��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$������C�u�e9Eb�����@��Ώ�C�LV���_$�﹪d�f�λI��U�'�E����_d�[�'z��dxh��o5��I����>.��p�����9���
���Ӽi��d��q"�eG����}5y�	$XӀ��1)��GUt�d`dp�3��s��;¶��NRnz[�<�/�>�2�ƏfS�~��n��T6�~(�q %�9����%���Xw~�J/�R�*��u3c��y[�O����3bEDh$Sk�RAGo��{�|.���Њ�"�!Tv+T&�f� �or��}2��L��"���B,h�>����
�xZ=,L�Dp��>��f�6�l���D�KǺf'c	�-�ŒҬ��A�-k� �����ݓ�ГD;�7[���)�l���CA�T?��_&8�>0Q����V�	��`M�j_5Xdah��i��{}�b��\�ms�����<b�8����*o���ҒN<�f��-�"t��x'�#�I\<>�Io��Q��5�����m]���+;�r�(��w����fd�׫K���ch�Q4 ����?�ɉK�����8�ΪW!<L��l.����;� �;���3�CHP������nͽ�D�"�4����̬�)�
Lm�=�G���n���%Dq_[��8��.Rʧ���"�|�&��]� �[Z�XVo����#�cT[�;���Q�r�M@K�%NE���q}K�A�^�e\����NU�C �!�\;#���_wh���e��l�B���J��=�r�	Y#J(�9[��X�8)���/�7
VS������W0^��I��r���g�%�</�J�#����C��;=��6s[]Ԋ�O�j��3��n��zً�Z��HEs� ��9c?	bէ��	xFA3�t�%:)_8�����GpE����@� �����%������J���2�t�E���]2�������kR�5( �;�>��|tt�z���"�8M�����#F��m*<M[ �n�E��w�.(��ʕL�w1r�"�~��p��Y���V��pT�a'���C�d��f����O9ҷ�pfˍ�7O���`4��̄�R�(.Z)�kaUJ��
��=z[��|��#6V����68�]��ɹ�$��m��x)sP��=i�+�٬ƥ�D[��zı��)/�n�5���L�����<�)�����.gS�]�cbh�g�-lH7�͎�ֲ��O۟����u�-��:�W��9�)����%s4����b���aW����L?�����{R��������E\,�D%N�j���}�T�D�z�Eྂ�-�N��Tɜ���i� #pI1��~GE�m���&?&r��A�\Kڐ�@�5V�VUW��+��60��^��җ�I�T��C�'�ٳ�	@+0��0�`-P3�K8���s֝JK^�g�'�R6�H�Olr�@��n�AMr�󠊦�䧁���n�n�q�~桜��LoZ~W��\��?ځ$�d.�XE4E�+���j��Eu\���s]I�JW��e6���K�l�~I˲G�+y��Q�G�Dy��$��J�wi�l����!:�x �J�?�o�X�@�E�h?�g�U����"�U/�eN���u��VL`fq�����<=A��M�S�LO���<�D����#A���v�L�Q�������Osb/�q��'K�桌2\�n��#��:Ƕ��Q�94�+�a�jU��a�&���?+Y�*�}C���c1���*('�}|�T�d�7[�`.�5?��t0����B��%�6�ݜ��Y��o*D��" �S�]ݗ��S"�K璓�TqѢ�I�%b��,&��KN���F3���8r�b�4��&Va���@m�j����C�`g"��[#��1y�S,N�bW[����+b��]Z�0��d�kp�ȁ{��Q�c�v&�~�sm�������dAiǅhT6�WG��{���ΚnG|��pn����A��V
��ѱ� ;����LF|�6��>���g�i2ޚ�L��"�����SI��1#�q���3�n�ZT�w�?ȡ+�D񤻏��qN��־e;���LSF�Y����	����=G���t�Y�m(B�L�d.���|�ܳ�s���a �q~��dhs�����9�W��Z�[������!a�T���O��LE$ф*�b�1tv���{tK:�{�C"_??|�E޻dS"M+VR-�d��v�$��h�\#�#��Na�`�+���%�c��N=�
M���(��"���<�><��4��;�q�og�I��ÙOG3��^&��2$]�B"���Ѐ�	 7�ZP����sM����X��GIRƖXX�<2��?�}����֜Lk6Á���`�W_�"��y�X��_*�g��$Gt�A\��������%�!D�;Z�H���{G?� �;($����.^r~;�O����з���^����w�6���^p��h����'뷝�6,���1M�w,t�:Q;�&�Ns��@Z�,��kkj�?���	q8��#=c�>r9��1��z�~n�/af}Ӱa���8,�����E��꼡19F8��V9Ɍͫ��v@qq	������"Ӱ0&��/' Z�@�۫W>	c��hi1"��hœ
0��E����#f��;��凥�9S�b�f�9V���Q2���#N��|N8�Y]%�;�^�,;T���rglA�C�k��N�&\d�`�h������ �-����:�&�L�����M�_L��e&��7Z��wuU�7�hE��Z2m ���|@�>�jF�--��NT���m�h<�b9)Gj/���V���ja/��
��5����ex��HG�	�f&�����I�p=g<��T�1li�0�_c�+�R5�r`�`_	�ρ�[W�C��P�˒�AL΍�7�w-˓��m��Sz�L�KI(i�a�?�������I���,�dv��p����<~ _0Ʋ7P�O���H#�9�+��Pȗͤ�$��ɒ��'��.~{��5' ���,Uן�!R�*X�{�i�o9��J�\(3c<"i��\
lWhU���s	-�I�<��C2	�n�)�'bA���FYexF��K�=��m�2M�����AQ/����"+z���A��R��JH T��o��YK��O,>�y�}������¢l���o��`�}	�Xv��$�dE���aiV���vo�����Z��X�~$�⮝�� ��s�p� �����<����Ƒ5R�06A�����!��f�טm���V�X��9����Z�޶AԪ9>q���D#�/�g��ߪd�d���G��5�"���Z'� ��'���")�5��[r�AY
��,������E���<i���$��l��8����3�l�@Y�'H�}����Nc�LC*!X$�В���!F@�V���u��4��ˢR��:=�����7�i6�O�C�*aݴ�&����Y�_G���J���=��i��zQ���8�5�X+�����. 6k2W�2���������=2�phA���DJ͒�3lr���K�&D1.�0k�3�; �7$QɈcʜ�䟐yhQ���
N炟�؜,�[��ڈ�[�GC��c���0X�
�sS��v��X�$H$��O|e#���I�����hGB*
�{�Ҁ!����r�<�0�zS��-9h���񏜼��I�~ShH��f��<YV���Ԃ���?N`�N�D�zU�ϙ��,���h�t��>��2s�J�9�`#���(�nkP��GpH�F�Kv�&O�ҡ'L{@	,I��T4���9x�
%�)�`���Q��F%!��+pA�`�߸ba]�/��.0;ƾ13���A��z��\�.����p�	�)�ZO<X@I@SR���s֞����#�?�e! ˳��_KD���T�J�b5����u�5WTd%�{��w���U�Xa\�{���/�8g?������q��i�lC�Z��DyE�ZnQc��b�D��VQ_�`]V����sD�&+:Cu[r`7Oܳ�ʹ9���:+��~�1{�"�(��Epȅ�=���[��6�Q�& :�
��H���� �����ׁ�-E�Yع�V�JB�o�n��n�_eĐ���zV��]�ؾ���V�p��l�Im�g����g@��?�;���)�d܉u
Un*�'�'���yq��V9ؿ����#@�:��W�,I�wN���D­�,%�j|UCƏ�G�+k9�X�������$w�.�9��1��'�G�Ch��--�"eب����Mܳ�g~|�p� ���Ň�}��V��	��`xGUV�=vpi�$��#OM#�)���P72��4���UX2����A����2���~��w�6T֪�g}��-��G�u'p���+�^u��Ik��r%�e�y��+�œ�@ٶ��
�|���$�o2I!�z�j���o/	�Q�ӏtԲ�*�3�R$�L�Fo��`_Ⓧ��d�㤼�[�B�//�BJ��_�;�Sc�r�������N��k7RW?3o�����@*�D�����~�3k��|��K�؆��
�)E�Y�G�|��i���<�g�}��ݦJ����;�<���׬.v�j�(��S�bG5������V���"�/4�*���db��d��_տ�a�g�O��鋼�d=gG�(�a�%�̹.m�tQrQE}2�l�L���| �G���X�V�n��N�Zԋoi��,`�.��+�~.�礏��z�9�]�3r�+��d�@ɀ͘�¶A!,��,S��$�>}N�=eSS[��ޢ��
�IB韞�	���.��"�w'��?$�#,�2���uqt���ժ<��s�2�9�ݍ����f*2�F� �>���EC�+p��=�k��sVLk=H�<�M}8U���*L�
d�#?5#��?��b���g�Z>i�#?A�����aI���qQ ���图e�B�έM���Hp����[�pPkv8<�/����˰
��Lrl��l���H7+�у�V��.8I�a�G��|R4��ע���l3c�o� 2<�ݥGw��J����0���ĳ��@������4�5r��ˇ��*w������b0���{ړ���Ap�xO"�B@y�1�9v>�pz�����E�e�"�m���y6�7�a��PK� ��æ��P��ð��n ٍo��A����T��F�1cl3�N���#�K{�]~Bx��˛#*�Ҟz���'�zڬ�-Ҫl�Oϡ�R�~�~�1K2-�)o+N/�$�"2%P��O)_���ɛ����4d�_Dt`������H���I|���������m��~6&��uHh�
	��{R��t/�&�	���K��pNjgTi�Q�C����|�8h����0�fRg��.ekU�p��%7���Cܢ"z�u����v��	\�v=�����p+v�X��O0I�܍,)��{1�)3>���ɠK�&]�:�hҾ�}�x�����٧�e5�ٽ���A���m�--~��jl����f�����M��/+�kT�d�3T����\
�R���H�h/IK��
<Ō�^��;�,��]f�g���0/2?-;SI+0G���/�	&�m~,��DSQq�F�uԡ%P��E�Cm����/�b�.�:%D�؊��JS>�Q�����ͅA�bq�ȁpS�i�1�hޭw�M�ᣵ��C̬W��S�_����nz�1u8��}�����M���0l�&���E3"���7`�ar�H�v�J�jn<���f	4���i�w������h��|[{�0���9�D2c���g:"�>����H�>�>�@8c�D�W>X&2�%|���Ӈݰq�.�3�܊m[�X'�dz�M|��ԞF�4��<!"���1J���������V�S�Չ}[r ��P�\F��-�l���m���)�M���SAxT���
��f3<�����l�0	�ݏeK��>��>W��u�c,����6BMS�-Jp�UAU% l����<���~Pi��ϱq���	KyeP����O)

SO��A�!����	�%=�U�|A�3����� a�s!��0*IC##ͱ
�Y��v.��2���$���4>�����ż���y��,�>����C�{rJ��i��b���Lfo���)\�O���ф�����t# t�򐊲��@�����&s�W�1�F]ٿwKw�'{F��ai���F����M�aPT�FJ��M
�;ß�n�r̱&�m>8#a�0r!��&���X���Z�Sd	�i���I�w(9t�!��cT^�|Py�m)�[a�E�儹9����1�Uj�S�=�?�v*r��c�U��r�Y2�%����	fa��W�\��l4D軘3�ڕ�8OT�x؎R�,�=�tcO��QG�k����I0���T�p�������nRs�������E+����aM8�F5�6|�� =�`��;�����im��� ݽ��ɥ�9w$��UQ�g=�"7�O\VCM
��?�'��X��(xE���]8�x�=I�0��5��^�Fۡ�Q�9H��/[�H��'�Xvi�]j��;Z�`��k��������\�Q32�j;?J���<�$0�`�!�����τת���h�tH�^��g_��3��?�
��յ@�26�_h����������-�[� 颓���2o�ޛn!�+u��]��kͨxe�>� ,�-]�.k�*�JF5)x���WEb � ׫0\w�#�T�[�ɏ���%JK&�Zw�6e%|W�����\�[m��F�����uce�*�Xs�Y�=5�!�Y����F&�;O�My[hhD��)z�I��������7�?~!^+�;�2�@~'��sa�����L�ӑaH��J����}�K���t2�e��Uq{M+�kyES|���8��ߪz�ԉ��y�,�a�>�.H+x%�)@�����k����U��]�{���;|@ͤ����{��@��KԔIq�o���;&D��=`�;�<��OK�<��5t`��U���9��~��_j�8�����V�����"lb�4�	�.�,c2��!~Z��K� EzIS{q�ҿ�����jY��s��_��*}@�mL���TM�9{o�g��E@L j�ҳz���`!o�5+�y�*� ���?^f�V[��ԛ��
���b��Dt�K�@�T�0�f�_���֙��st�Jf#�5����e��r�QH��)>�N̓N��в�P���DK�������{�{H�Q z���[��E�LC�GW��=e��H�%�a��k��E��X;L�)�;�=eUb&o�s���f/��V^~	�~9�N�����V.���GJaQUz�K4�s��Xr�~Z3D����N3W/F�}S{T�n����d��cr����4:��5��"R����]��q�&q��ˎ�eȡ�k�d~�����>8�+(1������͕ߏa<���;N&V�m����Ɂg�tܒ�u8`�ݖ,��(�c47�o�<�@X�����D'P�1���Mn��Y���/�stQ�dV^;6L�/J����[�mJI$�������fF��%P�����n�.#Y�3X�aZ�s�Mz�d���V!���G�Q�w6�H�1^�B�S�¹�M�������8��U�n�b*ӡ�+��g#ܞ��+O0"Ƴ�_wd���mU���5�2�o�T��s�q�DO��R���a��(Y�IU
\�,���@M���ӄ�k[S���Q���)����$PDb��Zqq�r������Z�|�������>c;�ѓj���P~6U�ÛF����?�����g��� ��)��ء9S�H�)�tj�x�f��$h[�18�m�3���7�rc;�Im5d�1� ��P��=��qzڃ}l�!���1�o~<��nM��gf��G}5v����YȝeULl�J�7���Ll%�	�l�QI��E�00��_d���'�.K�9���)W�D �M�Xj��Qۑ	� �3�z*��7$݊�hni�a�v#��+Qߠin��M�:�iLn���j ̔a����o�tGxZ�9<