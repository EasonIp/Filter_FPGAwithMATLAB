��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0��`q�M�'���2&��Ȯ�W�4��д��|�6�K!b�'mY�`��L����TR���x*5D~8��VP����i�ҭ�������Z�F h�1(om�?9�x%<O��=��F���3�a����_��l٧@�S�B7��K��ܙl�0�o��n�l��~�ڕs�u�����V���HG�Z����TD��6IC��W2@����86��ӂ��j�˴���S9�иK�|!�fg�Ѱ"iJ��S�4Uc\�:�H=���bGE�b�#����Q�n�T�0=���X.���v�+n�Pr�u�鍡��6��{h<�o�(��4�$���^�ߘ�21�˩����W�����o,��[��GW�H�hF�#��B�xh��U�� �d�e���=�+�bk\|Kc4���N����};N��{�1�}�+o/4g��wή��4B;4!�c�OP ]�e<ϔ��a�+|�{,���H��1�����6z-g;[����T�q�s2XP\�+���Mx"'�@�[��?I�;< <Ҭ��z���8��=;8)������|����2N���n}��;@�d��&r,׹����;��N�K�Q@W4�W���E��iv$ʁ�?������'�R�ם�I��in⸂�@�pɜ\�v�Ndqꐋo=iYF��˸Xo��Qa��v����"��>C�<�+�?�3	�9u⧐�T�0t��\d�1O	[qE�{��(�ݟ��!K��[׮���T)�].���� )wyy?��]�9t0p�ƻX3c��qf��:Q����݆I��b~:Ȑ[W��Ck7d���af��QZ��J���<�&§��W�������oPT���`�_�^ىr��J��fX�0��qX*%���XB̽���q�k�p6�Q1c�i0����'���I*��:��Y%�o8�����	͂SY��`({�ݺߡ�?�}����7W`��&��r�}���(5pɵY �����[7$��3L��G�|ҵ�A���Z�Ӥ�]�E�ǒL��4��J�tV�vN�W�s=��]��x�J�5���$#@ǃj���������㬐���ط�����Xn٨./0�q(qY�>�ʲ���Ό��ĸ���M��ih��m��2����[�0��(,�"]J�`�ɿ�ƌ)<jK����7ˎ�����h���������'Խ����T��6��V�ྦ�Cty�V/�����:�-��2��@Ea�� o��I^z?l�x�NtV �K<Xu���x��y���*5�Q�T,op/)�OHv��Tͦ=y�i|y�ٟ���t[�j_7�*{lq�9~��ʎD�#�~@���d�ѐ�]<�P���Ý&�c:F�Aw�@͒u^��_���E°ƽ���$�t1�Z+M�F�36��� >ٴ��P./�݈
��G�H��_[h�oꏻ]ň�k�g; �(����'�5,#�BE��Z;��t�<�����F�m0�L��pო�;�����b�f8*W�@X|oH"> /�G�&�'����r�}�����|���X��[;x����x!���Y��O/��!�����&ķ�i^alїh]Rz�\�Q) ��R�?�����﬉0wդq�3iǂ��%g���Q���	E6�&�0`�!�6*'2��հ�E����k���{�NeX͐�/�c�����2R��Z5u�6��2�5�dp/�{4��&+`�L�X:!x��K(AԆ-��4�K/�6�KF��B��z5)��R����q�G�?���%Ar���R�.��	w��5�AJ��3��S��n��w`�y3C�D|r��L�ڸ���`e��$�@Yܦ��zO]�,�^�ڈmYr���"�:��M4e-S{)�k�xm��0�[]H�[pϫ$��35��N��׉qF,���tjo�A���I�����ɐ;��
���߿]�Y-Iu�A��y��-&�7|8�}�tY��`f���;�,7�#ŧ��%��+��{��.��3`@����⋱����p|�^:Z�|���%/!��&S(�*	��9]R����E�����Ef�d������0L��h!4�:.!����CN�`�A�$�a֙��Fff�$���$%�ވ�t������L��_+$O�χf�8��n����I��s�[��Q�����X��a��Ī
/+7CPx���(��9*�4P���3x$zZi(y�F1�cYF�s��*���'��J\��ui�2�W0~����«:�c8D �2� /I;
�w%�`�H�i\ȉts���m��(��}�oT�V��E������(K�С^��@���M��у��-���!'�f������ԗ�]ke��O�`o�#�nkV�N3�怏:ـV�1�]�.�Ɏ ?��L �F��vqZ�b���Z��-�L��P����:N�n���
�PF.��T,��nS�F�ڿ4$d�M4>�r�I �3�8��]+�mX�F�I��"�X3��T2���( A�H�ִɭ�<��U���q������F7*�}0�b>��Ah�\��O�d�y�����>TVQy(�b�Ĕ���z%B�������H�����/n�pj'��1[�/��R���3��� �Q��P#�
<��$�;T�1�	���ݱ�1���~�^P����5f���U�a��'�k$�t�1�6W+�_�+c�J��Z���.1�'�ܐժb�S�̈]:],��o����H�R�V�]G��-�=n��Y�"{��֥<�*�){���eSt���b��R�L#���9AJ3�v�Թ;I�3Ǧ�ǌ��a�f���Au�4.��m���L�$���y�3�9N��Y`|}$򔙶GDN5r����0xb{�
�#�>7��@]fu�ge���S)4#-������9Jum�C�DGu��W���0*Em�\2��nU2�Ƕ�n��"v�آq�psZs��?J��^}k�K�{�ɖK���I�mh�����W��]�c#��cS_X�Q�Oބ�&M��;�64��Ad�~Ω���wr����O�B�͇,cZyv��
=o�2\����=_&����ڒ&°(B��i�:2ċ̴L`j\�`�����lW� ��rZ�����#����0+���I����F��_" =@ED]��gV� ��諃� &��=�����f�
4�x��l܍	S1A��.#�b6��H;��b�D��rP9X����?���,�0��!?�Suw�Ob�pTF���QN��;8�Xz���GJ�ȜIȓ��J�"&g���A����Wj��T�DǇ2�Ѻ�.q������&n���_;�Js�Hd�z���&T%�>�O��&����`��� ���߬s*�`����`C�BVE�.��R!�Y,\�ҤK�[��S�����ʀ[�`�� 1��Ga,@1BNU��8���M�g��F���"�}���~=radX��}�I�� �xjѲۄ�	�.�0ux^=G�;�}��q
�|�'��+be^1��E�чm���7��R�O(���{�B�nr�'3Z� ,�l���й�\Ψ�hNWV�Pn����
�qN�.��w����R:��2�4�P������uy��=VD.:�z.���K5�D|-
Ɯ�v�r|���إ-�~'�pà���ȉUó��%J�̤Cm�8D���%�8u�a���yb@�?��Xc��"�|��4?�ux�3@�l:�%��~>}Ҿ������{|r�B&��A�"��7<O,�Q;�s9G�о@�~`Ʌ�(�@�UO���9I��0>������p��Q�Sl��o$������o���~��u���.�Tm��DG�@	��$[n�T��g�Ӂ����B��7����^)X�v@����B����[��5�>�$��?��y�2��7V����Yܑ,���v����RO���e���ʗ l���Ǔ�:9Yۤ�n��z ,7Ո��>�B�I\�*o�QO'�
s3�ʲ���v(ܦ2��gӇ�~��̉�5 ����i�p7��l�A���#�
5D��=LXk��+�~j׻��^���óIR�,�a�t�d��l����C�0�N�W�`dc=���~���
p��-�pv���Z�ޠ��|-Xeަ�A4"di�O}��dg�*x+=+�@ٔLx0���`Ġf}�8r��{M�j`���%CLn]5^<��<� �ѫ�5F���2I��?��&�l�{�TsJ�,:N��x��ϧ.��8)����\�N$ˀ���k�
ʷ�(U57�C�=�o�LG��,��_���ȔY�QDA�ö$����tGL�:?$���1�:��B��N2G�A_PcL�K�@>^�y���i�=y��m��[�Kr`��p�J��T�R�3�Dڰ��g����Z���4-N�c�������+g���`s�3A���n�+"�Hy��}��-@,߂R@��#qS]Vp;佉u�Ǘ�ꇬg�nU�U����g�T�zj��Φ��tx��z�m4{��]6�q�����b������/\�ޒ��<
+��S�%��29Ii��yxJ�ewn�G"���5�)��@Y@��B���a"Al�;13�/��4����� ���� ��G#�Ke��痧��6D`��%�g�RM��feզ��X�O�}�)FY�t5�� �x��1�$�%i�F���܇c�3c�k
���̄���E�CM��S,1�#{��C�C�u	��=@����	;�Ut:�ס5l ��?C��֓J !�Ar�{L�����k f�R4������[�`� �h��4��+�I����9�m��I酻�;G�б8��-���6�Ey�k3�	�,��/��a�\�d�sJX�m����H�A�r���t6Uވ������˭�����d N.KEF��;D��v���Db�=�Cϕuԛ�H���3w�w-l��J�X�"7��5t�]�H��=3����1LE�&��������Aʰ��Zr����*�u�'�E���ix�Hz��/7����ݨ�Y�,��F��!���(�>I�	�	��8�1���]3	�2r����ބv��heʕ�y�|��?jx����=`8�=B/ߎ�[�@�o�k�GuJ$�Hl;ﷸ���� *�Rk�@�Z�ZMI�g81єio�H��-�g�{�s�_0t�CG��!&+��,@ѡξ���1YIV�
ؚ��W����\E��q�߅l��6�|�d�1��&z3�A�,�׮+���P�08�iχC�j��|re�R�w<�t,<l����^��J�d��sA���]��p�����jZ��
dxv�]Vp2J���#x��R�A?�Ss�U�Q.�&�$�X)+���I�4��E�<��,{�y��q����:���ƈ7Q��ؾ����������C�J����H�;4�5��j�*���{ek�4	:���О�ݟ�M�mnp��)��RcNr�]��<����`)k�폸|��{o>��d�'��*g��AΆ�,tF�P�w��zF&�E#��y[�6�?��(�g6X�롗�q�CQ�>Jˮ)WOaq����K��v��	�<�o��7h�
�xr8���r_|��[��I�D6H
�a�<��P�u��+�u DzB��J�x�M���}>Md�ࢬ��Yk��d���Q���uư�y\��6q*SW�\��������+ 	�⃛$�s*jQZ\d��)��Ks>�t����w;|�Q��-w�g��ha�,q�����i ��	����OHo!g0$� >���B@qx�h�h��R��3g��F}M��X�X/=l��T��Z/NE��XAMQ緟S^����nσ����AO�2�C�R�V�a�薖�	���#ސWFG4�������dƆ�g�嘁[�����E�^�]᭠6��!t0A�l�,���󊐣*�c}@!]��2�"� '������)P�u�I7Xa� @���@�I�}��ʩ�;������)�ZX�'��{k����ο��F�opC�wv�J�I��H�8�wq��v+H��/u��6\\�;@�猏��M��~
�d��Ŕ�?w�|���a�y�"�,�y��!�fUWs�
�;�N���"��7l��JY�F��n� zH��dU��G��t�4f{E��kޞV�3�$D䟘��k���C�����L��2�i�N�ƽ�os���Ԋ`=���Vs����kR�