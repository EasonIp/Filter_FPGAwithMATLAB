��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$�ʿ����Yo���n�y�2���l�(�GE�$t��tG��U+��n�o�ע��%fVC&�^~���=���I��Q�A��(Vd��g,�y!�UlrV�(FI~�9ao�D���I�u���*S��G湹=��g�	�ĝC�����\sy���ն�^u���^�.�"Y�Ť�V���̙����3����㜄���C�VY{�!��t�
�</�gC��]��N�[z�㿗tt�W;y�JM�a���1^�R�d���^�Tۻ����!��>�4�'l?+&Y������� �܁I�������1�ԓ� *��;7_U"2�܅p�e�^Q���'�OG��t�x�q�|蚧/�XV1|+7g�B�qk�#6K	A_���;���I�o\M��Kp]��}Z�o��"B1�JB*��R�Ŧj����VDأ=}�����MS�2��DP��|�y$�W�oc?��+8t���+(����t���?��b|u.r�	��!=�.�����=(�)�չ�����1+aKM��n3�:R�۳�%��a�p�$�P��@��7���U���U��ݠ��4XΪPI���0��[�L�π��Kp �/6���%�iέ�º��L�Yס�ϧ�T�V��C����$���"���ַ�*��~�r�u�K�{�:Ѫ"Rh�k'j&I',t� ��S#p�i9����;��	k�h�i�2���]ea<�r�\z��/`���I1�J�Bp��0�}O�NBb�n"�n�I�Ώ:{���7^�笠�8�� ];.�Si�U�,�`O�}"�D�]�-����mߣ>�"�]Sl��e�Y�e��}�2��n�Og��O���-aigF���Tr)���u��7���Q{S��>?-~k��5��0=Fþ/��ؓ�4K���@Ku�A����ɩ����;Zc�3EAyd�R��y��ܨ���͋[��l����l����h-�����Ok�Y:(9]����:�q���#�Xct,��Q)_��m��Hc�2��PC�jh�~�qNI-��{��Q}���jG>��f�zh�+�.z�DÊO����5��Cp�`�5�4��pBL�>m���<Z�'�W���R|�K���H'��!�t��ч��x �.	�sO��aB.�3ӷ5,����i���������fX�y�ã�4�ux�%'�ۇ�����}.�'-�qjR��o��i3�O8<f����5���Ykpӣ=�R�峯(��+֩>v1HLt�.��&c�O|/O��?Ao�"�:*�?���Q����V�Ԑ�y������ڥĜ{���]p��&
�js��|�Ȫ�\����J���]��x�3$5n��K� d,t�7<�w=�;���A:��"�Q�v9�������NH"uX����Ka��d~ ��0\�Y�.�S.���o�T������o oE�Eg��� oE1s�F��;i:+ ��T��
���	3;X\&\D�!FJ��}��L&����U�qŎn�;�vɾL%jso�A��l�D�kkܘW�]�%f�ҳ�}S!����<vXf ��Hӈ�l)%ﰧ�5��g�T�;ds��wiJp�~	��OU'10�}����Y9#c�������=�$C����&1�xjO�&�J������KD���� ���Q-A��e�I��'˨��D�EOpZ��d�X�pv<k^J�(~���͟>�}�����A)j�{<���'	����z�n�����N�ʊ~)Y�I���$�T�`�v�b�����^NV�|���Qj�EXq��+F^J��0Y��D�j�	����Ş���f}��#2];x�i��t�Tn>�/b2�U*�g���Ś�Y�r���q_!�j9���7=��T�i	T�ozi�+3fL���l�������B���TG{��lE�%3Ȫw8�#���U���Uz�ѵ���5��`�O)��|��/�r����e�NV�����3�]$��񬓻q�|�b� �h;U��5�n���j��1G���=�..� �{����+n�6Ý����� �� .�Y^�	-VG���@�[#�%9�^���f�9��@�J�)(sV�Q&2�s�b�`���fN��7'xS�kw�_�ތ��OW��BN�8k�\=j	�8٘�$hcU�:��g�t�JgQ��&tH�����&�f��?1U���n���ZB1����O����^��,�J����K����o0����쿌�U�˩�d��h���
k��92�|ٗ;|��֖�I	��0�1u�����Wg-��3�=]��H �#Y�5|�N���9�
4�Nq�����ϼ�^@�ZώC���X�0�Ƌ ���ὤ#��S���қW��?��?^�ǎ��ic�����>Q�3]U��/���ȍ4���Ew����Ⳃ�(c�(v�^j��T�2o�#)�ew\��by�u������ ��R-�઴�|�H�Xo�W�w���)p�8t��氫��!&���H��-�	Ĳ8�5���S�s+7�X�Õ��6�5���z�߁�n���OV+i���!X{!�t��c��ۍ^_�BQ�Y(A3%yP_�|���(����8��Fȅ�,���@�<1��#�-o~���x����
� ��xR�t����6/�O`�0A/87
��a�1�ȶ��lr����M�}����X�X�/9���&�W�v��k
~7����7�C���1�����G����8���'�B�3b�V3�;B���1-d�+��,��4��u�-�p(��	���c�\e�s,�d�YCA�a�b���2�e�׼6��]��̆�F�Ҍ��;G]�
�]G����Tt>�rM-��E�:�|���o�QfuM�L�kKVU�K��b,��c�|Q��YN�ILRB,�Vh�Ȃ�S�#P��P��&iV��Ԙ���J9���X�>�'�<~?)D��F͈��	�	�uVi}^�.����~���Q�����`��ŕEoF�q*�u����P�`��x���`:���/~&@�_��/��K�� ��%$�=dk��v��jB��2���͓�f��y�L����~�1�w(rx��[���5үs�R���JpA��@��f�r��v\�L�6ƚu͂���I[׀�	L�x�-!il���
���\�S���IE��Y�Y	�M�@>y��!T��e���sQ��!b[Z[����d�2��s����T4q��Tt�g��a�W��.�n�W�9�%�k�>��AG#�'ow�u�V���[&D�H�D$��)�.7���(w���V;�|��ٔ��{c3qf�紝H�yXrK����LIHΜ!L2d|C�ϸ֬�)"Nw�V���Ђz'6�D����3�,�|��ܲ�q0�i'x�6���}WI����{l�ڞ(���қ�{X�]��Ѷ^V���?|X癎;(�����@�o�����^����)��"�w���یd��ɋX'ʷ�o�'� ��P�" 0��Y��%���S�,����!B	
@��+C�j�Wnh�ܵ�(�m(���[�ߟ�"P*���j����]���Ʌ�/�T�ՙ��6���X��B[�]�0+�<�0�/���~z݌���i�9.ӆ�sÚ�D�E�/����������x���X�=���:^�Mqvz\���N������3d�D�z�����t����	 8��O�<�e:!O�,���-��~aʌ,�=�zlq��4������/��"���e��J�*E����9�������Z�K��H��CWE�;J��J�7��X�G�Q^�4��L�:������97�z~{����o�nI<4�ҸՄ��)=%t�]*��LZ��ܟ͵:�6�h��m����O�L��L�2TpI��UX#nC`$�
Ɩm�Ťj�񠹵#�Oh�fi)d�9��	�f�;��<F@)LSnh���#;(ο,�w����U�kc�z#�e���)$�*4 ̀+��;�c�_�u��s�u"l�s�~��nz�w�
����X�4�%��ن�V����G��+w��@)J��K}{��m�V�d��n�4d�]v��!F���qZ�#�;>�P�|���T�m9gK�Î��!�I0���28`KX�L�#�N �lF�@<�2i�=C�U5q�䉶l�o��)��R�XLY��`ߢw�� XP�Cw�c �놸k�n��ꢨ�5����;�9��U�YD7���9�ޏ�1�v������>f�V�k�L����(}:��y�˵�XGȸ�8X2��P!�Qw���/Y����oK ����Ȉ}��Կz��i;F���X����!2H�P:-BG���$��0;���r�w����A����sqw���n��P�b �-	V��ü�Ӈ�-�O��6pF��Ipd�A��pWz�@�?Y�n}���Dv��x�� ����O:"B���_M�+q� i��a*��o�U�p���CλrA5<��:?I��h�m�&��-���5�pf�7A¦t�kP��/�H��0��5&(�]n=��Zy�L�nv��SN����/��Y�Qx������#*��v����]����׆��60ϋ=��)*�#�8��Vh���o�������V�5
�k����L^��=&hT�r�2�n�r�8��.���1����w��u��W�~a�"zt�i.�L32�>i{�U�~��uW�q7r�~m(yR�d��Ȩ���3�|L�Bu�P���{��;�	Ǧ�ne��)1b8�{-�����C��{_����=�N,G�!�@�-�>�"�L����>Ϫ2�~����]Y�&��:+����LUA0�m_.�g�|F���<C5���]u��+-a\��V����z�*,��5�Du�� ����L�����ʶ���Q��*ef�8]=���ǗV!�GI�o�:��f������t����hDc.i
cBW��9)����b+�b/��m�3^��Sƶ��R
�:_+aV39�ڏn�V�lj�(/RbGR�kL���d?�����?�����m��Ўt����2�����HT�q{�;�J�i`:�5޺D3{�s:W�p�F��R��0���9 �����$Oo�k)�9)}�ܐ4ΛT|'�̮�,mRҮi�W��`�f�t�?0]�(8���EQ�҉��*��c�vl+#zΓ����!/f/V��(�EAo_�7�%��<R�ItPL+9��lp�:sy���17@��T�X\�p�(K��pBj���0ł�L(Jd��E��_u��>be��i7	�iP�r��Ʋ;�����<0�űh�ʀ�&J�������V.�Z��T����!�&��9��%�������_��,3h���Q��c���ϥ������\7�$�|o ��.t�s�30��;͗�_y�
w�&-��1��N���b�K�w�_�O>��������3��>��c�ʞ��䂢�075[�-e�z�8x�0��x����[�������O�7~�� �4����h� D���m
z���Vo[�W�z�MR>_��׫�@:b����m�؆&9���By<����碡�������y�0�K_�:���jW2��t���R�$@�"���?���ĵ�l3��c�ϩ��v���]�)r*K1��9�I(�=T\�=�*��I�,����Aw]��"��A"�n���.�>?!�PA��)��~�`���m�\� 4�v5�(K��V4n���P	
��+k���/�v_�`�?x�T��v<�v%�vu��Ӹd�mF�<~*���@��ǃ�%�ҷ�.����P�@#���m5*e��{���3-�
6{aׁ�$�{�
hI]�L�?oB��S��>��7ˌ���s��
V��N��'���&�|���P��2E ��z|��s��C��o�g��QxMI��,��9�DL�~_K��Jr��e��~��(��g��kCr�-qAc��4+���RK<Q+3��>c֥@�A��*M���w��.`���^Al��J	P�*= V� ��Y��0�3o^�������ќ��u:7���H"�@-���8<��\��)�_���r�	�|t
G
��ؚ '�mt��{���E� ,Z��e�dI�/c�t%X��gޏ�g@���N��S�cA�L,U)A�����DtV���GN��� rQ��r��E�#X����։~�B�oᠣD�x+���b��]�ɚC���>]N�dԇ���K�(�'F�z�����50�d��<:�F׫a���W%���Be�E�M�߶���� �F�����ik�(]*r���(L�D�bR�@$07P��YzL���y�jڸmїD�Yg���!�W�S�;To��tp���C"=,�X�bA{�r�����A�4"%9�M�j}�[k���N���Mh5�`�޴����'$���� ��p�?#y�o>w_�����Dah=�=��!�@l̲0[� cF��N���)����1�(�7W���s>~�[C���mj35�U�i�9a�u~��Q M!!���ѷ+�[hs�ٔ=!�Z5*{�`e� ���:�r&F*�&l)$`5]��H�n낁�'M\&+�3TFK$��E���{XZ5��9$m#c\��ߴo:����L�޻5���8(�Y�V56	R-� �YV�S\n����ċ�~�H7_R�?1!��<�<�9�r�niEx#�W��Q�U�����i\
�=q��l��b�Y!�e<���5L��rJ'��;MS���5�d�/�QیN�(L}e�F����&�1��D�������6��������ω/<�����ݯj�/w.7@(�O�-����!1=ކ�&��Pͦ�n�y<�N�^�`��c~�!iZ���~�iB���9�5}�x%ϥߋ�:�o~������U�٘܉hH�P�`���>�FX��%h��v(k
���_�V��DBDk�k5?��&����5�3�)ܪnʣ�T�u"�1')�)o����&v�SX��>@�4��rHT���$��;ͳ�)�"NK��'��Zz��Yɂz(Y-��>�M�Q/4���3NN��z��g���*���;e����:Nk�~��:�����<E�*�W�;�|���s��[��q�b.7�-��^iy �KB���r�y�:w��<�PI!=��py<=e�u1 q�H��m>�d�&�{�I�k�j��
�w:M�4J��Ѐ
٧��ͣ�/��K��o[�0��9T�Ֆ����CŚg��D�F�����Ĕ���&F���թ�es`���	�t> �X��m�VzM�\ � ���t�KA�i_�2����O�@�W�-��^Z�[M�M��Y�1��C�'T?9�$�b[��.�j36�-F�#8���Re �̠�0�E���\��=��D�d3��B
4F�RdQ��j�qx�^�V�K�L�\��f���P��b�JV�?|{���d7ÇA,
0$
{Z֚d��l����mB`Ye15�]�a�Pv/��]����ܿ~ ?0m�XFj���Ӵ�-n��?�GNu{`Oo�h�����k�[��oVyߢ��}g�ߋ��2
����Y�{�BV�xva�ҏ��~G�{/1DG�� cA�D?U��IU�#q[��xѢR���q����M�p���O:�8IV6��u����~z��H}���ڨ������ApEn�MX_��N��D�&jI�I9��Fn%qCj���M�_�����]�_щ��8��}��>�%i�����j�r�C�o�UnyJh��%����<"�/n�M���M��=����>��}!ٯ�*�1����E�<Hͷ�{z��e�tK�lՀ�֣�	̌�1!� ^e,�?���&��%�M���<�b�����(��ڧ�s#�Ws���x� ��sK)+Kdx4
DQ ���z�]� �:�l�w>��/3����$���ӌ0��]f�4��Io�>��sn��T��[�_U��Ĥ2�n�8��xT�?��`�b��c�>�Yŧu��	�/�G1���r}�[G��[}ϋ�9g���s#�#����$F�5�� N!߬���h���WO@�@:�Ʀ��k��N��T����%ܚ��e#����� �k�/����Qm2��*b�bWd��ӄ���f�6����0vz�7��ߙ/��
CΛ�ȩ�"�B�&���3X6�[�`戆���{��S+<	M�'���(��$-[_������sn�{�g�U�;7$�8�ד���YbQ�0:x`"�F��J/TW��׭�8�Rv�(�By��#?�&���P��@Q��dO4�E�%s�.2�!��8(e�ْሟZc�]2F�XҦ��Y��mz���m�\�����]E?���gU���?햕o+fvЧ�m� v��]�<<V���P�����?e��h�O#�f9��ԗ�Ǩ���%�;/+��6%�3�p�VSWh4T���{�V�<b��i�#M�t�ə��IZ!&T�i1��kO�H(�5�r�^<\IC�8���P�T�c�^�
�B*MT`Sv�|^�c&��K8F���WZ�Y�b*�&iwe��#��C������9�G���˼�G�0^�O�Cꭼ���]�b�}?)G��WO�y.n�{zw��-�2�r�����y8?�hK�y�	��%��m���tP�n�:>~������J�>;�����0h�D�����Kb�O��C�?�sL#�T�&Eaσ<��o5�1��<��e$�q���5��e ��<���<Q�9�y�9��1z�p
�A;5���Mf�cO0�ѵ �;��	o��<X��OV�����S�13s��7��� .`7�K�K+{�P�$���l�A�a&A�\<T�pa7*T�}60���u�~'���K[�/WqM�ت5��{�4�NO�XQ��Y�[p;̐��{BӶ���~����l0� '�HX����V�x��(��v-o�
J�[>O��PA��
13��> 8=az��z"�8]����:��f���Cl���u�I���7S����I�� �A�����W~����H&z~*q���9���(�	��M�A�:�%$��H�5�;ø�O&�\�	Y���l'M|WA\x(�S��|��j�/I�� �¿�q���-1���4��
�i�,������
�Pc��|�X	�>,3=�|���E_(�G�N�#�u�I�Mf�U5�:����S�?�*�uT�DE#�[�A�C�ڌ;"�.DU�Zsl�]Ǣ���8�2��"lT(:N7r���bR
|aR��tE����"�N.���/E�V%������[I�r���F���w����s&�c�O���Г�B���7c)%5m./�*Z�X���|/�̥��L�����:�fُ�d����ѝ@ѱ��W����c{�(C���e�a���fH���M=��X��xIz!����ULO�1rv��q����,9h;��Z5l#�n�
,O+x�OJ��^-	б�"�X��z!s�j5M���s�����u�ƶ��
���⬲5an�r��P��˾gC�����
��xF�f��G7ֶ8dFb�{��������`�a*����?9�}�6"@ӧG��H��/R�0K V�oד�l=ư�z3땶�dr���H��k0�y�������\x��%܃�e�Ml2A���ZǸk��N�*�#�Ɋ��<4]��=��y�٫����ե���k3���z����4����p���n9A�q���V�lx�)�BD����'�&�zͿ���L�F��&�����Ek3�06��5,���)�'jk����98=v��&/[s�t�pBG���H�l�A�Z�e�)o�b����/^��e(��ܓ@��ϑ��OJ��l�U'��0� �%�ڻ�̓2����h�ߞ"�k�w+y6����6iw�Ӌ��8P�Ӽ��,��":�lNJ�5'����{7���~����4�稘)��Yu�!�Y ��b%l8� A��V\`p;���-�s-�(M��<��8�E�a�͐��!Ƌ �Dʘ(���CV�#�_����a���?�{�Z��OD����)	��?�QQs7�{#�ĭ�r`��e�`z���$���R�>��F^d�}/��iI�����_9�e���>�?�� @Ǐ��s?�A�p�+��i7��NR����`�m�	��Tq����� ��u2��!�>�BTwvp�	U�!����1����E'�t��{ ���B�^N^O|"�BLS�5#B�=���@7�~Nz�e=�lc��"Հ(�@�gO�5@��6"��=���Cv�_ԝ:�l�Ψ�8S�Oƴg�	�ǯ�dʎ��*��?��k���I~�� 0q@��k����P������tG4����a_��$یYj(À�s$	���J���Ӄ0�Ҟ����?���O���ٌ}����E��\�}g���H=&�D���.oQ��&�uH�9�d�R1!��Kt72 9��p,��s���L�=Cvd��&��O�}�({.��'�l&;R��,�Ye�+�p����v	�LR������v�q�/>��0���N��
y,�T�F?߸�cj��,���
�Dw���[
���0@B?��n�_V��u�h��cM��in��o@Xj���2��Oŏ-)v3N�9���-�{�Y�g�Ҷo�D�ĵ�xl�T(Li�Q{2]��@{�8��@7S(u����z�[���(���6��5+��mY�`�ȸh��]���W)�(ȶ^�+P䏨�X�G��a�G�u�ک���}���D~�r�]���9��?w-[+��_�~%�=��"T�M���I�)CG-6#�^��FPKD�������W�c
H�{5'`�v@��X`Ö�'�Rd�<	���Y@��+��[O��88m�"����[�,^Y��maϝa��)4��:���i��X9�f�L��\v/�KRD�$C�V�H�u-mSS�����.	f�L�PX�S��}�V����aIB����������]� A�LUȮw���iӚ��a�/t��%�F�U
�	�'��ұ�_��-��QxD���t$��m�%KPFb����#�\7����0���\�R�ȸ:OZ򞱇Z�)E�+㹌�A�p�������X��C�bI�[a��O��N�E�l� �Gtu�ڼ�����^��f�U�ū��'�]�]+f��d^�dl@"�?g��]&��ƈ�da�z���e)�/l�>7�_̀
�����W�V4��'\�+0
�_���_�u��^@�����/1_�"J^����?�Zg��6�b����u���������MHBM���?����tF�h�X�LAx,���݉`������*��>�󘵿7�yz�X��⸇	��a"���� <s@m6
�gO��j��B�g�V?���b���5����N��"�.8��d�LYK��p�F����\�A�9��4i��ȅ*�ᤱ��1�ϳ?���e��ϫޑ��_Rz����������q�gM��b*<1,=e����?ǵa�}Ļ����ö�jE�Q '��v�q^�%�K��x�w�w|�t�HQT64�xoۚæ����J��˯l�����lM�郱�Y��������}U�?������I�䠘� /��(� Xe�/�{d �����fTw�Ϯ�J�&��Q)�l��5�` ��'�q�WO	p����b0�F@��grl3g�*�J`��~��b�%������2��íS�S��PZ�͌�|[��2h�t~����2hB�|��B�
ș���T�ZlPb������
<��_VE���D�;uj��P��Q�� ]L�?�OV孝��9�>Bϥ�� M��,%���c���<����H�gY�܁�?���+��p>�fT����)�@-X���:���(�(���u#K�h�@V�G�&{#��9$��D=�Q�2��l�<\}�.E\�d9�r�Z��9�b�Gu��i��i���;V�Y��ڠ�O���(�o�����[F9���r�"]�U7�%�U�G���&������U��S=z��el�w�w�]_���)$�n<u�tN'_��ߙ y��0�FuAZ�G������ۺ�&o(�~D�U9��ŋj�����ycUa�e�ғ`�Wf͂1����|N�ڭ�rϮ B�Ӎ��f�V�y�N$՘/��0ܣhvGR��Ef��r�(>��Kڐ��^)��d�<:�*�%�i ����+��k�����`9��q���=�n�)�'.��q�	H��c��8{�0�E���C��y�4_W7��]V��)���E�(��P���v�&��s �!�KJ>�R�s���4o�v�xl����m�%��O?S��1� ��:w�-f7w~�n��t,�C%8����3ߡ�O!I�l�71lA�!��n�V�lkIY���Ua�3G��[��kaGy�&:����|���k���O`n󚝶� ��2F�,��<e��
k���TT-�`�� �����'����}�O�kE�Q���+�6w~	��@Ha�����~T���<�T��%%�`�|��)3|<��QLpPS2��!�j���>B�5�k��? O�_d���r�f`�#���yee�������՗�g}|�:Q��M87I[F� �Cm���B8��OG�ͪh��q��H@= -�W�q�3k��q��R��C�6a�`���p���� �D3�p빧��8�?C�u�a[&��|�ی�#疙ronl���V}h�t�2(?9*��+����D�N���?H��M*8LT�ڙ2�B�� �xc>�<��&��wro=�Q����vꌋypG�+U�(،;v����t� ��s(Y��v�Gh�{�2k�5����-��~s��R>�/��B@s{�h��� ,�o�����i]0�}�R�����]]�p �3[c��y.|�Q��^\�4�ܠ����H���py��%Ep�C�&ړ�5+����3�]���p	{��ɖ�0'Qm����8@n����К��w�����:iH�T���?���"� ������<ʺ`Cr
i��ajS�$1��j΢��f �T�!Y�n��Є5nA���k�Gd�{�bL�[?��ߍ�"%K35��7=��>�4�r����ز�.|!e��[��+�6,åP�˂}��p�@�����s�LL�`)~�2��H���&��9�α�c�v֚a�^wω8�0��(�F�������u�6
�E�jN�+�aI��}��T��ݦ~��S��ԁU(�������c�!�X���Ѹ�2	�'3Ι
�*�4�e�u����'��Q^X݋��|�^ �ׄ@��I?�(�zr���;KI�Q��^��3
����l�B^��^eWL�5[��,T���5�=\��_���ոQ΅�C�Z��/ .݉�R���s\a�>��A�I�_��?��D�S�ӂC�pT,�'��r�oMm��|;�Z�yO!�RC�D��(9 j���?0_%������̬5��/ΣIy.*8S�
���N����*Hc�(�Ö�M�cH�P!�L���)?��t��@V!�����I�Ø�_�S�P��|X�ޘB��	m�>_^��u��aq'e
��\lj�t�4�#4�r~*� I������\R!`�V{�6c�n�D�T���a�溈J�*ԓ�v��+t�_�w���'��OA#k��\�mQ�h�2�ĺ� ��]aw5`4���r�H�� /h�}��sr��K71'x��b�&�}~�
��K{K\�e&��M��^�c�� E�O��[���P��()"[��w�M� ��eI��ȉbGZs
"և#�VM��p6�gn�~��(i4���do�'O�"ѿ�H7 �����Y��v��G�_�8�:�aq>��{d��.�lO
e�J�	h#9�����R0?05�#<�>Dp��}� 1 N?�<��x��\�X����9Еȶ���$�L���U7�{`�"���Ҋ����9tr/R=e+���a��9KS�3��)�8���JK���8�l��~)nw;
Гֹ����7q�E�a��AQO��9�cEܬ=���f��9�<����]�G���>ߛTh��d�7����2%���m*I�fl��;�^ib��'����D��Ax}�h��f�/
kz���K��(�� �*��M	�MQ��7�q�X���ihǭ���Y��hf�aA+J;D���Gk��X�	�n��r�Y{Jt���D���\}�#����:O��g$�kK]O8C�m�w�B_�훳�k�]��|�>� ����~7���U�M1#h���a��#O���J��k��b���z���� I哖�2y� <6�,s�D���f�<��t�kS3;_":o��`1�:��z���,���N��2�5sD�gL�3��k�܉���R�\� ��펁v{6Hג
UC�L����˴c�~�G�'��K�'n��տ�σNT?��R�Vn�<[q�t�+B�a�1Ǝ����q~-��:��=�9^�l8��M!/�@��j��h���4�t��L+�1�O�⫷c+���Q��\� x���rV�H �R#�t��;�!I��X1$v�=�V_��6=Ȼu��$���f��G�\N	~@��CӞE����*Y�����>��=��r��/�ZV��X�;P]+ǲh�����u�!���11�^7l� hz�ׇX�QK�5��+�=+���2�%��D4��?;���9V������F��3]��}�[��P,�B�d�A[=�hݳ����п��&w�Ɉ(�][�'8���+������R���єj%��LZ�V]�4�w���� �2si��07_ ����g�Q��y��t�X��1���^�v�1�K���uX��8S~f�F,kS��U8����˒>���	Cc��4���'o5yvǕ��]��'�)�� m�j�n	�c��o�k5]���_;��ї q���U6�.�^�d��>����;��HE5�&�{���\u��+����a[z����o����]�N�l�  �C��u��Tܴ
9�ʚ���E�{�1W'��b����_����ⵜ�Ӯ�<KP��u4w�4Qn�^.�`�sݪbio��ņ�x����{���ހV��l�Tl��>����WЗ�b�H��ʀ����e����N�5�a��r����M~�x���NS��ᱍV&0G���tZO(�sۄK��Й�c��ޤ��s�����38��U�.@(13�L&4�%�t+cD��%.��4�H��G�
�3�qM��k������8�=QKjи�C&�ތ���%$J/��u�9i��e��<< ��?�>{�<�W�)�$�n~1h����1(j��ġ��k/ln��4�|��<Gz
�Ш���}�ur#.�����ϕji��%�C������ӆ@��S�#���N������Q�R��w$�g�����@�מ�4�y4*|:���հrg�Ⴟ�b�>����`��\�u���!(�'���Cv���*����[g^�����w�����d9�!��]�o7F0�IɋA�$S��/U�R%sbɡx稪���H�g|��屉�v�D��x�s�~R����OE��e�J�����$��ǉ�
��$��ЇE��w��U|��d¹:[R��A��X!��Qn�@М�(��'랍0j=6ĕĥz���n�L�?��7�����X$Է�3B\���&?�Ա�R�}m �U5�y`T;HUɍ��-�o�?͊��߲�Kl��V����T���e	�f�Q���#\�_ ejs��(�it|%%KFE,�Хf�7N�<q�Xk���!4���Y׃�l�s�/�F:��	!�Y���?.����x����!��DԠ�Kf��A= ͣ�y���?�Y&��u���,M\��i-��=6�`�e��2Ý�4���ɩ�	���2tX�2�lvg	��E6\���H��4�K���3%(u��l��h�7��J��'B�;K���k�2�a2�({�iS~tY"��\�q���2py��H���1� �Bۭ�k�L/S���CP;͂�iT�hn�!e�3�N\z2�os}��Vs��#��!��C�usI��~�E4��$��,��/�Ȓ<�#�+.C,�C,^Dq���X1�?1�(wlv���gB��˦��s/T�kqr���7���g��)3	���BJoy]K>�	�:���b�'cu��@�U$Z�a��ݝ�(A파Ϗw_$�A�爒 ��2��]V�p�t�sUN�P�	���]!�`�d1/����K"1�hO��F�￣'����Hi/p�vYm���'��c��HԸ�wg:{a�d����?���Z�6Fe"�#�|}X�K���r]L���zP��5��C��/�LV����X�	���m���s~/���!�(��u�6�����Z��% sZ{�6Q��u��P�EB�IU��p9�cn}.��S�p%�`�ď�BU���n���Q�oX���v�AkN2�>ƍrV��6))ն�G���(�'�Y2�;��\c�|f}۬�*�lG��q�"A��{	>QA%p�Z�y/Zg1�Y&��)���Ǩ8��{���(��5�)h�y(q���78��aϒvw,��� Q`����Y�6��u]�嫐k���Xdݍ�uM�����T�� H|�s���ʎPLsc���(��:���)��II����[W��7�+�
Ľ?n��%��}k��.RǷW� 8!�F��0�U&ڼo3�>�)��s忬����0g �m7�Ӑ�����|�p��tlE��~���+F|�����k��+��P�90ZiP� ��]/R�ES�V��T&��C:]��geyﲜ��^Z��~(�&�P��	�յQw���v�v�y��iGL舞I�#h�>�]Dc4QuHC)�Ҝ�tM�jF�7� �
�M=%�-���:�����d���RE�J
+i�� �bm� ?ۘc�a-*���4�G��g�2N���=1q��I.�L�����J�L2疊k�*�Mn�d��:�M��Sۿ�~�c�^���S9�u��P]o]���,=�aP']�)��U�D�/�Ls�0Ȣ$FD,
�1j"�>��y�.�����s���;i�cY�]O�o�-7���H�M���i��H��H�c&�6�,�N?�/�0@�l��B�:�I�#�Ͻ�����bal&��q��4����	��\�Z�C\�ܪ�,��)�l�"�V��l�n�����OW|��ƫ���� e�u�ڸR�M�8���n��:D+QΘ6���Vqz:\����g_|\�f#��u�Lg�L��K�6\�r����E����?D#�,.]�X����r��x���ǎ飩�6�� ����=�h�
���r=�$}�0`�F��i�ڦ�zI'LiNSpo������T�3~~c��#2!�%��q���#N��l��5d��`G_RNSqNA�>��Mr�s��]�������]��P�%
��Sn%4`O�X�բ�c�A˯>��4���@y(J�`�c��NU���^o`�Ϣ�TM΢b�`hݲ55�9�J"�V<A��yQ�o��zV3n��x@���-8C*Y��%��-��	͊�WA�U��{U�Մ����9M��x��D4vj�:��a�8tiN����ƀ����0��Hjn�-ؘ�l�i䱐�p���)���J�t"�l͟@X)sX�+��+d�M�ݪ�L���%�;�-@�D�f�Qe�6y����>9#�V��z�9�����5�1���sM_j�.�	,�y���:��	��&����� �X��ch��G쬒����<���"��H�kiG�w�>Gx]��lB٭_!N��xo k`��G���I��fC=n²��b��F)ygш4a���)�X8K��ň>�u�� @�%g>��w9>Z�9���aG^�I�2�LH���?�{5���O�w��0j�~c�Czޏ���%a�`�}6����9qٴ�#]Y�V�����B��`2p�qS>a��("�a��Qpq�jTNX���ټ�������D�c�����o�w-Ʃ��:@.�#���t�0�ka���u!ʠ�!C�1.�=z$�V�%Q�����}��Õ�ܨ> ��yjp8�����+^�:cFvHN]q�6QU(�bH���a|C!�ArPUwe	8�7�O�>拊m-��lL3O�x�^H�ƍZj��-׎����q�/h.G���.��՜M��α<��ц���"�.��ZF�ʕ�HiML��b�C���u	)���[g8�v��m�+�ok���������K�$���G< �'�<�R>�w���XH�� �>	����3���� �H�K}����Xz'��'!_ѯ��foK����l��!R=���k������k*4��OU%�=+���$֔��^���=oD��/���ea"��^�,ˊ�y��������U��}�I˯���Wd-��{q9I�PB1ґ�B����d��:���:��SI:x� $�"�e���^F_-I��7�ŕ�->��A����D�ErF4]:������1g�w0D#ٺ<�n���,pj�pEK�!dhy�����hțd M��'��bG������ÔR0KSV�o͎g�K{D[��3�S�7/�+�0蝠8�ϰ���0��c���oT��Z�(q��kj��>Shϗ=�F2�'��-�<g��hks>Epy{�̰e��������P7��O���裐l�#��7e��+P�a=!�x��8�b&@
'ϛ��&�����~�[��G�nԬx�l7�Ȧ��)�
��0�w��]��
����{�DEZ?e2BLZ�kqˡ$c�`�j~q4̳Iiy�|�L{bP�	���%�Di����d;U�Vc�VTj�&����M�=K=�޼a�.�b���G��ka�����L�‾���>�B�S���c�dhP̕��f������:�7�A:c ��/tJ��ĵZ�[A��ۂ@*�����C��;��|!�sT����h���y���]4���Qh%�jz)�q:9�{U�±R�x�sr9���DA��W�!+��e�1�:�wl0.��z��L�15���P-ֵ�!J�/9�/��d�E� �CN�r������8�jVƜ�	���tɟ�0(�������ЍuŌoq��P)D��i�=z#���υ7;:�7��
���?���21��|�h������u%����F1��"uwi_�&5Dz�(�����L~7%�5���p���+'U9��>��#����*$��.�i��6�� ?:��O;1/���'24�W����ƕ����ZM~��<#��X�z�,4���X%�\�#�K6���h��21�W�u��R�AJ�A�\O"�\Uo�1�m`9�?�<A����u��_�
�YZ�)q���q��\����!(�Jzt�p���������(��z���*^�a��(ivH��Ʉd���B����q�V�e	1��Awƿ}r�T~r�Ț����H)�;]��$�_Ǖ޽��_Jkd��
g	آ�کE��Ŧ��B��5֪��k������۩��_jn�m9���Ʊ��\Z��(j�~'���Ϙ���LF����/$\A�W�A��Gk徻�w�P�;�g�k��WC��x�b��E!>Jy�a��4�9��!A��,V�C*�Z�&o��԰IT�uf�	i�8�mT��H��e�}�T�?mngd0��?D��:��s�8�ɍ�
A`��s�x�!��Ӌi�o~�yRH�['���Ozi�M�@��%���D7�C��2�C�Dl��s��S	ϱ3���w;�*c$�&S�i���C��MQ�8��p��Be$--�3 �~]������������l���N�pT'9XP�S+9�Tm��w �L�4�Xb�SG0��k���u��G���ژ�0�&��̋���)����#�k,%̟,G�=��00bNXX�'�5-�,�p�H`�A��W�{{��X��ri���7t�j�i,�4���B%�z�=�u?(r��6�(��br�mi
�A��̍��`��0X�MՉ(���ݲo�����O=��G�u�q�P��T��6Y��)�/}x�l<pw�ۼ���i/�N՚-@i�P˕D7jXGWՎU�t��w��߆/Fȼl�⻐��8a7HI�W�~ߩd�=��G�7Ř�=Q��9����1���r�����=PhF���pI�5��{yHk���/���?�*H�"m�sC��T�-֎ג�"��[��/3J���Uݡ̑��N^���?;$WzǴ�ֲ��P���:7��HW���\�xEsz3�\��L�Zz�>K}��P�93E���������4�c�d�εF�^��4�;K����+Gշ�,�oE�Ep'`g�����=�"�Ta�=�u�]PX�6GI��4�d�B�Й�qXc��_��>�����,ސFK����6���%���С��^`��QUS������g����0����BE<)M����_I�w)T��6��ɺ<���LLJ|�8�A���9��8m�}v���E�W5A��R������[}ޭRnkSLq#z���� s9���w���篖���e���Pw`n�ڄgsge�_�f�:X��w_ଝ�7�ˠ�v�(T��9��1K�vq�\Kl�[�������j����|/����x�@�/�ݹ?*���j_<I���p��.�r������p��Y���E��d]o��B�'��z�'��"⪗Zӝ?_5=�^R;��A͛�fV��ǹ����f٭��8jà���2A,+Y5�Z����s�/O_����ߞ���aiUL�q��i���.7v��=>ݑ20O�ޢ;+Nן�ь�KFjԅ8�B�P�z�'v��$��r�%ˢ��z�~Cp  Q"X��U� *�Fމ���L�iir�����wt�W�'�U��xKy 7hs(|+�P�tw�zɦR�܌�����q�c���)8��l��T)�E��o��H�@��X�m�a*����O
��hڕ�(��/n3!�K�I� 0���n�=�y>�?^歞���@��M�\�D�ޒ�Gg�t	���|<x�W�..�TG��
'^r#03�Bx�Z2$�!`%��ư�c��8����@�,uGy.�yآ���Vl#Ɩ��6�s���������sp�h"(�9�Θ�.yQ���O���ђ��ew�d.Y�P��Z����;��_jt=�OX[b|�75J��E_�ϴ����ᗭ�k�?<֦fCc�\�xvA8P����+U�����)ش=I�#�(ӢK��v��xx������x7�+]FX�X�o��4���m������Ɗ[�#"ί�ċ\�w1	У0t�4��)� ��9��qǜ��Di�'6ZV�������[?�)��0S�'M�C�vB����J ����Wяaz���~2<���o9�kE�d-�T�J�zE�p����tU�_<#P����y���s9W�*;)����8��nvRV���ju�?�E荓L��jkuʴ����¸��y�cy��:����NW�<�&���
�[eg=�I�qY[����r�	,���ɐ�����z4��`���V�!��G�o�)� G?�sdۆ�ai7kr���$B*.	l���I{�z��3�m��i�S��=��	��s��fY�=_u��]����\�jw�9B,?̟�Ծ1���F�ĺA�����l�����+n�`��'{��Byo�A����j�7@F���o�7ٙ�UY��YD���1M$�\�"�V.���������}E���*�#��J�T�� ��"��:��[��;�rl�0On��ٛ���	்=�4��(gc��&���1-ڧY9ឫP�%~����2�4�7F?�>�)=F8Q(�/��b7c��l0�C]�})���G�F�&�-Sd�����Ki��݁�_	�jRxa91�&�/U~g�Ju�����|\��ߡ����T��Bj��3_j�*}��Z���`���Y������蒭��u?[����H��Y�8�6�~�R�^�}����J��B��á�/U��(����[������2���u}ã��4\bk���c-�,�����F1��6� U~���. �O��r�?��-[�e�`>*.����Gm�)KL\�:�J�N<�"�̣�������k^f��,#(���%�����{q�ZN�"7��2�����lV,0f�"E������IdB�?���2�����Ojx�P��@�GalY�]�r\W����D��	=-y��{Mz������`�$����}��gM�-$�{�|$cZEy�O|q����op�x	o\,�y�r�@
,C����[2��4ؖj8y�=�[�3�����y� w���]�bQ2�`"7��C�w���2�Y)�ל-��H�+2c�
���X����[t'D�^��9d��+� �ѩ}�"���=�^Ba:�-$��Z1JqY������Oi;I��ܤ��ϕ��\V�<4"�<Fh����E`Lj�ᗍKH�=]��n�1���f�q��+{`
 ���Q-��������'@0�F��I����x8(�H�l����!�[N��RX�O�J����-ɜ�tvI��67z-�`]1�5Qb(���V��w�X8��gLp5��T�N(t9�|���Ы��ʈ:��/r,��2�v}So�}N@����DH�L��ڻ��2˦�He�	�3�Fh����*{W���lP�h�NH�0�5�k\���yCww�S���%��j�3ڑ[�c��#���Kg�|�zK&NL���:����H=�@m#��Lf�5�`L\�X8��~~�|GA�ܽ���d_PYcz��͎�&iY�)�"G�<M؉Qي�>a-���z�����r!�ѽ@��%8���^k0�_96h�9iޗV�����A��9N>{�!>��v�y�J.��?=�^<����'7���Su�����G�GaZ�Tg���̒�Q�H�w�ȶ�������h��1�K�:Cx1>�o>%�
�&'�<}�)��jFI4���,E{T^���1�&)��[Z����G�#:&`�~=Ԗص ٺyj�8�#�<`������7L�"�2�
w.��<�gׁb-I��(�5��DϥȒ|��@ ������N����@�éi݅��z8L�f��y�pdO�J�0��w�]<�'Q��do/�T��˟փ�W�)j����h�2��[Y���
C�Z�/40s�y%��
*Z�����I��HU��%�T���IZ^1��9��?%�$�F�lX�u��îs-�pga\Z�0�F�o[��wT:~^$�.�M5��@3�Nwۻ��_���R��c�NO.�Q@U��	�i7ߍWuB�2�7Gf��t���O:ڣ�����|���s�@�p�ؙ�̂��א���Z�k�U�{��E��!5�o������]�����ɇ�$g�F��E�O��l�k:0vF�on�DmT��[��s�߁rB9eAFۛP�Ą�������3;�氏zz��c��*�-�d�Td��ύ �"���)d	#f��*��R;Ї���!����_�+�B����c�$��lL�'/o�.�B5S8g&/�o/m+B�Ѫi��-�v8�RP
�^���w������ɍl=��ϲ���Du�n	U���"x>�T���7v�lhab�a&��2&0ˏ}���Y���#�t�T�����
[ �}�Ê�Xpn
��7�N�F���R�}Q����6�N�|r!�I�]$ba�����u5Y(��q�`���\k�C
�hqd�6>�ԏ�;�B��\V�Z �;5h�SS��y� ���k���ٞ�yd��%�:���K�&�&��[r�bKNEqb�!�O�%��q����2�3���V�gzo�0�h�(k{h�*b�YQ�}��F�:��5�~! 8�z���f�3����ӝW��ˍ�_T�k.��j��o�IF �ɇQW5.3��L� �&�9��.i��� u5�=W�e���=w�Ɯ˘8Ɛ�̵Cҫ?S���C�㸚ZL��ó%6��]�����CLY�\h˰	'�i����Y����^��;i21|��b+��卺�cp�-4VR0B�v�v$F��� 4��3����nj;���4@�QG3@��Л�.�h�3>"�P��쬯���ҭ�3V����eK!M,�CA�3]�^4�0"7��j�z��?��������'�[��N>�+���p^�p,Ǆ���2���S�2C��)�;`lt��@�30���76��K��:`h����q�b��x��,?�Jvّ0��f���KIw�#uU�o��3_��e�f鶝�����5�1t�R�Y]?v���Y"�`%�*��:\ύ��<&8u[Bx8��!�ɪ�p��0e��Im�g�~�"!�b▪��-�=���ԡ~ ��ύ.�4>�^��K}�-���|�P}����ync�h>����`p�h��yƖi���{�wp�-9z[�y;:��Ƃ�*d"19��@t.�WG}О3���.\&��Q�y�ı��LX�9�dA��0���p�n9���b�i�*QPI%�?(6[9�p������=O��b���>>��8|Q�ސ\���j;��j�W�Jg��!�s0�K�����A;^�HsH�py?Tq�|������ѮlG�GE�LK��ܙ�j
Ҡ<6Wf�W*\#w$dfW��1�z͈��	�X�(;G����Yם'\�n0x$����f�d��i��Nb)�eܛ��G��zh����\*��M{���a�GȠ���||�(�T��}Q�ܯ�{�Ĳ'|($
jQ	N.��Ӷ���/�/� Z�+HU: H+�t�j\��c�p��#\E�z����D�;��	�u�4K=�j��i��Ɓy���J!έ��Uی�~�$�m��;�8tSv�C寠"-x �9�O P�R�bh��Hm��h����e�̼�q8��� �����d��f����/���ҏ��)�ɉ�".��|�:#u'��t��!�������u�H�]E��Jy�RA\=�M=
CdI���&I6�FgNO[�_�}���{�ڬ��_��R%��\-3������+�h����,��<$�&�_�_�ɾ����×�x���C7
:��-���=�O���ȩ%�k���h��[�j��'���X�n�^���嶫&~q1���䳾�У|�hT�Q��xb�
9���~�ϐQ�!|���U�'�A�#yJ-^Ŕ9e��zm�d��k���j��@x�˲�A�̗͟���2�`3ALIp< ŅÒ�A&��I�a�X@��&�!�!���z�F�w��Z�-PM����K��l�pv��
�ǽxGGF}]3�\���h�om��&�g,�ԧ�
�ƶ����m��<�I�+��ZwBϷ��7N�H�xtJ�R��6�V��k��
9���@���Ѝ��K�� �B&�p{��m�nM��G�Aʿ�l��.��tW䢈Y����m�wO�-� @����&�=������[��	�!7���0/����<�:<h����o� ��^�-����Ģ�{�����L�(���Vk�����7���+��!h����+���S����9.(!Sc��4Yz2��i���2ݦG%Ԅ�xo�>�)��w\C��[�&T�1��j��{r�
�Җ�a�W[�����o�p�w��9JPv�*w�<콍�I�U��,&�<ֆ+1�%^��:D�'�u�����I�c�$������ЁΨ���m�Y|&yD���4��?���c�HŹ/Q�a�@q[*zu#��6�6�О�l�/<�q��Q)�Lyعl�h��F@���um���5�+�L!�K�^*��kO�X���ϩ��|շ�T��Q�WW�r�\���4�����򕴁��� ��	��	����P#�8{�Sj�>�`���[ �3g���f$3���akXYW�H�["�S$7}O�iA��6C���@?W�f��HCњS������u��U<Y��w�9?j���#0�|��f�R1�v�}CҜ���>el(.B��6aGV}�ŵ���	S�Ju�R�L@�}�_����������:`T�I�j�Y���i���>iK>9�_`�8�!��U�2P�m�Yi&}��	�����C_�3kf���={%Jg�&�g�W�f'��ztm�+;;4��o!��O������x��1oQ�y#��*�%��?���W </�z��~�oHY	,15����ү[���O9$\s��a;|�w�^n�5���48镚���C	u�|����}Z�pN��%�Mt�(8l`HS��+=�"���Y,g�}5u���O�'1N�<��G_N}����!o��)�jYn0�Úqw�Fg������z�PΩ�"�؉�e�x���S������ �,�X�ɅX`k��/5&�xo��aLs~JQu�)����m��`nr�+z��8�po��Sک����������~��]V��4��nΆ�1��G�)�8��ޮ�C�� H�<�)�9�T�V�D�&B���ɫY'��4݅ŤaM|�����L��׶I�V�=�4�_<�L>Ka�~�>v�/�gF��U��}[�~<����	�E� P��M�^=
�^r��ٍ���G�S�D��(oB�t�b�J�`Mdcy*CeH��d���`٬�&*P���o�|��מ��G:j�� J;�`�=�������M3�����D(� Ԉ0PeXu�@�1��x�	��S��~K�z��Я�,{�G��y�-$�峏nGA	��$�G���z47c��9Q��;�X8�
�|k��ւ�H�O��Y�`���:�����iд ��v,�w;�xxpo��q SF�A�G�Ԫ7Y1�M�;23���Zy:OTU�����@z	{UFJoT�N\|��'nJ<���x�
�����h{�|>,�Z��e��M����g�](�a��
r���	�emD�� ��!�1':�35�S[Ċ�0��:��m�ù���t���{)�b�V���J� <�����-d�����pq�	t��S�(�Cː$Ke�t�%U9/<ֵ�m���N���y��m_S���^�!���A�fC�i�L��"�e�\2</j4�*:��l�-)����Xu/�l�1ΉZ�5b-<�3r����p%.4��^���ݺf�f���~��<�͈BÁ���rzAAK�7-���"��D�����KV��1N/ѕu��+��~R������F�p#��/�b�zG{��d�JĔ2R���Ļ�O����sL��D�(kO�@U=]�p�ޤ������0`�k*�}�QCӦ��5��J�P�k�D�0Ne���*�����
'x�'
uv�~�t��Ϊ��q� =K�8 ʅ��ޫ���5ؚ�oNQf�tp������*�2�������R���gz¥/P��<�"� ���؜�b�?��4�F��������vߏT�P�k����_�R�z�,���ƺ���9��P3�h��}%v�S��5s��ϳ��iqN�����Kڰ��;�\�]�↪��Y���M\M&�.d�B��=,�,�ñ})�3���N��M5U��}x#}�?��$��e	6�#zYB�Y���B�๵��\Kv5�����keD�b��9��W�>��o��0ceBQ=�Iy#;΋i	��{�FeEQ�����a$�]h�,n�&�(�\��A��/���x@�J\��nm�㓌�m����!-�=u�4��Q�jƌ�ʪ#�RF�[OLȿ�Ӷ�����0��ē�x"ο�I��wA���|�׊�{���+V�B{��۹9l%E����z����z�(�Ԑ����$r��C�s~�ˡj&�u�J�|1x9:���������W�_eh�L�X��Bx-U��M�BG��_\�E��j�	'�:�R1�f�`ek�4b�;���P���J����Й4��J�+�!�QG�s�Ώ���2�%�/��u�R���.�Q��9Q����2<�o���9�0��H4Z����@Z��E���2l�_�0W��f���-��¯+�K��#��	�"�8{�[:�0��l���k0V�Ƿ1Gi�{AB*���X�z:/hS�o���" ���R(�!�+���&��7"�!فD��D�a�.���hۼ�!�K��O:����PT�z������|�V".���?���$>O�%�k����%'dw�80} �	�x](<�Y|"�a�1��w����_�1�阾A�����@m�oӈ:M���vP�%��j��,*��*�w"-��V��"F�d�9d��+|�g��-tb�~�V�ګ�wq��"�v˸���h$��E	�t�榆�g���b{Z��UysG,�
��5'Zi�7VD5�{]���]Wi/��ך�V�C�4��~��0mw���(iU�i9����`(O�'[��H���6qH�3٤*��?G���W����UXR�೛����'8��Hh��#�a�z=�m*�������YH��+)��4ߊ��+��L	X^�Ť(��i�[�F�נ:�Vt<��4ǜ�У�����W�O�T�wb���|���\��&ꓒL\th�ʣ��D���jo:H񞵄Xj�d�6����v�����O��=���K�ef��6���ó^�[c�:K\K_r{�H%O8�rf�N�:�AS�����>8
3d'm�����x��3��'h�t�	Q0��v��@~K�� �\.NyԊ ^�UQT1T֨ށ��@P%r��:}GU�0���A����:œ���۞�a"�C��k��	!wEq1űE���)��aLý6����`���E��X����=e���d\�\��wUm[�қ��,0� h~C[���þƐ㲒D�n9m�A��"���+�~��L�ˊ�/������Fڇ}�G��Q�H�"_V�H{Nt�Cɻ6�OK�cE��@lE�ލN�D8�(з+���Ԝ������q>�M$RlŨ[�$Òa۟�!G�oL�b��dd���C���gn�4��w�.t���iUU�=I͵2"W0p���/�9��6����0'W�+�q�j��;FY��捵��!"8
9KN6C)!��|AP����WH8н;60�����I��$�(�?8o�$:�Ӧ�h���l9��<<V��58j��XB1�ts�?� �؆Q�߿t;��\�x��n�aò��&��{����(�Wh(�KR�v�X�O#����'o�P�R���m��ΧsL���QL�Ιv��6U�R��lk�\+�x�.��,���K�D23f��%�Ζ�.�YE�Z�	iZ�ŗ*�mF��z���U1�;k�~Ǜr��/ B%u����3��ҞBQv�Y�����@]k�~^�g�����g�%s�yC�0XK�ys�h��WP3:���oʸ֫����4;��ʘd��~p}s�2�B� �j���M	6�z4YJ��wy2l2Q�m�c�~�C2��h<����@�]��������D��E���(?F�E���K����\XU X+��R/dHD��1��` q�섢�%ϮP�*�����%�:��Ous�"���7�fv����� ?�hr�߾��M��
7 V�Vg�\�Za1�u�ri�P�͹�_��5n�/��u�n�̹��� 
\�ɏ~��"��/�K
��e�3��p�ӊ���\����@�8����:7�IT��+�X�i�pO����jnqP�Vv�k64��<�؞���_��T[�|����V.uq�ꤵ]��l�(�&�nJ���RqKfo���c:��
��"u9O�H������D_��A��6�Q���i�k=��Zp��?ß��~S�BK�2�r$�ցUG��o-nO��s518���Z���\�'��N����H��1�1���9p�[�_c�;��k��fG��.�X�Y=/�A'%���P���*sS�%{�㰃r]m�	�*/��u^VV�8��t��d�%���B�������&C�]i����V����O���kN:��,a�w:����p��`,@j�������"��9W�c�%����r�
x�N�������j���uz����Ǩ5�;Kq�͗�ZO�T��t3�u���3W�S;�����`j��B
z��?����$�
0�$\�À��OA�0+ơ���b$�&�0��g��-W��9��佟�4�Ü&��Ј�$^���w�(D�l�e(<&�_L����Rz���CT��6���~��.���|A��D��w7�c�˝(����PGU4�$����H�bd���95��c&��sU�t������L�jD|���g5��cDw�u�h��ӕh��IƖ)���R^82����"��2������w�:���1>D��e��OG==W@R�m20K��Ėy��bG�y���]��B�w0{$�'<c�2};��b���Z�Ǻ@����! ��	O�� �:rl�Ø=�� �5.��A�'GK$���z�C�J�u;O�����LDN�����`m&�Gy̱�0��yN[�G���i����r�� ���������xS �X[��Vο����Q{���P��4���2~��-�;�X�t�x�ǡ�� ���q�S���v�0��K��90����>0W�wfQQ���q����qf/���X�Z��`ޡAJ@���HXT����]�������C��Zx�ZɄ�lM��<{���[���W���#��9N:F�Bڍ�D��Ҋd��P5:�U �Co����W
XR~��ku��l:�O�N�~[N)G� Us�-]L�ҞC����`��G�������ݸݮ6%7�����N��{��KXv`JA��9`�d�/�lvoB�S��/���>�+�Oi�Fs`~VYs7�먶thf�����I]A�����V%��K	�I��M���r�E�edy��9C�?����"�<�8�� 
u�u�����_�����/*hq�;������I�7](�r�̅�O�w�e�Ĭb�x�}M��i�}��t/���p�Kt*e�g��]-v[�C��/��]���࿧٩�t{�����0�q.0!$�lI�`�G�ny'���fJ���(I@�*@��ٳ�(Ya���\�*�oD���`��59U����*.��q�����0�aown�y�]��]C�I)f�UZ�SH�����{�6t��Ƨ�ݛ��;0����9oVF���~�m��}Ovw���f�Jn.o���X�,R#$�0��!]�0T=�W�@�r7��u���[O��
tkg �7��TE�R�Go����Ud�;n�5>uT��HV��d�;W(����>��c��A|%�)9Oh(�����I ��1��X���hZ� E���8�j{��$����4�J�}�n�����dCȣ}C�,"1��k����~�.�8��t�y�<b��RuG.ǴԿlEh�5�&�.����q��9Xi��L��9	�^x̬{f!S�q�h��5T�s�S-��dV�������漟��U��G/�\t⇘��M]����F�x��< 	+��T�\~2�ǻ�*_�-�%�'?�O��i^0I[LKp+} �Q�C��5D�R�D���@}��hC�(��ʁQ1#����溚v?��V�����\�%j�f�$u�}�o�	�\�L*exZ�<}jQAɴW�� �����FЯ̉|d��J���r;y�W$k�LK�-�º�3��!.|0>�/��xaև�GrC����6]#0[�r�������<�h��\'ֈ3Ge���&�k��������C�6�Km��i��+�r6����3N@S@��J���/�2�D6�S�W*�$r�Ӹ�Z5�RD|�����km�wU�e-~�7"nW� ����5�Lk�٧�tv�c����Y��_���w.�Zo_���?��M�������sؘ��=�4N�/�K�Y<��v^hY�ڪ��S*Ufļׁׂ�����ck⏶�7�X�ɹ=�@�=��582W�4�*�L�H����}@�	_yZS��3� �����0��<�<zwU�{�� ��l�&�޻"�<���x�V������ic�qg��8V2jYmz�)��B�j�.�]�o^���@K�pӖ�mR
^�6�����.u�����E����):	�gGSs	���@��{�ȯ ��"TH[��԰Kɳ��I���@�aE��Iz� g�8f�C32�5U:c�����%"�d'E?���m��0�Q(���n���岂���d��ؒS�����-em�8�u�nkS�W����(��[Gض�D����������� .�ն���FG�i�ct�-Ϩ|X΍=F���ZFlE?�wY>��l�����]�͐y�*Ύ.�V�!Ng��žm��7�� ]8@t���#�L�߼���:�3����δ����ƩS����8!�Y���0H�[?�Z�������#����1x\�7�1x�+�M(�p��h���	Vi�}����1���bPT!Mfr!����ʷ�k����8�q�R�X��f1���:
�ߟ"��
2��إ�pΌ}��+���+�(Н��px	��"������.Y�W[|�@(�B�6�u�������NJw{1�]�R瑙���RuB�]a���%%���Y�[�j��b +��5kwZ�p/�ĺ���@b��:��cO�T>A�G&y�gw������@�#>�/���o��ۯ�}��,$%�K
X�-Oh<I2�q�u���?qھǣ�����\�
�񙒽���Q2`fi�g�P��}��Š��	�c������ƫ����tՋD�L����2�zAs:�Ƕ���Y�T\�H;ܖ[���t�<�g\�i����(��`��������u��q�Eu�5/�ޯ=�F����/�z?c'L&�)��.���DX@���v1K��t�sV�g񕓎�Y���	�'�j6���F	���/Z*����}�l�F*S�ŀ��G�L��b�����4��Q)������yL� ͐1��Fy��ă�Ȃ3!aepl��B1�9�n�pZ���!p���:�?�t��[?+��.�t��:�yk$2L���K���um����Q[9E��88���c�r!8e�"��y�P:YYV�k����]�u�x�@Yԧ��
�"��T����0�������� �P�	I��s��Âs��a����#'˱��jqm�/	<��Y��2�e�J�.23ضً�ǀ,�������u\��m�u�0�$�}��#�M���� E�aVgb�;g��ʾgc�Ɉ�t��rM�i]��?nY��
��&�k������ �
�=1d���~u��@���'@*D��,}1���L��������l�ߥ;YT��1�zb��y��0�[����ڻSH�P\��u5�;��3����֮�����EV��]�_���UB-؈{���J��V v���9��8,.~
H?0�E�b/ɗT��g�$���^���߈��=�&&�k��f�^�M��E�-@7!�m���O���"x�m��Z��ox/\�kb��\˪�^?���e���esP���椡�
�ӧ=�_�W�'	���iJ�z�]R\w�3?�wmrv��<t�4o'na&|�k�e���(Q��w�*$���L�$b��3L,��Y*��@��_�Iv���臺�!�m��nv(� ��3�G��>-�ɸ�hcHY����o�������}�A��0nao4b����ا���IU��>��{`�����5�y�~��f�=oU�K��+����Q��/Ca>�V�z�S>�����5�����O^�Dp=�K3�0P�[s�g����b�,Z���4����	��e%��<�n8Ĕ�❻��q���6�;Z�F~�`O����ITA/$S{7�z�����2�mn"T����92���O�����L�^"���l��>\d��-;�c���|��fY�M�UJ�j���ZuF�J��6�^�C^[IƩF�S]�
��-fг�R뎎<�[8��T�ed�?a����x���,,��̿ �Q�x�5������F�o/^��Ar�r��	�fN+ζ�� nηVse�&������O���G�����$�
,D4iR�j�ZX M#Xi2ZiI����i�!Z,21�i���I�.n��`�g#�A�v=��푶�|��9��Nl	�����T~xor��m2�%�\ā9��vQ�j1���:�U�#z�K���f�lMp�z�ܜ0m�u�co{����ܣ�NN}B�����C�m�����9N &�(8ڨcj�}>Qc�H�<�y^�πi��0_ꮕ�+�����6�6��N�(� �0uC�=Z��|�W��rm�����?�׃�#��W�m�V���#�>�y�JIR�*��r�����m"P7wq Oi����4+�a��?�aq ?*_�����3�r7��d���a���=�'��x�:����C�%v�U��H�נ^�5-���x~�Xj���N(��i��d��c54ă��=4�!����N�\���/,�DۃT�k(�.����ۚ�ӰT�US�v �')#�f�m`d��ʵ�j	ȭ��� 4����na�jO6_���emR���P\*)��i؉ЭG�Z?lP���79gS���������Og �M&������ά_���gG�'�ު�����2��n���T0�$q��X"��x�a�'������a��&o�G���c$b��-��hV8L�4�>I�cY�^�a^�OX_og:���CB{'�
�L:V�7]��4��2~O��%�,Be�{M�gU�c�Zԗ��Q�˔J�5:�B���/���M��uC������3����R��w<����v��y#N%�eO9�eR�t8�����/oh5��t1J_�߹e�6ҝ\Vv[M��R�4�&�9c ���N�}��-����I�1$\=�e~RO����)���tI�g�~ �Ql����Ч�dN�K�2g@z�ÄU�4�+� �q�6y�N0o������o���ױ\�:���co�.h��^b��hٰE�z��6�xJp���Y��b��snz�)��3`D��e|6���/���*�~Z+<NW�m�Ne��}�@ߋmH�Z��13`"?�춺o���I7 N]t��sz���n��p(��1�p1�qzxY��}Ak7�r�����?Qt!�D)q#��I�+��T> �6��I��<\y7����������i�j��$'�[��Izq��"�D���񌏄zҐ��|�4�4�����>8`v�g��E��2�pAZ���1c-��tʳq��c���& �'de\�κ����a�6��*##��#��H�x gD�"�2�6��Y�'aG�U%�u`2U����$���ћ7���#�����Q��2��OI`��q�!���+"A���L�FLN	Hٚ�o@�c�p]�ڡ����?]3~ ��2nr@�L'��yUbK^��yh8�E'c�X�	��ٺ~]e�&��T@�\���3v�ێ�v�
$�5���P1|O�\�G���~��Ze֠�����g�bRMVx���p6Ƕ5��-3LA� ��'�%��x�˜��[x� KM،�	�qc� ���۹�:�?�Y��m�78J	�Ƅ�5T0����Q���f��s���x�~c	A3��@K8�C��]u�	��r)qߙ݌j�Öu�m��`����-M��o	,�Nv����Ixx՜�~���<�Hj�1ؗ%1qXE��a�Xu%x�,��V���L,�O���d��� �94П��#�x��3[�ɺ�E����U�w���DB#3`��|�
\(�������T���%��k��|�����FY�sJ��S�^� &L$I��Ԉ�=����qQd¾�J�1� ��՝�Xu�D`�HՏڥ�hL2�$V�cޝ����!���'������Z���IG�CZ��*F�R�6t�� =�R��cﾱU��s.��˫��N�c��]��>av����(��e�{���@2W��\7r��C]������0���E��Xr���ܱ.62Y��Ӂ�}�%�>���y�YR]�J4���d���Ί�uPbک6�f�d�`<�fmV,OC�uC����%2d'J	�D>�	#@�y( ��z�B�'q�/
�̴��
�I�1g���[��@����}׷�~M�0/����0��|���tԣi�����z�]1��Ȅ:A8��J�hI+��0����]�*d�|�Z���gWV-�NP�o�\�56��(-�0�K���S2;Yk�|`p�'Ox�/Ow������Ex<�o��̑�j�D"a�2�L9�Ȯ�������b 2£��-$)�Sc���;��K3�*ˠ_���_��uo�.�oJ��'̖�Gr��`�.���"��M�Є�Dly&9���'��fNx8=Em�ik����#��.��܊�5�V������^~�f6��<@���}�f�;	��_G.c��9#Y��
���FN�� �v��_&.ۢ���7�2�=��82�/��9C ���a�n�f.\���H��]�����{֬Co��1�� ����'��j�M����*�(���[�
�ȤqQ��<,�|}A�LӜ2��^���Nƚ����-����k3���MD��\�ԓ8��U�/�|ǫ=�AU��$�t�{�ˣ]���>���r�c�U'�d�-<q�n��:}v�{`����=�Bu��ؠ��eC����6~V����<�=��S��������$�
���L�"q�t���_�!�r.~�.H&r�ʣ�}�	�<\V���K��V�BcS�����Y^dJ�B�m�{*�,��A}�@���y��Hu�_*Lք=���F�H{?�O�
��ڔ7����6Y/
�����xͦ������/f7$2����t-ܭG������?�.����O1 3_�Ō��t���k<l��f���7�\;���QV)�<�4A�z[��?�6���I�vZ��5)B^w}�Jn�!���^�6��qI��QO��������
�nޟțw]-]��lMs����*�Q�����[���묬��?�u)a��0dLm�t	���D��S��Tj��JH�0}��ު�i�=�ao�����%��q��-�YR���J�ݲ �3�k���W�_�`�X{ȞQo�tG�v����_�,w��,��r�fΒ��|`v#\�*�:��8���u3�r�G�h�6��~ׅP�n��!W�=�3�V{���R������zx|ܮ�_���1`�F�C�5���:h����)L�$��XR�D�u�BP ���mF&DR�h�B��]����UO�\��
@ߴ%�s�i��rD�'� �z���*���딛\�RV[����0=�k3�;Y}뉂rD��Uy�������7�)�cc����A��|��ގů�Y�d�R~�p{@R�>}�8G��yT{�L���7�&<������cw{�?�� ���	��>3p>����.j�P��\���\���X8�`|�S���T54��q����uJ���k���6:��@8jU�Aܝ�:���T\��Ԥ<�U��Cc+�{��:귺��m�T�d£Gc'���}�Õ�F0�k���T�>?����L�6�K��(�w���!~�cN<���3>7�gb��M�r�M`G�|�8ܪWsE9�~��^��O��;���71����)}���z!N���"H�	fvT�s�>��|�Q�Il��PM3�'V��u�rym:���^�-��oL�Y�_��M��C�,�~;�I�|���-�����w]��;��IW5y>��j܈�ǺPcV*I�Y� aV�������]�ߛ�=,fU�3Z�P�`������xj�։t�,�!+���i[]��!��n)% K��H��A���|�a:�D���(���I�qW�1�En Q����K�rC-=�eu�T[@����np;$ �E'2М�����VΥw��-�,��j���A!����>�����Υ�EP}�j���11�J� �'�w��R;�J�5���$�c>�|q�H������"��#J��m���)k�D��O�Ǐ^�������`2M�oiX`�y/�I�S	e��j���3(�˺��d��4�rJئvA�:�C��Zu�v}���C�s3���{.���OX�Ҵ�!�TK�8[n�@p[(�L�N�:\�k��N?v{��W??��9J1���aJ7P�`�4��1X��fpSܯs��c4OkH#S�h��v�o�Tf�Ul/���k�
c���]�"�Z�� R�>�L�%���k�6��Y\~SQ��T��a�M�i�
v�i�Y��Ղ�El9DԠ����A͝	D����R�B�y&��P�����EQ��u�џ�?S��<J�Fߣ��s'(icDՂga�7\%�پ���:iϣs�e؞n���{����Z��t��"�C'S��Ǣ��LJ#g�ak�����+D���0b㽗�hҸ����a]~��)�&\�(�����cDd��\����tp�n�g(���MP��c���<%��.
E�:}�c8f�ޅ���f����Q��&��������$��{�m��03��3�9�O��|E��r��.��5�*�m�<7����iS��C]R�r(�=g��ݍ~��X��W0�|
���9�(��y����x!���W�&��yG>��	��L���D?h��Ո9?H�r�4�ji��͔��&TMI��L�j�a�B�·zq˳���?@�|��L�J*,4�\9�e��fH�8C��8IlXLK+��sޥӲ�ϱі���I����$)�����"L��"����c�ut5x�JB֜�Շ,NM}��CH�v�+�j��[W�,�n(� ����pP���3ߡU�27�&���֣�!%iQ~���'��3ɨI�'[�� T�[6�C�n����E6��Ow!a����[�Ia���/y�)!�t���0���3���������:3���+.曁G�3��y�j�4�	r���2M��fk�Npd�=p�_沇�Ģk�N�=j�4KS��3��W]����%L� �z����v�o&o񾰐���GI�eI:j̶'��ZX�ȭ��؃U"���s���Ŏ:�y�~�#ή������������tP�~  ���e���)l���E�2���N<�?�4���[{8jmi���kQi4���w���ۧ(>�J��Jp�_`6.�*���_/T��-��*{3���Yu]d#�C�wE��'e�NJ��S�n<��Y�,u�����\V�`
~f4��7�\��u-k�^�W��d%2ΐ�1��nǊ��qA��o���C��}�@qI���,@(����-1��i ���&D�)A	�=ݫ��u�|O�{+S�f�p�TOFNF����]�v�m�N��W��lg�!)nF`W:���qw�a��qJ�InH { b�)��+��u���\�V?�xV[���@p�A