��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$��p��@+��+��S�x��n�[	�^*��'�����r��c���(��#�8мs���g���{� ��c7��z���#d��H��h���Ys؈Nyϫ1�Ĩ�C)U�;)���N��I��r�FR�lK3�H�K$��p����=\=1�	�ِIFR����l7���y��mst�@8�����W/C�η�؟���{ֿ���Paqx;{��a�v-� ��4��YB۲@yK�S]oh>��ل���K��z��=����(�=�X�IٓH�-�nEi�a�Ɇ#&��}��a���"���+⃀E�6�D�Y�38�6���Xl�rF�+�C3�>Uk���us��qL�pl1T���v�>�L�u�j,:`7m����c��ڐ̬�ߜ�8k(5��'_�%\�c��.mVl6�مeR��^
>߉��T�M���b���orF@�ؠ���*��@����+��F(�{I'��`�x�;�>z񽿷ݡ��n<j�/�L�:x�0n�\s��:�Bj��E~��uZ:�FM22�O��5�0��iZ����U��p�x�8r��M�
��z3���K�^�R��k��=�+���D�i6�j�9WoW���3V�k�Ԇ9�X��Ma'�1/eP��7޿�Q$Q �|�h�[e��W��s>t��xꊺ���54�5K|@�N�^@Xw���:��IX�o��z��S���7�x-s��p?�����"͹┯���~ �!.�*���td]a'v7nl��+�4����j��zzZ�WX��}�n���=4�JX�I�GD���t�j���@UF�����?Zz�rv��&��`s��w�BLX�7r�&��-r��O[N��CVN����JnS�D���	,?-����)G�*
ԏƁ�6~-(*�s���\�Z�����Tm��wMne���F��II�Q͒�t�6%e�XE���%�������X�(�b��#������.b�����)�/d�o�^�):���'����)wi�kf(��M�^��+�O��)*���0�\�����w_�~z�$�Wb���z��Qj�ɖ�,s6��{�!BE�>�o�`�۵�1��m��R�����R^�խ����:=��,}"�!G�ސ.ԝ��,HI�27{�l���Yq��g�Yy+U	�B+��>�	7�W?���1�˃�֑�{R7��gK�R��v�W���������O���
C�eq(�n�zqfs5=� ����;� �F�S��H��H^�,�Xv�=RW�`GW��D���H�2�����Wi�kM�R������A�I��?�!1�r�i�?�Xq�I�1�p>���g0�3��ߜoWȠ.kɼ��w��*�zc�i��N/���Ƙ��%����hC4��w�wͰ�J�I ����������Մ$��g 3�m�d�ϧ��gJ�_'�b:C�.�ST�<���m/e"E�������0/[V!���qG�}���`G RR�3B��	��,��4���sJ��Z>i�O�r}�J���3�
<���@�I���d:�c��Y�2q�����1�om�}�`��B+f	��P���ʙ���X"������g����O�a�"���5'�'Q�,$�2ǲ$ ow�.�����",��Wߧ�"a	U���~ƭ�=����(h���Lphע�G�W:0ʒ��&����b��o����%�pB_2�&�t��5��@�E�g&����Yx�eOq��b	���K��7��f���U堃΁,�[Z���n���pbD&��_\Y���A��~q1$)�Q�W� ���{ȓ&V�#�HU�s��EJp�.��6(�v�C���N�=!z�<ǜ��1/aooaZ�p��}���:��d �y��B�0�Pŭ�����z���Qe���X5�z@�2�jK�C�&�/�'By-���K���J�-�3�'�b�!�
a�2��:�j�R��}_��r�Kn�6�\K��{�fmg$5��c~��ψ㕂���W��Ƕ~�"��Q�iw4HQ榝6�Gy`��R��Mk3��}���J*Ej�_T4��1pi�[9N13�_�~֖}�0�M�Rt�(W��O��In[����ۉ:,�	����j[oLc�S��X
D/�m�K�;x�;��=c/�S��Ʀ?��40����H|0��qg�=?���Pak;�0q��d-��6`�dWĈ��H�)���{�qZY�[�]C��-���>2aG��*2�Ni'�w=(d�
��W�s����i��%��m�-�&2c�Cg�x�
�_��uY���s�څD�[����>�sј0�Ӥ�O�\��f"��4��*��{��q`������rY=d�T��Ĥ���oxt��S]�WLH�f�M3O���Ra�y�����.��4-?s���!78XV�\������L'sO���������s׵Qg���/�Vb�",�
I�9��{�J��o�u�ŦiL��w��6-�e32B�)�X~G��Ij��P��4�$��dG:�g$��^�y��A���	hf�%��'v�} �뫡%9���T�����/�g�U*�����j�x������:j�S<��^63u^la8c)e��f�V�v&��U�!�[�#�IJ���7������eC9��D>�(�>�O*���6�Z(��Kd��he�n��ڵ�iB$$��T���]c=��uɣ��MxǛ�z���ƮaU���ZZjWy,p�?u�S����]��]m��T7�:nҧ��M�<֓E�LO9W��Gc���j��OA��D���b���+����������f�#�۔J7OV'F��I�9uA�(n��A=��nŞ*�Z����6Kk��s�q`](dht{x�^�,��x-9h�N��2q��!x ���='�ش�e~�*wb�r�*��o�U7����%9�t�P�Or��2E+�`�E5-Ǘ��<R�m�ⶑ��~�i,��T$17�_0e��i���V����nQ�=m��v�T�x�o�$ˊe�rV#�[��Zzeڔ���?K�n�잏>�z���������Pʓzl�/q<��K<nh��T�ȽKra3��� 9L?4%��@��ڶ2A��%"���۳������nz\0$P���+1��*�X��Z��V�4�c��t�������(k(���h���gʞ�S����/w�}`Y��HF�o�tpS2�,���0�!��w%1�&��Ѿl����z�d\��
�����Fg��g�rfP�+���m2� ��r�#�k��*�m<8a5�v)_�)�]BðK�򡃱wjp��R�@�O_�A0�4��P�˷x~;�7fA���p̻�����7�,�i�tlc/�2�5E4�5&=��5��O.��Z=M���^P��gJX�?/��9PU-ظksײ�3tŒv#~p|F�x��_�G�{
nK�H�:�1ޅ����lє�d��/�&����z���0 �%�N���ٖEQ)6�M M��D�� I6��쿴��+��a�MU-$=E#Z�`��H[iV�[:�`Rc }�^�d��mh�@X���C1��[`sP��
V�Hb��~n8]�hA��F�㗉�
;�W��xE)]^����D4�e$��Lc�sOy�0Q�Ϧ�c8^�4�(�߬j�7r?���G,'i��=eB2,n���:i�x�T��+X@���
�9��`1TD��\4H���V=�ǣk�ii9�6���.��_9ъ̑8H���c0'ԍ3�2'<�f�b�f��Q�S*�t
�D�{5c��W������[���=�4��IJ� � �	.�e<�S&I��OVā� =S	��f ���+;�"������`��G)�A��D�Zr���_�l��pE�Q��G������4V����'����$�*�ѿ-�=Q;Y�Gj~[[������P�(���{v�Ҷ[E��aj!���,��<�	03������B8�M/��g/sc��Νo�Ax���J��ht���}�V�ͯ.���ա�ջ,&��>���<`
V{,_�gF�D�#��W�y�N�)Y��]�B�-��� ��*Ć��	���ǅJ��q�m?R���^��8��r�Pq�|��]��8+sIVih�]^΀�� �<y�1W�'�g�݈$���)S�Å~ylrb��gN?J�w�7I�#}��`�y"nZ�v�ox�LJ����@��L�z@@�������x侣!0��S�������>=-�nROD��"���od�������{p'�PVM�V�;�=��m;9U7��jCS5Th#?�5�1ɝ�\ϑW�;���F��՛�,葩���	8,d�����U�1�������O9r�潃n����6�*Ef�$��M��i�2�Ys����c5�.G������p��4r7sT$�s���@uת��~��S��H^Y"��������Y�e���O�95�A(&e9H���-te
���9_K{�V��vffn�?	V��U.�ܦ��ʑi7��nԄG�׀$�+�P�2��؎l��$��p�܉d�����В{L��<}����D���Dy��'�.�G8w�$���������[f���������CӪ�[KC�
���koQ�)�1^X4�gj���&]�i�M&Q���1�c��z+��/8��8B-f��/��WV�Z��hI�,sA��|�_�@�E�F�,��mk�=	D�Uܔ����3%\��I��*��� 1�y��@�ז�
��bD��y�WZ\����V�	I�9_��"9�@���Ũ�u-�����E�hxZw�h�Q_��'㝜����;����vr��?�_.�Z/��+'Rϒ��mt���g5����03���R��7�CϾ'b�qI�>6����| �	(S���l�@��͕]�V�o8v���;E��.Q��HxY���`�G�f�8�XsYH���&�;�l�0;R�P?�cAʮ_j�#E"p�eL��7/�nN��
G��r�zt��Bs��_]��'M�@��^�9�Xѡ� ���a�QMB(�|֧|�5,�����s!���W�;"1����*���=�e�� �Q>fHg���5�v9ٸo��s8�$*��M#&�D�j�D��SUG:�T��1�[�Prg��U��j�HR��p�hm�������wV�V� ���ֽ�Qi^��!�9�h��|��	�֦�2�~�CL��J�֦���ڐH�b���ݽ���i�4vpWcQ�?-�~�=������/�C��u�F�N�����{�P/ř�
�ͷv��J�綈�u��ww�C����T��n�.1>����j5�f[���d�v��s��ǒ_�%y������^�0���4Ǻ㺭wj�N�}�Gy�MxwU+O�l�a�,]Q��6C���=N�%| \�Y��|�G�E�j�d�8p]��}h|���$��;��S|�]kO i&�d�%"Afevx�%�k=Mu���t�~��A�Op���o�1:��#�D	�G�_�Ӭ���Gfya[%^�;�{��Y�ߒ*`�B��z�/�{�,txg��cٮ�V<Q���Ⱦ��Ѐ숊'M����q��٢���^��T���g4q�Z03���-2��l�i�獚᳁�_
 �@nWm�+��n5�l��ٝ����SP��#�'sn�n�|{G��U@k2b,*�"�l<��&��v'�C�T8����Į,�P��7$��!�� �`�~��"��KD\4{^��H7h����iC���^%~j������b���60��Z�	*�d?�]Q��j�j��{��oL��4@}���M���c�K����;ã(
�>�a��,x[ܿ��U����6�G�9ts>�>�:JoG�O
���n�J���kx*_���T5`I�!�L2 �u�KC�=��r�����o���[Fn{�z[h��v��P&z	�#��JĭP��5R�crO��v����"��~0[R9�y��>Y��<~WĢ"���'b���H��N�>b�{4�C]]:�8��f��%� ?�=������J��0"�Z��D_�d#���4����[�B��Mu�P�6{��� ה����jQW�o�6�T$�}8Lْh1n�*�����x@P�1&�Jh㿙�E凜�:�r��+�o�����);.�kB�[��lH�49Vaz��8|�w|k�9;z-����ɩ�#��c"����~���B�S�a9�- 0�7�܌��]�6�*������p3-�i�/��8
�1�~���S�,n@��m���DS�Z6���(����A�`��/�g�BLHj��~!P,����h���c�9Hbk�̨1��Q�r�<te���49�C�|�����H��}z?;Ç1`������-}ф�Z%���O��IJ
a�Z4a&-V��J"��̩0ݖJ��$Ն�r��� Ja�^��9�:+��,.6�}}��]u�N��.��Q����K��r���y��^� ��/]��__@dJQ�}�j��
�`8}{�IM|��?Q�k� �/|~�Ƽ|-禔
O�/E�K뭘t��-�]��Wlꋓ�oWp�.gUN�������ަ��I	���m�Z�0�t����V$����L��:�p�	�KuPj;�UuFF���8l��[�1�4������0*?��+h�?�Y<~#+�'6����
 I����׾&���F|<�M��R�'�Ǌ�/�(T �l>=�lU�΀qNf�>�J��GQF�tf]�;�1$G��ٹ߉��>2,_�.���zn�}e�K�:rS$��!O͞�E�g��1��T�u�����L�Վ!�����j�Z��� ]눦�&0�p�ɣ��p�H��fn��#^�5vB?I�v��X&����3v�'�=G����>��ӯ2nGX�'�o�p7�$����J��y/����d�<	����Ip{r�T�p&�m
�N���aK��u[Gy���u�%�M�P�����{�{�:@����-��k%
��ρ�pyj�R	�_a�E���Q�@�n�J�m�Qop1��SG�������R�sd�:_HfU,�}����8^���R���L�{G ��Ŭ��Lz������g����u5�e|n����&X�S�O�T���&�HW�(�+ar�y=8���5���
(nQ	���	|� ����ą�-
4y%f��濟�����I�GB��櫾G9��*���$w�{�{��0�g���¾`��x�$�T]�!�Ѯe�I��S����kS�u��ƝN�gU0/�p�ßm�{�ٖ���uP��DR���eb4]> a�@����3�j�Z�Ǵ�!��2w_q�Q%�yّE�����}��<}�ߗ��s���#��8Ѽ����aK�#�;pQ�\�r�kf���rG�\�-�d�_��KfV�
J���&�������R���!@L3�U����wX��Y�XWSmz��(?�k�z�V(1�1�6�~��:�?��,��'#� ��N�|P�^���.���Yg[?tf=�%.*��~a�9+�D(��[E5��2�J�����J��)r,V*�ʹ�k?���.<���×^�������;o.�hìr;>�	ͅ��+30�}Kĭ��j��]ɔ��"�J�W�
b}�7���׺	�ZRk	#ȩ��r"�	;?�����$��N�K]��y��]�)�.1�a��L�II¡�D|R�����s2�|�%i�cTwWߩ�6���.��>-����ҧ5.�Ҁ/��C>b��-� lD�����q��
�g�'.i�t��Z`m��Z.,���d h����f]��'%�e|�'B���F���$�#n� \��dv��A�SS�K�nGٞG���L������_���fhZ����y�v�\�i���D�}�(��_���!n)r�.��$�$�,�u��69�;�ዲ��B��cO�ơ�ى^�4"�Z�"P�=㉹z���s��j���	�ѱ&"�>��f��Efx�Ց�Z���Wu�|�����(��x��z��kim�'�S骜?x�ںl�*� Cwt"�D�������DЂ6�r�=���$�c�#X�@_-����=���QS��nE��\%�)/�.ca*f��n(��[`�����V̆Ju��!F���#2�ё,�0]�]^�$���9�h.{���	R��0mS{��aiD�lS�����B-[�
�{J>��s+��	�2���J�'�T�l��FL)&��LE��{\p��l�G��&�24��E��T��B���]�S��m��e-l79�]l��f]�7\w���m��,g5��?�����`��yv��,;P^���o��!�`x��R��- Aھ8�<�w�$|^�G>oS��|�aԾ~L��rw�<y����D�|X(Nǝ���|ewM�}3�{�|��L���W����yF�����3���c��ą�'�B�6D#�<��<-
�y��K�*� ����Va����~;"������/��iR�?����s�,�.��v��NV��p�_��N�J�uJ�f+j��)�|I��Zr����1���$j���Շ	�uԼ3՜o��Ů�T^�!j�K��a�	���"�iH(�?�d��Sqk;���/�j""-@���-��v��$è��Ĭ!Ն��]�D�L:i��kfQ��O��l�ԁ�M� D��I�yw���ŏ��g��y�0�u�rM��౔�m$,y��^d��4@���3�8^S!�D���[��j@����Y����*��~E��,d������0�h�۱�@e�=������-�e�7=t2���;�?�;`��Zď�ʏ4��q=g<�[����a�(���a�+S�;�nvF�j>��7�b�P0��H�n ]��rR��TAa�h�VL��>�'��n
9?��Aƽ��tN�V�Hx��P�����w�X5*��� ���k*�>G�m�P�D�S����/��ͼ�s�����	�0�o4G��iVE]�Z�)��,���ݼ꥜8r²Y�@JI�>^���IB���t/W�3w�����6����j&2qN�x�2�7wi��R~h��������~7.HW�����v�3t�PSc\����0���˓Z:�xb��N @0���y2 �ͽ��y˹o�:(ɟ��̔'Ȣ�C<I�X�})k�Z���@w6�nm�

,��3 ^��'v�Mۦ�X�O����Q���K�l#�#!#)��1KP.�X������eMV.�Në0�I+����I�����)3Kh� �>��=�v-�Dm�[~E\
���fT��V��E��nm���s |
���]����MO��$	^<�t�=�z:�ڋ��R��6�.]�@J v�Uf5��`�/��v��|�	�#��P||#��*���v�;ά/3{�G*��8y�ؿ��m�8����|�lOI����<~��a�:���l���-��O�/�|' m4��~�cPKB)�x��G�l�~�,HI5�����b��������M/�ˉ�� uR^������͹�J,�sU��,}MlC�R2Q6�hOf������D�a!з����o�PP˥ӈzF��\h%k]gm��<S�(��<�LA��!��^svڭy�`&l*=��G�3H����D�k�Ǡ��K�Y�3U.�>������E0�$0��m�B��.��Z;� ���Uxoa/���'��'X�����f�
�6�1�G'U�Z�e�{�CT�m��f%���:\�R܉�A�x�e��
�uJ}���
�gbߒst� ��1�3��G'�DX��p*P\l�	Mk��O+�gU_>�u1��H{ �q�B���g�LB��K5��)�#K���2���^!�&�]�2`����O0Kt}N�D���:���$�-�+	l#ǳ��O&vhY^	21��S`T]���.��ޠjч?��|��~��������;���+C��Coy�3�o >�}�@��z�0��:��LX��LLy�r�8�26�IY��{��MՉ�4~	�����d6���7�2������.{�p��E~V�H��#���V;>'����o6�M璚����I�z~�O��Z�D���퓁��M��������E��e�d�n��������}�D�U^�R�֎�{�����w5D}u��Cb�m4T貎���iB�u'��=���H�#ɏJs�׌��J1�q����}����<��p�t�����#�p^ܺ��l�8�z����B��9�Oٞ`ƫ�.F�˴���hTh
�(�A�eI�����<[��ݽ�Cj��x!�|������ש@�n�ݛ/=�����C߉���O��W��9���D03qG�*�E�S74����APCV1�s���[𺙥H���4����fr���W
J�]��!z5��Oa���t^����z1ݿ8+��	�n��`�Y0tA��'��N�8�p�g�X�HTX|-����&ρ\�w��Y#���܆С�����k[y�daB�?��NԳ	�Aq��$]�)s�6�R��i�T�R^�mA�O��̎���
uOK�Fh&9�\�l[ZЀɽx�E�n@�r;��zyl_�iY���/�P��0����O���4f�]�����4._�Z�������^�|3TkĐkq��������Q�}��L/�\z�״&��e�Ħ��jh��s�\h�>�����H���RvVȶ���O�='m�ʻ�)o���O�/�ѷf
���ì�,Yd��yIJ9Pw���.�>`,��y=�_�<�Vr��|v�쨽WkKG'����g�9�
�~C]���m-��j
���.�� D���/�)�a8��$���8���皖��E�և@���d�0��(Q>���(�*��!�dL�����l�U�,���%�I���o^ ��������ЧT[\�e��!�Ɂ����� �Gf�c���K^=߀��m@y�7㳃��y5�>�	���pGm9SEp`-�Yd@_P�Sd�nq0<�I+��&��w��#g!Awj�:�`-l��_q-�H��0�8gm��� ���4Ӳ�M1��r�/����b���Ց}����n	�|�,-iv�7����O�WU�M}J����\4���ρ�0�e�Qx<�M�;����包o�EI��0U�kg/����<30�)�}�_7�ݦc̑�ؓ��zZ��6�~����r��P�P�:9�E[���d�>����O�9P�e��p��dd�U�*c�ʴACc	�M'Ber�{�����\𹹳}֑u��ϖ��?���Κ�5+�1��d���y�⨈T�Zɠ�][��;�RbJ�k�Ґ֦�\?|[U��ɍ @�R�r�XnF������Ѝc���2���Fll�7�(Ld
�x��~��J$^M���%Xxi��?o"<$����E
5�_b;�ki���|w���7O����4�S�M�I���-�"mdh3b#4�*a<"���֠���{G���ᵰ:��7�E�/*0DZ���U�<l^ځ��ܰcjf�y�mܧ��͛	���f-&Q�֒#��J�����*Y~;�%1���0)ָ�L��l�6��8U/�w�y����`�K���O���#����=���w��g�()�� <g����|�>_��BϬ�'�x0�}���痫��2F�7�@�$�ۗ /y�~E�-��j/�i��J+�BrC����=9�Ob	�ϐ�M9
�p��1w/�-ŏ�I-b)h
���2	��Pɺ$�P�s܄蜐��4�-#t�hS4��� �ha� Ve[˷�;�����6?Bt���H=��w�m�x����EYWw"TՋ~մ����K���H�D��Z��$�H�������g������xY��8Fy�|�UO\!�.F�_�0ꍽ�X�n�<�q&,��%��a���7�Q7�6�j������ܵ����wW���r���CPJ5�C�XXԿ��ߤ[��1�s�Fg3��5��j����&r����Ffs�<�c"$?w\�`n�${����2��@r�*��;���A�8NgN�d!0e�{'���inN��d�*��f��/I�mJmfPӷx�3��*W��V�+��ha�"6R_,ɷJ��Z�M�B �|��v��4_�'D!�������8a���}��ܿ��R���������#8Xa�թ$"C$��U�����raU����Bpf*����Ss���>�� �f�Q�$����������D���3��D6��w$	_��گ�OL��gMS�`D���X �ql��*񆀥�����cr�i�r!�2�����[9��X��7�C����l�����lfcW;���1�؇exj��,�Ys#U*���:�	g'X�-���9�)��rQ�+��$��f���6�*���<��O��⼚�_�	�#'�>yL$�^�K�ٻ5y��j�MD&�&���*t�V��_H��Æ��l���q$�b�m:x��àz#o�wt��N^�(#������,�?���F'x������s���k���0 H��,��N�Yn"�9d�q���%��S��{^�r�ک�
�-"]��P��}q~�2�~���&�j���QQn�?���wOD�w�)����Z0ͥ�Ko'̙���/\�B��������6�^2Ԟ�cB�z>�]�Y�G�T���� l�ku�+	+2^���'lg�L)��s��_��.�*G8輪=�҇�ؐ���^��-I��;�7�#�h3@6g�N���}��Ya���rps�����,O`Yʌ;C���k��lÔ�:n�䍢H���&-ƿ!հ��I�԰��_M��BU��E���Z�T:4����*�8�MƦ���Ko���m�nX�� dcf,�a���['��HJ����/�m8����>��"��=!�ˏ��Iفa[�O���Dd[?n@���Sޓ^�,+��y�Ͽ��c�뉴��Y�5��K�a�В$�Z3��}���>�{���
?��땚�
�{׹���۫��ҡ�g"|��I��x����ExE���@��w::�����?��f���;m��i�M3C��A|e*I��x&_MS@��ϐwgX~�kn�{��B�����2��!�"c�ϙ�e�|��XD�j��Sf"���|��_�LCXK�G�j�#��sa�B�lc�@���x�����(�I�69�f�8F|i�D���ߏ�1+ �ʾ1M�m�^$�����%1�_~C�,�%'楖��O�f瓯Q�YM�kY��u�	��8x���ř0j���1�$�J�3�{_<�i�2����,����?�@��D��᱒	$�U$���U'�Q
�,��2��`�H5�H �d���y���k��T�G�����C�r�uB�b��=�z�E�9��*m�Wjj;Tf����Kh������?{��Hu�_��)��S^��a� �8M?�>N5Df���~�3�#�3�z6���A�����'�W���������["� �G�.�H��,�m�.���cW��r��brZA�`6�C���X:*\�RJ]��<����ǯ>Y��8�؊J�89X�K�*����u ��B���-�X��R���"!�ɷ���!��{�w��֞)H��F��LB�C�ޓ��ag�/���J�'kx؂I`1kd��
��*[z�PU��eF�3�
(�`?6�ģ���cm����$�9#b���0����D��Z�0D���m���4��z�	$������'�.��P+@ae�/5Pr�2�߂CR���C�3�F��A�	��BO��X���@��u�C����o���%�ё3�`P~Q!����;i���d ]���4>�����2)��x�>#]�;.y�>#7��}�%��7×�7�b�X��ȅ����y���jr�k�xǅٙgl�;�1� �����>���T/q����	�,�{��I$����B�Wk�vTo/.�ca7�c[��P��Ö�gے6��s����6���\�-��)MBވ������ыC,c+����3�"Q4���S%�|�W&|	�,���8^{��jS���nO����1=�Av�CP�܃��_7a��x�6����;L#X��u��7���s�]`�p(
)�K��X�X�uK{�K3a�G ��ȏ�?�#�_ak�ș��J�|�$�x1���՞�rҜ��Y��s;�+O��I��b�|B�M�{P4l���A��SH�&}W�b5)՛ew�	2�.c�&�o�$��|E��Kp'�~ʞhGzZ�-3DH��	�k|�f0���i�����Z%_���H�8�-I��H	�2��\S��+���&!6�)3X�V��u�]�c�<*&}��j6-Enapf�����0�8��.H��={�Cmq�ze�o�a��!c5[���Kw�3x���n��` Ɛ�(/���LWq�i)��h��S��N��eP�ё`���ifR
[sM$"5�t�P���n΀?~��UJ�"v[��c�M��SL�u�qP��8!w�,��^���� ��=ڵm/,5��UPUsR��ޖđ^�xd
��i
��?[>�]�f5[�r7~��ų���i�&0F���.�)�u�>Y���ؘ�%T�s���3�ǦݝT\�:}�L0�չ�ƛ���y�˶~O\��.^N���py�V7�L�c�$W��6�������}+�B:�6*Q.��MQ����1�xS�w.�]�i��V`����*)K�Ų_�K_	LQc�JQ��<q�