��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�J��"4�=�7(�T�JѺ�ő��,\��s���ӣ�F�؏�+S���B�g^�h�[�;��Љ��P��iԏ������~����y��UU�MΧ�:�a�[��m�����Kz >�[�z1���y��L����G�j�ɽ!�v���?���k�3�����+�D师k�;�!� I��߇$@4[LVY�����22��fav4ߢ$�2�u`oݗ�{o��,�`-?�:��!�x�Ė߃?S�a���6Kɲ���
�$���۴�[���ҟZ.GCY}�A��ϒ=A��{�H��L�SZT��a��cm�HI>�ŝ��H�֮�/+1{�W��.��Q��qm�n�����\x8��C�'O�s�������e�࣫9!c�СJ_y�E�Y��{��h��÷�c�W�b��2b뮲d�O�����]RZ�[�7����lM��u��X9Q8/����h���o�(l& ᶛ�8��˜P�'��؀2��3`�'Ѓ�z�Bl;�
7Е�fϵ����a�G,
ݬ���߅n/ȜJ���nW�ؙ���q��ߴEr~��faP?���/��Y职�x)�TTX%;�^�����7=o<�U�m�h`�5��F��5��im��C>s�(��O�>-\�\! h����*�k h�M����8LtJ|����&�vބwS�T<,ia<�A}�.ut�ڰ���.9^�br�����R\�k�u�4���/d6���d�?떩�
/�Z����hޟ2�O%�^)��2�>}�>�+�s�n�w��l �Oz}*A���b�)K$rI�ρ���Lb[;%���k4�f���ॵ5=���mGբB�`yo�O��	��O=j#��}w���32g�œ_���m��;�U�y��O�_I�9|�z��#���u�S��or�:��|=RjOF�����@)�	��>k侃���b��Γ�?����m��O�:�Z����lڔ���v�i�gc���[�����d���Kh���h�IDO�I0���I��d��k�G`�֯��b���~;�i��|�r��B8������σ�ԛ��������^9i���^�0�[�����\��H�}$Z5#4�M��m�R��~?[���P,�X��V����(�H�鶞�w�:;���[���┺��j���͢z��g՞D�R�ú��-ß�K�C�Q&�wM-#H���Ęb�ض�<ڗ;ނ���!�W���2��%�`v���n�[����t��.��Z�8I8���F��80����k�<v#/8#{4��hÛ�]1���z��J�_	q۶��y��-0���pX�"'^����lj��)?��IނK�a6��L�g�*�Vb�g��u<�{����6��T�0��m_:�Qҥ_+�����a�=��vM����y���":(�V_/lB��=2M�e�d<�_p�}��.WګL"�7��X����qt��:���!�4=z��Y�x�i�����\p	L�����!����"!�U�-Ȣ#�]f��c��$i u�F��[p:;=(�܉��H��{�?)�����ّ�GH8�@�Ŏ�B:qs�1]Ֆ������&!_]үV���k$�rb�'V�'va��&���-�V[�(���6{�:�/k�oױn�D��W��~�
���ނ��?+H,��.ce��b���:�G�=�F�{�vy]%���wH�3~�Ai���Q)aUl:s�}�<�/j]�u!v�Z��􏳽-N=��o��N�~cob8�b��k�;/�b�DN��x���I��;��>U7�U��ȤM\��@̻���0��/E7G�����g/(=��Ժ��h�]�NY�#�t�����Kv����E7���x�*�3�����B?O|���S�"6���s8?bm�����]�$Y��ԯ&1rG�������7��!�Q�V#Q$b"+��ߌ����I��	�Ҝ�!r+��`� �~݀�S:z�|o�ƊF��Zt�=��/��pR�����z03w���ؿ��,n_�e⪈�1�;Q��Y'�`�	E�P��ٕ{MyM�R�����̞�[Q	�zV��dJ#J�P,8���h��K���-�t���t;����|��❍cN^�%��Vr�sJQ	e�͚��,��u@=(���Kx1o-���6Fd1�pOB�|�D��Խ��Ol�%��M�9�L�n8^�E?���8��'�<���{��WkS�ڲ������ʲ\Nʝ�+�c�u �L�^�\;!�H.�q�!F���/{Y�e��V?1s���!L?��d��[���*j�����Z��D��e{4������8=�N�I�슌�F���(��^Z�t��g��{14��<����P[/�;x a�&��Xu�V(��K*�u'�Ը�X�W�_�	��9&�gD�<苯Q�֜5G׬���[��ς�J��)NY/�X�W��H����Jݣe�KU����#_�x9�IC���?l"��6M סy[�Hz|vp��8]sm����ecOSu4->Czwr��{���h���Lr��K��*�W��lG#�����K�0�r�
֥��$��c&�/���㍔�a?c��]����rЗ��.�JQ�+�F>�ʹ�R��e5�2���M�Tb�7��H�#��ּ�F~Ӊm�o���_��M�{H�/��NJ�b@��<y�(`��X�*��JS�;K��/�"�����n^?�[�Z�����ȍ�
�I�?�=��=��rb̹o�tx<M���ܾ{���T�/�؄$־���{1a����K�n��Q���3`������w^}?�I��x�RE�v؄M�!��2*�X֞����TJ�
�]S�2,L�!��HPڂ�u�Z� ����-=<�44�R�=m�C���I����hw饟7c{��R�־LR`PK�n��.�]����>�Al�m���TC+H�?Ey�ߣ��Zd�����U110�e*�6�#O�0���9�(�"gm~�%}��,�F5�G��C)Q������C����� hW��F'�
��𭃒a�v��xi�q��Už�����~�;6uN�/U?�j�Ř�pR�����i&�֒p���b�����UǨ9�$\��}��q����""̌h��"/Ӓ��f�q��/ш�0�� U�a���:���4+M#��V����x5�T��?���R��B��7�$�E��.sK݋��[�y$�g{�x�^���uG1X���yz�!�}9�?�֫W�� �}��N�F��S�[�<�\v�6�s�֐�\�{]�/E���-���h��vk"��^4��-��3�o�J���j��Ө�F�i�8�2l� �.C�y���O���Z(�Y'}�j�h�]$A/"��IS��C��s�D�|��2.��;�W�~�P઒(.�>IM�&�H����^����L��9IOT�������2���itq^L ��^S���',f:uG��#�I������s���Q�%�x�́�X������e�<�)\�J�Cls��	�Ȥy�q9W��2���c�$�Ö��4_��D-{0T*����2�)S-�ga��l�&�i�����;4ʄ�_�{��������á��
���
�3m<�n�ii�$�����ƞ$���H����X#};\)sr@&ӱ�������ur��(��9SdA�8�3��;��Z�'�*�0D��GiJ�<x�y�{6���$�=��3N���1�X'�����s��망�2����21��¦������٩���J)�K18��i���O�,e y��w_i�Ɨ�ӿ�OD��s�=G2P�<XSq�ɠ�B~Pb��7��s-�^�o�����U�}i�б�5��:md�sY���	xW�L��> ��<��|��g@�C�rd���-[�K��R�g���\�f�b}��I:�@%Ҽ��b� 9����e�}+�-dN�W�c�B��ފ �HST����xw�*x���09G
U�8u�C�,/G0�
�6��2y/ث�����Wǳ�c�i��z"�#-z1���Eu��?��C�����G�x��j�߻�)#�>��������5\^Bؽ���3�fn�.�2@��<5���A��������h�Zw��T������L�ɟ�g�S����ڎ�u_�a 'B-�n8�;sl����5�>��,z����?�Z��g��#������E$Z\�>d�%ԝwϱ��(�'f�ι��CH��6�Zx����궨`��S�H�XP��b�+Vt�+QHN�"N\#�N¥.'��Y?m���"�jr`�ͪ�%�>o��`r�|%FEy�LPyM?U.��x9�='K,`�<p��V��NP��[p������o�pR��n���m�:�G����g�����3�����iuB]��$vDⷓ�CK^�T;v�fU�q�#IQE�͘=�U?
�1edK<�e|��9Ed��l��]���)�s���B��)Ô��+���7�А%V�o�Y?��e)��I}$��\�����`�Nf�ɬ=@��g��P((xEU/À�h܄c�$��Y:L�ťy̣�x��Gr�"�U���q�e�S����o�������␺�� P3�S��x�I����y"������!�&�P�|<���:}� l�/��I�:�GD��(���1�m����#��^ѹ���O�k*�6#�=x�^������|Dw_�^w��ƨ�6'Ȣi��/hA�	��j�0Z��Q)Xʄ�Ӟ�삮VSf��s��R�o*ݨ�c˶�v�HJ������6E���0 l�����Vy�~W��u�-#��^�2�?�wL�A�M�&��I��E��o�\��}!HS�,0�W��:e��d�|SnB�%��x];�CE�g��K���\&�6{,�ْ�Zt;��f� ��tM����͏q���adi����V�ŉ�RUy^�W��޷0���:�OR;	�͋�|��L����G?Ԙ��:�W0�*�ȑOx`��2t,,X�i�A´DqZ��c�'U@���`���hhN��Y�4`J����=��p����9�=��J5��m�Uz-�b�ښ������<�_�kW��K�-�/Q�>�����L֕S}Bc�����|SE5�d�9��a����^]BW����~q��F�j��UZ����y_֖K"Ը�����q���;�!1������s��?�94���!����9�G�Q��0%��;i`��Fge��c�@��`R؂�c�7l$ $�<�!$Ӭ�8TF����C�����W��E��g���}J���.ɤ�}������W�O�ĩ6d޸���E��'nݑǌΕ�TDW,õu{$�ޭ,���#�V�+��	3��c�QF��oB�m~v��}�8ڀ�7	�)�W\�"MgC���a7�e�l#��|�0���"��$��B��N�� Z\�-�������n��!���"�Bh��n�LJԙ%�6gqR��h2�9����y���tg���'�\��T�;�}wk�W����uv�c���#�[����@kr����82�����5E�B���;�o���!�]�t�F��q�EZ��v�ZP/��C�L�h��d�\�X��^1�#Q��u�n�����ɩ&��Dt�u�.$Qf#�Oތ�q����A'�]���.��x�1;qQM1�q�B a�e�%������(:C6�ƣ��+�Z��Wzt�?�4�c�!q|-��ߑ �5�\��b�3�|���;(��L�͜o�%�]Է6M�iƞ���́j��
x�Q~������7��2�mԉr��?s@�p���>��1����x[�'~���H%�bEx]�d��x��5~����ஏ0f8Ƈ�|1�w�D�Ī>�����F�
:�$^0՛�:�@��l@Ϟ�o$8�����°"M|�#�7��g�B=Q��x���o�^`S�[[��P';q���H�{������a<ՙ����}v�����a+���s�k!�if��6|����m�����G��$�h'c�X�w�Cx�(�j+�����ܓ�\8��<����T?�=���l>�����W�_)���u����ab���q�3��x�[�Cr���'����kq��#��~�*�LRO	���) �P/Ҋ3ڪ�{|,Z�e\��8�#�C2$�[W������ӬJ�$z�vN�_��u�m��Iw#�P�N����t�%�{�:�2*��ع>�q>^�G/R%ژ�px����(��V�m�r�D����2�ity�`��~�-��oAO��C �"�~+�q|	WyA���\fk��d���S�jW�<��L3&�B\�a�;F� [s�#Lc����BEA9�4��}�e�<�=f�מ 'Sw��qϲz�~L��~���m��3�ҏD� x1��#����}�?�|�ֽ���Zi�
�����^[�.�]��S����)�#�J��=��嚬���3օ%-n籫l���PRTu�[����No�-� �8��)y���;2T�	���M{&�l=��ғ��N:��nտ��H)]�����ߔ `:���6�/�ʝ�B��C�5�[0i�L? �iY�I�gc*z5}H�?`��@��ԨJ��$����;Z�eH�P��FN3�$�2�gft���IY?ϻ���4&���<�qI1�:�UE��#wѵ������^�x&�Oދ�E�鍭�<�x�������U��u�
����q·��������ҩlk���$q4&�W�s��pJ q`����1��i9��!�#��\\�$��ǲ���?\���@-�Xg���0w�
��'�6��?�+�V��*DrB<�B�'3I���~01�8U�A/�T(/Y�Y�������`e��$3da�4=V­�ч3�68-*����<�wS��F�%Eg�iH�Mp�@԰�v��aKV,��T�2����Z"ڗ�3�g���훺�î��`&��.��B�0
�Ee�S��@q��B���Q������yh�ݧn�2�֞��ҷ��؏�gk��<��uV�ϧ�H�X�Y�?�,��#���0�AJ{�*rJ&��$��:��n�AFL|)m�٪o�LVj��Lw��JK��[����X���r���p�ٛ��>�t�a�$��:�Msr3a�`t�UN��+$a�-�><�Rϧ�����w�Y�jB�g:o:\�OϪM� (;oo9t�a�v����e�u�0t@߬�0GϜ���v#��b�����e�o��* h�yt�K������`��C?81K%ݰ�pG6qi�7�G�Y����=�SU��~g���6���ٯ::U~�<�i7X�ML[��x�I�t=g�D�ve�M��'���+κ;1�W��Ȑ`ڦ���>�d;�0�p�����gl���;Ja�R{&ɘ��%�(�<!��굩Z��|NI�Y�χ��|]��Yٜ��B��`���K�J)T+�b�N�4%qpZ���c��%��D�خ��ڜ]b��o�����t�/Q`O�`��Cg_��5*х�P�M���w�N�Z�����͛&��R�
�tOʡl+^�D>���Z��`ߘ�8�:1$h+����;qT�_.�m5�����cE�N�u����̈B3�j0d���_��9�"��W���X�� Q�|zW��	Q�C�.܆�����°�����AcByd��P(X;��I�Y-����T�N�#�ؠ�q���I|E��^E����h�+9}:�V��\�T�^ 'i��"&�a��kP�����NV���9ź��o:A��y=U��{S͘��G�V�[QF^@{)�P��ʖ�{�]���x�s �57�k��\� 	��,ٿm_�Lz��8��5���;ѿ��(9^����`T�P��Po�2�Ig{�gpbt~%Daf(嚌�MB�HU;�u:��7S7ә�������O�(lL�aC7���,�́.���q~>���N�]A��^Lr�s�_YJO�o���	�k1�p��F��5���س�E��'��ݓH�7"�v��(�H�3X/.����mc(������cY��4J��x>���h�
nD5�N���ѧ�z`u�z~7	��aU��S��Zml�Ԃ�U�aE�\>`\.��n�Q�N1����$��	�1���s2�R��kJ=S?�J�)�Br��ߦ��q*D�mŹ_'I�KফTE�9	���g�����:)ǧ�ޅ����8�s��?�����-';$'i8����-<�K-�@3�x|"R�#'R�'�+ĉ��Q>��"�$�	扸`CB��W�7����iM-�lf���h���u'�j3�ƱHr�k����Lz@�_��i�v��F}r��<�U���a\@�6T�k" mr�Q�X�j���Iޅ���|D��߲ˀxT����Ҁ[��rrO����	�Y���T��̃�%���I���,B2�$���At�\�t�[��J��V}w��*{td\��!�R�?�U�=QoՎ;g�K��|�����.���vf(�O:�� $R3#�~sB)�l.6TX�Eɔ��7p�����!/���/�)��<��r/�g!�Ac(������g�Y	�R�l���Z�Ɔ��逛��l��D���-<��]R2������8�u�6�H��3|��Č�@i܀�Ir�<�����N�K7�eE��S��9t/����(���$f|��d����qȧ�&�حl1oH�5�nj����Y�(v�k�{a��5m�����`[�=_�[�iT��k/ˏ����<����u���o]e��yd�Am�X`��3bg����z��ˎ��hV�0$��|*i����&�:. YU\��Ӷ�I���j�j�:'\�' >V�*d�� ������Z��&ҹa8��DL޺ ���ij�|4��aͪDY�*�����KP��ѽ�y���S����4;z��~"���� �l��ԩAw��5�	>��-x
n�7x&,���u�s�ٜu|�{k����ٮK�~="���B�w�bm��㲊����vѷ&�'+COx_>'�9�Bx!�$���Tm��S���{�(����ɪ�T��Ǭv5%��qLJ�4�߀�����2�qF'%�|&�b��'�� ��=�"n�*�oX����T����EM�0o��)��7B�����kYl��:'��qߔ��_I����6�H��LE1�,���'��?�*Kq"h�ɘ���:��o��ն�B�&nV1��3��V���q�k�׽�O�tpw$i�(a �V��'����Dm�{\۞ٖ�Ь;YG��	ٶJ��f��D��8��T�i&��b��Ȭ���P|�9�m���_ū�s���=�[Y�C��H���W��J���ʉ��嚓MC/�Z�l��7m�Ln/���y�N�n[����ȡd/� *?U��eSm�{�>EJ���5��r?��`�fC���s�8�d����(���N��H�ԇ��'(����o�df�J}pm�����%ao@��������7���XI$+������Q�jmP7M�FXj�
��T�����I�c�+~N:*���>����2��� �wn� ������_X~:��8o�Z��bM[��4C�m|r�/+��ZQf�B*3�.��������	G�=д���� ܒlYRM�a��4��3�a�t�QQ�CP��f���Z1���%3N��O�l���[MS��`�B5@��ϡ����� Ճti�D6�b�fۗ�0^Zl�@<��Q�5���U���m�6�|�;{pt�,�	G��D�&3q$����U:?��Ȣh�`õG��Nhh S>�X�z}��M:Sj��{i]*�}�t~��nZ�[��Yh�L[;ӻ�:5�� 2�i���ځE���|]$�S��G���d�ub�)(�+#�kbk�i#�X(��݌����>)�f��G������?���*��sV���6����r����}D'�K���l�<:���a��z����'y��\�)=<^	��h�P��?�N��6�S���UVW���1��զ��B�[����(o'��I��}ˬ��$���wASv���vB���E}!��p��T�AŎ,-�u.e�8=�Եi��v���I�?���y�������׿Nb�Ǵ��0��9�pu�>�&��'o�C92�d�jJ�ȯO������E��J̓����^o�byv�1��I��⌜�Μ�`�=�XB��{�CO�gj������@�xT�=�Zl����ߙ*�u���8Er�6X�}��R*�P�e��0��W(�갴�)��MP>�%Vri/}�a8!�L�3#CW+���q�E=P�c�?*c���M�wy^���]���?�c8s\�$�P�6}���xw�������b����}�iB@E�o�+��W�#'��|~���lN|c}������j�ᮨ�|��jЍB���H�-��$.4J�=��y�D�)���̾M6ǫdP	~Xa����\F�Zg�?�yrp���.h��د�J��W�W`�w�r����ᝋ����e�k�Ͽ������͜S.����b��c��5_�'`�����M�|L��b��o���&nR6�aD���A��c�����3|��X@ʅ¹�Ofc�
��G[����l��<F3�k�o��UBx^���d����Ч�֖��}��g8�C���Ɣ𹛔��3�����H�T��垖鏋�l�g	�WD��`{��7�ܰ0� �ܙ��w@�kk��
�6�V` ��F��S�ht!%6_	F�*���b^?��XS b~���D4M�}5�!��ws��J���>l!�s3��`.�_�L�θ.�������X�
�
u�X��7]tt0�7�'{Z��v�{#?9����Ñ� �)	��Iy �n�1Hs&�X�滠������u6�9���E�`���/p<���T�FѦp�pQ����̶��hz� ��V��� o����I����Q�ɢ4���v�L$8#KZJ.�9�X�TH�J�����+˲ڣ!�\0(�tK����ƳSV�)�5�W�0�u��~]��1�AinD6����"�Z�K��\�9Q	#­(��m�������p�Q��^�I��y�A>�/
)�j��JE�Q��nDl>7B��j����F�P��v�uC4�����'�nm�={Y)þ|��~�[j��u
2�P!�3n-]��21���	ܩj�N�E\�Sl}�.���]ύ���>��?�sNE�b���VPwE2��Q�~�ԃV�L�ma�4<��ye��uk�>]�PGQ�#_���:�v�߄���3 ��qٵ�;�L��'�H�pE�U��]�����y��ڰYtZ��l��ϔ�yc'��������ŁlD�9���29PtD�"��C|��%
�)A"�<���M4��ev��D�bv�"�"���=�,@��5)&�a�Üe �����6߱�����-%B�si��.��=�D,Py,#IV����}��i(Eݤ�z�f��].�����O�}>�%�^�og�v*}[�I:�:I��;���� P>�B������T�z���[�6������_2n����������$w#Τ�Ët�I��X��_.0��thx���yNž���E#;`a�``���=|ߴ�?Q-5	�?Ýb\J����(x>
��5��"���UpAK���kTՎQ�-!}���ˏ��+�(�W`���M����,e�$�Z5��7@>�p�mNЙ�z��ϣ�f�dH�oy�[u��j�'��J�x��g�kL`؊��RԪ�Z�bҷR�H�6�]+�h���u=`t�?O�ʞdH�L�Ӧ���F�'� ���h�`�ޖ/��'"l��~�wU^`b��?�?O�����E&n-�OP7��v�	_؊L����a2��b�Б�ݢM�Aυ-��
�`���Uj��'jx>RY3���q��G�M�ࠌ]"���≎����9-�L��1t�;�U*���qs�4PJ�k�_��7��I5~������Rw�_���(�V>���%aZ�~��� �s�!~(� �^��}R���I8zSj��F|rR+QuML�n�T��	
�?&�6�&��C6k"��`��9�efZ@O�`�����H6���,�!���n�2A��x+k�M�Ճd|@�qĮa}�yF�Ζ=�.���C����CT��No��rj��d�U��=��M�u:YAm�(|�F �`Ɋ����yrR�TY�a�q����qˊUF�\T�[��NMB�?ܨ����d��N�.
���:��KcOX�N�Yl굔V:H��2��`k��a	?ө7iâ��g|���v���Mmg�U�U�M���8�+��X����G���x��~&�w������du���ژ�/(��y�蚜����|:�*����kˑK��a̖�_}�ض����6���e��uDVۀ!���_I|8 ����ǭ�W#�\��ϝB|���_���@.`�dI��|&���.徝�`�kQT	"z���{�^ʜRG˶:\Ͻ�]i���������� �ʑq�:B�.�o)���0���j���Kmo��6�I���z/sd�@Xd�?s��h���|�\}�y�w2 [y�(��e*{P�X	���pt�9�s��v|����U�_��Ry�]:��cK�A�t�Ϊ����5���!
��n��(��a'�xP# ������=H�|�R��a��1�`?6yUЙ��/L_��������2�Q���$4N[u���=F��"���*�Co���3犎�����F�9��H���/�Ү����-cօ���!��pDet*����O� ��̯��2M[|.RL����w���F@�{�n��X��뾲���BV�иjР���5�*+���K�7��q�̴�9_'�֊[-myvd�R!ĩWj�-�2���w����䲷8�I��Z_�Y��!���ӿ�f�5��!q$�
p��׳�0��϶�wm|�|I����V���/�����E����}CA�H ���dUcֳm�Xo��ج�k6~���o�TÒ���'�;|�Ğ{��}��:�J�����k`�v�Ӫ��9�ܖ#�U:K2�#�x�R��#���oL�>���1�4v
M��0����}pJ\�?�O*""'�@m̃j�;X*?����&��8Փf��A,id�O[����D?S�X�o��	��ĉ�z�U	vJ~�T!�y������m��ͻ��#4k�a�Sy��m� $���_�ݺS���b���)�S���R)��n&��	a�(l����'i�Fy�d�/��W���DI:������7�>�� �Q�Z����jl���H��k��C���Z��\�8����4�2�#�.�ӯ�4t%� �q`�����3����}V4d|��i*^.%R�L�ʈ�g�n��L�L�C�L�0gq0��2�p@�_���Ȗ��V���,a�^�����qv���:y��g�X��@K���ո'�JE��S�o5Ey�sܣ(�'�J�P�K�}GaA�� �V�V�!V7�3�Ѿm��NU8)�
�=uz�D��(����5��R�)�u�i"���O����D'9v͍�`u��?{;؊�6�r&q �ZR"d���X�޷D�͚L�W�AO��'���j����7�;��]U�oS⡁k����D���cq���a����Mѯ)���|�uO�ƦLhI���.=�@��zP}�?͉=2�΁�Q���;%
�=�'
��7�2�N)^h~ �4���C�������=��1�#�KZ�Ž`�{����+e����A2��+�a.P�`mP֨-G��\�7ǀ.%sŴ�	ʕNח�&!;�_���4�p�9"x+k�(Tt"���V%0(��wヒ*6�	)�ڬ�;Ϩ'#䵃���^�Xud �:3�M��%1��՛�����Y�ôY�����b^h>R5�DQL+�-Li�.�I�=����Y���$�5��i�#ZX�y�)F��kIu�O��m��ʐ	��{>Pt�]��Z�0�� ��%.�<���ߓ&�\��w�ox.��>O�x�l�1@w�BjDs��b�4�an?��+����q�Rކ��d�/�d�"�3/ɿE�NT���8g�@YW�"#2mG��ws��>��W����u�}ֲ�.�.���u S?)^s]*!M�����R�~��~b[4�E������:d=fB]�nXj߭�ȏ�Ċ����1�_�r&
xj09׿4(M!97e)ЍW����"������R2	N_QdI*��J�Kd�	3�pN���rb�L��lG l#���XXJE)cA��Uf�}�M�2�h!j ��ۛt���6��H���2��-��a�׸��~c[�j�r���J(�����ˈ��:uF��R���Ef�RgM���#@%�����g���f8Ӱ!�k�"�*�e�	.X�I�]�m��R%A~�'M�ަ�3FhF�-8��(�s��:�)=�9������n��{8�f@�Ʉ�|�*%#j� |7��!�����iÉT���*[�����F�+R�~'�D��/�WH6-ѝ��
�V��)�d���fl��P+��k�/�Xʺ2pNdY�X�����R��k[�mH��:L�E�.:	;���]�j__�a"�Q�*�L.���&����{m�U�T'%(dOC�=u��&�3����*Rqo�������B?S<J:��^r��m��iU	�?*so��_�n��{m;]�����:�z������%�������C����TD$�$��n�����s�l�7�uXq՛,#+wOf�t*n���9|���͐���S�\E���<���t��P�"���"��G���lz�Aз���\�"l��t>���~am�.4�������Td�cp���C�i��4�˨R��װ_Ƕ4Z*6m� �nIN�b:B/ɑ°��7q���Gc��G�rK��,/���zv�?~�U���L]2���D��Wv���P��)D�N�����:o�C�3���.�b%G�=�9
��R�p,��D0����c���+/y���N����
�}����~�9�������h�$�K�Ǘf�[���u.U2Y��;�����Ǫ4o#mȵu-O-�p9]k�Xr1�F�cc���H'J�pU.T�X��!>~���՛��m���<� 8`^=w��F�jL�b��E���Hz�6�Ā�_Bo۬Cv{���#^��%,��2b b��dy�fSM'qUs<�,>�U�,р���!hg1�i�ўd�\R���%X�S`�U��='%v[�ڪ	�����d���I.\P�H�����>��`o�(�?Py�+)�"�;�+�4����-�rYn�d�}5�D�/��(���3�h5]��Pm�,WJ:�I�+Qs�~'�	��ߗS6�Y�ϰ�*�:-����K/�k�� 9���T)��}�r�>TK��4����d�rHK��	liCI�|NЪ7�2�R�  �k0�U��=(�W0?ڹ.u�h���x<�9�yպ��a\����3�^����z��x�_E#��>1��d<�����Ƽ̈�.j�����+�x���$����M��+i�������6��Z\�C=
"��_A;�O�&2y����R��B�$CE
 \]�m[^T�a]�A�Q���a8��Ӊ6���m�Vfȴ�8p]�3����^D�;��$ᔀ�5����t�t�WN�ݍ�3g5���j��_'��ۅyı�ϧ\l�\��>��q\o~j߽�Ϳ�4�-`���k�L��k}�4[3�s7��
����fՅ��١�?@	
,D�#�3z�*	)��yҳ�nM�J2@ys�f� I�
��\\�V@a��8[&��Z5��㍻M�J^��<�Z��!�魨�~����9����]g�S�˛i-H��5�o.`���=7SF'9� 9:�3��K��UK�ߣ�X5�u�a��8UBo�5������d!c,���h$�#7M�%��箼>�_`���p\g�"tz�i��Z����Y�6L�Ķݚ�>����b�U��v�	G�np#ɁXv��]�s���ޡ8"���Q��ɍ7ӫY��&���89bϨ�H��SW�oO,�y�g9nP�$�{Z����`�ݔ������e:D�Su��?<�$�KC쓾@1^�Ԩ�.ؐ�6����(�ZA�O���e��*x�Ɯ�y��=���8�8�fj�@#��k��U;O��64�ܜ_[�q�(�>���|��?F���z�U�	w��F?q�^6�L_�x�՘�m=`�jQ�8���~}+s�����3%��u����s�M�x�/����O���i��f����Zō�I�QVр���������ڤ+g�l)Q�Ģ
c��{�v�g"x�@.x넎)��w���Ux`�Rܽ�^��q��H��9�}��lP�x�i��uB銲|��5՗���>Q��:�s�o�w^��"�y�1���f��
J����!U!��3rN�� � ]Q&C���˴A�uL&�~T��EJ�,��x�M��I;�qw�W{��s�$�k��s+�"���<�3�X���֩]�/���u$E4�{ה����˾]��Uz��y@�����X�0��&GҔ{p���m� ,��?��=9�p����
PC;�>d�-�������1R֝?�`�T��	�L��yꖒ��~��*���^D�e'&�ΔI��(���g='�w'{� a�D�7�i�v��-�_Й���SC���TϘ-�84���?��V�[V�g@��ٮ�Q����/�1���,{�jfH���jX~!��g<-/���S,7.x�W�b�����}�T9������D�?^�d�����+������`u~ўG7���߷�</�X#<;�D�h� r(�>��c%3�Ô������n���O#���$��,�Y��]�up��#R~@��O���֢��e����03��˚#�5�'T�*J�|n��x��|����ǆ� Ş0�p�R?M����'i�l���X�8��[�و6H��Su q2��PK�wtC�`���
��:�TGЗ���,Qb'����蹻7D��x�{c�|�L�x���'���9�ّ%֍	�=C�j��S̍���oӂ�ށe1��W�P�t�cCܮ2�^<�e��<��! 6��.�q����v��j�ؠ���M��*k���v��h�MZ��,g��뙛�ZtLI�?��%����w��ӥ}g��L(�v�o�%v�]{'U>����L�/e+=��*;٨�qt����iA���j� "Q[|�T��0*�,����� �Q��tcw�V�"%R1�]��C����+��n���ї�{��4w:���z�e�Ab�>�߯޽�ZJV?��vuȾ����CH��2BG�Ax#�m���}� �$RP/�kz]��?�ڑ�I�,�Z��7!x.ei"�x]B�@]`���J;P@^d����_�=H�����5?��`��#��"�u��u+�*
&8]�H�3p�mR���]��[߸l����2���ųҹ�����C$����F&Ѡ��H@������]��@v�L�J����Wɯ�1�{L2W��.}"t�N��.D�f�����څ<�nT��Bg��j���&�����
��|��n�/b��y��j�3ZkH�+���1kN����j�Q��Q�AL%Ŵ�G�q�c:�Tb�z�e˿W���І���������Ѯr�5�H��_}�j�[1�33n4Ĕ�z�F�H�:B�4b0O ���������ݗ��t@�RK�6Ϊ��^\1;��4��V_Z�8��[j��q�av�VڸwWI�<Z�9dg��D0@`#�3~��,��$s�����.8����n��j$��K��8�Ȁ������������3��<�*^zu~F9؂��?nJ��e �n_� }��ǡȻ[�!��/NkX&��C�Z`�%혜k�-vzu�ĕ�+���.�|��5�K&����Xg�X9g�TǛ�d,G]�jK//��>k�A���A�iw�Fyc�V��/�2ɬ ـ>,q'�º�׺"��F�i���-��GtA�D�a7n��
D���  ���ljr>;�	j��?b��TQ��U!b��
�����^Wz�e���/�UW�0ӽ}~hcAg��W�g\�`��]&x�̽ݩ�/`��Q�F���BN" �P�p,��R�����缈�*��{����cX�I4�aI��djzfy���vH��},��)	����2�;��������󼼣p��+��#Z���y.�
 |�^o��X��h��"Po���%[ yT��':��*���C�Z�߄�`Bߠ�s�	�G�T����*\��=����"��,�f]��"��d
:�J���t�Ԡ��s�$�u�3$/=�s�/l�A�\F���V�ګ>b�hl`I�s�{(�#?	�Q%��!�o��jАY��s��;o�00[~S���U�o����Ҽ+�^Z=y�Ue6��czDX5��ߍ�J����@˕�^�p�'�ǎy�ͩ�*���O;"9��S��P,�B�Z�+����n��<�yV�J�E�A�)�!	� �M�l�ä�B�ĥ�J��̪aVҫ
ć��LE�3�=��|Y�k�'�d5�c=gnWkw��,S����6oS]�_b�.T|��*908ڳ�@D����_ɳF%v/�K�[Ok�pV�*'�P	}n-igG�^���U(�<�� ���;n���>��^|{�U�ղr9;��H	e�Z�K1���8M��l�R��|�)��$'�ҋ�bvju����=^���ݪ�-�y����q��>o�i�8�ɫf��:�OH�3#�B�UC�8x��ꉂ#���}2���a$���Ҵ�1��ՂI�zs!Վo1����� J	d|�u�'������Y��1�c��g� Ln�4����y�9�ꍻ���p8�r���0�WoV�Џ	D��0j�S�7��.�ݺ�)~�\�Z�Q4��!�fX��{��3܃�Ua�#B�ز	�{ө`V�;�����,$�B��w��w�G�	�B{�~x�?�@��G��=Yf>t�[I7܁���'�~2�|"��C�08�u}��;X/e��y��k�Fh��UB ��b����d�	:U�� a����M�������,�j��{���kǿ�dGz�&��#�-E�$r�+����ۢ�?��p٥��+���٣�+|�0�����b�=��Z~2e�7�ҘEK�ųj�M�zH�Ǎ�:3,6�i�;8�Xso�����e噔���+F�f��d�Rp�v������vRt$��o���YS��Q?]�F;��׈�յ#s7�x|L�J5�/Q�ʁ׭���U��5��(�d2��i�>\�1��yn0XI餕�?嚗Ħ�Kֿ�+x��
�b�Uz�?f1]��y�J�V�X>��<��I�A)a��!p�my�L$U�mxc��{<`��TΎ�����Qt�b!���x��M��֮�LV��)�dRC5R���y�w���B�ZuH�)97 ��;C
�U�;z ���3��y��A���:�uDǇ��5���)-(,'G�9Ǘ���\c����ٯQ��[�R:%!_�a���+H Jt�0����K�P��y*2�4<�l�8O�\e��/C�|
�4��}S e��D���y�m>F��$�7-]��F;�6��Xó"�c�����h}�Ng	`	w�$bpI�Xl�����~�L
)�UAj�D�`�wC��?,��`Ծoq�?3Y������Cf�)d�mn���߀ ��xM��+�@�����V��\LNz5h?�]v��SN���3�9"��"\���S7��Α.�[{�ϥd���dI=z*֨����4��ֺ�N�Hlw�}���*P:����1����;����������Lf�h]��
c��6K�]y�M �j�M,�T�����e�^�[�u|�(�3DqgCm�0�z�O�|:��E�߃ê��ՒٟuM�ý0o����.%�u7T�/�RP�~aN�C�6YAn(��JYgb����?�K�yy��C�3�����H�;��v���eFWڹ��U\N�������8�f�����������������R?�3��b��WѠ.=lG���P}�����q��}�����}˶[xn��@l�jKI&��ķ��$*�m�}��x���eьa��9i��2�8�QS�:�n��浼 M6��-L��e*��/)E�A@�F�6�I��+�"!p�s�.oU��4�4��P����_���G�C8:��.�7���?�x8����ῧ@Q z�Ny�����*�}������> ����]�NG��u:Ĺ��fH�:>%Z*{�$���+B�#L��I�K^�Hk1V��c��p��O��p�i��k�zϮ��T���\nOysB�j*��t�j���5�����44�s%2OFOEjfb"�]_��-hkU�!n�r,m�NB�l���6�Q��$�8=�Hs����ͅ�n(L�.p:x���DA'�f��sv	`��/7[?��%\�� ��,�dB5NrRL?At���x�z�C���z����M�7�� }�0�G��dnl�J��}<�:�O�V���-��V����}�%[�Z6H%�Q�*0�V��Q��'J���g�tP�x-�%x��{�\�pk!�t���MسU�RLɪ�C=�5`�"ʛ���ƭ*6��5N �<�3[�މg��}�"/D���p]A9^�	3��o:���x�	���¤6�M�r���wی��ju�q�E-E����	$G�?2o߼w�6E�&A��q=�/{k�b���AF���!�[�|JzԶz֯���B#݄=B����6"b#(�C�v���ה��$�$��{/��d�-�	��tn�%��b�ʻ����#�~���j`>�I�WW��`NF���4�5O�_�Q �}1����MjaO�[�
��Eu�W���v�j�b0�D����_��嘞~uqXKؼfl��{4bV�Q��1_|2ykK+$�ϴg�lo*���2����7�?�L�@�����oF)�@wMp��h]]��p@Y�1���sH�I}b�{C��ü���Aw��쁉ȴE�0��|�q�%x�	oY�9��N �:��(�I+�M�L�B�)6��4źӖ����vr�FE8|c�W����f�'�9��8)-�r��j�GQ>��o���V�#��{��܃[����{I�Jw/O���֛[G��������r��jeq�/uY�SD �)ɢ��	�N��w��/T���xm�)��[p:��ο�n�B2FpAS�s|B%�B��[���q�fԑdg���/�pB8,?q���.��Xri��7����Ⱥ�f�h�m�)��6[����D�n~��^y3�ή��V��%�s�1?2W��@����Ȓ���Eq%kw*�(�Tvz�(���ǳ�OM��c��dj����o1���|�"�X��Ͽfa�tH%��я>[�}Ib���gz�xA�w+i�#������#�!�� �3�UҪ�-חǨ�qK�mf�#�N{i9�r���q������e�9�~8�F�l��\������H{�$��ܹ���t� ���C��V����Ys����M9�¸�T؉������Un��5�]��o:�5H~F�]�4Z�AݫuB�th�����ێ4�&~�V�����  ̩�O��!�W��V����<J��Bo�6�a�4��a�Vt8s2��E�o�2�t#L%n����pE���/�~([�#��I���
�*7My�����ӥc���<?1^�u��}נ�[ H�479A�Ǧ����#a\�y6y��,U���%4��̨NqL�;qv��eݓ�C��vgx��k�'���G<�y��B�O�("��.�TB��T	�:n߽	m��4�Z����k�1�E$4[�S�OZ ,ptp�Y7�B�mO�ij"�,uM�wI_@� :I`	�����N��E�JF!Ro�-��eX*�rL���U�J5����za�nO��ߴE�c�o��$ZK�4o�b_�%�FB��R��itX��?���Pu�d�I��vm=��qXS��D�`���oB�}�4#�<�E�s.�b�S�1s;Q�@7���7��/���h����� ��~�v�	K>�о�;�����	nY�{c��K=~�Ì�ȣK�{xg�^-��Fg^�|`��;�?��m
~o}B��EY�k�c�U��r�38�[��e�m'�/k��魽�1|����M@�s1���Y��������lq�I��.#��ͦ�A���s�1pVBk�n�e-@W%�%n:}�o����i�sy	O�Y���;
��P��3{���t�f��5[>�e�6��E�{N�з]v9�&���r�f���Fvr����0��
��5��-n���A�o3<f7���O`⊺����e�m0A�b�oq������Tm_��_�R�7�d�88a�+?��T��#���>�����^��W\��#lw�p����OhW;�K@�^x��x�����NQԓb �v�c�<g��a;�G��;M��[|��`{Iۗ �Xӎ�5�31y+�rU�+��׷*"q�a-�Wg��!L�羛p~��oh�i��%:wC�ހ_{kǵ�}�dV���c�+�IN$@��a����!ن������,�� �\�H=� �ڋ��0Gw���^��%��A��7�d��a�>Y�L�3u�ʢ�}m������e�ql�I�[��Ѽ�[�*��S���_���ӞE��`76��8G�ŉ�5�Ǹc�����,w�Fc�� �'�a�QQL��r�E,|m���)P��ў��J��CܩG�o�[z�XXA%-�,Hw9+�K�c>�y���(K�,�Jn�1���vh�.��j��Lr�H��/#�M�[:%�PQ�+!�D>����4��ʽ�4�:��]�jJ˽1�a�	s:����Y�K��P�kӶ�!��X��vU��/~���I���]�����B�a�<L��>�������ֿTQ#�Ee4�@Ka`�"�4�P�2�}V���-�,GF�@1���o�2V
�
�Gt�#���SrGz�Zr�g=��!N�npK��@�J]�fH�\,�#Y���rt�E�]n���=E=�S�[n��n�*��wx��b%�S�.]"�n]l�B���j�=�+VF�?
�7���v��0�����ҕ{��LJ,K�':f�T#~3�t�{�� �κ_��G��̚d��8@	����q�_HdD>f����U���f���X_��?�0F&�	��������6�i>����t�q	�ߊ��B�Ȼ���d	�Ja�������Z�6��&7�������ҎE���7����욦XE]CX�E"���@"���ReK!���)׋4���c�cf)Ҳ�(8J���yg� i�m��؆n6Yw�(�Mo܄0ؒ°����S�($I� �r)�d=�����SD��GѤ ӵ0��փh�/μ�>�=�d��@��i~^����h�Y P�������b?Ǫ���&�cB��y��R~����PP`_��F�E��	%���%��:����"�Iw*W/��1�Ur2�'\�g��d�w3m��2��J �������<�`����]k�ev��<�eT�����5[ Bw��\��5���R�$^[�J6xi������4�݉�QJ�`����~��Ǯ�P��dW;(�K��Mz
�!C�xY��f��X��Qh7��Ϗ���� `���&'��E�힉j9bhE7�e¹�>��-0�\ı���<�� a���0���x�Td�t$�gє @�;u���xK�/�*4�&��?�>o�S�H[��'�o	πG�0�����m�GV=���[/��~_/���^cv�o�c�p�1�4��F�I���w:��Nj��c��2���w1"�{ji���x쌯)��	3�	0�B��)DM>����TC}��(q��0	h�}��J�$�>���O6[y �Y]���w=��s��$B��]CLǼ%��~�L��f����	۹�m'B�e�XF��U*r���r������J�n��_�7�z~�lLCu
Q�qv�
��=�j�'����F���{Jv�����%.��u���݇i�����(3��J�uc��,�9�Nh(�8������Y��V�q�m�Wg�]��n�;+[�X�����$/��5�B�M�F��J�֧���o�:0S��~�{�����I6J1�9�1i�Q�ͅ��2��/N�/���K�&��L�,���u��4�/�I���D���g|C<2:��T��^�G\�3�g�'�"N��ǝ��b��tz�ݯ�9d�[�D AQ�pHR�v�����q���c���ذY������+���9���JS[����g��S��wZr:��>�{P�U�fn��JkEa�aR����r	�O�����t-�@���`|7���l�O�\�	�q2i2.H�������,�3�޶��.L�nX����5ã��`�y�"��1��EA.F�>wSɫ�,�$��0�ӺfF������?�-��-;��/0r�)g�･�u�����sr���uH��5N^�V	ҝ��=:�%�|v�IA��40 �s�b�ٗ.׭�����w��C�r��S=1�,gR"�i
v���upnp�ؤ9$��H��d�ހ��r�j�k(��}`	��oF\!�/@�!f��p��_�u�/� /�7gv̲4>`�`�9�C�Uc m��=I��1�J�"�M8�q��FV���|�kA[,I����eL���-���<<�_�Cxﲞ|ۺ���r�����m��+���!Z�e�x�5��t��>��:9����B
�n�ay������=��3�-,���ެ�+/��׸z���y���;��E�A��/�'��[��\��ƅvR|(̀o޵�Ug�o�7�صlǛ�3B���ˠ9��/�xtq�E�Y�<���,�����3�u�Z�抔��$oj���Ǝ�Eq�'���}�����t3����/��I��9&�m��/R�F��}+z0�&|����iʍ��f�-�9q��'���

)	�*RL��|g,���M�M�iV�cuW�KJb�M�"Q�L&f7��H��	q�"f���D���XH�ϯ�&��;B��Ȅ�7 �:���Č��6e���k�h��V�����hܺk/��{��/%��_0� ��5�V����E4�e;�_�ig�����]S_�C_<�Q�7���w/�3#W6��zR��C�=��K���ʵs�9W����8H7ދjfb���z�t���(��.�Ɩ���X�}���Y�4Mgj�[��qKgl������z���_���m�}\*��ռwt�$}�T�qM��07��kDNg԰�A�ѐ���|r�D0@0�b!(4�F4u/ō�N��rN3S�!��$/��V�׺�DC��Z�~��H�uᲟv��b��FG]

4�!�������8���\G��ٱ��;XȔ��.h����*0�D��`�5E��<�[�m�΁����ޭq�	ɤ�3Ų���x�	4Ïx���g`��Όɒ����s�鏍j|T�oY�1�ν�?2����܄�5�*�r�M�����ܠ/Rs�(�c`2��0�k4 ��\qLd��_M��}֔���4�>W�s������l"�ؗ~��^�LHp�;8�/�)G�&��-�bu�oB�>"�#���P�{�^���I*��M����>�3���Sk_�� �M�Ye�q�������o��CG��X�3�%��C�Ҝ�u��|קa����}e�|������DxV�s��	^ؽH����!d���ƚ����|
)��M��� �W�wr�6����|��:fC�c�b�$0�s\.�
�!�ʶ��$��D�KX�8{]��fI��M[ʢB��c5���C"�׫����Q�_��Q����3�>P��H0,�	�m���0�P$"���~��/�i�x���Gxp��>��HE�B��ɩ��f�!C�v����gA"\�ә�0���.���t���ԋW�H��O�L�8�j�6����IV	�u��G[����[�����W�9���h�eL�N$?��߾/�cϛG�wZ�xyi�W~1<Ú�^�$�$�I :��:���Z�����1uLd���5i1up�{����ze}]xz��� ZT��l���} ��Ԙ�1��*��"��0Uۉ���9=r��z����eOS�ZQ:����0/�����(��ڙtHfe7�3�q���g��*�ˎ�`�9}N2���+)�y2�x���~A�%�ht,CX�X�5��
74��4}A����W4Bo�įf�2^�.�"���`��Q%'v.�j�1#�8r�(Y0���pA�����-bE�hA��PI�s �0�J@d����^� ��������f�Wgwh���{[χO�T�M�ƊuT�i�U�����
��˞$�s�Z^c�3�ּ�9��C�O���	����+�;a+Ks��23�2~���{;u��џ�Z]F&�})�$$Q�V���H^��S;@�;ֱ{�~�P�9�2TLwv/J�j�e@5�_���{d����a
8��z5�g�$��5�mD��P�Y!���&|QG��۔$���4�R��3a*P���/��^L?º�Z\��N�c���w�P��,��E��o����k�FzI���8cKR��nB�od*�AZx6����ד˜Q�zR�J�J�i�3]�$�l�TS��J�BȱU�;�6s�v�[s�W%]_מ������F�7���n�y�%v�<�*W��e�O.dD7;E)��*�!�5c����P����?ȉ������_'��@��w�h���m�T���"�Y�����H
�$���R$xl���0�ɾ�vO��}ՓB���yq�O���]�^���p�\�K�]�ϋg�#$�ʓ���^g}���&&��]�mU��d�fzg������[�N�_�s�q�T��x��%��%"��*���?q�^2*�6�Ț� �	]Y[|�&d�<�ܫ��g����бʇ!��S���`wY�c`�H��W�\ :�� �l�gp�>���y�5D��Q�'� �����f+!-Y'�}���������f�BQz_x�_��}��)E�D�o��������rY�Ee�x%��(P#�Zy�[@R�p�|�8hq�oh���F�O��k�-1V۞+oۆ�K
�K�� :��|���p�>�� C篺�Ǫ�KԗI����V~بE�� �����	�]�\�w���[�ޒ-7L�rk��Ei���Kr�Yxe	����b^"�ޛa��;�*Md���j}"Z��>4���&�Y�v�q����s�<*:Da@����P�x�ؑ�*	�K���r$9M���xV�0��`���t}����?踧-$�ަ۰�S7�;E��M�#R�m�e�3׭��� �U+R���[��Sܺ�����ɻ{�-"'��#}A�i��!m��P�f�ʳ��wfT��*����.�]]k��Vɗ�v_�r�ͨK���u���p�2��k+	|���*���ac>n���j�m�(�\�o��O`����90ͤ���#�Q���/�Qt,��r�\i�C�G	v�mU�-�3o7]a"��e���J{B���,�o3��9Є.�x�����yy�׏5h��㙍��'�[�Ƞ�g��H�T���_;I�I�������k8T�D�y���d�x�,���3��?��R
�ux�'Nڮ7����k���#�Pr�t�,YV������`!�͞k�=�g�A���8Z:�+���x� )�%DVf.{�%�OP˺��ؔ(�r�R�^*��ъ��@��f�a�r��lx5&�MN�0�3'���_�U`�|\�V��{�v�e��O��sM�������	(�&`��xД��N�3��x�Kȸ���c]- ���m^dz�&�y�/��ݢx>O�̏7ix@�Ÿ���?�Uh�n��l� ����d<Ŋ�d���
����d}
}�R�����; ����y�����7k�z �,�f@�~�8V�ɫ��O�`��C�cxt�@޺��*�Ш���Vn;�����?��f�EξS�������y]����R��@0���p�zG��`
j�#��"3G��N)��C���4en��+J�!��H�頌��v\#��\��Aʿ&Q�#rٸߋr����x��ޭ�|M��YyĿ��ֽO���H!��θҰ.g�*�'���R䄧�T��F��{K���]E�*Ǐ ��z�J�,\����ҕ�_��|�r�P]��*	c�~��;~A�q�\=��c!�-����Ԯu9";��K�_l��5��z��ʤ�/ ��~��Z�$�zb�������/qG�rT�og���h$sfZ�L���L������~yBm��nJ�{����p�k�� b�6��񌣄f-�IĤT�C���o�s���Vr��%9�s�)1')�'����PCsj2q��
�˻GWL���^��Y7�5��|8�>���%垒�������ڂ��B���fe���@����`�V�o�p+�'_��� �o�����TD��Xo����My�{.���J��R�NIu`I>��t���Wh{�<zf���=�������*�&N@�Ӡ�8=�����!�����\�`�+&�\O�Q�4�������o�-+u䅠���fYF�{m;3�w��-?ً��*@\�jb�Wj#M���c����3ڡ���F�(El<;�����?~C֊��f,?a,+K�y�� ��f�K�����T�
`�:����溲�A���
	| ���g4�U�~�*��ҟ�ey��W?�]I���2��:��d���V�]�h�k3X�"�TZ��8<U��٦P����He��.�y�٭�
p��%���i���묩��Q$�If�?��oW��Y/B.�uFy9Uuc;c(�U�~�4�)������MШ�%w�H�%�S�`rqG��yl=��{���M#�;e�s8
�ץYֈ0�ߢ�
U��t�oo.,��`��h��3�}vy�������J_ai�4%����}�7B�E@2k
�`�J��GV�I�}P��7gǰq�}�E�n��?��K/"s���~.���&Bj��0��\���O���Ƿ��5�L]/��@�瘙�|�=��n�;�߫J�j, �ڱ����g
��dt�w;�����^����\˙MN��9K/#��a�+��v�A��4w���Cpny��J�a�[���@�7#��((6L$��q@r��ȥ��4�5ѭ�oQ��ty��ۆO'��G�T�W�;2�R� ���)L
qu` �8���K{Q	LG"k��,ź���k6�w�\w);���%�i�z������ঙ��ʷ������Ա�|3��<��x.���#���"*Y7or|�+�!����W&� �޳��;��n��.����n��ɮ��UW���@�S���BVIn�f����1�=u��j\��"��+�y�pigY�J��︱_�}������%F^w喃��Ӈ�_ }���/�k��H��2@y])���I
Mx�i|�L0���������yP;p��[�����;��sG{�]V=�6f(��q���H�ʸL2L=9��(철0��E��4[�-Ȁ�.��b&C&<���9�@=�؀s���
>��ax�B���&T[KV�m�Ȗ+���=t�ʅ�+�)��$pQ���!+�w�8�wXD'~����?=�gX���,����!��~hO��G�U(x��f�H�u������y�ȓ*n�[��X�Ϗ4��$��������c��˼����$,�0P� �g����r'KGv��HM��
�?���䰉T��/n9�h���n�b�}UE����_�>�@),�+?�y?�����ɉ�z�b)���f��5IBƎ,[�WZ�L���$���r�M������\�o��l��Fo͎�6�uC[���	T&_oa��7 nk^[f	��d�E�f��A�֚�,�|�i/Z�r�r��Us�_�#K��
���T�W��l�#cV��K��b�8zM��K��8"^����j@�0���������t�g�G���j-���36���SƯ��%%���틌W�FvT�����﬛�-r}#���@H��W�Y��a,����P���4aH��ڕ��Q�@��g��N{���]&�왑�*W�4bY�NRpl����LB_V�����{�-D4+�w��"�չV'�4�xۈ�T4·P��MGqtR6��e�e�!��7��fX�mS�ؠo�R?�|�?I��},ݏ􄗩\g�*
�TM�/|�Tι/?#�ϥ�v��)cQ�?��/K+@<��t���ñ�g�ۯ�t�b/6h�ۈZ;b]�,���*�x�ul��g�1u��Y��q�Q[����!��Ā���I�?��&���Y�R�mR�$s��U1���@�CO�y����$_%1��		�@��k�[�tez{�³�tG�ɒ�,~��e�p���y&���vT����A�<ńQ�yȺ�Q�T�t/ ,YLs��'A����ܕ75�,t�VB��K��X��'*݄8 ���ww�l��E��m�Ɔ� =&��Ә��۱s�����zn
D�wt��jS���Y.�-�q�(}]*ws��!�̑H�&�)�'� ?9!��(���W�_��؏Һ�
���TS8��+mTOl���z�"L#����Uy\����������_)�48O�]��<�>���1���޶g���/mqF��Lֵ��ȅQȳۤ �7�N��S,C�'�=9?���O���Q"�Ǳ�V��3���n����i��7�8ݟ�fщ�s�H�V��t��®���[���1_��B^q!�����Ñ�Yk��j1�*{������N�4)N��*V��W��䵊`l/,AL{��$�1�i���ξ����C>Y��b��P?��x=��c0���S���y'I�c��D��|���� y)�����Q�� C����|�Gж`(]��A�N$��e�->[ɜ̯�,ö ;�����/�ӔX8�<"	�)UB��,Nа�����^@�ݨ���$(���j^ I�E�֕ފx!^�+�DEZ -`��e��#��dj;Gy��C]�N�j��Ye�frԏ��*�����ȟ;0j(��ށb76R�&��ǆ�����j��3,(b	��ӧYwE�Hr������l'�������xF맕�Y`������)#��|�hL%m�e��7X -2z�Z�C��WK.7s[]���A3VK�bL߱����
�r�yR�D���ѯ�=DJ���T<2��'�2� h�;S���d  �"u0R�ۇ�� z׫"0I�e]GZZ� 'v�	���ԑ�!*GrA�������}�=/������k�Տ��vlF�1�#������=Ʀ��� �aT���Z���2��"q��f�ӗˑ���I�U( �U �#m#ޞ�[ZE,��H�F�ܧ�O�zM�*����*�����
:3D��C*`h�"�A,[L�G��4�������(���JUq^6b߮dkd��ţv+E�-��x,	&��L��#͒��	�Q���m�����h�{>�I�����%�ۺH��-,_��^�FS�����_&^	�n�'jl���t�[*Ҍڈ��
�լ����M�!1�(�e������X�ƣ�Qݤ�&���t���$��~��+�>�,����<h�T������M$3hn����}m>l�Vt��R����YT���;�i�h�6�Q��L)�Y!��H0+�}}wx�����͜�0֋�����h��/��I���l�s��q��%*�.$#D�(y�&~n�����.xE;���ƽ���EPPLqU]B�8�+i��)M����dr!�`w�s��b��3F��lfp��i�!��T���V�����L����Ԇ��dU)a� C�w5�l�Cy�@@Y��_�Q�;���K�� ��Uv���\�jI�}����?R��m����	]ZcBªsG8��� V^��V:!�G0�Y;���v��X��i`���Be?Kġ�c��v���&��E������|A��'�-�+�N�z�.������qn$���x����D٣��a��]��|\	���  �\�oY�s�&0гfp����� �^�{�����i�����m�RO��ԡ�G�@]���s��B�K�ij�����}hȮg&[�����5�@d���n��6�|lɋ��L�"�̬ ���������|��:���6��7=
R��)��[��#��Y"�&�\-Kru0�B���J}˸[E��v�l1R�� g�)�#������i?�cҴ�b��xhjpv��;?6{
�@��~�sdu�ozW�n��� �����&S�!�W�Oʇ�`�
��_�fC�Ax��:{�sfiC��y,N��%?J�x���1/;�'L2&��ϩ֦�D�H}��ʛ�̿�n,��Jօ!JL�IK���0F�ͅ��6��Q��c?;�8��#mw�x��Q�܁��%=�Ul�̊����8,s/ѐƈ�q畚�L؁l��J3�Ü/�s������m ����,�����iݸ�t��tf��?B�>���h|5�8G�g�3�@�����ml^z�O���o�� E
ai�%��!.� �m՛3�@�� A9A��(��0�j]$w�f���F��~>�g" ��^"˿���U9H�c�-�l��ٙ/���]�V��}�q�y�O���Ѿ��.f��O�[���QunG�
���	�TV�ݯ�k����D��N���$'
��&!��vW"�4���u��/eS�|�Б�] �^EB�Pˡ� ���C˴�q:�2�`���"_L@(U�Y�݆l�غ�R{��U�jl����]�$����y����<�}��/$B@�ja�-;�����y�E�ȓH��>��>��kd��ӇDYQ���E�ПQ�-:.�M��~�7��Jqf�=Ͻ��M'"ڳ!��hg�&��i��mo.S%��^P2M��'��f��@���A�m�A�Y�k~�֦�\y�������h1���������]� �a��*�z`�g:���سi�M�v����;)��i��qV�� �:y�n����D�V`b��5�RB���X+C���S����n��<&^_�Db��z��Lnu��n���4�-Ō1���f��㉓��x�M���K,�{��rk ��Nx/P1��9��.��� ��%�O�%CE_�E'�*�r>�������_j�]#]�l�(!ύx02�0�p�ІU<�.C��=�&oԂq1�ͼ�}�j���u�UH/�������'��/��� �����n_C٥Xz-K{��F$���	���)�}����Ҽ�Ⱥ�zN۠В�w4���U�=o'Ӡ��A7D�����ؚK%��7p�'�r�19}J��	�Lٛ_έa	pf�=Emʵ��Ñ;~�#/8���e�(Z��U<�#��:������jS���TB�<���o�s.^�zh�H+���$�K� #���l�r�%ҍ�~sN}���ͻ�J�c��t�Z��r�5�x���~?�z��h���K(�e�.�s,&>�� ��w�Y<��0fC����_��#.}È�w�yu���f���z�Y�Z�~>
�o�(%w,��+�0�i������[-�^�8W�S[9�������)�B+[��D���6��YE.`&�u�&��]y�����z`ne�T���i��גq�=&��,�@�w{���g��D����iٟY2���Eu|Mp��_����i�!W�->9���3;�r����)��5C:���
s��h4���Y<�Ht�Z�Vz�2�I5�H�Q{��ɉI�Z�Q)���.QĄd�v�����o��c5�*��)��t�'>xHA|xU��q� j��
bֆ��)1��~9���"�7x�f��<���d���YV<W�}(�宸x����&�
��/F?��P�A:Y�v�.�0t�.���k����vԋ1s���g�����6ik�)-�ukj���K��րQQ���ONZH��ٱ��J�a��<�������O%t�},��0�0�e�be~P�#�̩y*�QŘZuC�^�sQd��ˆ�/Tp�P-��"��@����u�]����H���3��Z�T�N�J?�Y�h���n�If���`���&�l�L��X���|�+\1��l�����xh5x�"Ks�䠉ΙK��u���&Ld�����$��\b�W�M�D:Y���L�+�q�|�d�n����#����*f�(S]]�� ��t���1�O�nQ���x}��r0}k��R��m~A�9q�U�CU�
��F��S�b��v �S+J�~����w�s��o�S���i}+#��Ȧ�?okm�N�� Q{ѿk7�GE�?b-��,-?�W�?9� *`!] �6��8~� ��o�L��ϭ9���T���w
$М�2k� �͍h����CH�u"�����Q?a�e]�X0d��h��Ι9O��1ָ_�O�B�
q�Mǣ�F\��\gLΗb3�)8���?M���${ݠ~h���6I�Г�ۮ�B
l��t忝0U�x�kV����D��Z'mz`�V��	y��A�q�ﹳ��ǫ�8BΪ��tJY[ˠ��EF�¨��6�K��m״��{�9������f���N\UhMQ�o����V�ۚ��ф3*&K#'l�]qZ�*F򓊇j5Q�(~K���$h����:f|D�'[k��ͳPa:��䭴��
��vj�O+���� H�b@\��uC���i��*ĸ�5�����_1[?@Vf��mO�@{b�P�|��M+�$�Z���j�Çg�W�/�����z��M �c�5n�()! �b^*�_ד�h��9���.b�C-�~}�/2;�����v��@JY|[���Ƅ4a����*SLT��_�6:*����y9��9a�H����\Q�Ӊ|G�h�zJ{��T�{K��a�� �}�/��R����$�>ד��fE�k��}~�49�B�Rx����y�Q�3ِ�#�`G�H�j's��п;�.n:�f�p��E���h������gn�p�8�p:��j㇪5<�l���6-�K�ߴ�Nܲ�՗<b �3�/�P���#�A()	�bޱ{����u}�(��/f��PP�|M88KG�c��:�
���>��֡>'L���9��N��� $� B!b�^���Ck�T�[Sl$���ye�i|�$�����L�W�H��m}�tY��	�?QI�Q�'�ޣ�~��R���}�v��K_I�7v_U;��}��fϵ��E#���-���`�f"���EʱΓ��t@l���9뷙l�wU��82'A���i��7���ꉆ5s� 5Z��d?��z����7M����R���/Vp6@�U�t(�ȷ�hE��ӈ���َ[�7o��G���s�>��H�� ��֖��Ch�	�S9�S�T�>�yE�'h�2�9:f\_�,w���H$��X�C�eL4��Y���t$����x�Y#���>��(�Eĺ%y���m1��&�DЍX��[6p�=%��r�� �)u�Wa�X�^Q��̺���Ӱb��O��c���⽓�2r�9��nx(�QT�D�lphۖ��&��@E=�ǯ�<�4�R�Hӻ`SU,��+X�-7� Xk_Q��К��?X���i�v$^֗Ͳ~��"�;�����8�z��U�M��ȼhH�J_b��T��>�{��x��r�����[���_ջc����v�Pj��-��W�wU���"퉹���?�:�V0=�C+m�A�2�@7L�P� BǢ!Jca�^��������z��"�%��5mj��5��X�f��I����3.�x�cȬ�ל;���Q�B>(�Ɗ���.
D�G�a�H�����J�c�+�$����?����멬�� ���7f�х|<u�\a�ei�+��\O?7�����o��)��Q�����5=Uy��X�!(0?P!Y���]-��CL@M�h^���x���Wd��9�B�cfs/�P�u�9��t?1�̓W ���W�s+���j;�����5V�u���HM�y�g��69�`�n��ەT�Y��3���Eȍ���G��Z$4���d�O�o���ؒ�u3H�22rq���-T���BM�s`/j��>�(�M4w�"ݸ����G$�t^�A!=��bO��gRV\�����������֦<Ž�*���3�Ė��*ݘL�E�z(�aD�u�A�z��k���:Kݐ���o�o�0(JgM���ܵ]._�X45�݅�KG����Ԟ�G���iBr�8��4y�\����u�Nč����kӆ��4�a5�k1� �9$���ht�7F�|���-�.��Phg��u"�k=X�])�Y�ڊL����3�l]�$j�%O�`c�������^=rE4��-��.��8Yi�k�vS�W ���S��'_�p]�S){�C&�P7%>�fH�P�t���+�Hp1��ľr`��љC���ivT'.@�wR['�o���%]���S//�ҏ,�A#�۠�6���1(oz�,��Ik���Y9y��Y:b��l�-�nrR$<r�7��(c�Z�gq0�����ń���(9�+ݝ�ӱ���0���Z@�)*[�5"Ҽw*|f��v�F�щpB8��Y^$���K$�e��-U{�F�X�L���a?��y������������*QvXd��������%
4)[7�E����x)�Chqʪ@%�jc���� �˕ �cI�i�A4�N,�g�����Z�N�5�']BSf/�T�\�0IT��n_g��0��t�G�<6���h	1����('ȫϤ���"��lKa��zܳY�^帖�ȵ�i\Ǟ�:��&�ٌ^�I&Dٷ�qSCڄ�s�ש���o�*=�E��;��?�;y܃��\Ď6}��΍��5��i�W�����\zJ��f��� �x�y��L �_��@I�*��Z�`B����>�e[��z�v+�;��Z�S���Q,�o K��A��L�?��% ��L��r vPX/d�KÙT��q�wk ���	�k1���_J��um �N5�U���{Y>���v.��ʫ@$�ӊ0"ܯԧ">H�a�?��E3��[�pB 6<mVq����MWY��I����+;�kp$W[&<�Lo�ԛ���]��5}@���A�Ys�����3�N*��E�m���4zꛞ��o66j�26�K���g�v�{]�K{ո�Ͽ��V��'Zf�;�֢o��Rn�Xl������.��4	��HzVwd���mM��q��.�\�
*MEʔ��Š�%h��Is�EFE��w�A����ef���|��b����S����3ӞQF �#���]a��1P�/i��꧉�(�_���`B�����q��{�g��2(F�m���W�q����:tmS�t����LS�t��LM��8_Iz�F4���tk��BK6�S�M��ig/<���.Z��	�^/�e�G���3rϏJ��l�W��|&V�f�(����;@�)b�Js~�_*��vn2�bn.lT�oΏvY�o'��jM��?��Sx��X
*��7ʹT�ܛ��T�I%9C��M�5s�/���(��K��<ͩ���`�Y!�T8~(z�J�_�;���ҁrrI�kz��ŀ�
�MrR�	hl_���d���18Ԫ���
��<�MƋZ`���ԵC��5�U�s�5h$FY��e!�Vix��HF����J�<b|R��������p#lp����L;�OP\g��M*v�u���w�ĝ]�����k!�!�\�o0�B�6�L�����W��D��7�,���sU�x�LK�鱬���?-a����+"���W/��ڿi�M�H?x���c���~w*@�
�Kj���+����+R�<���-53փ��������������hIې����Cep�?ޮ�����F��q��ĳˢ���ne竌˭�R�X�wT�5&==��3K"�0�A�?Q�ҼWT)� hC~.�Fb�}VY��aO0CL��>���������xHxӗ$���+������G�o��I
� �asaiA��P?U�bZ���l�-+$Tq��q0��\�`xS%;{cf1�yS�M�����֌�w�Ɲ��<��4��U�7�P'��[(�*�A�md�1��c�]��W��T���NO�1�e �!+�ݺ��d�i���GYb�ߥ��cy��c��0��!��'#�`f���2�K��`��;�i�4}�V)@:GԈ��<n��/��LG3����s���ܐ0�3�Ӊ�ɸ6s��s$@�씡¿��&��+nĳ��ș�m�����S�0Qj��[^�<��)���^fLh�i$�e�E8u,i�j�ho'qF�Jr�^A���^����Ȋ�a��T�]#kOQ!�O8���a�NPEZ>�7��9B�|�}���}؋��<ܫ�}� ~�L����F��VU��,ȃ��'v�Q�7�J-�%u�J�F�>��8l݇5�=q-��ln�༦����8����Ϊs�(�m/D!�0ɍ�m�rˈ��&�A�Z��`R�����(�)1��4�ߖb��gWw%])fS�BʔĔ�x s�0�}��8����������&@X�R���8}%����Æ=�U�1ͱ�"B�  "�"�M����\h�f1��1#��p�x���>8+�>��Һ����-sW����[�Pʮ�u�3�-��Y|Lk��z
���V�m��Q�z��{�R��h�N��T�s+8���}/:���㙾<QGl��PT��8MA4iV�rbD�������4�5H�)��J����!J<,h�R����Y���D/���<[��q�Az���X�`��_�9`+Nk}m�|�T�z͎<�cڥ�\zbO
����rʮ0�O�]Vя��|8l�0�b�0�]]��ϓ�F_|�	.�&�W�*�uF�A��M��`S�S4��5~:�g�cY��U���,u���P�T'���6�3p�,7E�K��E�����:$��zs$���\���������(�� �X���hW:G2�?zB��T����8��]X8�"�I�H��Tb,�.5����UT�7;iÒ�:�k	����W����`��YF�q��!�>Ր�h������C\��x!/R[��P X�.����Qn
*K-�
��?�p�*Ģ�r��z�ѷ�x�Lrٌ�\
;�U���UqC�P����Z�k�}�=otT�Rx�Y�"���7��zO����P�qg\[�a-�$��f����Fouгj���B��R~É�\�#F�y�H��J��um���
��0=?��y�v�U�wd�GD?�هEs=d�x|-u��9�g��T �<EY�$X%e����a������6j�Me=ߙ[m�hI�a���0aY]��� ?��,?����E�;^�0�ֻ9Y���yoSi�>"�>�2�R��-X��v��m@ɲgo��n�Q���N���䊙�2��g�D4���s�U��K�����݅�	� 윁	� T�ð�7��bI�Q�a�[�c������k\�q<��a���h����n�l��ÑQlJ�I�vF:���j��P�#�1=D��ɮνK��lu&B|���"�&J��Aew�=����rFSU�l����{���o���в�*�Ǽ����kQk�-�5�u^���4��Rp�M��<��nX�%M:I�f�W����=!q�����Zf���$�J�DK�3�m�:�Z��.�R����}�Dp�+ŭwGZw�7e�Y����=�����|R��Qq��,�~#�If1_�L����;� �z�RXX T<a��R�M��A&}�heQ��@)0r��kl��cV���j�".	b�[���8��b����/s˽N�$?��O�Ѳ;ɐ"��5����ů����t�Y1b�P���Iƕ��K�\,�Q$]D8�§�%>�^���n��^�i5_�!�xP�-ϕU�Ҽ�e?E��ym(l������<��7.�ʆ���@���u�v@RS�?������o�-����ݎhw!w96	�4����S� "��Y�/F'(�{��HK��X�/� ���LL���p5:�N���.b{�6��'�iKp��.8��d���l;Lا�.%`�>�~�ӌ�½Գ� J�dh��,G�Xh�`�E�f��Ƈ^��t�i\�}}���#IZ�P ��7�����{{��(���1Q���8L�-��2�yq�ܑR����Y+#/�9����&-��и͟D��,:�L�"W���⣵�$wR��W�|�i��sG>P�8b��e�6�ʣɁTϑ�ܗ
f�E��Pњ����}����S�<�׷����c�p��Jr��A_5�n��j"R}D�6�����h+?�AZ�=:�uR�I����^'�툗:G�i��> � �CP���,��gU�r�?�ZoD�����r�/a'���
�+f��d�Ps� fò�I���.�걚�C;�1ڸ�oi��T��*��a�c�P5�sO�:6z%nv]>:�6붱1CݨSM1c���Q֌!�|�h�]���-K!�_͒����ڀ�	�"5�Y�C� ��¡��T�v��.�W_���ƛ�!�+�@K��zS�y�kz��ZV����0T�� #��굨@�r�~\�_���֬��_���ܗ4��z��ۑ���#��Vj����3P��\X��}���!S�N��R��m�q;)��_%k�H$BZ�un��J��֊�1�W�6���I��nD��V��e�o+;��m��}��\�<
��JJ�Z� �2��y=db4L�3���r{��x�p�XS��a�������X��i(E�tt	��1���W��3�Ϥ����za�=t�ɣkI"軚f3�瓰5�UZ��'/�Z�I�~<�kuݡc��
�I�E�s7W�('���:oD��h�@#��sJ�����,W�2�q���f��M!��4�U�qP5�D'%�gY��ċ?Z�V� w�j�
�]ܖ��<����HZz&_ND^�-�����c��*ebX�M� �xx�Th�C�8D2F����c*�����o0$	D�K��\d�ǂ�0Lv���i��Yk��ʌ�u������B,hL�F�RF��)꘥$���x�	��G���U���,��	��&h!D���N�_�E�G1���k�0G'V;�բ|\�xB�~���6>�.�����7�G�T�@�.�Co���n�ਥ|,W����^D�x�o��*�r�pΞ�/P�+M�B��0�ۢ@�D�kF��cp�<�i��X�M��@�|��
b��_���,ѻg���xN�/4.�59���� �Nhke"
G=(x�0���ػ��',^Ew}3u��-�wI�t����~��Z�/��H�3Xm�5�b�Jai��a�G��o�%Y��O�C�*���r�I�i�<!��N��f���Q�F�O팬�:��z����^N 	B
�a{0��+������٩��X���%��ܕ���"]�[31,ʁ(}� vR�I�s����w���ķqՀbZ���Ik��>����)4ĥDmG��;g�Z�������Yh��~��N9�^۹tLH�,���A���6�o�+<�KU���bQh�!��;��m���]�y]��(���d).��:�8C�{�	!�\��ܛn?x�c�����84#�F��@ጸF�|��્!��M�}���$��꺚���%�?���Ev�����n�'��_��q8�1���]5ғ�/]��j�C�B�ĒF�X����g�3`N����\��+�V���a!�J�p�~�7E�Q8�R�t[�b�Z.���i��?�L�t,�E�K�]��sA1�A�j/����ώ�#���Ay̚��#��2��􂏤���N._�]H���J��Q�t�#�_���{=����-��d+���`�i�y�΄����X��PA���,�.we�a��������+`�C�Wrz�F�sH+k�b�Ov�����o�4w��n���n£.f�����j?-����a$�ufe6߬�Oɡ�DR_��$����^�U�}��H���f="#��0|�r�3�_�1�D��B�������/hu0�b
�e����&e��64��9�$��;�����65�.R�f��)�GɆ��=�f16
鑼�2 Y4/��<C�y�
�����n�C�R�K6N\��;K�M��x����im�\u�0P���U}z��au�@�K�}���&j=�p7����mk�^��إ2�	*Q��,Ҫ�*$��b)�^+�ʑ�)m�m�k?���BBY�$�3�Emv��B|���}w��ĳ:��Wyb��@(,�����q��e�����^����|�	�&�}$^jy��ĥ�]�S^�S�nR�f� �k��I{�"�@��aHɁ���f����-g��7����G�\�O׽�@��
�)#$��%_�Չ�+UnG�����1��Q����u�m&�T��p�Eq���ükc�!| �*��Z�T΅��2��1��ǎt� �D��Yl>�1Fg0�v�ت�w��E�����h����'F@Iq��w��]�~p�������I�߈
:2�)C��}�����I���
)!����"��B����^�<�0�MV�C鏃ygY&]��7��x쁪ܧ�`s�R��
�tʕ���9�,J( ��.`K�F�h��L,��f�N-���������r��"�Źl>�$�H�m��Y�����`�>���v���������Q�����v0l)_�a�G��y�j,��lgg,S,28�>�{���L{�t��ȗ��^=�a���}�Ne��FkQOA�<��M3\Ml~��\��v�/K?�t��`��	]�m�`h��U�h�"O;���3���ޝi@š�I���G���5J~��&:�4IxK�"�`�ƱMի��:*�q+��8����7��=��Fc����}����s��!z�▇�fѫ�
aBt��ebl,�9��n�O�~(=c�9�8}��&��Pku��/�l�A,b���nCb��Z0���O�z�&
�fMKG8��T6A�à���#WF� C��� ��;����>}'��~5`j+�4t�����A�,�����U�AIg��(�R*��z!d�7Z<U�E�gǱ�C�[%��?WX�|w��G[���`�.���34O�NoI���A�7�E-d�� �W._�]|�J�q�E��c �5��'h�����+U���M�
R��O�<r� �8�Jy�5m�F�w���y��Q�N
8�2%jF����$R����d�U�}sL$ccy�I.A��_ʃ�R�K>T�V�[;D�z���j�7jŇ�$[��6׉��T�-�Gn��`,lW�:O��C9a��j�� ��c�������~X �T.\���K�'��1�7K�o�S[�vZ�yb#�O�^n�P�bu9� �&P��]
��S�	tyQ_<8��J���&%3|�ȱ���V��P��v��!�aE\��njm��:��. ��R��jԮ����~{��?�jjm5��kB���a}X,�H�Y�f"�U��cd#j9�[2Fn�!/�te���Ta2��C� ������O�[���c��ߏ7!I���C�/�g��j��>�y�,�1{J]�}U�/m�K̿#�b^U\g"����bgE�f�sN�����0�F�M�C=�gz�����9޾.���Q�H�?9HlN�g�N7'�/b���_��+Gʅ$J�R$���ت9��-Rl�\�p8���/#�緓%օҨ��������'��������]z��%o�DX��C޾�\X(������o�	lBq篫ҧ��v�h,M��V���k���_9�RPʟͽܷ�s#�r=�GV��\hƱt�A�G��O� ��c˵���Y<���F����ReB��S��Ĵ8�R_ ے�'�bu���"�PW�6a�!��)R��?���h���7>/qB��HB�r^_�J�*<�v��j���T��ə�`>�V����\y�,�̶#�C4�%�"Eg�YM�
c��N�E �E֨f���R��V�������,eT�'����U�B�Y �q*j����L����`��9��D >�Z��,ebʍi{d	��ʞn��39�1�e]��Ӳfl��3�tn.� �U��-J _�������{kܞ�,�2��ީ�2Eu'��	7y�B>Ҍh�L������V1�nD���;�K�� ��&���d�a/ Ϡ�?�����d���B�h�l�A�&���t>�� ��G�����63�qJq&�����a�ɕE�S�$]�J1���7r�)S	�F'MOF�/Hpg9�?��#�FÁwj�=d�\�?#����k��l&�JDI���xa��XK�U1�2��4��wro+�@�A��gM&��/�
<	^Q��c�Ϥ��;�1;!�tfu2�2�I@���;o�"��rk��֮A]�Tԋ��	[p���#�H�XE�eH���zAu�{	G��mpe4U�H�zTV�����(g�9�$��g.��wj?-����������> �X�.䲞O$"@ݒ�thݩe�������^g�q}�6��y�A���>�'F�:���Q�-�26Ϣ�w��9R�	����`+!u�����䇐m�ȼD�%��*l�_S��UL�D�Ŭ*ȧ�0��L��&��T�`Z���h~q,�������ɩ��nS�$���z�����!{Z�i�� S�TR��Y�0N��Ju����ChU�8BhP���70A�,Hb����n��-��3YE�G��3�����(��]�q��
��P�E��y酢~Gh��/H7+������������-u�9*!�ް�ܰ�Ϻg�c�|5;�M�N6�q�;h�LtW��4<��$U."��D�	߶�N�O��4���voH>�/f�H�H��W"�.���Seު�!�3WPGI��6=�%�( �����7m�Y��?^;'��a�
Kׁ�������y�}D��P�}>Ȃ�h��b|��P�X���?vv��\��,�N��A��/ cL���襬6Rj�`�!p���#,N�" �����C��o(N|�ѻ]n/�')������Y�/���l���2b)���g�����X���x��b�l�}���&�8Is� 1�=E{��64�H@�?�]F�~�K�������|�.MJ�R�r��.�8J)!�#�\�	����a]^O��Rn�����o_"QHx9-�<{^}���^F��i�񌍟9ztx�D�E��{$8Ut�^��K)?�j*�Y�Ip����S��S	�߬ FҪ��;��Z駬����y�_�Jo{�I���q���q�7e��>h���?��A�b���QI�+�϶����;:�+�}6T��E�N䷷K��g	���J!�ƖSG�� B�1ח`ň5v��!�볱�Ēq�H�D���,	���HT�������iY�*r�|W�Ni�Y�����:t��������� �I�u��,�}�V: ��3��#Y�|˽%е�-�bw�J�")R��E�d%o��S�?u�4n�B%��;���Y�7�Q5L7���h�|��6��P��@]��`��p�NՔ�7�5DS`R��Ε�"�5,�ڴ�9�@U̞fӊcos|Ol�,���ĳ�}���]F�[�w\?��,�DЃ�1>Bh�^<R�� ����(:b�|�3��bJՖ�7w�]�˭�1���I���v�\��8��2���d��kn1�:�IL^,�͇j��n�`�_`������]6�-D7�X�s<G}C��7�� t$��Xg��t�"���l��m7s �� �mJ?TO2K��I��R�s�a̾Q�h��W8�B�0g�2��_��ſ�q��B��5E�I?p��쏷��R���[=9�c~�6l`�ʈ"70�W� ��j�|���#)��r:n��k-�����=��)a?)�yr��Wk��5���a�Y/��y�4��#Pģ���q�o�;2�m�7��з�n����!E�������[
s�����%͑�'�D��･\���.���KwC�.Vc\H���̗������YہT�!�w_7J� �q>�v�F�T����7�-�*��o�I��7��p�hϽ�����Ny=���"5�����:�$�Po�P�:���~ұ�}l�aR'��۝���P�t���z�'sA	�����u4Ξc~��<�ww�������s�c5��G@�I#=/S��Q��*�SS�0�"Ӑ;��5������X�D������	ь�e�j�S�Ń:��I��%�m~p fEQ)�&��/��d"f#��Fr;�������~�,�'��k?�{�#1	v�|��"�u��q�K������ku�N2f��׶����E�Q��Y�����O��ɳ�4�����.�'QN*[j���,�r��T�=�{Q�d`�C�Q�3�'wjK���SY��ҕ�.�5i!��w��!��f1ä�x�V$a8�W��Ey��;!�XV�_��^9k��;�5��kЁ����?�{�\ܸ�����:8�c�Ы�sH\�r��Z'�6C�ݺ�i/���F[�I�o̓���+G�J�[��2�,����%��:�-�� S��،ÿ/8 8�ɿ��\g�O�;h/�{�tIP4�X�4�-�7�3]�hhyw�G0(�-������U�Ņ�4� P�C�}l��Fv.��jl�7gZ��}R�er�(Ƙ�q���V:�_�p�:����Û�d7Kn/���J���0�![�U���R�dS�2$(m[��@\�]��ebo�]�^�lX[Qq�)��� ���,��WD�?	�>�C���hUam�����`�[�L-a��`S��p���dl5\��.Hvt��E����Ԍʏ������@3A��@v G������I�/o;��V�P�ʯ��.
�K�R�R|�ȉ�6�o���L씩<jV�������lH���"G�7M�)�S2���ۚ���~�Yrд�V~�<!>\���/Z��1.�nF��m��k�N��k|!���>�x*�<mĖ�<�X�AxEbA��__c't�,� R^2���C|sFea��l�p.:��Z�{��:�p��[R��/�	�ݹ"��t��>_�_&r���ez��pv�F^��a�Ew,+Ζ���l<C�~<M$�2G-�46�b�.�x�Cf%�;�["+-��KY`��Z��k��4`-r��qlawF32*8Q����VWj�s��{UcF˔���|A}AC]ov�1��KEtAP U�.����0�`��]�B}瑲II���oz�������ʱ��GG��W�rQ�^��R�31�_l;O����$����Z\c��$�To��,�F����G���FjF����W���i���HK��r�7uOy��}��/�i�����=�E���2V�-�����5�K��$�~%���0k ��� Y^�����U�Yϱ'n���k�詍MA�t�J���:���M��\���M�������M�f��[��f��".���Ƭ��!w�C���^P����R������ݲF��I�������	����}��JU�nf^�u����q�� ��#kK���������5�b�7vr��֔@�#��J����]� �h�� ����ǭ�65C��aџ�&�N=����AG�r��r��K�7�.�p2<�z4<J��殇�K�lT��7�z�;-/j���^�}�K)��A�֫�Դ�ʻAC�D.�u@@\��[�~�r�))m��B3a�������=�-��z��m�o�2@��"��=��[�mN)�m�H��q��vY
�� �R��[���'V��eJ��p�B��m,ep� T�	�)+m�E��'��"��Ƈ5�RǛL��������R��6Y�ò��^���g�[}�^�crƅ���("f�����v"P��5�+ �	��No��ĮjW�@r�uY$��_{4�<�=�m���#�̽cֱ~X��E��N�{������i���}��
\۩]�zԪ+���_ԅ,�`	-i%4��Z�t��w���5F�e�(�>;��ʖ���p0-�:?���'a��������A�x�jA��ǃ'��z�^�/�{�������NI�4�������A��Y��%T��|Qn�'W�� �'/�^[�c]�(�t�I2��g�o�O���:y.��V�-k|o��D!�	3,����U�9���鱗�X��jE���B�b@�ȮAzZ�������8w�\~gtu�?R#��p�/�9�FdB��eQ9e�������_�|�1��~+D�x����q�ߊw��4Ο��Gj#s>��`�U~��hQu�oG��![0Co
S�Z�d�t�B�-d�"/��Xo�so�C���۰�B�>�E��W�$�%��i����G�Nъ���V*���9}X�m|�S�u��7m���O#�m�*�,٘�Y�3����t� �HK�w,}��b�q�{��F�*��B-�2��{�� >��E����bN���T��ќ����|;[4Y������$�1� �0��,�!3JU����]��0	����d�z�,h!,�:����)�E��y��
'Dn0��O����Hc���*˹����hce>�EzAsQa�~P��,�&�0T�[��B��O��-�*�ux�U[�3{��k[�v.�Ut��1�	Z�e!����Wn��M) �狧��ɓ��!0/
h	��/��A\�G@̩@�cg���T]FL>m=$���g u�O��e�(g��O�'��@̧��D�2f�8SLGE�$����y�߽�j��t9W�U���	H|GT@�͢r�^���9wI�p���qC��4k�0����=�=H#�~������󞼀��C��'��"ĥ�eWqb[E�G��/b�R�t�
x"G�.{Ac]�AI�����@��
ܽvn���� D�_h��S�I�f.<g�����Y�5�#�-�=���ik:6�
�aI�Vl&:p�l��+��6���dy��,���"��s���V�@�a1�:�����*���\����ֆ7�ҷ��c||/��O�Is9�~���+Gv��]�v�/�r�%�",�R~���������I����QӇt!����3��.R�>|Or�(�y��[P�a�k���BF�C���4�Z-t��qjR�Bm����L=��g�tSH�⧤LѦM@{��b�3�
�5E�;���T��Fq�`V����E����t�|��*&��疉WO�&��=mS�K��&�iP�֪ɠ��R �2�Rb�F�-���~��%�>���y�SakTpr�rV�u0(_�C	c��{�O�[��u�SB�4�(}����s�w��q�鎴g`p�U���o�&�"��WP��d� ��w^���k�E�߇�� �]�9y�ע]܀'+;�HA��?��-<����݁��f������ػ��P^�9�mu�l���J��%�׮K�v�	:�R>��g�`��Ur=/l���~�n�G:c�Σ>l��QitB��r�ո�'#��f�[�_|���_���v�І�%�"�W� ��W$D�4ƚ�c�}O�U��z6��)�
-+(�:'�Ǌc��A��vo��c�Ҿ�o���Ӌ�G	�l�.����[��7����6��Bq��P�Ųǝ4cz-��|!��0?N	Ze����jz]��{a�PhG�X�0��H�S�R����0��ƃ5/��'v&���Q��ֶEj[�'FKg%a�Y�t���CF=k���������!B�}ХnE��]�B�9���~7�ճ{�U>�R2�xy���c�<KY���lr~C�6;�����T_��ь-�/��&*05�Kj���Qp%���}�w��,Dͫ\���>���{>{�x=K��S�J���^l�ו�"��8��(�0 S���<�Z��U}�(�����i�Ju��@�XA�[��"�J�O���"���Xs#�ryu�$<ם8>�MR�� ����w7s#�)&I���-`�&ݠs!p�ɒ�z��Y�9���O�t��X����xh_�+�ȁ����_EY+0�"�^=4��}�[X#g`T�'aV{C��)��"�1H<Q݆6%�~���<���[ Pq���\�����b���u�kQ���剖��
R�~?!8��
��)gZ]�"#p7ip܃�������ӽ<;��b����5#O_�(F!7��w4�۵9!e��8@E��l���wm�c�#b�4��#?w�p�(��IHCc�
]��ABD1� �a��tI��5�\f�3���N��q.WRQ	�Sz��4h��2�8���L҆bw9���4��N��xd3�A7�z��{�".�=���v��gq���.`�1�mT�-��b:������Sѣ��� ��4�h���Ͷ%���L�"��v����c'P�OSH�Rp�@"��vr��Hf�A=�����w�IH�|���fPk�DW@�LZ:Z�<L�xaˠ�a�g��A���EJ^�Exsb?�����g�욎���y1���n�"��0fƃ<:��քH!s��ڬc��ǭ3`����JrN�P��3���Ñ�}�g	$_＼���4�G�v(��0��4ԯl8��>1yV�`8t��V}�.5=���N_�%b��^0ip'U(!G�g�Y�-��54�	���	���<���f����!/���������7���������׈���Е,͜��q�(	a �l�0X҅`��jKlIM	�Dri�D�$g�ݵ�VP�#g}\S#{ykN�A��������s9T�lX�MX��1�Z�{��\E�F�i�����܁�l�������i,D3;"\�/˨A��T��Ta��;LH�,�>VarS��]9�jn9;����	�~L
y�[�����.6e̺:���v�BߍMm�f��ߜ�}�rw�	�&��|�T�2Ii��zt��aҫ��!:�{ك���/�;ψ���4n���.";Z�=k�@�j<��m��a$�0���^H�aX����3��-���7�Νk|���J����v2/3]�8�(ծ4�?B�T�
1��n����U�mm3g���2]$���V�)��nww����x �[�h����Ϥ����ʞf.�2i�P6o}1�R5�[�"�H�e�%��Qү��k�@�Q�O0�����'���ʿ9��ɬ�#a��Z���ف��
"ir�`j_���#���:��jä�#f� �F���E�[l�Y��>���(7W�L��bm�{��չ�e���b�Lv�G��	*zDs�l�����Iv�A�nT{k :�2��c�����{�n]�;�(|CQZ��zD8�ě��v�F���&��t-��`B�l�oV�[�UDQ2c������᣽�(KRF1�,��G/�Yߩ��='Oz��`�c�!���K�����&�t��R���#�´,�V�`�o�hE,����e3ò���S�Ӂ��R�.ջ�o�;NU[�hj����@�=���Q�������C#­�1��v�/�}�U�q�҆Ô�Q��ɣ��E㹩�p>>cN���q�m�$�^$
K�*ja=ƀ�|�w/ؗ\�T�bϰN�(2D7~��$������g�B���#��|�J�=k����B���ۊF���hj�y=�9Y��ZN
M�M�Ը�;u���Q3E�Ep_>�Rp��٦�i�st����Qz� ��IJr)�uP���<��}��3�r��d
f����z�C���E_��qRl���E.���֨��U��`q�ĺ�H}�ձ/�����v�^^�A��Ϫ5�K�7��;�-=��3��TBD"�5'���c4on������7�z�N+�$���pݠm���g��K��_��4;�����ZY���=��I�۔E����B�:���t:�FS�Xn�oxc/�7�8k;�6yUgЇu�@�
Y�w|E3�O�DS����3#e��k� �5l���o���@Uzո(k����0�'�eݸ3��������Z0U�����#T8�i��4�1n[�d�{��B<��֎�]Y��/�idN�L��q"q-/8 EWÅC
h�ϻ]-��u���+0V��Q8̽63���I�b�I)xh�9��ܸ2���8+��㷤������y�Xʁ��ϳdĀn�a-�:�b������%�5�S�=�>h� ��4�����pvd���m���4��ڟ�e�P�J��Mb���J[^+�g.��'�n�����N/D�������Y3�C��Â`�/pv������#��1=ؗ:����ъƵ�����@v7��x8h2ҝs���U2���E�S�Sz��g�@YE�S�H ��Q�=07��r�8����6.y���`�7����g:�	����j��(�ڨ�Z�'n����/D�w���w��>@!Ԁ�lU�Pc_䅸��(=�jt���z-r"~�	�@�������Z�Eb5��?���ຑ��fF�70�g�ud1���oD��y�
�`��?�g.`6���]*!y�]�6@x���c¸�6魩�DDm�|��6�u�Zl㜽A����V`H�4��W5�T3�o�|g�ޜ�U��h)Os�O@���)��= 3��s9��I|���9x��~��(!���3�T��b?���p��ç
3� �\n
	4��sg
�%2s֐O��R��ņu�妄�M�N�nJ$�c-����?`5˓ �����o+�*��-q��69�҅)���ź%me)]�,T�C>5��C�Ϣg�RU?vw˩k���
.��IS�d��U��]��v�5�ek[�.Tx�w)�����oI�Ϣ����'�o�4�n�i�91������pH��r�}k�֨����,��`�[��m��S�B�'�Aԓ8>rM�Q��x�wQ���f�lp	3�x�O7I�\h�P�h��5c�:L�D�f��m�k7	�t�1GR/ӪoL�_q�&�V7R��B
M壙�H�ł{E[uPGF#D�����=\k�Ό�em=?v�9�C�'���&?�ʤ�Ӗ��1�O}#��Sa�)/F!�6���-roB�ǀ`�ec'����?M�§�I� ��Pj�8�WP!��j�Q�ӵ�����ٜ�7uW�Ph�F���;�X�v�o�1'Z����QLO��Ik��0-��8И\#��Y긞e�B�횼_J��PyhGH-��}���d��f���F@�7ܝ$�e�K��n��=3#�m����h�2�������&��]Qg�$@Jڙ		�
��a�]ͳ�eU�)��0�B'X��;�SuO?%�"k郓$��"�		�!��hh��_���V0��5����3� �m�.o�V��	R��S�����d�/�z�'�O��8���.JC&ĥ.L�����T7��=��Q=��B�؄~l�.$S®0��vaǽ�Ŭb���x>�2ź(��+Y[���W��fMb��v����U�E1?���1]�5W�� �UL��m��N���
<[(@�jN;<RO(�*GpTm�6����V"��fq��w%$��6*α֨zMKq]3:)�ȭG6L����H'�_A��<P[�$��6��|�����q�� ;he�1��G�÷!f��rs��X1 �8��@ ������4)r���)y���5-�>V�ݛ ���{)�d�A�|1ny`�Pln>����I������~QZ"�ED�6L5+�W�����]}�^d�S�u�J($�Sj%������Oˏt�{�9�ЁR;�Øj�w:�-9F��i�x������\_��cVZ����q�>�|.��9�&�u`��|��?��d�bz~��wT��ND,�N�1P|#�MN���!�K�������HO�=V�N�g.5��ψ�f!-y~0d&�ʾ*��*��!��F�j}{�<��:jQ 8+4���.a��#%g�f��b
k�	Q���s�Hi�[�;bT��m�t��kW�ƒ�2��`�eƎa�jPY��H���@H��M�
��ܿ��p����_�����뿈b��BK����ϵ$2�c�8��Q^��d�^��������X6�/����1>��"J/y�R���?�<��ʽ�������+Jh߹{���i\$���[�`=��{�0Zy":��� &
_��y��'xu*�������\���Hn�=���.��F뼣L���.�ڴo��E����x xˆ*�(�(_��DLy�h���^�n����ϗ$��L��F^0��@E���Xboh�2��}Eӳ]8Ŗ��7wW���/��#���#c�i�K#i�v�HF�{���ǩO6��=[rdt<B����˫;jf�j�j_9���KR3|�~���-iA�[:%�����%���s3Xd����yρȬg�
��ΰW|��#�,��n�X$˚�!�W���T���+�|�����me��%�T�ۣ���a�������#^��G�	e��6���h�ݜhܬ+�=���^4�"�����s>@�}ҿ��:�e]gNtV�k����dg��P/��]��)(���5߁peռ�X�U	�t��ǯO�5��̒�!p4�� z�t��4B��<��W�1�̅����pd���1ĵ�"��&aWvu͞��ċj) ��g�n�\�#�%��J�\i{
�ʀ�}Q�\1���3E} H�L�o>ڣ�n#�E���O_�
!xY �^eѝV�2C�j
��?�t� ��X:"�Ky���x��f��b��~<Y(�j*r���/z���8���{N_�ms"�2%�����#{���
�G�Ut��~�CAe�#���HH�y<�p 沈��?$B���m]A����x��䇹����M�H{��F�2X4����Q�g��w]k���E۹��u�3	����τ����qpl�9:�;��n�;�h#��r�|����`F7�@�?�$S�v*�4���PE��z~r��:���%'W�}�g�H8�^z�v�S�D�:��n?��U��7�	;��?D�� ^�ԭo��._q�_?H`�ߨ���1�ꊷ��=��-i�Hkˡ��#b�i�/SX�~Rq����U�m�J�H�B��ޠZ�;�R���nT�8Ԟ�2�89�7�_���{k[�D*}��c�ި.�E �ޣ�H�x���N��d�2Ç�Z�3 ��S�O�	w��|)��§XV��7��������Tu���U��myi��`��M�%�e���4��{U�����]�*�:��+l`��?�ux� }�
�gW;Q��D�ν�=�
8��}vD�l�ިK͛����0�R�5r-��Ƣ�N팠��(��J7�sm��'w��Q�����?���j���5������|,(��ķ'g.�� ������<r����m,��v��tp�m� s��D��޽mD�I�����3)�?��t��`Z3��bYD��W�'�Y���~�Fro�m���9���]`�B<�z�sZq��-P�G9ҿ^�3�(Q�����
Y�K����ذ��wC��nLl����g����	���'pI��#��%|��N*W��ԶQ�ؖӏ���D�^D�6z��5܍�z��نt#�֚rR��W_p֯]�N �R��/�H@'OM�X��t�.�o߂E�E�D��VicEb���U���?Cbi\?�9�yl�M�B����æa�l�A�G�Y'��_��7���).������'���S ���oj �{/�'�:�0��u伱^�������ƒ:הa�ښv�����{�䰗�i�#�Mt���
�����ƭ�G�i�i�n���5m	0�~��˦=���
�NT��7Z��]�[�o���տ�(�J|W�U���f�c�-�΄I�:y�u�o@��k��Hz~����Ěɑ�F�@ԡ{���e�������ʃ��$�'[��j%�C�۸xt�q���cz[�v���7`L!�p���\�|mėXe�9�q��K��ЪB���ڇ�c|�Pyo��uz?n%���yq�Y��b�Q�U�>�����h�d{J*_J�������Ai�(�-
s�E�����ࡐ�����y���E��l����uFؘG4NR�� ���~ t��VO���i[�S�}���⁅pt;6_��|�-ң��PK�V ��)��f���b�tҲ#]���w�]��� j*Cޣ_u�{&��je|��-����b�2��6���ԕ�����/T���$T��ge�zj�
4��%�aHn*θ_�"m��� )�ߤW����s�u��{:���A�M % ��p�>Gɶ�<'b.�Nx��_1�'��1f6�.���Q&/�v�=?�M�zy:�[=����'` �ƴ�c��C?�br������8�t��=�,�z�E'U'I�E���6;Qo�чm����B��4�`|���/�e+w�}4P��U��_�5㤜�N�x�����*#W��s(cN&�$"��5!����u��Ku�*�Ѵ'����B���r����Z_ڦ����zѽ�К���G5�!n)��d��4%�~���{�-K�gK6�v@UsN�����pV�f�����V�L��'�/�:��͊5{�ˑm�M��br�ߏ1 �_�[��M;��N�s`mk`Օ����¾-j���<�>���g��1j�3(��S�j%�k�O�'�C�0����V��_m�D��TQF�h.�y7A`�{쯥��"89e3���J������K���;n0q+�]�d��1$+�6�Oa:
?u�j�֝�%r2m�>H����Z��z)�-�Ұ���c%~�N���iҚ�L�ck����(�]mG��w'S���!���7�I8"Z��Ʊ ���O~�X�v1h%e��H����'���9!-RzQj崝^�h%��5, ��`�u�t���h�ft4'����W]˟'�T�!���$�����ZUή~��]b9�b1=l��9�b�K�.��f��4�r�)�c ��H��j21��|�NrE��I��%ߓ1|g$&=9@���G]9�P~�3%���U7_�a�8�o�`�sr-&� <��n˪?����kr|�9�
!�Դ���.��O܉m˾���=�:����L����~�;�
��r��O�|�'0jͺl�T[S��@ә�ߟuL�j�-#x��ܳ��c��"R�; #X+WZ5ɳڥZbǴ���rʺ�ފ������g��$�.�_�=m��΀�;�/��svW8�BqS
\XR��Eߏ���?���~����.�����D��}��$�K��� Z���bй����>�e�'�f�`����Xp=�
�'s���x��ܣ�#��H*�-����ɳ%Np�B�z�_{�qb�I����c�j1��æV��"��K�Ԛ�5p��iصQ�*g�m����g�����"	c�sǯ��L��Vt�{a���X��k��\.=��pt���G|�A���'���i�־O���:D�)p���𛼸�PTO��"�a{�j����8��A+��C���>�u4\`hr%��rj�>ށTY�V���L�	�	1o�O׃��̾��%,��1�{#����^դENPCv�Y�)�\�h�c��f��)���6�Q���!�}�]�yx���n����Χ8]٣F�W6����7A��S���x:��|�S,W�l�*/�Sz`��<�b�Dj~��`V��9��\�r�Ll��<ĵ�N���_���(�<�>��%M�~#��o@�zQ��F��B�Z{�|��lW�S�{ۗ橠U�n�
�Y�3G�$����v�C����)�V�i��)	�]�N;|����sVG�f�gE]0�b��k���Px��\��TF�'�<JO���8��A<~��鵂�}��ӥ���MG?�)�W�	���lk�,�n��r� +�"�Nx�0�~�����	��M,�g�Z`(kr�]���F<����Ɍ�L�ut0�����k]�hf]�S��"bZ�G�@:��Q�
jp�Ȏ��u�;�-�pw�:P�)�NMu���s�#�:�2�Ⱥ�ҀzT�V�t%�X��������?���""��$�P_M�NRڠ����W�Z�"��s��1�P?nm{=W�dr5����9�Bd�1��u�h�4: jK�4�|����'u�|�ڶ^n,x���'��zH�E[k���5�j�Ϥ������̚U��T��ߑL��_��O2V<s��J�N�=զhf�4h�k(��U|��W�z�e#�͛���0iP)���m�y�����̈�=��"ة6�.�N׬ZԍޓZ+�E]���m���>)@�B��m��#��Z�N5e �_o�)�z� rJ����6"�v�n1������9@��Ԓ����ֳ52Ѳ��E:����z��l��G�Nݷ�=o�n;i�H�& wV䋉oK����l�6g6qR|�=	l��hGF���~�0��+ϳ��3�(�r���Q��ۺ�
�6�6����ci��!Gj�� �1�w���H;��`����h��.! <L"�b��Vw+��'�҆֨R�7�Is�X��J�6 �LP��g�-{�6`�x�fvoSE�W1hl�[t�ƍ�US���/�$X#E�Z��\�k�o���ȴ.uqn��mI}��B��9fV�
_�����D%��<���S��3%	�X��Q l�r'��\�g�vR��D���^��^�� ��s� �������W�2,��X�WT�,(�Q�T��A'�1�G�!<1\��a��ey��~����VL��A�T���Byd�~tz�%��T>g�Mp��7���V��i\���V�����A�� �c�@i���'��Q����Tq����0���l�z�,�	{�]��;"x�����M?����k8im����'���RU��e����/Hj�Ed���ӏ��U9���MP�V��r�m̊f6�$���0�{/� ��eҗ�䏞*�є�
:���s^��g�{<Kw��
Gc�U:}�R
�m>!jA�����gx�Mwܤ���y������L�,)k6W�������h#w��Է�52�꼢2���̩�kE���H�svB��\m6+Ю-�pE�=�8��4F�@&J� ��I\�Ǒ��o��@Ggx��Ǵ�ᾶvD�`h�1i�AJda�-��Ў���6H��o�L{���!W���)_%T%���.����m��K����m����E��$����� *�����)O�� �`�#�{�BW����x���Ȼ6��f��Y�Nrc}9���|*�l����ɨ�GV�*TpB��3���-�F:�S?Dk�l��e����u:���{�4H[}m D�d�4�9La���A�"��iҥ>�Us?C����|�#�����0��TE8P3d���T/�|�O�)4a�S,3�3 ��[.�
-�/?�J�7X"���GN���Y]��u�&�x�LJN]D�'��P^��T����7�/���[��P�fv�dz�Ì	�Y=A�v�Xt.��1�'spe���&��^��}Wi��?�;"/d���L4�_=Z���}�L�t�-�e��M �!#^�>�?�Kw�9r.�K릚���Z��,hce��/�*�����X����11�:�y]�n3k0L��Řs4U�X�1BS�-�d�&����ư�v�#��g�
}���H�`��%���"X�N�]<#DHS����� 3?_}]m��b�๞,)L]2��@���=��6XP�x�뎋 ���wP����x�v�l̿��똊4�R�`�EhX�.�B��X 9�}�a!1���ɜa�;#�@_�]t��R�>��O�$�����!9DBf�3�[̿_�8,e����r?s��B�(��<@8����+X��������NM~L$��}�]���8����Ը���Wp��+R9i;���p*�!��C"�!��������*�I �7_��,m�����j�L���ӣ��t�)�wC�)���.u&ࡏ�$u�n�p�����_aՂ�ijoR��J f�zj�aq=���(*-	͢H��"�4/����:���Sӭ����%��g���`�|<KH��-�V���h��j;�k��ш2~٭�S�Kjw#��5�h�1�'�n9�,S�S��i�f,Ll5s��ŗJ�g]��UE�u\�OC�NYY���2�z�����n!�Ea�ո򂆛t�����޻�t�._�h�B`교,5�k4ſ�+��B&L�� KӬ*���e4������
��P�'�o��%-S��Rr+{����9�Ѵ&����7j� ��� �u��`asrb�8���;�ͻ����UĿ!��}��`C��øC ��N8�K<����cӠ��O"��AE�Ɲ�#e����v6^��|���8zt�fUJ8�M5�W�f�<�k�k#'��c��	^��l�YʻGM�{~13�N����nd�uEV�|9:
;�Z�b^f�1�;>���,�`��Þs<�]�P�՟k�ϡ]��!A�X:�� �PG4=%�ܞ9�9N����Ȍ"wE���|7"��|�122�# d��'��:ȷ�5��f�^�)��L�>8M[O,(�B�y��#.�$͒�+n��1da�����C���O�������>��@u�I����bw�Ϩ�ia4)Ôk���|FߔvV6-�i��Q�	 ��Vݳ���|�;���a�xTׇ+_p��m���;����c�G� 6�om��׬7�m�+V����(��b �0�_)FrR�db�С��BM�m��� ���;�o�������!��^�E2��Q�<x���7̯�T��'66ߚ)YtFyk���Q�T�]u�mD�ۆ^F�kk���g�\*֞�c5��KʙR��O�J��揎a��8:b������&������gػ��] �Kv�UN�_7��z���]e�;{)f��L%AxOg��3d�
�#V�B��}A����	,݃ QQi�]p	g�:����3l�A�4[A�a��Tr��k���/:��7��)���!Wqr�]Ui���W��u����D��*Bo��J���5��"�!���G�! PԀI��'e
��s�zD�z��`=����ȷ8����0U�Afۦ�7cįO�3��!FUA[���EA����@lL�X�F�9L�?g�H����nMg��Y"u�O��S��F4���TW����uQ�e>7��S��!�?�� ���sI�ߡ�́Y�o�6�	�l�E�������&@�J�_X��F�u肇�P�����HOؿ|#�K�~�T�*B4���}6R�����WO��� ^5#|I�V%#.ɔc5rϿ2��d��@&�ؽ-J�[~�}Њ>�zpY�:��b\���[;�`�����E� �
'`���BAٌ�D�+���,��g�'��`^���|mu:��9 ���$e?�-1�A��Q'N�Z��NΠ���40����3�8�7IF �\yc�ga����7	s ��}�iz�^�:���Ɣ�^���^~s.��ߜc�;��ď��{6�,����=�O �8�+��f�Ņ�'d���}.]9��=�}dފ5���p��Qz�G"ɘ��I1���g{]�����$M���ݼ��<�����i<l=iɧ�6���n펿����i��m��Ԗ��i��|�A��7Pc�s�☮�f�q-�1Y;�H8�7����K:#�Q\yS�:��S�M�9�>�[�qV9N'9���w������v�))Ke�K��+%�S�#Q�R�T�ܟ����t7r����`�,�A�GS��yGǂ/E��ĭ*H��ڂ�5&��웎���<c5����ka��M\�m�	|�����b��Bh�'-!ާKU�h�(*���"�j;����܂V��C��(%��Jo�^�8�e���q
*>=�8�}6~�>��ԃH�ֱ�E5��\�@��zc�47PC��C�`g�U�/��������ܔ����2~L�:��O�>�=�٥��X�h&ź:�S��h�j����l����wJf��~�
�i����B ĚY���� ���#ٖ��ͫ�R��d�I�1��Z�N"����j���S�4�1n��ٶ�����[E��#*7"���$��KN|��դ|35�ܹm$�>�X���G0m�yM%�u�`g܈��"�����ܟ
:9�a��DC���ضl�^H\����⺢^�ݣ����,�ϒ(������74�y;7���?!g<�5�#�K0{n�UOq! �?<It?ϋ8�0En��x��Z]��O��I���?C�'�J� <a�y�ڐ�nZ����\�W�����`%0�F^���mx��i����|��5#��<�n��Z:zZu��y�'O�I�֑ĉ;�#��C�vX:��C�л�W��O�^�EḚ����h�b��f�`d�,Kಏr�ao��oⵯ!`\#����p��(r�x�z|��.{܆ؽ����d2�m>������I7�v��1EX��y�׭��H\�#���]5S^�z�~*�^��5 i%� ��p���'g�w��������g�0���m�ZP��g(�ZOW�I6����
6��8�,�mU�j/���@���0ܵ���.V'&n�����>�"|h������2U��6�D-��I������B�:JpboBJ��_!�~����lK���'"nUs���=�n��Ń܊�#�ȗ� S���ٓ�O�)�I#����љ.���Z�֯,ă]������{�>�ds\�)
���T9�B(�~�n�c�f.Bb>_X�Z��{=,�I����	3X��ܥf��'�͌��2=���À���o�7ό�����N��QlzjCU��_h!/�09+�r
������ϭ�����3�,�p�s��\0��s�-ec�에�������~����q8��~J�;u��8�Q�w(�ioL���
���;QI�}�|=��;�W
���4��H�(�J>bTux��j��E�L�Dm}�ڪA��,�h9o�3!9X�!hϕ�-
_�Ʊ��?~��FO�$@�8{�6s~	�C���t`����7�W!����[J�}=�)���5xm������~#���Z)���lY):ݻ)��!K������9>����!��6�
�9Oj�����^����G �삨"Z��yA��Ů���8�N�GN*�t�
@�-	�x	��������ZN� t���+�>p�NR�+��*��%�(��:�h�i]������������[s��b��p���$	��¦�'}'?`Z�}�����6�Z.nXB
�d%��B��ZD���{��dH���3#�S��L^��ZlY~����!M����y��·(û����ǸjXr�l8-ƷI�b�� ���Z�V&)�dG�rE�����棤�F�*��P6����Ӹ��9��̗�@OA�U��I��#:M�&
T��&��eeQg�r��eK	�����@%��ca^f�ON��} �ϙ	�t#m��i�	1�.�<vR��y6*s�6~��� �������σ˼{���D.�_���Z$C]�J����͉i��[{�ڀw./[���Q�fV�qM���{|�t���3l�Ѡ��!@GN���vl}Tj�D�vL�������<"z*ҧ0blg/�t���R�k%Y�S���{�*
ʥD����U
�D�q��S5|p�T/{�r����*��j��YPo��\��Ph3�,D����'|����_*�{ae_T]�a@N�G�����(��i�	
ܨ1�j��)�x(��/Nҽ}D�?x���N���[�.��1�]=����b�k|	�3����[��{9̕!J�3���լ�2�5�N  ]�B�c֐����A��R��ōg�*��gW�8����S�EF�B�gn`�4��]h��O�t@��w�(ӗ���T�(����8v:�O8�)��ҳ��Ѣz��̝4J��$w�^�B|H
%G�K��$�P���z�f#;dJ� ,L�7�ǰ�,4JQ�=��K�Ԓ䞩��	�1E^�|�|p�+³���U�0iI���p� T�� ]I�edAqń��X�d�o���YN��\| ,�rZl}����D(`�_�L� Q�.�Hw������Gއ�2Q;����: ^�ݱ5׼�N
����j�/��l�Jk)�5�[�a*xo�]���Vdm�(�s*�,������6�w����'@���H�Z~�>U�5�#
�b؟Y�CnBQ\��������t.0���YFT�i�P��i�n)!��ߌ'�Jm�IBz����gO*F����Q���ק%�7�Y�HP����Q¾E}y[N �vp���N�Uj�Y46�Z����N�1p(u-uE_�`�4�E��;�=qɇv="�R�ߵ^��i���V�<��MW�]d��<����ߔ�8w���M��:�o����`g��3�pG}�:�>2E7iB̋;�(���OǊP���Q���k���+��$�*f��������%dP��V������	��e���>L6�J�$�DYtS�TG�g�>�
8#_csk�2T-���ϘR�K���d���?��szV���'X�)^ީ� ��i{��$�$�}=֍�sx��SC A�������D�UxQ��
�\T���y�;��%D]�7
y�}���K��8!��`��Od����P-nw�@H���p���^Sڪ0jZ!�R~P8�2��<�v�0o��+����Ӹ[���J��	��?s=i�������~�w뚜���:�HZm���I�tOd���t�u���iL
����,-�3�W�d�����1VfQ�f��(a>��sh�e��>��� ���![�����(��55��lv��S�|Z�(��Ǭ7%$��f6����t*�K%"ԁM#,�P!�6V�X�wvv}�gM��G��de�1���I�m���=3QP�T��o�@'g���"� ��g0U�k�uJ{Nɹ0щ[���\/����s�v�ʑWL��و�]�SOu�D��ݿ��¢M���zg� ��J7|���Ɔa�\��%�q���V���bH�QmJ�P}�~@�O�4k�0������6�r� I�#�7'|E��DÉ 9���Y]�r��1��J����s[�i�܅cwI�����~��ϋQ?yz��&<�������[�&�|q���^x"c�w\�֩�B�ƣ�l��c���y����������	��z@�U�;&�u�=$�b<F�Q4�V#��$���&����0�B�e�	�4Нv��Y�d�^F�d*�EN��ɼ�^�@?��E�;`c�d��$,�i�����/Y����o5�JI��2n<�Z�n�XՁ��.az��c.wf��PgRc^1T�=��W�r,���5�~��9��/.�y�>Ӣ�I�o�*��8�q����o�����1H{c [���{��vq��\'��R���_��<��Z���Օ���xܴj��m6�j�#�Ϧ��<�����`�e^ᯞ�e���4��=\�^hN���j���:7��;�����P܍��8�5_�s:���`�u��}�50q�
ʎ!���6��e�|��
pa��rA���;�:	������K�m�˺��l�7/�rrsit�%�C�&G�
p����W��C��� mv;�!.���xg������U�c���˝���N{�I�+ �p�d-a3���P�`��I\z1 ]x��:5��."6Z�دyf����$������4$��* �F���l�d\�c^k����vM ��$�h��ލ�t�<�N�n�Q��SBB����`���R�l:�(�n�`dIÏ/߁k��|/�K-��B�%��ou�v� !g� 9 ��m�s�.y�D�uP� p�� �'p\�!���*��s�%���F�Y+�����)� A����vjEB�d7zE����nu� �Q#��nɌ|y��`	WFD��X
d�ln}����Z©�%�M�S]p�n�j���V�LG�^�G�0�KP+�in�V4`�ݑ-ϒգZ�{~k��+�[��Z��s���o�`��c�G�H��ܣ�c,�z��a�=L�R�V�s���Oӷz,qDr�Oߞ�Te��A��+t{��`���y�����--�(E��f���H�f�bE���%����YU.%"�R}�0Z�i=�/�8z�WĴ�,�K����II�̯���@(t�jB�q|�kٮm�A,*�P�Z�'wɹ��V�r��F~�<Fg��Mⴷ4ct�V	�N�����X��*�K�	!�W��ٺ����a1�f�uî�k�T �:����6ԭ�;}'�� �8qӑ��&M2o�s��KH^���k܍�u� �[qܼS��ĳ=�ʿ��rn�%�z�s3�odT�&�p�g��1'���#, �R���3U���n;�cb��he�C���u8�&�>-|�d�U��6��،�g���ou���6��5�3Zx�%W*�Kl���4�m�h�_�Qgt�j�н[\�G�S<�1f:6Yo?�>%�o>���9i��LwֹB�Z�k���}�,R;�b��r��݀�M<��gē��X�%h �����,Bۄ���A��riBߣ�Rz�����g��1�V�c�u���m��-�Y�D��(l��o}7��3��5Vꩅ��_��[nu��B��CW�,"�S�,Xh�j��@ȿ�1Q���̠�쨷�\�n�lНs$ȴ�#���v��>�~B�0��e"<EKn��Hk�i�	�����~� 3N �1�B,I�"!�ݬF�;���#CQl�ל���l���\A���d���>il�0X'�=��'Ґ��=�`��b�c�*���dr����
%'z�E<J2��ib�b9��ᕝ�Vl'��$C���x)4^�چ���#�P����EB;�OWe�On�%�QE��kD���j�ੴϢ�g�j)Zj�GAE�8��:�����6���x��eҳ��x�g�9�E9���" �y�s���ҹ��~�U���.q��MZ�q�����y@�8|��ҫ��RXg��<�P@��د��?��#��$�~C���D:1(r(��îݾ��u�}��t�1�6�7�qڼVYH�7�Ft�����k��W=��B����{��x��0���������A)�� 'K��T�d�v"{�oԁ�-��$������sk�N�L� ��2wοR�WR�O�3��8����9`<�����;	�3ڲ�Np�����X�yw�Nx��M���9��#�t�H�{���iUL�<a�>�̃d�^~�]�	�]a��]��~�zA�V��f�>w9������ר�$L�h,���@��i2i�S��H�h*pA5��P�c�L�0�~f���l�+�
�q����*M2E�D�,H�~�
�)��-"��F��7'%~��|%�rE�,�|�ኑ.B]ⴽK6�NG�bZ��ս��,�	 �o����)4-��zH*��%s9��^D�d�T����z\ �����߾�cw����VoǞ�tuR?���V�Yk:䊻�Rky��ҧ7LB���e��PN^��5T�tQ�)��k%���|�
�׺+/\��i0I` C&��G���x2���`i���t��Ԁ '�n6��U���4�
�p�Mے��<�Y"�"wҁ���_%��ko��;H8x�ms����ր�+�@R�W 8T n�����Ȟ��������H�/|��8<M�_���e�G���w��G���SR>�|uGk���5-���N�-�o;.��c9��Зo�Ar��+z�|��X��Z�-��è���]kߪl`ҵ��oeN<��Mo΁��BP3V�����BW�G��~�-V������r9���J-_av�(*xR6����6���RT/X�f��؉�H���C1��XKS�/
.��Xm�RD� Zܕ)��7�-�S�>5��PK���(�/���*K�mv�\��?���w�pܸ�-㥄��z�#<�5q���Z~D��~h��y��Xo'i�2�m� �r�W�@_b�������zGe��G��s�컢�au�E�w^F�f%rn�+Р��l"�/h�cտ�Y�E��K�,�a�x 36
L0C��d��9���y��?�� ,���2��o~\R`�b]�R�bl��b{�#�t��
�T��?a����p&��)Pƌ��k��ε�%��z�-9;z�J2��?��
i[�yE�����g�z��q���>���Y��ժ����X��s,���@���򾺍�P�У_^��Ќ���N
jR��8�p��3���&s8�:�VRxK �"��i������n�绨�ŭQ՚&G���tf*t+"=@�tm8YG����:���M�z�\�l���CV"t
N�1W���Y��v(p)@m��*§ف.@��f
۱]�(�3��I/�R��Y�}�h8Eg
}�=���1	'
R�L0��x��N;}Uu���_{�7�/�N�8��^�]�{�m@��h)mg�}]��>��d[��\��N*B`hD9�`G���z�Z �*Mב���u�ʫ�ҩ͟_A	�<���[E�w]Ŏ�5�|b��p[�Pl�iS�\���|g�)��3m�>�����S�<KU�4��p��Ӆ��������^ww��>n��������@�͵I�;ܼ��N�ܡ���Pna')���y�6Kަ�!8o��$s3��^�Fq��<!��M@�٬�?"�?��<��BG5��3�nY��f�Hɺ�F�QƑY�;��ß�̱*��Ӹ�7D7|�"	��L߄ Ψz#U3��I?����&I��956J������`~*ӟo�Z#���8m���i4�ؽ�\k�Xdt|;@;�>z֕�$�ܺ�B�Ԓ�߱���Y%�nS�h�������6,B]LGF�7�{�o��/?�}N�$*�,�[��=��5�Jߙ����n��SO���`�G�N�;��=.��/��p����j�' ?�Z���)��н:��f��������t�G�TE2e�M�v������.�j���0�t-��[���� ��xޘA~����Կt`�}� CNom�w�c���D|��S��ނ�p�����Jf�����Q�E��_h�n��_+3'�g�D6��g63ĥ�yV�adl�KCo�}~��]�L<� �����Z�)d2��j�6�]8��jW�A%G���yC �u��b2���j.�����)����\|y�1'6�����1��#���� �պ����� �֋��,K�hWUz����i:j�Bڀ��@���&,���;3L-/v�����P<��<���7b �b�������� �z��qA���0f��Ƨ9�@*Y�I����a�|�shr�#�G���|~�g��]�7��Үt���1�$M�:QY=������猭�p�q�
�<��r|g�3�~']<�'=�G�ML+=]M\	w��͡Tp-YL욤A��Wע�Is|�j!�h�9)��}|ֆ�.�~~,W�k�*���穚�D|�kg����H�G �.�{B(�W%\�4UT��b�9Z��[H��bN�>���c|���j��lk�8R&Hω��׏O�I2��Y�f6r�T��GqS$���X�'"~�<C;y2߯��L�@w�HtR�6��f�hx�ߔ�'�5jt��bkz�ى�uO�� a%�	<!�(��f�r�"+H�\"��fU҇��]�щ����&�I��G���a�Ky�\ƚ@*��_5\_�:Z� ��.�u�eY��NYC���˙����Zr�ʶ�����ī� �eo4�W��>��wp<w$uI�`u��/9=V(��zow�p�_y�Rh��5DHxփ�x�3��i��n�z7�aD�ʶb}h�I�AsXޟaC�;�i�X�@`����+
_��> $R�pr#���6�-�_z@�|OA�ܰ��j���8[߹8�/ӹ��D�����ܳl� ���(���ў�<� ��!�G����ϓH�q'�o�]��8 ���8$�N"D/�2*����ܩjO�+k��������%�1�2d֞t�we�yp��2;b��y�?�<�m?�$쳚ǪI�H�� ��bMx�dw¬)� ���_۝O�
˘��ލ�Z�B�EU��㔓�p$�Y[]��a%�y�]�6"ۏ��Ԅ���i���Sv`�W|���˄��ٿ���B�m_�[qN��Sj)�.���%C`�nV�3��[,J�P9(��}]R'���[������_�����Oֵ�� ��ߌ��ZQ���ݳ��a@�]�w�����7/$����8����N$� (s��uG� ����4�*����~����O�."Ф����/�N��h��8-r[~U8�Y�V6��s;пY� 8P�����<s
Uq�?ړ�m��k5Z��[H���H��WY�Մ	��~<(7�o��݋�k���6�qK]�����4Py�G~皧�N
4����雴���oH8b�K�]�R�Ӯ�1u)�'�`��*\z�Y+��2��n����S~�EZ�a�d�c�U�E!B�p)H���JtB���=��G0�x>��p�N$��^�d��-���f;�&�P��&�R�9��ݤ��
X#���,���H�NÔ��cd� �a�:)��=���i~�[:����굫2�Ϲ2	���S;|�au��/�<�:mn���(�'�I���2�Jv�J�b����:?��y%�a�x�&_�ވ�,Vp���i����w����N�)��_v���X+OQ˙��\��c���a:$�Q���%w�~�s���m�O\�)5����L	<'7�� {��ټrI�TX_GD�D��'p"��k� ������������d�2�T�5>�b��:����l��nlW�Y2Lg�<�0�7�9LbQ�yj��tx�D]�ukd)j\�����b��Ҝڥ�f0�j�~-8�#5rB�)�D����m� �4ד�޺�L�@X#��Ǝ��Z�7��`_k��G� �����O1��	!+ʠ������-������$��_-�J[/t+��\��r+#�����/T�?HGga�e���r�����?�jS ]���O��e��Bn�Iî^8�D0����_H_P��0w�7����� �)`�ɍ��t�y�����0�����tIn� ��ApG�!�	�@,��yO�!x*����p��	قRR8�f0������ɻ��k�ie�
h�g����]�>�����lH��i"V��-��|�s��z�1j��3K�cʯ��9w�C������V�)��&��[�I7rj]ŉ�g\z���\��}�3k�=�r�i)[�
M��20�ܬ�G��	�c1wr�8�ѿ�+�k!�+�3� b�J �g�I�wJo_���A��r�tꠚ����{��i��C��iL��g
�ƒ�rc��4�P�p�	���^����:+W��&�7ʳͮ3:�壟����f8�V�Q�c�j���;c��
8^?�ч<1����0 �e���i ��,��X�!=�JHV���^')~���%p���C�������u��J$I�ģ�d#�e�Q�S�r<ڕ]�U�T/qj�F�nq���_%���'��b�n:��HR�B\;$ F��� E]�A��.D�|��G2���8��c�]P�Qq�T��e��'�)9(����2��S]ƞlE'U����uOԦׁ���X*�"TW�̞���h9C��0_��VE ��tP���x�{���F��w�P���$<o����
m�.���C�|Q 	Qz˦a�ɗ��)q����f�q@-h%��ǞN�o��L�!-HY���Z�ݭmƲ~��Dk���Rv˥�z��p��-�#yja(��CC5�u���������W�G���%�3���Y��;g(�b��,�)���W���5;&a�աY��4��t-�?�!
i���d�r�l��g���\Lw��U��'����F䍯@�Th�1����q����i�b��ͥ�`���+����ѫы߭V�0�7V�z����en|��M��G�ק_�3ڶK�񅎩��|�y6��N%�&��߷��;�h�= a\��l'�����z�=9�3[�ӓS�e;tĦ��Нm�c��qxI����RE�~G18]��썿E�ֶ>��R�'H������l���ˡ�⋛��0�З�R
�U	M��<Or�6��^:��-����.^���qq��J�����O�K���=�-jT����d��Y��㢜&NOs�K�S� ����Z&�A󎳙Ը�^��U*qڴ�
��0yc�?�&s�**��3�}��g����=��"�V"��ZN��Τ��M�Ѩ}om��(��\&����+$�����?�
 �/��5"�i��R�]���(MrBi���\r3�o�&O�ѧ��j ���HY<�5??�]H&l]v����K����DPփ}�*۬?i�@C�"x��B��χ�e��+a����V��{I����ȵ���?�0�V��6lf�Lh)W��ή,�7�d��t��u�K��l�v\/�i�7m�d�z���ʞG��p�a8q����䋐NYߨc_���L��&�Mr��o�4�jP��5#���8nMUiY�̸2��!I�����f9=���n]m�y,H�B|��QI�*��l������9�Oێ���B����w)�tǍ� �^�eA(�,zVu!P��즘�?�9�&�4�&Zi7tWT$�`̡â�cW%�dkN�"��.%�� 5�po�4	� 9+���Ag
^�&�}gh�p�5��?ݑ[[��4ӏ	L�=�Ȓ��j��w�Y�pX-�2O����p��!�Cs4�>9�\�͠2���Еl�_���=ܐZ��0�P���LDĐPhf�)`(���~�Y�P&m@X���=�衂�0�/���a��Y��L�NZDW4l�hu�������Ծ��(X��$[5F�+�Β╍r�a���2	O&���=/�c�s����YE������A��vy�¡X�b�@
V� � � U'>G��1�`���_	/��l�yu&K�Я�nQ�/lg���U���0�\i.@��	挅U�%()� "��t{M�1Bᩙ|(ίnq3Т�qy���}]��C� 2<��+�c�P�ky��kr	�|�-eQ5��b����>H�9�[YM�j~ќ`*~�ȒN0)������xe�9
�{�G�fLD�	~�/n5{}��Y����w���'��Xe�&��a@Xw�?W�a;�=<]ew`Vw`�Al�s
��k�2�u�:|��	�}�_�4q�>p�2R����S�E5��&(kw/�J	�F� D�Z,��^c��կ^%������b����A�L �:)u?���̸�~���z�>Wa$p�M>`<��z�֖2��F���l��5�=��p f઩�ʜ�CN:ީ[���2�f�c"@M`z����K�*���J�k{�e#N�o��L�'(�	p�DG3�h*"xEc�zI��z�jf�f��VG�l���g�b���*8�r8�<�X�S�:�u�N����MsM}n(�憶��K
s�f�<k���5�:�6g6�$�r�Z����/��-5!Y/�u�sK�l��+�,�Ԏ�qԺ��D^?��W���j�H|f^^��+g;�p�@G�w�4�1�@�8z�~����\��a-����ARV��?��bG;˩�▵�܎��HK��:�_郜4UЌ����9έ�D]1�e��oZF�rL���ԧ_
Ϟ�n�Z��P��_/���T�b�^g��"BT�9�1��!���(,s���!K�/u%�XX����1�R#�-�#��mţ�̻""�_���4��i�|�_���+�F�d�bd�#��z_r��~o���c�~�R�:�Z+���B���f!�7w�lP}m�d�ڕ^F4Ar�,9��1~�ma�oi1�N�wo�ć=6��˰�aZ�u֩��1��8�$���g�=6`I���«o�>�B�P�R�S�7��p�ş�������������sx���1�E֋��K�:���l�q\�I��c�"B��|�����qFh�)�7U�O��(J�2J�	�kb�O��q��]_��%����%S4`p�q3���?�3�\����U�'�<c��p��vԼ8�=�p�@6xK������BC�MjJ�����6���{�J*����/�������}�ر�8c����ʉ4p7�[����;j�&2r�1*���q]䔤��z�$>O�BD�L!,)s�]��pNڷ��}�A���|�L���=�`=�-_��k�lh���-# ���<�l�.�zʓG��j�)�_���R�f:�=y��U|hˉ�!O�5:"v|�����CK�V�q�m���d�)�sqL����ɩ�
�߸�^�0�ɴ�l[9���f�ULO��L�W鰚�:-��s,iC�>��?�8w\>�_�L=��?�N�����q�R�����\�̢�.��ja��_�S��X��3̩Z����\W�4 zv����|���q��m}��m�o�i�Q͠�`���Ě��^�����A
!�A�����%R�VkDp�V@��)�{d#�my�)��o:�������t�b��:��	�"r<2L�ٹ9vR��e\�w�9�q��B�7���Z˔j|�@�&>��C������}F�k���E�,�p�Rm�y��_:�q{V/+��徢�N6Ux��:�(�+�J���\�,`Ҧ�	���)m��/�l�&�_��tYǻO§��/��bh�;����S0ʿŵ�G�>٢e�����T��Y=]�	C~N�ԇ<SE	�-�>UiYL�iQ�S��A��A$�-f�eqޚ�V
ggor
�k��:����M�0!YIш��$`l�E����>�H���}�͌ˍ�I��j�/�u��i�h�rr"�P-E�}�6�}4)��C�E�6B�ٍS`{�; ��?�2�&��Ə#�D"�N/{I:��������D@��`�K)"w2[&�j^��<g.W��Pm�Y��pT+<�B��&_dU�~v|��mC����۳��ri��L�4�����}�q��@j�����LP�w��'�{)W�SE��jxUs�T򑠪溃x�ͦ�l�9����EI�oa�A��*�j���R3W�P�I��se�Bt(	��d�p-�H��z��9�;�N��ՒF�^�J��M@fAg���I�o��Ty1 ȭM�x�*m'KS��Վ�:���@.Qhh='�QI�Mv׭�k�6x�� ��-�>��"-ݾмՅ��	B>>B�,ů+F%����fU�@����%H��B"�$� �sӣ�FW�fޗ�M����P�t��3^\���n���B	���U�7^� �u�R���XQn�b�v�͊S1���o[[:T:����%�]����R�Q��X,�$�1�H�6&(��?5'��N�s��Gɀl�U���c�����>&C�	���ǰ]��p��ᾌ�7�kK���J�x��<����9D�B�3*fy�ҀQe©�=�D
X�dp!(����$�懬j,� -�1��%�T����i��~1��YJa@�2&E _�^��}��8�7fI7O>җ3.*R��L�6��#h�:+�D�[�5\��z�3���6e �H)vS�y�P���X���&Z���|SN#3�tezC��<k�"?(�Bױ
��J�l��!&9�!k8೬sL{ˡ�^���7�]_�	��0�]Uf��w��\j1}��R���-���D ���k���#i#4�V���y�W���0��M� K~��<�Fp���
T�i�W���uM��6����H��A-M|���O��^�U%����> ���Gn�Gl���`������+�}^�z��0�PKo� Z�)�K��Xt�RC9� 뒕��dj�Lz�T�8�+�/���tQ�}܌�bY.~�'<��˿.���c��(���BQ�	e��KqBm�:	��nԁk�����Z���;�t¨�-z9����X�&
��)8Q)p�.�NG���$��5 �	$خvǼf�`��7	~���3õ�B^K&
�w(A��/V����iP�ϵL��u���Ҫ����FA�����
6g	��㳮f����E�^gBB'��4`�P?�����3dy��-��R�Be
��d>G2�uH�����u����)ҼS(��MFze	���6]MSv�*Ȉ,G����,����Bu�H����f-�_W|Z�G0F"ӎiF	�ڦ��z�8�t'�sN-҉�mY[�u�s_��_|����-��g`��'!*���@��n��c�>0]3U�h�B��2�J��ƗƁj � KV���/��WYI�R�)E�G@�Tt���r��Cĳ��
0�� "0��hV(���9�����r�m�H$���݅�3��v��������t� F�1�A��]�|�ӭ���j6� �J8��84�4�.E����Z�O#��|������=&��k~ m�r��h�!YKrT@g����'2��rfcѫ��N����)PȎ��U�S�yQk�7.��ķ9a�}��L��1��i>��i����� �DB�/*����q!�G��h�3�|�Fb�Ž��T��{�7�����O��)�����K�D�����E�F,�ni�J�4�}�POG��!���F̾��Lb�be�q�����MV��XA��؏�؅5�n��z��V�qN��A�ZX�3y���^5�I��a��î��p����ψ����2.k�ݵ�OYp��h�,l��(�)�zjsBBCd�B���@j���m�ޮ�Hb��>
�"E�l�0���]��U�}=�eD�����޵e"4 ��>�& Tw����;�;�(7�>�DjU�����G��;��W��y�]!�th�
�
u�:�2��|C�/�=��	���J]l�����+x�����2��g�ܣY����;v(\��M��8��C^fՀ
��K}�1��Yg���u��ޥ��5 ��?]��/�nkG?xJ���K&���fHT�xx ��4�g�{��3@���p(RZJ���=} e{���3L�+��p��R���l-M�%j�y�2g�xr�ws������8�Tesw�0�6���NN�.[��򅺱�-����uj�̒�����p���kY�3��)V�T�l�����jEO��������K���=E� i_:���n��6�;}[����MPG�ЂH�b7�f�5��fy�����bj׆�"�ŏT �.�p��Xx��jM��<��(�yԣ��`gÕm��Q�I����j+��z����S���A*H[)@�;�~��Ie������]+�bT�g�%�1_�v��.�����f�e��B��$����;���W�S?����T�yk�Rfj`�TY�w��+�}߃ʒ`M���a��b�3�1���cig�"T�r�
F)�Q� �53j·�.]D5��TDV����5�0�y�dھRe��`-�x�$�,�ߺ��ǔ`TB�Ϯ|�3�K7o�lc�?B3̈́��2�0k�����to|r�H2�OF֓k�cf�A�����.�d���}3D	�N�J�#~�޳�5�tA�ϼS1�*�8qr�lk��gM;^����+�0�]�L�nT��[8A��Y�^�O\���$��Km����^����������N�L�4�y�.�P�ټ���E9��ϟ�,a��U�h�p��^.����5������S�'9q��4ʯ�ɉ�NRĂ��k
��U�E���FЁ Չ��k�u�'������r�F*��; !�l^��Ӈp湎�߳y�AG�^ͷ�8.�O`UF`?�k�['`S13��,�nǽ����$�-n�bǘ��=!�#�/����el�v������zQ�AE�U�٧J���QxC�aA�b�A����y�x��ЖN(��� F4��_(�:�R?��IH�E��w7yP���I�f_N��[��\+�)�d����_:T~�/y
��t�϶8����j�1%��:1�Vg7Vi�#���E��j-)s\�0<�����o����g��޸�F��� �a�Fø6��\f`�\|V��n���_��,�Cn�Gd���$Gͷ,l"5����뜯�lQ�zǤ&ہ�l���0�\ۊ:/ͭ���l^���c���'��jg~靖�@g5�;�����M�ba&�_�f��Z��;��9FQ	�0�d�c�@�t�k�H�1��<�*��O~H^���
��h���C�=�K(���ύd�&��"]�Wn\2Y�c�kZ�]��C͇��G̉��������������a􉛛�%����T�9Am�Z����l�_~�����C���49�p�e��=��)f�H*��*=��	��
*m��2gZ��"ʉ�A����)��;6�%���J�aXq#xx�����czml$+�`��Uߏ����_�	��u;�������Y���&�v�V����(�}��wj3 ����d&H��%>��UU5�)+]P�A�ʴ� �e�g�C�	�?�`�DR�� �R�b0���P�\ܮҙت;���B�0n���Yݢ���\��g#c&��T�3Y�y� b>����`0PY�E�E��w��z<,.=߄H��/�`���{V7��y�8+*�f�$Gt�4��k{��B~J�h~
);��%���ܭ�a��{[�B�ĂXma��@�H��#��-�e]�\��ɚ�h���nP��,=6��n"�zm�1A�/v?﬇$w�6�r;���3���|�hե�A�Z�ߵ>g���ja�`n�zj%b2�� ����Ӏ�K�
�Η�鈰�)�O�٣�:ʎ�W�(�N��^<���k��`h��e5�0��u!��2���I��S��K_�Z�E�ޕ����K����k�Q↶���'E؊��u�;a-��þ
�ߩ�yW���o���YU�@O��0�~ǿWq����T3�e|ж�<��L^j��8F6<n�= L]yP 楤6���A7<�]�Fʏ�DB9y�hDe�5H����P� %�9�D�֐�[�狎��t�:�K+2�NO2-z�Ð*^���S�w;�]=���.^�j\�蟓����r�G�)��0�6K�
G`��P�>ϿPl���X����f���� h`\AJ�z�nG0�
�_y�u�t̀CXE����P�ތe��E�L�u�dw�����a�\�3xE����+��քd4��e%e z=�n�h�G�b��H�I�[" J�ʘc_�!|zq�>ܾ��*�_�:�f��
"�̽=�*�າ8֜+�6� ���X��x��w����ӑk�Ɇ����_tU�_Õ����ժ{��'�Y�P}�
0_ywC�_ۼ���[� �N�u��������\)�V��M��q�r�vf�#^�2������Rц��Z��� _x���-$nxX�:0���-�2��Nok��t�-8�[%�z����bt�蘆^����ɚ�7O�.�H(\���R���	�}�L�Y�+]{�x>f�H�!KIe醂��|�)�PJ���q�}�D�ր���芞�M<���.?]Z�R6�Fq�_󃺝��B0'�Q�UP��Lx�)hQ�n�U�UJ�s,L��+�핤�N�x���F��+��!�8��9�10�+X�����?PjT|�.je0U�Dxe`͙�3��o�9���}�̾g78������<I���c�%&�ae��f�h��v	s�P���f�A����/i��݌`����_бt���cW5�	$ˣF|Rb��0͕g#f;����]¯���p�ݏ�=���O�t�0��]��o�2\�]-k��H�&���ED�@���9qؘ=�<)�F˸bⱢ�����I�����/T��s�73��>=rs����>S�C��F�M���)_8����z�w��l���HW�r���r@I�H3R��CN`D�Q�U�WY�Z<E9�&;�����|r#����+��D(�4�9�Uw &ccDB$*1�ֽ�(��"��(��'���I����T���ɫ� �m��9x�h|���T�|B�����XW!=YL���P�����_�"��'�!�M�����:�j�2�N)�
�=�%�]�M a��@�Z(�y�K�ݎb��T��5[��9I^3�d����������N6��3\m%5�9�E0DX��e&����1^��o��泛�K���<�ǌ���Ŏ??_K�#��Y�r)��ߣ�\�jN���ǡ��M)�w"�}#�m`�sx`Snz������_<.p�\�C�7�F��2[y����0��h���k��개7�9(��j�Z ����y���6~��Ǡ�)${��"������d�U�9���m|���To/9z����/yi'l�Nl����*|�<Z *+}С���m��J�7��9fp�8=�4��|Cp�E~�[6���p��!t^���0��h�rz���J~�EK�[r�5eF��Õ̀=*='�4>r��c����|Qc|gr� ���`t�(ꎱe%����*��h�^Na��t�Iq�7I�o�(�Ԯ��㤝RۋϢa��
37�f�f����vUґ���Z�d�H�=�d�D�ǒcv�I��������O�[j0!ȡ@�w*��M�D�N�~��_	�,�UT$�~<_�N}�;<K�s�Y{+'��� Q�0?��Mv���0g��9K�����?�'M��ŵ������mP?w�e�͆�����.zϨ�F�n3�z� כ��V�e�e�?GMф��E����7�ɝ�o�_RS^Ae�����J@DU�!�C����sD�n�ILͨ�Sѡ�x��٨F�X11I���U�޿���kp����1ղv�8�-�	����C�Rk<Q�됅�|��D; ���Cꆃ<5�A��EZ�Qȕ�-���]o��D�*	��']�����H�n���a��f?�;�����tR�?[Q[9Κ�?�P���q�La�~�z:���p��?|��U'���1��&�~�E���k����Z����>xp�{l��w���)W �*�*p�:�#=@��|�r�n�1�s�������� k��-��E������M2���M��P�}7?���7I� ٕdp�t��(���� )��8-ג����?��8���7���E�Τ�
{���ibҫq��yG�y|�\O�;*Z���HB��@� �ܽ{*N2C��V�⏘z�#�r�OB8�H�h���4���C@��e�<̾=�f����9wJ��C2�(];�H[`e��N%�Ģ��� l��Nx�`�$�M{,����!wU�,���e8�g?<0��j���>��W@���y4���v��$s�ȇ����?:v�P;���r+쇾�Ӓ���J��=
"��$k�P�g���#:�q?����ϻB��[���]툻)����] L��K �o�k�Pp��bc�I.e��N�$�b�dc��Qωj�6T��~Yv� �[�D6GS�2�Tj��*]ZDT�ĕ"o��=�Gz��ɢb���:�mp툞���YHUj�˻���y|�@7������}6���i�����]c�͂��"ԧa��<у�e����	~���w����_�r\vȀq2�����w}��o}����Q=��ۚH��jaUo^U(W�eW���|�5V�s��)8���/9�jH�ˡ>�`j�>��;��iq.D�{�:�{����uC+����.��I9n�� �]λT�M���ng�H�+Q�Ý��+zaf^�ّ����AE��?�?����4�v޶p�BJ[Q��0���q�ܨw�c� ZKz�����d�&Qgl5��MT��p�0s��5m3���&�ѷO�J|��5eL��Osp2�x����ś���3\.4`gئ�m�����I-������*��D��^iW��G��(&�\�];��f�B�aOm1����\�c�t^��Ќ	Y�z�w����nOqM�0��ֆ|`����T�>�d��0���1f)�ZqP��7o��vR�_p�E���Oi)[�͍z��W��) ��Q��Ě)�dʡs99�h�>aG)��2��%Y*��˻7^��C)�<RT���Y��L��a���N紮�C�m.)O�*��_��˛��m|�ٱm�Ly��^��>��W�x��5���k��+�6ݠ�C	��:��x�p�L���P��^[rK?��D�-���V�u���=	��	{���կH��E�u@O,� �I���I ��њ���\P���D�������Nh�B�B|�kuׂv�W��BTF@�Li�z@���I|����'�r;��+�Ӥ�]�����%ݓ9�&��t��/�O�*rmnIn�[��e�lJ��+j�`�P�E��j��C{�-��%�B�4���4��<@����bW��3l,�ڇ����#ٹ��J�|e<0\��E��+/\�ىQ|�h�Ѵ$���VD��h
LնR#�Ji��pb�,FIͽ7�Q����V�K�N��Ԏ���c�ӊ�ה/&n�0������q����22��%eHL��y�o��{�%m��̊0hE��N�C"� 	���N�(2�젣�n��¶d�[�ŊC �6�V@*`�	��#|:��R����`���Y��1{��k�s��j�G}�{�b=��k�ZmZi1
���j���A�J�?�_IͽI���K�R�CXL[�O 2ª�ɓ�}���=*��beQ<b�i�nA����+��v�.~���H���4A�U#X�([�b��u�p<�ԯ���5I(����RE�}�Roz�>ID�>"�z����h�g����ӶB��9�:��O����*re����_��c-�gs��΅q���.�����"���߃x^GE\	�\�G�����)�}o_������w(��$�&[�s���
���"<�p�M�$?��>�b$q�}�� �H`w�¡}���6�ٳ��;J�i8��PF�@����.T�M�2f�������K_D+u����fZ�@�(>G��/_��#}ô�IU%Npo�G����t>�6�ţ��4����/TA?gn����}$�����
�Ky�;/����{X���)+��D�JDN,��ӨJf[�:�"N���S�F�T�;=�������]�)s@G𩦻�*R�(-��r9��J��i����\9�0���I��wR�?k�&����$�QJS�r��T4���k�a�y� ~�.�8��K���Rf�e.��~�ԩwJ!��̄�B �dA�BH/Ĩz��U"|��H)j�C��b����৚Z7��%�\Rh�=�b�_m���|޾k�.����N�4�
V�/�kˁ<bO���M�i�e��λ�;#�$��� ����l�@��˖�dy����M�zh�jc�`�2������"|�m�0�o5t�T������v���:4����=��H�(϶��b�O�o�����&�i�DF��1��*Ҷ�1����6�����spT�`�.+���� '\����p�0MȔr��:E	��MTZ2�}�ELv�^~��>*Z��;/}��u��~���CibS:Ki>��2��$
��6H���h���R�_��J�}�3��ڶ��Კ�[��S^�op�(�K<]�P�����s4��r�(�s�&��	s�DG�o��'a���J�q�1��A��!#:�m�	 S;��y�}ѐR��:u�ȁ��Ѯ+gI6ϴ6,�eB"����L(t���|7�V��ɗyE�JR��;�ќ �+,�����`ٕY9i8^[HBŉ�W+��#s;���&�j����{s' R#ø6��1��íF;S]bE�=�/`*c��g���*-<�㉅?jo@��u�]R$�WZ�>�ydN�2�܄��\���̲���[<�@h�_�EW�ג:���sy���ةHV��ѭ�d"�Oe�)Ie$�z(ޚ�j��Q�:?VZ �Y7���m,�{;�\�p��{*t�*�����G��#?��7�	���o;�+K��R��ZV;R��̧a����z��2�7�Ť�d�D��	����@2��?mH	���`�
���pT4��'B��q��!?~u��K���8�����Oy�Տ��B�>Q(
짍Xn\8�Rk@�:o<�r��K0��ǵ��g��7��)n��#|Q(P�z/%ֺU�4r��o��,h��
�5�7:�Y�nX	�6����J>�}a���X�~� �2�{�t,G������XY] �j� ꠙ&��%��	|�DĮ��ďF^ɎE�q����3�1��H��a�.h�k�X��g�$TZ�Z|+fD�����H�X̗3���s>6hg��X�����w��|�X$h��&T+����[k��� ��[N�5���:;RqM��g�~�K��A�9/U�(j�,���Di����=F�`��\b�I3�N�6�<��>��ަ靂���o���B��F˅�?��
uI2�g3�lG��l���bJ6l�&��������f@��)�~@� ���Uo��ʄz?�6}9�*�ݜz�eA�Wq��Kgoa`D7SH�w������/.b��`to�o��úh�h���q�5�~�I���T�����[n��-.y�DW�	�:�tv/[�>���R�`\�
#��A���;���`��}tXg>԰{R�Z	R6��y"B��E�=��@��ȬTImf�FyKf�uD�4����^��@���P��kW'�$�;�z=k����5�՜yZ�#������l?Jӣ�ZK�QI%W�yN�g�Ux���$?8��r�%�S+:NJ����u]��(�;B����
;:8H��(u�ͅ���aɥ�������~���C�Ɵ������̖�ç���Z6*<r���[s�؂<^&�͌���G-E}�QqG��˜�Q<�^����.Yh��M�Iid�����ɟ(;B*����r��K�#�.�f� �#ο��9e�9Rd��z0��o$��w�Nl����OM=G�� �n�9��KVE���U���YLR�M\&��ȜL��p�.�w��X�M��`���/��c=�ʑU�5�3Qz���'������0�i��!s�I�"8�?l#�D��ˏ�i512mM4Y��,]�!�b�����l���a��G���'!St
6K���b��k�,���Zҹ����ȣ65:�r�_�6��`�^`KV�������7��Z��wE,��O��~t���j>�jW�
��=���jSҨ|�������������v�Z;o���/@��������%F��P}dڻ�Ld����9]-�;F�U�����1�9��,536Tt�ϲ�儝@�M����5�l�y�`h���K�m�%ț/y����s�e����E0�v�7jQ�${��0ٰ��_�G��
)���,NDՃ�=+�2d�x������jVV�A�v1:�I�)�������f�~/��{��vf'}鍇]�(0���yu�O��},�K|e��=q������D��C����w�s�C}{Ӛa`����w����M�{U��m�ڴ-�e��z��mX����z���6�0i�N�Pb�Q�~eM�����g御{^v���<�2+^w��P�u�j2�&�s�[A��$���h^/������x�� Ps�����6��R�*ٗ��A2"�b+��4���:�5�޴N�y(��ri����s�|��߄�.�`�1��a
�C�-t��F#Ԍt��6~�;��]��u	8�I�R���j)�����Wēl��������J�~#��S�ܓq��~v�?2�F���Ǹ�z�����V��ʎ�D]��	�?��_N4|����g;��..i�P�5.�N�+�5;�%+��T}{~���;�F��խ������i.�������:H�9��ئ8�+q��?dغ�Dh~ʬ^���T+t�(X�>l7��I�6G� ݃�m������"R�D���w�J�	�X��=tsR���F�R����h�a�*�ؗ%O��*�B��BcTM����
�5SM�)��p7v-
q���8h~�e��ch�_��`�X�6�U6�]>���L���d������]��c�m��ÐQ�k���`L��2ydQ��F���f*::"w��q�4������]q�sid���}��=N��T��

���6K�3�ynP��f�7�1� �y�'�C��Ⱦ{��ywgFn����f�Dc�A�/>Y
��mjӪ��J�쨳n� ���q#���5_��OoZ.����"�jZ�o�M"�9�J�,�4Cu���f#�'�%Y����� ��^�Ԍ6����,��4��z���_c��\��S�?��|t�����HO�����c�0�&�T�qIt;�Y���@@��o�R�C�3�Ir丯�k^��k:`4u��з�����N�'g� _��V��Љ|v���(C��hU�����P��a�_I�K�/s*S-Y �RĪ�-攌@%���[����-�݊�U�\�챨I�r��ӽ.����a�/ k�i���h7�Dh7��8y�5*R�e,�����.Q�;A��.<R}1_ES`��)}��{���,��.-�C�V8�U:�����Zk�6��I��o��+�^��º�Z�j���	���ަ����"3�%KO���dC��҇�N�^�%7� r&��qznl�i�I�E5z!-�۵��<̤HzK�&��E6u[yM����k��1-h[�[��A�j�D�1]rU>�5�Kz�P����ȂS�_�1��Щƞ�jo�� $���rv4�x�aP��=��a�0�6^u��-���:��L_��X��Ѷu�0��LB��(�S�@�g�;��u��Ɣ��gt�<���WLS�C[ȫ)�͑oDGz�m�#�Js�C�@,�G9ؚ���b�Wd�4U]���k�p �$_��0���Z�mt�g�|_*U���b�#��~���v�V�;��L��m�U71��[� �e��D��xx��s�������G���r��J3����z� �F9�|�i��8�I�g=D��6N�Lq�h��	�S�ޒ��~���`T>���u����h-ԟ_C�=ߔWOxh4-M������8���	�>�%�J��c��t�=7,�P�Ɨ��*?��&)�0�V��iֆS���m���m�}�d1�w�I���I�����;�������v�T�v���t�󥏻B�b�7�5|���
���
Oi����öN�Z�ݖ��s�>���0p�_�?��8}�W";\+�|ު�"/ ���E����tW�{`mj��f �u��%��r%�9��)�� �⍍&)y���K�^
�����&�J�	2W�X�@\�Q<���s�;={oF�d�x�܌MK!�Ğ��,�o�X�1�E8�^:E�!%�h���Wx�"�%�g�g)�=E\����*v$g7��f�wgX�	��Y�=���5aOV��L�ږZ�5!y�
au�L��+wd˦�7�Q"�"��￷�DBt1���ѻw�ڸ��_�I��R ��O�+��鍆�/�7�.����z��)�22�#R�<��T鹺�J-�u%�GӰ����j�
��_a5�E����w*e�a� �S�d1����#"����"[I��	Tk�	3S�o�J3)��`�%��B�}�9C�Z����о����/�[����Rav��&m��j�p�;',,�K��x;�)5��b�5�l�5C(����*��#�!��ޤ�[�5�N��W:��DT����6�&�f\�*Ȼv&�����״�hH4{���YSD�p���Ƚ����O��'����'�_�x�V-|RUvZ�E�%=��{�tӨ����1�K}�^+�
^ZC��O�|��d�#�s����O�!Wd�{��D�2U�z���9�;D�ؕY�t����Zƙ�}z����_�_�;/���8����$�;{�I�wKmZ�zx��W!]���pf�>蘶�q7�j��2���5�:r�L#>0	W���Q#�7b 0-�y�+8�0�0�o�m��]�۶\\�\�Cb{ݏ���>p& @�K���ߣ��c�
Zk�7^��I��X1�,^}q��N��7�����Lsk!��.�<;Q��c���eV,���w�k'u#��U�uZ_e�f��x$�Q��H�Ń��;w�W���B�M��+/h��L\V����$�к�@�8�c���kѺ�R� -c���be� ����A1w��"��Yf��q��>��������0sy,�gZQ$���ou	��bCwZhFf����P��t�+|ߖ[����T����%^4�61+��ATG�ּ�^%�����	1"48� T𕮰�Q����n�o�y��� Z�*�c�D<Ld+1��yo�_�"���4���4�P�X!��1�3)Н9#���_'G�<!?r��M��,� �d�S������ܺM�gu<�!�b��g(z�lP�U֔�}iHC��{Pus���p0�Yd�S��&�ĭ��8�B�8+��W�R&x1�^�Db�	���u���?Q��v��T����eK�0;ﲂ��	��}ŧ���W�̰�[O�&��s|+�|8�0��-�j��� 7�־F=f̥���Γ�����!�\Q7}6VzA7L(>��r,ǯ����~�b�6��w��xK� ���T�L�g%�9���K�6~���8~��e��;ib�r
��ī|����}�@��Q�D^��>1���U���Λ�S_�Ԫ��`0x���|�X���8�p�����9���᎖f�jF-�/�+�w� a.]��9ƥn`˖�Ѩ�i�Z*�ߟ�"��t8�-�W�Lf�Qo8� �|�'���A�{0���`�&�&� ��1!;8MQ/A�`���� b�~��H5˅x<^�����R	>��\ zXZ��jtce�q��E�݀�E1�k����A�2�;S��Z@6��g ���g�՞j{�j�s����۶:��D�H	����v߯ӭU�չ��ik~|y܉8�kt����Qa3���4���
�l�n���x�c��抺F	04�Gg�\�'}b$�w�[��J�ͩA���f^���+p8U�����/��Rt`Ɗ,Rb��������rVQ�g��^��/�?N,$�AU��rȋ�@�x�s�xp;�� `&e�VaI�3C �b66�A�����ȸ�y2��dme��c-L6C\P��ܴ�x-)�DbZw}y��3�jɹ(�����H�l,iV�R�M���Dre����+}tr�ұd�W�HIr���LD��8���'?@M�9���f
k$�!��!����R�ѿ�?�M��x��h��lWv9�[M{*O�J
�6�<.����M.;joLB>#o��A),7���ظ��u��Q_�zq��7~�U���"aK����5�FW���ޘ���Ph�&c����v�/����m}���7o�w�+/���"�y�/	hc�=���H�\��
+�*ϟ�n��x*A �y�Ǐ2l����2E�y��7�B����ؔ����IH�� ���)���у�o�!;QB*�L���t�si��4 �ħ��`n��0OQҳ��������<z��\x1'�5���wk�-k	�<ܟBi^��/��;X������"!t��ϊߣ˃���
��@���=�{װ8�C�Or���P���b�=$]�>%��K��IB�5��-"tp�����Kz����������M�$���(����_
Ь;�=��Ѥ�]�
`} �/�E��9xI�b}9��fF�^��	��W'��?��nB�a�Zb���}�y�"�/�t���h���>�|�]�"�<���������*x�@���m�`��x����T��;e꾈&eF�%�4[c(&i(qu٣p��-�22"$É��?�kZ�؃�`�"GEA��w�-أ<���#��#2HC#X�3h�N�V�``����a�Wf��I�C�\ӊO�o52B�|���N��V�/�ԷE��#��V	��r
N��DS1��܏��1x��R���}=��u�m���hbj1��J��|S�n���Vfw���@�y�PhW'@����FdvO�z���M��?M��nZ�[�3�s �5����"T�r�M��]����Z����+���w,PF��$����Y����[sO��Sٙ�A��G���bz�#�0�㊠����v�vm&�V޴�a�SԮĆ�_����Z�\�H( ~82��FhxP�0g�w���y|�����N�<pM��Ȩ.V?UKg���CA�I�_�[Y7D�!Z�0?�C J��8�<��tj��q���iew`�������Nq��c���q�d0J�/[�6þ,u4G݆��u�8Y���R��ܨ%Gf�Y���fK	7#}�5x3�+T���	��D�$Ax�i�\��UqijY�"�!.J��O��jG'�ը�|K�j�I���b0��Sۙ���r�M_���X�8U�9�<�RB�;9�T{u�nޏ�=G_���'��Hc��/�6�Y7`@�#b��+����j�H���i��XY׭�Y� �
ގ]��?J��h�=@��tV�[����$�^�]	g��<��o�QIɣ�%�v�XO�B��q�v^ �y����-yZ����|p�v��ۚqS�U��0���Ǐ�#��H��2�l�r���vW����
��Z��ܬ����ތ׵�x^_�)�[��� �ǾYw:v�\G� (;�ԁX!X4L���Tɲ� ��ٗ'�h���}���K�� �$�g�P�'�r���]me��mV�=Yr�D���L��G�����H�.;��$̺��� G9���mo�i鷺s����a3�I����0���T�S5��j-�HX@�@-����I�&�O�˅�[��ŭ>�Ku
��E	��_�����7��Q��6:זr�=�9zu�d'��y�J�f����]�}8�}R����Zjʌ^�4����i�Fo���s����F��O��^����M%�ߐh\Qc����P���0s����sWA;�a*���N�+�~~Cq��rw�.�r�������ev�zm��5��Lk��@H��r�����F�Sa �����]T%@���s���D��Bj$�3b�$���s���USs�e}je�c��8�8
G�JT�`iV��2�N�����o�3|{	cX����UZ���C�q����蚆x���'���5�c�����S�	��b�����0����.eC���uJe"%
�?8'��.�O; y��:n�s�)_���^�ze/������cb���IU�Ş�=}x�W�����Jd���)霓دh?t�gi㆔VK��kn��86��hlԮG���5A��A����D�V��΃�9%ň�Z�j4zv���#�S{��f?�I���H�y>��.`}0p���j�H�ip�!��z�^\?%?�J��˝�,$|{�J��k��Teǰ.6�C*��O�ړ��_珞W:騏UI⇰�gc��Q{�w�3Avl�缅T��a��W�e�u�O��>8v��!�-�Yˮ~Y
@��
_;��W-9PΨ Kn��2���+����������N���Z4��k��j��Q�j&KH�*���ϻv�`Di����(=�F�6�ih�^�VH m�E�|�����?/v2������{��E'Q�(�,]}�4������Hi��Q�d����wZ�QGO���7�pi>�:c�`#[4]��6��Pܵc*Hn��P砛�#�B�����C:���b�PM�mGR�hXY��S���H�"R&d�M��:��Z6+���u+��Н�cM�!_��N�_>�;�ȏ��f��*��Z78�S�W�UM�KGA?��)����2�>�ZH{eYg�*Ŗ?�K�>��6ˉ�THn��	9lpL�0��,�����ݽ��*���3��e/�rڃQ�j�s˅�k���f����B��f
�S}�g	]�N���7���� �1_�⳧z�hO��B��?ծ���$���qs�.�]q�m%����MhI�c���F ҤY+��wd�)K��lݢ���_#���&��E~��c:߱J���Hʇ��~r�L�9���;*?�&�}=� Qc�ta"�לNᕩ�`�����vzU�*�y��m�1�9��9�GKΐg��<���G_����4�#1�_wL]6�N�7���<+J̘�:av� ~��� ��K9�[IH�k�$K�7HQ�5�&�������C���~�����q��a=��쑓S�m��+�j���e�r�o	�3�l%�%�����p�,Mx��o���kz�^R����q�[W1��>ۘ��<dL��4%cm�g�;tKx�@BF�	�(�{`����)D\_���!�d1�?K����]5�pS�����|̻�g�4������K�^�ٶc?��(���|�@k����O��Y�x���\�L�6�R#�Ŧ�q(���P��`I�3ow����A�W�4!Keb�,��,C�C՝�9|=&��k��-�'�2�Әy���y3n�@����l}Vtȴ\(ރP���N`e56C�(�x��G�����bɫaa]V���@�x�>�I�~��2/_' �k|6^	�-��������EE/�sh���+��H͓�ǆ
l����<�x�
@[0�hթ����[P,��4Vj	5	CF:|�T0�8 }'[� 6�1f*��cؔX���ehȯ �z�v�;ˢ���\��:��vt�+�v1��y��y����2���:���af#�N��8�3�?�����i~�㳗���hp$��B��O��*�����/'�x��4S�ޘM�CG:��1 �uŅ��p��O;��Y�_�Y(�uB��Wx}�~�����u�#;(,/�ǡ�|�!����(��5������(���	s�'�Xޢ��n��"��u]hBFa���"MU�St��N��b���7z��}j����? o�}���*�Xl�s���4������Y�b�8=�k���i�s�ZZ�b��=`J&?��g��r��	��#��ZӪ��eG���لjL�(=��m�k]���J���Z��B���z�7�����뤐U򉝊�8K�"�ڨ�T�F����W��7�9�5�<9Ò��/��]�	y"b:8XV�KU3�}"��м��_�+ȬJ���U�!�H �H��뀓���eZ��Ymz��Լ	mN��U��HR[�E�*=d�	P9��Z���__V��2`x��y-�o�b�I��ߪ�����V�܍�AS����.�Ж(4�b����K�\*�a:j&9\�0ןNyʾ�*kx�����EtH��Z?m�i}�<ј�����
[_ʀ>,}��C��5�v�QH�A���yK Jz%���`d�!&��m�θ lG�ji�؁�
�8Q@@� �,�y�c�R����[$~�Pս��w�G�O<�=	�c!��o~�zBt�!�݂��ywjf���������s%�Vԅl��5�A�>�j�S�RȮKDZ���{Z�mz�bl��%V���Q_���Wͼ���S���U�K	 �ʢ�m�\%�K���ॹ��mϝ@r��L;�j�A��̦G^Ҧ[�_���d�?�������rNf�j�Hkc=�o��A.}�hK=^�$�������;�b0�d��M���&k݌ Y�\�?��N뼑�R�+�������,1$<��JI���Q���_�+:���w+��Z��DWSYװ.�Tdp�,"
:A�3�3���y٫i��Zt�m"r�њ�W$���2�y�C}C�d0��n~�iE,�k�8^.��
jQ��m�xjTc�ęw�/��_(�+�ͩ-Y��UU\VVg�yH�]љ��
\k�NYX\�@���V��ȡ��k�0�Q:�r�Z�s���]� �iDW�?l���d��m7Rp���*�Uj/S�L�����b��@�T5	N���Wa�4?�
�ա(^��V^aA�Y�!��:5����Z�c�,#~�O�!D�SYW�<`Yz�3��	]����}c߱�Z���g�{� �?�X�r�&��8�M�t��٦$��,�������A�[/xa�y��R�����=q���)����N�58��j5��`�\��g��v2�F�VtH)���۝p8��:O�͊%}<ы�췔��l��eu�x.����Xˏ�^�4-�h>!�)ˤo��C��0s�Qrv��[#�&w�$g╄���JCn��FKG[���ʿe:���!<��<ä��3L�5EJRK�`�m��,}yK�}.'H��L��i����\������$��>
+�MN�.ɹ"��١L!!ӫ�>O}���5ΐ��#�%�8�,]5�G��=��e�i�����,H.Y�����0����<jp��L�ૹ #�A@��w���ؘ`ي�K8���p;�BRd���R���E�B�����иHӣ^��(�n�F|ኣ���.Bz�V��� �@m�ܞlP�<��Z��훷ዛ�Fy�j۽7�*�@��{�L5g��+Ro���a���j�2"�_����#�3����1�K������a*\u0�گ�T���x�b���K9g��3��J�0m��%���+�qeЖg��l?0�~�z��W�p>cg��bñ���UBĩ_ec�L��_g\���r
�L�߯�Uٳ���f%*Z��F0�V L�k����O(��u���~F��ώ��<C�����i��{]js#�6a�7���9���,媯��DZyP�`sv�œ���W� ��1���@��5aE/?�����FwT���Z���@��ڗG��G�	���N��"��8��P��9?�2\�&���K�����'���02�i(QZ�`9��f��D�tS�3uH�G}�
��w���	?���q5g�e������5os���b���%��ǳ&
�\Oҹlo��L	úD�*%^f�U�qvמ��ry#�����������ʊ����c�k�
<^fa�)�������X�L���ܕ��+�X?����r'^)H��I%��$+wv��>5F��� O�2��A����,���te�t`�U׃�Ϧ"i�`YO<<0~.k5��n`����R.2��}c��Υ���"���v����3\6߆R}�B��SǢ��T��(
�bY�:~o���`/���L��3��G��l+�����K0�����YG��>ۛ��Q7XZ���l�ZW����S��3�����:No2b܏���H�q@�vG��p�J��o6�ƈ 1f��9#�^�3������x%�I
���Jml�Ea%O�%ȪIY&��ȯ����X�)3�M0�\�h��l��/�-8O�� ���� 5�|X�ʆ^���|h��pA`�M��6f8�o@1?C��E�����rVH�n�d2�-���z�$w�.c2�GF���m��Á'� �n���c,�R0�;+��I�u� �I�)���>��`H�R12�<xl�{��� ���I�9{`�^	)[���`�RH�8��۬B}4!��:t�=A�A�m���YM�}��N~�=c�bm�"p\Q�]��H������
��</߃n���o���S̞e�������/;Z�0"��k��<��Jb�]x�.�1��^e��� O͵�=� x�S�x2�����m�CO�v��t��R�;�}UU-�1���J!�(���˖�rX��u k<�'�l�I�h�e��+����=�<3�����gĳ!]���}������`�0��%%�.c[��x@�9Hv �.��]�#&׾�j�>y6%�웏��w�ba[��dJQϢ���W��2��N����S��v�zW��vZ"�K)u���^ eަ7�O��Y�3c܀>_�E�*�g�.8��󊎯%!��}`j����K��K	�M)�W�H�Ku5��� 9 � �>rx�O�:�wS{�_���6��'��z���챆_���GD�]7��
�^;v�V�'j���:�QĄx^6B�лO��MP�����O�}n�1��HH������	M�o)~=���f�˼�-�+}EMC�ț�{}E�J+�BuJFfQ��_E/9q_+��5lz���\�r��1�8;&��:]�6��M����˫$�kpM���n�͐��h+5YUݱ�߁i�"5�M�{'�����2D��jE�*�+�q'0$� �!-��/ ��|k.lv%M�Ճ]��Z6��IVcA&D��	Ŕ�m{����5��9���7���G_U���\߃	����}�x�\]/<RT���h�����~	�h� �SZ���,�-�.l,���
�t6/F�Gj^�kW�#GAcB�$�
���?�eTuYY}��Pt#cCI��+�35p��֎i6c�7H�⥧�uK+I����Mr�*2�T��;@� hUi��耉,��vdB��كJ�c��r���Yw�=��X@zE \uO��T,�T\��;D%Z%�/M�n��N�Q��Sf,����Ql�o�M�ѻ� �u���S�Ɂ'I��;�]>a��]��.Xz���PTp�� ��H4A�^���(��
:��^���a�y���C�ҩ-���7��������Ò��@>�6��}��a8�D>)��s2L9��.޼��IW�K���������4ԛ?+c&�h�"R�<�"���2�!Ok[!�ڸ�ǚl/�<�?�9�H��v)�M��g/GH�"a>N3߮��.�����)q-UMt��W��*����C7O��	Љ+�9@�a\��a�Lm|��Ng�v�![^��a�y�kz�K��ۧ1>�}����j"���B�����%;xL,����U���2��'*�нc������"��t����Ǟ����J�-��{g�[7Y6%M�o�sK�ʵ��mu.��24R�i߳c�3%�j����&�b=z"�Uy �@|��7�/�z`�7ܷز�L��uuޖ�����
�f��٧����r��^���%�R��(�X��dr�Ĳ��մ]Y�R�T�>���ѾK� 9���rNU�CWߢ�w�S�bO�kntc�J=!g���U�ײb�b�;$BP�ϗ�6�6���>,~��8�n��M3�
�O
=�ٛ��Q�6J�8�3A��r�Yqp���#S�[��O#�ȇ�}��]�R�O�˖�)�8�f�<3r�.�:D�I}��6d�x���O���@!�X��S�!��^�ڞ�7�GB��ԁ�����J���-,�dN3��2Y_,̯�74�T���-����,&�t4�H�5x{K8��˃�:��i����Z_�e#x��C��&��S��{nv��L�L�]�рu,��%;����l���mI}�p~�J=�8Z�{����7�L�����y<K�e���b�Jr��%=/�sP�충y��Ù�[��[faJ���#%�fMu-^�h寐}�$S( �Z ��x��|G�?*/7#�����G���5Z����؄~K�h��y��(`���&��ܞ��G�ʈ���Ĳ��$�{�Q�{iM$�k�3|�
���i�S���6����Ii��^�r��@���Y|mh��G�-�u=OA���r4�$DC��������/�7�-!�s�7����8����zV˛�W,e��SI2^<2l��^O��]�?���V�2R0+	G/�̽���8L���!޴�Vn����:Πk��z:\�ޱ�K�Ko�0��^Q}��_�ߵϊ�*�����1f���(�]�E��źlX��&��(�t�ٸF�@���"�L�3#j�R���@S��{E�9*�ăs�0󃍷!�`&SBU�V��p0'�rcv�#���<岪�ff�[dI����ګ���0��8P4 N�������$9qDB$�̤̉��u��!q\��b���h�:R�Nz?�#:̬�Cڡd�g�q�#�Iy���b'�D���ŵz�~N0�~��kF�M����ϗ�tid�Y!��ae��*!"����md�^+)V{��{��/B�Z�����I!f����x�4UL����/�e��%��s�v���W}��t�rGo�A�=�@��jͺJ^�w�����I�^V�
3�A�MYA�I,��8�:��*z,nDƣ�'n��o��1B��>���G4m��ػ� 0Q��+Ex�od�]Of�3�z2��c��A*/�mzEAKĦ�0�YDA��x������x�	�H`�^[��R��#P�'jˤx�Q���V��E��c��Uɰ�������k��	�w�������"��P���+9� ��Z�:�����i��u⍝�f��{;��uU�r�G40x����>\�V��	)-121m�)�L�u�������o�)ԡ�0hmKh)�%��Pu�X*�ȣ��h;:_w[� ~�3 6�n��QuR�L��1��Ao3��8���|�2�"<�J�=F�B~�����=�6�3�_l��]�6���A;�J�M��4v��pQ��(:s������L�׋�	t���@ӡ,��ؕr$f�,�+ͺa�w�'��H�iJk�
��T~�r��L��av �ӿ�kk��Y�VlWD]� ����n�ntyYe�o|�F��И�m0S�IBa�X�W���v���d׮ΰ�9�?���L���� �ɼ�}p94[��X�g �U^F�	|�a뎤��Y�$��n���Ȁ��^Qrdzfsj_�X��?�س�\�;'�#��� ��M���������x�Hco�A%�_�y?1�����|	�R=��x+)�}�[U�m]�׷)�P#�/���̝�M�������)��5?�J��39[lz�����}�����֝�*�ڹ]gj 	�m? ��tǕ�z�!����N`QO��3'��uL8v�5y����z�~���r}b9���0���m�n�c���3�he�W]T�(XB��,�v�������F4��-��|����I���S�(A�O�S*�3h�������p�t�p�s�iS�6�j?pYQ� [RK�f=���\]�W<Ҿ�� ���9�n��F"�{����1���8�e!M�30}�� ����t�/��G�s_�^��ܴ�3�:)��@r](wS6�~��7��e�E�j@���K*��eTKY{�5�\QK#�����*���[E�	{dn�T��B�le���v8���2�P�G'�	�܎�-����xSy6.�N�2H��XH5�g����V����,vc�ed+R����pS[��44���m�C�c>��%�"د���g�����-QS(�x��~F���嵯��
X�x�9��i�vI�?�@ŭOK�F��=�����A�f�����b=�I�x֭�C��|����BkʝV�x(G��Qz���C͡�_�:ɀ1��`Ս��pk����5q��z}~Ft��y�>�p ���9��oT]iNfQw����f�l�Ũ��Igh1����� �L��""X�*\�O���H����\�Ǉd~+1�X�܊��8�;�#��H��r��x��(���I��#8)=���e҇���`1r(�j�>�+�E�"'�"���8��S.�v�kr�5����X��ˑ�
�7J漣��S>�ė�)�s��P�	��>oKI���}������f��YI�E�k������`��h5�ϫ}�]S�Ak��D#Am�\�7�i��T�i���U�a{��9�F]f�"h�=<T!
b���.�W�W!1G������<�6���ל#i���4*Xj���_��J�:5N�.�.Z�b�M�f��G���*���*���P5�G�����lۙ������<�[<*X���B �D>�	[)S��z���^�.��A�� `�DL4�f�G�+\Gܓ"�O��*w4��;q,�,��D�bo�����Ҍ��>H<��r<�Ucc~�M lw���t�iw9�zXc��6U6�NXe1r�� +�4Rh��cݣ�|Pڲ�\��e�!St�L��i���(L�[���4^W�2=X-�S�IqP�/�zK�"Gׁ�Kz%�Յ�] 5���<�����B8L��G9��:�hd�Ī{����>4�r�ZWrgkQuo��_5㵸��z��KB�+�Y�G��f�UJJVMN;DS���Z��_��Qj����B.@*��:�O���v�F&Cv��,���-��z��ma��:��	jFTlWCD�h�>���w���F���ȏI�"k�@�y=@�]t�|t�t��~f�T:Ă��<Ƌ��쬂�j����_���evG�+2��r���I��W"&�k�Ofj��d�o�D(\����S6�OHtϹ���Z�4�
�?O?���#Z�r[L���~9��xPpJ���Ve��5%j��̨+sKd��^�v
e�*����%mSml�?��4ro:X�4���<I�9͍}�%&����R��{D�3��Z�*D��-�B���
���qD9{���"����%r�x�Ѡ�:A:�[��Y`��/�6��G{y��2�e�ϩʌ]%k3Z��FT��(��*x_��G�f/L>y
�٭�����@wQB�SΜ���}�`���hv����W�	c]D͌�%��Y��(�3ٌ��1��6[�����RL/�JZfXj��\7����[ ���/,��<���(�{�K'JŽ�yOZ� _۹��?6\B<�X�r�u|r���%��nh�7����إ�AYՖ�����:�]!ϣ�����.٬׾ܸ������t�.&]a7#���,gȄVc��zģ�
:��s�r��9�FTFg�f�Z��!��EP5'�1�@_�ǂMw�Z�Bq�6Q�]Z2���&]�ژp�,-�,,|�~�D21�\�h�?!��F�a�\e�6ҼeP2�-�̓տ�-���N��.�T��:��f���?�>��FG,{=De`K�h���㘼BY�������\).ז��ؤ��N�]j~�0t!�i��k�G{.�P)8Ŵ������M�,���ύ�p�Gp�Qy�#V[�ɥ��� ���2:ׅ8^<��|d\@Ld%�IZT�� N/���/��Vt�VIx�Uu�����c8�;=b|�G+Q�����9b}Rٲ���W,6 ķ����'�^�=��~K���5�&<42r��Z���pza��v���p�uʏ��-��|"��j���'
�`��m��H�A1K[,yR��S�n=y=ғ�QJMw�b������9�	:��5�OhK�i�����O�WP�K>Ƥ�B65�ڋ�=E��6p1ki�/����:�pL)�:��_�߸���܋n��k ɜ����B(�C�8�������8@G�){JR}�N-�{Q�����"�����&/
h���51��}��q�?���:'i�l�����f�W+�F�_��^3��쐠���}�i8�*q�5$z���`��B-�\M��:	��L2���Q
5m����ekt1�m���"M
H91��$a¬
�3{P..4Z9�l3�f>�u�����[�z�L&ʽwf�ɭ�u��m���CH��Ibo�o-�z���+F���'t�`���0�S��e�ec2�pݓ�;8�l쩇.���'�I2���;� ��Q����=,ѽ�N�Z��ƌˍ�� 6���R�/`Tv��o�z_� �����t�����:�l�� ��œ�*Ww�2X~��lJ6��r@�5�,w�ݩ҂ⵥ�f��Bg�{8`b׎�
s����:e����� 1�V��U*֝���������!��n����r�l�`R<�:n�7{G��4����C"�KS��0
۠��E�$��F�����C�[!�<LI�����I��$�G�,��Xo�џwԑlK�ޏ�)�J	TՂ��<�	wIڛ',h�6eTIև�lk��m[
�ɕb�3�6֌���2wjۧ8܁�@[� ��c�S����է�9��w"(5��Ǘ�`���}l�b��E����{��|(Q;�AOA� ��(��+AY��1���b#e �4�4 �%�����`��(Ĝy��̽�pB��]?�̈́�/���*}�u�U���S)�'9�n]6�.;_�ی9����U|·��[�a�'gl�0D�\�Sb��Kq-`��(:n��?�ɗӚ�i�$�+�h=�ӥ�^s<<0�t�IW[1l���x7<�@���}*5�_z�@��$���(e19���u����0�A�8��/�{�B4�^RT�F��{�"UגQ�{Y������t�[v�Տ3�}�0e���e���E����ڕS
��qi��3pG�M�2`��������DD��.�F��
�������g��J,�7���D�h.��,�`]���c�D�육�a�	�&K$}�ũ�� b�"t�}"u:gո �+�0�絰"��789o����9�m���T�BI������E�Y�DJn�(@ 蝄��s树#r�{�N�-2���?�j�M�[�4�w��Z�g|�\uL�#]S���<گ�*�����5�zb�+�:B�Ҙ��"����أ_��ؖϘf����B�D 釅��K�:"��y�2�]�w�U��8ģ�U0n����FV�$�y\��J���S�
��Z
N��h�)��h�m{��[x�b��~�)E��	^��W8�Pl�$���щV�,�-.G���?��V�tk��^�w�(��M�L�l�TK�mP؝S����7$��.\�r�S�Xn��NWĬ#�����m(�-E^&�?�������k��&�Qc]�{�=J}
��l��XM��I�d���R�*��B'�O�уJWe9��f*<��.�p�04�3���R�� ���/ݫ�n��tr�n|���l� �S �j��f�5ět��?���� ^l�SLb�ճwW5�J_p��������1{�|�7��3����I���Y�a*�E7���R����ښ	R��Σk7�H��c ߮]������Qg(��j�M&礼ˆ��=���У4��4/��hV�x�}��[����t�
?%xx�4
��XIA��yd���s$d|����֌^/�(�~"S�T�O�-�Z���ӂ�)(v�{t���ȧK`$*�W�]Zr*�XiU���� �/5���H��LqC�� ��<��W]�'����a)�f΀��O�=aY:i�VA��r��i̝��-oo�O�&a�o�@D{�L\�f�Ս.:�BcV���D˵�%Ȍ׍\��������5�r�ŅAƟd��K ��{Jڿ߮�Ƹ�z�~S�M0���w�I�lndt��
�ʙ�h�V��l����Ι�����ꬠ�"[U��ҽ�$''� ��U	S��3�u���/;^�L��Խ�4���^�\�>�뀓0f�"И��bԔ gx����cN�)�U�3���juA�����lJ���l���L&��IZ�tF�E�ߌ+�(����9 �[k>���.qJw�?��Ȧ��!�Ŵ�*�O�?�N���>G��$7�o�:{w4��x��F�rP�i8J�#y׸s.��{�ݫET��.&��>J;c��&�M�C��x}x�'��ъ2LG�u`��M��GD�߾�1�/�����
A��eKoՓХ=�V�|y$������{����B �]��e�wɝ�kr���V�ڞ0���g��}����c��5�}�yn�ꧼEd�׉���!N�6_+�)7{"�i��}1�@��~�0���d��CeΐS�>kF��ڜH2�V��w^�x�;��"��<���H%���f/��&�Z�A� !0�Q�������m��H��v.J���62y蛺�qw%0�MH,���m���Vֱj0W��2IǓ�A7&�٠~����H����/|wף�A��%.�*���W_��nn�W��AM��wi���ڳ�<⹈�24�t�p����Awb�x��(k���U�~��CJw�:y��7��]]Z95��N�7�CL'N�cm�HbW��rb ��۩��`xQ9
��syP��)w^�,��Z4RDɁ��Y��$�Ɠ�+a�Q� :�^��@����$a���� ,�Ie�I�XE�s���N�1*+rS��h�%�MJYK:�*�?�fx[�L?�k��U���B:����x��`�T����r^|��0N5П���9j���m�Z%m���=���Kg�VJ,�{��hY�]�;n�gD�����Q����P��!���{���1�9ag>�w��SmXk�ڝ!�v5���4D���z�Th������ �����*���6ه����M?�B��b����˚%L��=��'���$�2-�:�J;5��a=�8�һ��DDa�%9�`���@�;��������hie��n��v��S]:>��S|V�r!`7��b�)Y1�g'�8>1��A�v�u�^�k�VV֪�4]1e!�i�^9���D90�$�h���R����[��$��?��(L�@����d{�N�m����G� �#o��E:n|,�H�g���q!�]���V���q:�SY��=�z�m�1�A�r_fMR�X_��"ֿ�?��2,{��#qgj��ɡ۔�W�Ps��R{����=[��A���Q������Ha����[}B=ՀH1d�j�� T�%�h`����֧��]P}����݈_�&��Qnj=�T�v1�w5� z���|p�����]O�JJe�ټ6�T#�kn�B)��.#��&��!��.��'�'1U�Q�P ���]��εR���'E�e�p�e��s��I.�8~m�+���@��m��i<���Թ~�5����\���U%xѬ,��ƞ$c;'���jz�X.�V��@�`?���r���$�V�Z�-����A�r��ps�c��"�����T?dMd�#�/��e0��-8R�(�構��L�q�ڻO|��#�J�i�*��,SfUH�KH�$,�o��%{���TA���y˞w��E��3������`�I鳥��&1a|[��{�"A�Yh׸�І��wN�$D3mK�y�mr��i`����7p���ތ������Z��j�T�'��e�����q����0ۧe[
��q"�Kڳ�_w�B)�s(:u2�x�������#u]r潛���R0jd���(LS��n�x<
�
8�.��0'�O�S�;�Q؎?��ʴ��&O��SFS��>��G��7x���?<*Q�P�I^��v�?U��T� ̀˼@8���������5�t�U�~����#*C��Q�6fj��9WD�+I��'Rk��,�?W�]u����Ø_���!$�vf;��%�����üZ�_P��ۉ��vss�2�S��X�D�q�*e���D����$1*j0��ي������U���ڷ��~�/�&��9@��\�1�"_5|}�P���0ޤh'�鴄Q��["K&�=%�b#�^@/�FB�ޔ'��^�+�i������6ʏMb�]g؅h��7�8�e��M��%(fe9C�-��x0Aj/��}+�Oc��wW$ĿE����i<J���|��$Of���V<��_ʰir�������N.��DT��uk�rs���J2	+,'��\@��M]V޷�c{���`z:����sмIP.�	!@/�P3����^޸8^�@G;T���#��~r{�K���(&U#G��]k��ag����Q#��U�O宓�>L����1�.�{{���:�蒈vڈu�{7bc�Z�Ñyb�Mz���)��0�]�;7*���Y�܋�R��Lc���J���NM
G���^@\s���*���}i�����JoZ�M9�z�U_���һ�_$�3T���M1���C>9G}S�L�|�����n�M����=�Y֣I���b
1t�v`v>vZ�� �3�-��i���8����g��ʆR��g�Is(k�Jfk�
�;R��{''�<W#��,�+_�8M�� ���:�Q�nZia(���h݇$��!��'׏C#�h����Ȓ7e�	q��L�Q�ʊ?�����E�#�${0��D�t8����&�L���d���?�����J�o���Ou>Fι���M��Sa)�Mc[в*��TE�sGI��xV8����a��)m���@?sj�ȗ�QV6VP���s�\���H<�_z%]�j��--x�;��2�6#9frI񫭇Xo�_�DУ����c���y����>��Vw`�a���{�Ϩd;$����7��f��1똭 Փ��9�<�T#;���C����Ջ�����i-FI-�Dҟ��H�>���=<���4>�I�د�W���c�Q<H �z��~�Z�%����
�0�R6�aڀd~0�>5��f�����2������d�"��F���i[j�t��)�A�#D��C��Zc�zI�~��E�=�5��c<q+<����s�����g�b��?O)�5)3�Y�r���j��ҳTQjSE�3���� G
��ۥ<l�z�	6~���H8��P� ��a��}�<8U+�(�Z�����~�揀�SR^�k�~��+�Z����n��?��+zO�j�!ܫ��4�E��߮�_��h��#x�'�����k���>�]��r_1���S▰�4jܢ�l�:s�1Y�	�9-k4�����So�T���� +�[u��S6�)
=�ǐ���Ĺ=0`9���P�-'b��7�q+<g+��z� �\��T��+!6Dcā~�%��o�C����N{���~���V��.Z���/��#{���\nqE��_�զzE%,��3���)�������_��r]5�Q�*fRg��U�X=��l�Zt&B2�({Z������#у_XA���Pl"v��{��ޅ1�}��N���I��U��l��
�*��'�1��3�nO'Ǌ��8�����c5��֥�D�鲸8@.�b�#@,@-fBc��Lkh��4Ul#Gf5_���K��ol�^�_�A����8�#Wr{�S�+`؈�]~���Z��R_�P񢮾�*ɕ�_�����{��E�Z�"N"�Ƙ�n�b$>����2�$�+�Cm���Ë�m�jo�Z�Y�п�������[ܙ##³dT[���Ih�QwShаG��bjU/h#��i�G�#S������Q뎰��P~�޺�S�1�l��Ơ[�O�炃.p\��?���9\GB��c��V+���.m�_'���*h9z#0s���4�lMV��L{�U-2_H	@��ߑ�:��,��NA�>�H�|r0�KE��Ů���F���("����Y��190ȭ=��a��O䂛s�ۛ�����č:%��KKFOE�1�ȔT�o�H��n~2��ʞG*v�rJ4����f�7��l�9���Iv/7�݆����^5P����_2�J;`���3rX�q�����"K�v�T
n�Y_�԰Rb���/uXy��Zi�؞��c�l�xI�MWrAT�Ч��<T�#rL�^b��d�v<95�����0����(R�U�v
@����0&��~`o-�i,��G�a�b@����r��eH�á�ho��V�sN'o
�����C�6e�Mb��nc����E2�����M#��q{Vvc��1�����\�\F�R������-Sd��8�=����w�#< 7N�3;�� ��2�S��T������k䑭#xxg���F2ɜK��2����޺ԫB[R>~��<�N�IK4�G�Gᔳ��-��mG�G"=�5P�ד�g��o��#	dQI�n%u�y���C�i����*�@��ۨ,�wb�fn���]`<��\LQ�"m���~�n���.��������%���?P�����1'�ԢWĐE�yү-rk��KF�������צ��1�!�-���T����r�t����䞷�t0��6R�Z���!_�I��k�`>�̭�j01i��=��N�~����z�e����Y�ʎ�AoϢf4U6�ם�����S�f�DҊ�I��$�B��L���l�Mq�W��%�2p$i���9�/��V����u��'o�͝9�I����D<M�u���W�>g.�.� �ն�^����&�,F"0�y볞C��.EZ�)2�d�&��{�{���Iz�fKP�FJW�³��w�P{��?����-&`��iG��y"��>�_��iW�}���%�i4M�
���=5m�)'M�:��B���Q�,�c�\��X\��}"o%��E���&:{�P�&F����k"���'���l]abU�s�!7`�ľO�O�a2IHk�E�	�����W�IE�y��/^���r�t��L��x�-�s�M�'�je(ҩ���6/M?(*�t;}ބo�*Au��S`�)�BUG�N�-ңsa�j2�\�'a�z*wVBiy`/[��>0�o%e�������B��$24��^ R�[-5��/j�~Z�'t���T�wK�g��^�;-��J/n�p�-�Ӌ%:E�P�o~u,Fs+�-A���^��#����j���:'��]׀<�f+�Ph�pu.���.07�^��P�a�m�9l�����/Nw�n$���͝�e�U�]���
�?c�fR�"-�tW�����0��X�1�B���eum��IL.�=4��Ph���L*V'M#)"k�c�s�깼��ђ���;q�/���z��$y��5�����,��7�vx�;&��; �E�UIJ����7z��CZ�����ۣƩ�خ6\
M�*�{"m�}��kR���S�I�'�|��K��̘���(�	�b�f�.+&)��<)�����F;|q�-r�'�x$07dNi!���{^\8�u	��̹؛۵ t�/ܤ�l�[@�V�DJ�=��l�X��LtS C����?+kvD�x�?Ku��Q�h�y�-��q��A�:"�K6��c�M9!�ϣ���nc�>�=b���XOe��a�˥��D4��	O*�HESq��Օ��� ��^W��#^����� ���󃆊���5����q���Z;P1���z�#�DLDG�K�ٙ��]�,��ć_.��㯩7��ۊ��[��\.C3��#�K�)��C=B��D&�&'��$"��\����v�R9;3��Kn\��BBΒ)u�ȹ�C���ޛͨ�؝nf �g���Q�?BI�}X�)̭�nmW�Ҳ;���[�5��rP��%�]h}��n�aN���+�*��+=q�uAI�T��'�,0*�]Hn��,U��*�xbi��$��2�Ort���@��L�~;�ױ�׿2SzZ�Ԗ�ҙ4�C\�&��?�C�?�+!Qǧmq��R�~��&�3�'e�[ц]\{���ֺ��Y3����l#��Sqde�S��i�IG�3�*�uCed{#`Ճ���n%)��Y�n/g)D�gi<[��1����������{S�2�@��Y4��Z1vTm,�Od���r��]Huϲ�����Q�_h:�N�������n9w|\�q�Ƃ�H�d1�I�����j��^	@����Zھ�ڮ���F	�5���h��q�"���䟺�����1�ǈ�wn9]�V�� N�0�/薁O�JL`x��8.5D#u֦l�����P�!���l_�
�n�Až۪�^�/���B�3M�����n1_⇶K���[7]���*8�8OC�m��y�Zw�xt��J{?��0f,N����H���T8�s�}D�"�Y���:��Q~�k��=SM��C8�%^�3 
���OV7X�=�y(pĶ���A��+L8䞘�KL��M��ps��l��/��A�JS����*U7J퀔�f�ۓ��1;��'���!���*�r��4�)�8Z"2�{�AY�08�`r�!Hv?��� ��D��`T��g����҃����~S�BR������+_O^/���qlG��K>�:05d �.�����B8 y�&gD��^��O�W��Pu%s��2��Ş�������
����,f�1��.�f �8�I&As���k�])YTt��o�_xRM���.���ɝ�tp� �D�;��]��.N�Y��	���܋�#�|)�����|7c�c�N ��3��=\=���ϟ�q���Ӝ�'{�WN���=�J��6��ؾ�\S?x�P"��[*;�}��>O�J�cI���d]I�%�8���>>�;�G:���C��D|~�0kh�#�2�Zj��
���p�]d�Y��x���j��"�m�!d����aNw[�hS2��6��Ge^{�	^{�����P󆪧��6���%<!)����*����Z�y
�0��9QZ�8	�L�u-�K˃0k��2�vcDi����	�5�Á�XWrᱸ��y�	��G�ü�dC���p���[!k>,�����(���$��W}[�k�*�>o��˲���Q\=�-�+�"��o���NW��a����� Ն���[�R�<6�u�=��9ؚ��o�,Ժ��ĀPC��3�|�3_��s�[U��3��L���t� ,�_B��r����P�oq8��y�P�h�ժJ���Ϗp6�¡e�C������;|�3�f�����1s��=5��Ѧ����C��Lq�P�����g��{���]ܜ��^���a���g ސ��a��1���F�o��9�Ď�#;���-w�M���]���~]*x�i~�7�f �\�����A��&���#�k��`隄�~�� |��@䋛̼�a|�$QՕ.�𶇬�ɪ̺�#k�I}�U ��V���Q@�v�G�F��gc�E�H��kW�r���H&ʟ�($s�����E�֚m���]��g�*��>�{�	���·o��$�)�����&TD���P[��r������:�m��YƝ
�܅�9��阠�����2��+�H�w���ã���Ea���ѳ�p� {Q�0`��O�l������h��X��gɡ��ӒԚ���) �3�3����귷}X���2�Ϲ�����C?%�K%V�j��hCg�5��X�h�Z=�����6��a��6��vPp'�z\w��>dgh_�	c�>Ã,�}@�����ٕs�����s ���i�_��C���v��(�b`-�Ӥqe�L!�q�[�?��~��")G
C<���1�34����W5�/A)�]��6d�����j�} MyIkHv|���S�䊧������I��-�?ï���Qq���6!4��B֫�+V��/� ��?K�M�?,�]%���	s�����O��U�����������/{���({�P�;��������@�{Jصj8�Cѧ%в��#O7^�d5����W�j�Hb�T�;m���^�7錄<�!蠴-�0C�ab�?Bl̟���>�?��H	T|$'*2�K�0s�Ȍ��MNH�����E�}V&x%h*�"H�@�j��<�0�����([�0���{�����&��\�����'���'Qo-v׵4g��=~�}��Ym��>Ni�	H�Wxu��Zj(��1�/#�6f����=_�]�D*��'/�+Շ�(��,zCys�ѣ�� 0�՚m&���lUE���	��F�Ʋ]W�=����&@�uK���08�lȴ��h���%��HG
��8z�����̀��C3l� �xO�4��'�]����,�wQ%� ���c�������|��b���T�O�)�*��%}\���ܷw�y�3�i!���./@ �L�R�d
�$���.�k�h?�V[�9�?p�S�'�'uIISNg���aeR�틢1b��;�z.k�/��y�o~�h{a�30p�~?la7&S�ѕ�x�!��Uj����y	�@���	$U�C��W���ǿ̨��Z�tB`�"E����Y�����\��m�ma]���U]���M9h���)��u"�������	�e�{���&,S� ���gw�Х�H3�U�����"s`�w��%e�v��0o���>�x�;cM����_��7COڛ����*{J}��f�4D3��G �D`��M	�ܻ�`��!�m��#���־_	/-D�F�Q����N_ϣ���a��e�_�4�/�C��Ү+�?>S!�K�_A�"Ro %�L��`ƅӱ,k2�q�) 3�w��%����l�3C�C�Q��W-]Ls���z��`h�2���)0���ґ������}f*�����.� ����|$�l2�$����la�	�t%��}� �a�oX��N XP��8ڂ@�L*�'�����y�k�Rw���̔��::�� ���"!ÿRH���&���b�`(��(U�֚����g�4�b��"'�4��m�i�t��<�P�e���|Z9�� �Ӷ!֖�	Y�M��~�K"7(|��)�%Hxd_rW���Y��l����(�����6r�9�`��x�K� ����J���s0bw��*Q��˷�0f�e�H��3te���i޸�6�q�=cM}��6蓂��j]oK��(א�R��g���-i����#�Uݞ�?��=��ף�yû����d@��R���Bl��/�ə�*3,_�P��)��[��|�d���Xr�����|�H�V�`��vf�[w�nGy�:����
u6�-�!�{dt�Ң�Z�䄊v��,d�c�L��D�#L����|�m�w��󺧁�WʑM�h�7�\���5�sKN����J��_"4�H�Ȫ���"�R���ÓHY��!�ͻJ���U�>}�=�U������b�������ӝ8`���9ܛ�J"�n�y�� ���0x+$�G�'m&����+��-u���J�/��%D'�̮r�o�`���'���_äu�A�$�N�~Ry��>�W%�-ՙy��Ap0��������}6c�z�������<�تk��X�K1�'#�.7?���w{e�r��2)�l? ��oЬ�J)�, fNT�����Soʁӟ�~�h�)�n#U���d��?�M������%iS!%�]�O!��Cx�)X�!̤a̜-�-ږ&���=�qˠH���}��GOo�
��8�櫺�0��K-h��3��E;}���Cd�R��ND����[��l:ч�M�7�M�y�lb����o�`S̚�0�ۘf�aE���q���	�~\.!��b��:@�ВuE�UA%���t	�{����a�7 U�,��p0U�|�Ѝ� ]�-E/O� [LP�W�������0��~���U��F�%�^��zmHX{m� ��"���Uy��1����@!�2|x:���cn����J���c�1��D;4o\�0�N�^�T	�&�L��J�2�~A��k�sP��F	��W�jd����7���۞��A/�y��.��$��ޗ�i��*�?Ⱇ�n}��}��`dXe�3d�m~���;��KrDH1 ;�I�s�@�y%(��<�A�B+�Q���k�R �%M�A�A �@��z�b/���h>G6��W�@���BGS�-]��a� �UaSK�<CK����K�*̍+Ȩ�}as��f��w@�w�[d��d�P�p�7xa�}��W��,e�q&^K�Y��XN�����EӒ���Ώ�G�����B�.W��c�o�0?�[ѐC�N������S����}�,:O��L-���?�Z�;t��$d<�=1̗���-©��G�A���Lkm�"�>��
⦯�����&>&�C��k��m�p��ڴȁ"�Y����`�,^^d�E��!-W�E��(ȹJ{���a_C����<��^2�:���"� F��uU�ׯ���,#��D� �hj)#+\d��֩�"�UB�9�������9���S�nQ���>m�2n/�S
��f�*N�cҜW���N�f�D��߸�C�<��/O�xi/,殄��,N;?A��jEB������zC�����}tR�o�$��(������?�EI��N���6mܝӼ����!
�e-"a�וPhN�y �J�i������,6�]�y�8�a�N&0V25Fku��<}��N��.~�����t^��-��m2c!�H�է��p�_���+�wl��|�8�A���<���T���nmЀ ���uٸ�=�yM ��ze�r�-o�~u�0_]�:^`"ic���\-��P�lX؞�W�{_8!�eF��̆���o�N�=�?����Q��hP�����]�%����j?�t�B͘7]�"g�?l)@yˬ��ݭÊ��`qh��>�jAp&�(���E�s�4�b�֬��a��j̪!z�Q�/�Iq���~17ct@%q���H��s=�!�ƞ����|��(Ny���{湠Ea�{����V(!��$#��,na3
��D�X�J-BVt���>:3�r_[ 1�z��&�a��F�c ;eP"�H�Y�">�������⏚�p�ܱ|���<��uH:�������B�����8J_����3���ڡ֔4�dA�e+aʪ[�9GE9�WZHu}��9����"�
�{���[����I[�9���:���?a�;)�O��@Ιn��Uz�U���&y�T�<4FV|J�{��H�1~d����A?]ƅ�� g�=hn�S�fI�,����ǀ�e	��=�4yMZ(���^4���D:r	���p}��٩�8�2�R�P7�Zk�Jc�P��?7gS!c���\?
�%*e�k��e�f�p�u<�୸�̕,T��=�������Ū��o=g�<
�OX��d0,M۽$@1��e��}p��`����Jz�F�R���`Z�Xy�-ŶB�J�����ݑ `��^.$ø�)����lľ2�G.�ќ_
��%�h�(97!_�����'��!�YL�T��_�x�È�f����� �Ƭ�tNW8/IWuZx�r�	u`���S�~'� Iw�[*�S��ɾ�{Sn2G���P��z��V�2A��gXŰ�����f���d����
�}�
D)Z�qr��/�|or�zxE��NB4�E�}��k����W+U�B�'�}�R��ȶ����O(��Y�ƙĳ�����%1V��~�J���27E�Wx�r��ϦK�� I^�2$�gKv=��
�R�������0��-Uj���[�wWr0�,��Ak?;\s
d��ħʁ�'\wjiΔ����HǙ�<|`��"�#��%J9ڭ�U�5[]�C�5�	��(�����Ɍ�����H6Pf��!�����I��췼y	��5)�]	#G֧�y�'�m�kh�pm{t]
�� ��Y�#�{���WT ��=r�i��`)y�����`�q\^�h ��й�;����l~T�C**hX�����8�w@������ϛ��OC�NjP�W������K�����{O��Q_��_��Nr�L�jB﷝�c����2��d�.ο��{s�:�vX��=ҙ�&z]z+^���~a�����|��rN�4Z��8��Any\~�w2_���.}��=�y�4%����9a����I��.:��.3f�	���$$�g �rBb�F�r����9ߖ7<�u!`��,'���)�_�x�~�7v-�T�-�C�u_02;�I��A^���ǆ,S�KBg�ɴ��բ_�vT�(E�(> 5�/���[���ן}���������l��d���
�2,�f�X.�`�E�=u��<ؕ�_�:�v��";n���$����xU�bR���9p0���Y����-��2O��@��˟:Ԕ�Ԝ����O�X��N#Ό���L�Z'7��7V���am�;`fcd��3�o~;��d�.���8-����Pe6��P�
]}ćL�x��/������ˊ���?��Á�}h~��P�y`Lp>���\��z�D�NHb�ٚp/�5լ$V[Ǹ��_FC׿����U����)�Z���/�t��3W��lK���m�>��v(�ӹ�^4��}7-sN{P����J��\����C֬�l{<&jR��,�ֵ��&�T���MT>�E8�}%�|Jr�z��!W��k����Q{��<���3�#�}�N��F��T�еwzג�qM�(Y��Æ/�u�N�
M��k��~�>4��Uu�f�W圸��X����w�rqf�d�C��R��O0��>���!��e^}������q�;r�{���J�;3Ĺ���+�ŏ��*	�*�:]PN��?�p������m�q��]����p:űbw)�q���� s�M�ӌL�A��jg&m��{��#�5�ҡ�ױ�S�ɡΎ�����Q�`�����|P�hd�K@��Y���4�0MR�2��C���>��;��
H=�gX��X&_�(t�z@.!�,f���L���+�B9A�8:'$Û��!�&���Ӏ�/
���@G�'F�����@~�54�7Ó%zR�2��2>=�nVs$��$���i3L�E%ڮ�r�a	�m6d�k�_�C&�rI>2</~��Q���ţ���C�