��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M��*����g#φ'����T��6%.^f��8{�^v�wK�T��fAN(.�oC�Yt���Ao�>���� �h�*��9礩[s�Tj˧��Y���oG� �'!�D!�#S��E3@b����}��doB۳��P����F�.r�Z8Bg��������K~�g\�l1�i����r`0���Sw����X՛m�ɒ��Fq{�GT���܉Ub��o#���;��V���
��ħ�u#ĳY���Ei�Տ�#4�P!���	j�c0G�'�(t�g�5g�O�U���H�x�{ؽ%�qT�ˡ���٫^�)�׶�rn�.c����Z] p�ֆ����s��b'��qw�3�Շ�O��)b;6��!dg~��ڗ08	��lQ����������ԯT�L��<�������Y��%�~J�i���vka��s`fȹ�����T����;[�sR�`Y����.EZ�e�!fM�J���W�I���!�u��L����Tq�q���T�d �� �>R����;{��z��L�C�D�){lx���A1�������8KK��t"1�����-�e��<,!:��«&�*6!�9������3R�ζ<���>r�֓|�Clp\%$�_�^�RB�����%���m�.�Yǫ���L�u���e�)��O��,�~��vۡ�0�.C�%O�Ml/m\�I�%��۩��/�J�Tʚ(D>y���苶56�(��wNhX��pl��2��1x)���,�V���o��?�K!P�Д�Oʆ�h��8�!8�gG��*��0���1c�����C������9�}ް�47�SԄbT��u%�cʚ�SGu&,�� 1���m<u�B���0����*��3{l� w���K�وx�'�Rx$��#2�)Z$��E�EPE��sD��;D+�L��>
J����ݓ��xxx��D��49�������kN��Q�����2΀^����sikV-��'���� �tJ$���F��H��ub��<�1v�0sQ��5�L>�C4;6��v�@�Z����j@���8��<�5��ܴN5���# /��{�n"^`"l�j��L�;�� ��fn���
ڈ��y�����̥ 3�οv�D��p.��V2��RV�|3�=��e`2:_?�~3Ǜuӳ�z�#��Ct��4��X0����D.8�x��Q5�҂�r���=n@bQ�x|���喏H6��1`�Ⱥ*"�<F������(ܵ����y�����eo���Kd�je.���*a����Q`�ƅ4aN��r���ȩ����{����v6�[�����a"��E���m;��,9ٸ�i9\����:Ig���}�2��̊b����ȵ��Z�`PN{1^�'1�:�4(ެ+-.�h>ѝ=��w��XnT�ke��,X�J^�oO��m��ǵ	�T�{��Ю�''ws�;艟�c����pR�8ϲ� �xf�ͼ$%��Hy�:�R��P�xXXR��W��`�y�ڪ����qva�v�W��{EDj�������3�RH���-Z8f��m�x�lpD1x���i|ʹ�\u����Z:�~D�+'����Z�o&K��(����8tȌ��ʻo��|7�:�Y^R�����_�D��5E����'�T�����M�p���F��
����w|'�'�"�����W�&C2������mK�%wשl�% ��Έc�X�n�+�z��`
���D,:s�����a�ըd"[�Z뙃��ܝ�������^bL�Y��E�(b�r>�fަ鿕x/v��ۍo�E�z�/��kK�ؿ�/�^��HY�~]�P?���0CJ߈��Dy5?ٵ��q}�m���\��O,#����LG���|�#@3�:�p�
3/ג-5Y��@|�է��*���E����dJu�� V��!}������:Ta�K�˕�Su#ʬ�������
������R_$���&7��p��W�o��|)���%S�>׵���a�TxJ�����|�c-4����ܵ-41�~	R�H�Y:;_�$���@U˭����� h�	��/� C�UF�N�V�
&@r�/r�V��2[��V�ݨ�n�͖��ߓ�u8d��9�2�\v�����|e�CN0�"i�}�aXd��c����^D�[׸�n��-�}p#s� 
����ܤ[�)O�HXƻ5hM�@b�hL�$,@����A8L�E\��>��9��c=��%"s@o�U�]��׮[\/��h���C�Ğ�N,�n�+�P�a�O��
���|�v��ks\����ý,�&Gs��<n���������xFoF����.e���9P�'������L[Ŀ���!*
R���Kup)*9!���%��21�j!]�,%��e/e�o]�iih�eLP��}$;��lݜm���� 0\���n�j��-L��V0_��?����K Pi��$Z:�d�,k�	{�L1ɯ餅?ߦH�.�D���%��/�>���ӛ��g���S:��^��I�;��PyJ�7D�3�w�^�X���gQ�����m}��n4�,�ƴ����v�Ó�EsEћ�hD��x4��̪t,Y�Nos�m�<���������8{4{��L�);/1�o��<:��U�u(%$\�R>�H$�3���͠�%�1/���6T��(��<�)5�D���`�$G�y�.��_w

mM��2��I�oΏ�eqt���}��T�Ün���w�@US�`�ާ0��R����)�f��{���X���V!�9�U*��ܷ��U���R<Z�&����ե��޲0 P��4PJ1�Gs��h������Q��y�� 2�,u��Ҙ�Y��3��cI��Ʉ�����$���Z��7�^���ߛ-xm0�Zؕ�����e+��K�LW{���+��gK����g��]c��4 O�z �)i�pd�K�����t����.Qo�������u�Ui^Fwҁ;�Q�d3b��6;�d�߃�pY_t4U�/hąH�׻��M�M�lL7/�8�j���ی��"�6�0^<�a�FD�3�����P	��ŤD���i��/�*�H)0�:�\MYIٵ��ʰ�ڞٶ ᠽc�COf�Z�f�O��E	��C$�A�'�SF��
����l�÷%�H�q�9:óL5!"/�\%��Pd�c���*�d��A��B�Nb S��I���vO�AV|
'?����{�Gk�O"���Y�pխ�����S�s�k�i���k!lx���CXr�>:��P�?Y%nG=ca�HD�s�ŷ��lU��*�C��N	`1� E�_'4t���0M����g������c���,2"��=�1�X�7D��.Tl�.v\H#��L��E��- g��v@�f`u;FJ�2F�j�iM�{���R�(Vo�;�h�xn�.�J��KW�;�1%c���|Q��	�J�*��m�4��K�����	b����0��|�kD���5e���Y8:<��
�
�zb�F�WQ�%�z�d�7c'��YcH��F��\�4�T�r�fE]�y	{�Z'eD�Y���w�`�=��+�+�G��������2���	>�w�y�ꐞ�^X/�]M��iD_�5{ճ:�M��uK����
��h�v�T�y$Q�;��lXh���F�-�P��X0�<�N@��  �G���UJ�-_�@r����^�������'p@���T�:1!E^��p������ثx�f�����k6P!����T�/��*+$�P�U�n��if�$7Ê�ȓx��rn��?t���P��U��%a�0��}U3D�7�b�*ͧ�H:�̣�dd97q�ӏRT�J�2���y7kzpL��ߝ^_n��1��ʛ5��a��������,�MS���iʔ��f�l��Uxu$�����[�A0��l���Y��4��^Z��dp@�����;�B�jՐ�aQ:��'���\g�4�NxR�v��@��*43vA�N�"�Oi���	h
7�\m��e���'�4^is�߮�$����8F�Բ�.�*�\�ca��38ۿg�ru^eGD�i����Ņx��0�L�٣/�G~�e�i�C
i����HLn�@������f�fX9�fn�`��Ӓt�ZE�H�Z
x�FȨ�ӸҀ�b��یb��^��8���}�4��<`C� ~؞�*I�ӌ$���R�qE��)�p#[�[��q�Rf��/�[	�)��1El�OP�jD�~Q���̔����K�`}N����;�N�����p�$��Q�%'���s��X݊�k<��g��z��I\�����N��)���j��Y";❚_Uw����'0_���y�0�`G\�����>UЇ(P<�;�a;�Hf%�_��yM�8l.N�u�̀|ld�+���C�*�dv+����/M�W�]<�t�Ig����홈|��m*�T�v��>�BMQ�����ޯ�%n��H(�D[�*������ohk��:��\!RV3��Q>����L�zKXe������fJ-j�0y�Jfs0w��C�J=��խi5�K|ZK��ą[\������٢�A'��#����?� /�%}���O�k���\\W+:�Gٽ����lN"��^q��J�℟���E}o]h����QE3ܓ�wD~�;�?졻���1����(�j�RN�~AZq˔��^�ږ�Φ�����uK��N���>d�Z00H�$�L��aU�@��Ts�dl��;nz@�w��R�)]]�!��<�2�e/w�Hx�;we8��m��� &����
^R�P3�Q��e�Û��u�s���#ܖ!�$��ʨ��,��\�S�����Q����h̹�\������y�|�����Z)�}���C�&f�m��D	��
l0��O�ȗ�J�'vs����[���%a�����ci�.�nS;�o��}����zo�Rvq�y��$xsC.�"+��1�7�^E�`im��oCA�10K�9��2�_�|��½���Z?�(��������E.�]|��9��퓪9�1/��*���S�#�$I*[Fx{f�	k}1)��K��轎�ya����J�jc4}�y�s[���v⨀7+���^vʼё�/*B��/Z��@��&�;�Н8u�����Sb������]x���g��i���Q<�4Q���a���kz߃x���1�i�"U�Q��>l/��S�F@����ܗH�������/�-��'K��N@%��C(CG�җ�6� P�Ŏ!扴�V�	�>���|�t	v��S�m~cP�w�% :x���P��!A���'7�(���/{�if6��(��|7*4�s{�w�$y�h!��s��dSiUF!۷� �(2rPœ�:'��P��D��J��~P��A��9��ݭ�M��jԿ#;�S#��]*�����f�BOA11x�[J�4�����C`P(�j��.���ϯ�A���Lؔ�ɟ�4�!�][U��BR��P;$��@�*��m6��)��8G`'����Ap�	� ��c�svF�^���8�FP�V?���z����q\ك�2�d"$��.�;�P�\�
��&��f7��0���i��u���/�������Z�����x��2�c� O:��s�н�^��`�v��v��_���d� u��!q�����!ܶS���[�ݙ3i��V���+�	�&�vQ�a�G���,ш���y����W��F���{?�ZY̨ѷN�~ޜ�tBH/�1s
�1�=��辴���05���,�y���n������@�H�G)�I�v�@Q�Q��4�J�_NH��_�����wϪ�-����{(�䦚�L��D��+I.t*&�����\B���
���	�Ic��_�i�{
"�/AC� �L��<��/�X-�G��"��c���q�?~qT�ya=�׺�x`d�eJ��دՉ��U�(7j��/�1�j�A)����u�� ���P�v�ƥ~7H�/G�6�X�6 h����|>�х��� �'w����]���n8Ð�{
�|�l�<Jh/#�o��7���|q�L����5�GH��td�EYʇ�ҳ�%��O���8t��S��X��U��|�˳0�`�d��<O��#�1��O���@��y��j�az�@BN��9�O��&�B�8�ћ�5����Hu����^�tw[|&����ʋ��mw`ΰ>��9N���z���Y�`&Ȇ
'��Y��Ԗ�n�E
I��"o��n�A�Xt%�FT�@��4%���`X�M��c���X�g2¸cQ�:~2��?+�!���Gm���'��s������,�Ϯ�D����p����8=d����v�s�L����x�'�{�upo����Gy�'�N6��G�F����s�\$�
�#�c(f��!DT='*�eL���M��g��QCU�(����w��������Iz����T�d��dʡ��k�a54�A<�F���'��1O�aEi��α��UI=��6�X�@Yj!��Vr�gD�j7!�H�����Xh)�Ƹ��������A/H�%�l��o�g��1���O�oT����/��҈���>�!�/��5��wx�+��R�G���x�u0a�4x�v�gq��1NZmg�#B�,ݥ���o�w���vr6ؗ=i5�$v���>ԝe<"�~^�:E۔��%��,��b�Dd*�(
��ix䗾��"Q.�!O+�C��l�*f/���"�N�v.�*�����O*�n���-�6=n�,� Z!9MTX-#��&	�=9��:u�:��� ��K����K��'��4�)֝Tp�f����O�_�	Ə/#��G��m �9)i��NP� ��6�\*��/K|P�\,�5:�9�8����
	bz�7�Yd�N�
�2�3Ϗ5o	���f�n��Ǿ�`O���Լ��#��P���Bj��K9(&��1<yza0y_�i{��_3v����A�>��b"(�n墽_G�^���a��c3�^*��d�\f>t�����4uk,�7��Ex�qc�,z����, �8R���]�ҕ��e��'@BP�)G�ƽ�[�}8�����H4��]O�~�ﭦj��S����6���ʠ`X?qVN�k��@�1��8��̇�l��u����F��cfW�����z�Z��@���.1Pc�,E�Ǟ�-@R���l\�(ؚ�v��*���>0�8��E���������Ij���1����41�5#�.MNg��N�N��9l�[\,
@��=�!N��v�9�b��YN���b rv�2-%��48@���6�MrH�<[�,u��lܮ�Y��{�-W�l^j?�`��jjwĲ��yZqf��#�6Sh��Q4;��.�7Z�j��e&��9?	5߹j�7đk,� ��+�������[�5д�*��g9ү�H�0��U��%Y%�a���;�x0G�.�#N��[x�7�
1�uTV�1��9w�/��d}+.����j�[ss��Wi�(n��w����]��2z��[�v:��%�b��~Ƹ�E���;73G|�̾�,�E$w
��6�%]�5"ˉ�E%.��,V��Iex�6����^�U�A�K!ȉ'd�������!~�a��
K�χ�_~�;�0ڬ�&�"f��6�� >��6��Ƣ��F�KR-#�giW]X���-�F�{[�T�wx�,O�k>���W��Ho'U�¾�hHsfVy�����!4B��ed"[pc���RC���ed'�'���8����O�M��F���� ��d��bT8��i�"G4{FL�y$���U�ͪ��Y}Z���*��۽E�	���/o����"Tԁ�PrF���[ 0��} Hh �2�y3��K^ ��b+H3�9%Fy�]-`ΝNNz���(�����d����ch%�;[WH���W�`r�v�T̻̾�{g�	��sߡ�"U"�Nb��mU6�Mj猆�1�o~��v|��9��T�WnA�L~B�a$��aI[1t�r���R�K���4�x4vo�*�ન�Ivs��JM��9F�a�����A@�#+|��حS3����1�}\��u^�^b^η_�g�}Ϻ����| 0~ܚzS�!jVA�[ӊ~��<k�无�k�I o߯e�	�����I4��ߟ`�õ�< ��L�ڭ@2DҘo�us�*ʼ�D�(X�Oπ7�rVK`��Ex�+�@��W��������A�m]�L~1�F����r�����QR;�$Rѝ�o�y�j�OM��D����](�T,�M��=����^���5r��K�����>��k1`����/���r��FZ�k���8���� ��M�<�/~2��py16rD�߃����ǩT�G�^�茴x�������!"�1�;�� ��W��� �?��L���:����r	A;R��~,�SH����ސؓ��'t�I8�9�}^�ڌ3L�\*u�Y���Ĕ�0;�cC��3�z|ζ��$8���+B������n�Od�k ��V
K���d^��~�mɋ	�/�`~��\��@Qƃ[\w����z�wt0�S� 1L�;�Y6���t؏ԇ�Ct�l���]s݊fq7o��p;h YhuB=�Z�כ>`�&�40{�&����U��3j�R����tfF�����&�7��r߅��������DT$�l�C��1�_nQ�#�W��d�Ϯ~2�L�"%6؋�v( dJ|Kv���10|j16�A�b��J<�j�F�B�GX�� O�˚�FF�g�r�-�����.�t��u�#����C]6O9񐁇A�+�vF�h��n �e�.lW��(FfvR��$���ň���,����C��+ݎ���ZC��G��ܥ�l�/��"��)a�xA�z�L:d�f��������_�F��>�2�\�KG�q�P�C��<���U_���)wB-zf���|Z�O�P��Kp���X���R:�tao�������� Rt��ͬ�z�u��W�f��*�f�⸓4)����smKϢ�2��6�~�.�:�?v�_��:�m�S��X�tA{2DdQ��>����LX�ߓ�,Z�3��� ������oHJQ������|ׁ��O�G6��ʀ���RؖNиx��l���g�k����٘El"���
1����de���*2dR�d]�+��A�04�JUW�1i0����Ǘ��~O����(8�����Ӛ�	2�j4΍o�+;mj��ĶT��{�������Y����֛��f\��V���
�$�%�A�9�@Z:3XM9%^�.4MA�^t�ߴ����+O��-I��N �_=^��;4.��언�[h�@w�1k%��4.d8.	�j��&����tםg&* N��>�`K�T�*O�5�i��df���y+�k=��@\?��$g^|b��V�8��^��o\۠�#ȏ�$Z�F����l��S�����-�ܳ&&�Ր����	�P�׆IEķ�opqQ�?/���3n����,�+T�6���� GA?y��eȭ-&�vه��p/��ި ��ʅ�"��>��2ª@���X`r*��Յ�(��,!A��N���Ix%�����{��:*Ű]~��p97�|�Iy���+r~���ݡ��䘁1��%t|k�9p��mٙ��_�4�L/�����VK�=���"��=h�?M彅�Z���Y��vOԆ.�֖[5@��n(#ţ�����O9�LO�����I�@{��r
.<�G'g� 2
�D�x�6v��
��6��-��˺��L�W�Q�-_��&DP{j�;�w���9)��×��Y����k4���+_D.����g����4�.��1��ܗ�*�mk/�tZ��-&�<�#����&@ߝ�79=ʻo����k	`�0̩(�̆SsS�&��K��6��bB��%�?�4��\�,:��Y��)� �	Ŋy*vu�t[�9J�ug�_"��\S|.;�Ω�%��?�q��@;��Atx�qr$�97á�@ԱxH`� �
ɷVo��qD4�/�C�,ś@�Ĳm��C���ʳ�d���K'�2֐ OS�Q�I��5 ��}���ǇXS�|��1�����$�ҿ�Eu�2R�;��CyKc58�#�,���gO.MC�1���>�����KdH��?��]q�864x'R��h�Nn�Km[2���숡(��2�n�Fg��eCz2��l$�S@��B�Sր��q�T��������U�^I��<�N�B�x�h�)@3�p��\��m�:V�=��%A��+)ܮI_H%6L�y����e���|���?�Fl�k.�'�yw::Zi�����4�?�/����ڼc��^}Ovm��Y�v��W_v@��8�m���P"�m��������W� ws��t���ta�NϟG�W�����v˷P��yHfi+�;F���z�~� s���ю�T_3��;3�璺 �|ʡ	��.I�[@���m�����`�e���%l�R�፶Y'�
4���"OmqP�s�T܌]���K�C�r�������	���S.�)� W(������	�d�	.(���tϘP�l����zS2�{K�0���v��r���j)/��q�o���B�FM�η�`ѡQ�DJ4OMuo�ͳ���.c���2�����$�����?u&�W�����v&{��ͺ���g�א��(���ix1������z�/D��g&�����i;�hۺ��/�;§�Ĩ:�x�=������h��u��2��G�I;�cU�p�B�%��&�z�)��tU�P����Ч�I�%�����F�Ă�,-��=q��4��/�X��9�> ���'Pw�$�{��De�C�ra;l[f�W�E�L��fI��\Q�y�lb6��\j��G7�;鱒�s`Q�m��@�I��e��]�ȿ�A����
�J	��]˩R���	P�+&UgT���	����e�����.�9�Y�7]O�*�|�Y~ן��crdl`%��d[A�:C��૒
VFS�$�<x�ǀ^N���'��5�*�gzlX��T���T�cB&��4�j��Y�U��3��^�}^�l��D�iL!��o��V�(��x�/��K�?�m�,����/�T�Z@E�d���O]èI>y�%��x{�T�F��E|�fٿ�`g��b!U��GUL����M�Pkť�)ϧ�D��p��
��B��#�	�vP��\��^l\�e��6vv��tl	�H����!q��]�_� K�� ;nG�!0�p���ҵ*L\�ak	�#\<�W���3*�]�~���⟯��:DRC�Ƒ�V���w���U���a�\��MQ<�>.R������DhR@0Q!�2�6��n>��!]�f�#"�[�F�B-�@�y��d��
�V�\s���ةO���]z�w@�&�N&���|�k��s�%�wj��&���Վvj�g����˫ȫꔯ8��s�c3��<'r��ó�8��A�䴂���4<�Yؼ`��m!6�6�7dI����6�0?p$��l�A��__#�Jx줩�w��P�?z{2��̯L~��{��s����3�WFl�F�B�nh#J�@QZ-M(Iu���^Ⱦ~�#��E�&�K�#,
�n�m��mk��������p�.� =M�N��AGz������f���d�:sd��ՉJ���g�SDI���\����VR/T�����)Z��ujݗ��c�if�{@-9{Q�p����\��V�������3UH�^�8�~ê�-�gS�$�̈.-߈�D���3:C+E�o�vVe�sR���1Q��$����y�Ä����,RF�I5�3^d����V*���ԯ����	Q'�x[>o?�l�w��a\�1et	!3A��(<_�*:�"��7U�x:�~s�*OG�s?Fg��09��D;��2J�k���/�D��� 6Tߙ6N:N��v��3�0ؕk�s�y����!�E�����:i���@��L�����(��
):�3�(tu��Q��e��~�H}�ENÌ' �X'�y�'-�.��W���Z�%���%�e��A�������L��aƹB��+��V�%O��#?JW�Pae�@���`M5)��Ø��c�;�����*2^��q���g�b�{;�ɐ�ڹ�a)=��ي.��O��I�]�c����w�%�/:9sp�B>O��4�ҟ���y6��IY|59y{ˤ �S=�	ŵ��z)�B�\�,"Yt��.���$��$�C��O���~��\Å�?B�m%&!}d;I'��M�y�5<q��(M=.^Mͷ:��]���l[���
�:�\m�So��*�fYn�����T��3�v@gڻ�=��KItH}��{t�����`�ˬ�%��Aa3��������~��X�*�f���!aӞ���/�Et���=��/>�L��'��b�
ts���t��
 �����1��'�L�^�n��S�<R2��FX	.!A�;.��z01'�9j&���]��!�: 86�҆�8��P�m]�t�H,�(�E�`�y������x���q��KoO1���qʆ3�!Y���/5=�f�ŗ�gd�3b�P�F)�\Kղ&%h_��$���)2[>�!����i�>�7ղ'12��ݖs�"��oR��ăS��&#�>MYdr�X|rB��X3N%̷�q�w�u�MH����箲�1���W�I����bx�3Bn۝0���]e��K�M,�kGN��/���S/r*��*-����0ʣt�=��N13мK;�kά��h�Nš�!:�
�ό	����npH6�,�Kq5{���6\6b�D���s��C�钔J~-y��Gg0�n���Ma��"���M|Ix�G,5a|�+�V��WHu��"C%p;h>FsN�x���L���@������w��H�S�8iuwi '�m�K��F�v�n�c�l��ݒ��9�|"�ޢJ3�dV�X���t���;�>R������5�"6)6Tf��ۉ0"�r��Oź4������� �F`m�(��d3BH�;/�B����<n����oqT`��o9t��Y&��d����� �'��+����.����S�	M��=d�g2�U�q���{]���i�1���L2�̣1�;MJFnz�E�p.�s0�]�@k��zk����!�l�a���(
xi��@�.����{ZC�H���QA�==�,)�7}n[q�$�Ɠ�ڐE�D��+�5���F&��Z��n�L���9�`Sd+?NF�'m˳����ʛI�����{*�mQ�D�0)HzJ4��jqOÅ�T}X��~{ϊ�fh���0�-�WV@���@�ZL|!��Io#0��sV�n31?���F�0	r�;{}T>>
���=K��%���ѝAdh�}�5���#�b�T���(��=��	�Hu�}(Jn�`��s��w�bL�����/�h�q1�	t��}�z,�vxD�ʃ�з��p/Q#��f��_�o�<�&��`;7u���H]��,������k"�Upe���Y�Mdɋ����G���eߦ◂d�!�aur���?>D�^����	su��YB��չ�V5�Y=hX�pѾϹ���-�ER�9ݽ*�y�5K�y�>O�p�!P�s}rm������ԧ������E� p�HF�3`�>��4��;��yI�BwA{�V�$��ڢ|�yy�?(�	J�}@X����X5k�{��D�c<��RT��s���Mą�}���I���3[v�)j�:L��fj~�IsJ:0hsg����G��+?��{�#�p�y)p~�"	D@��C[fs�}���b����ȩ�Ȩ���#L �Y�
����r���[�Д~��Sy��K��`R@������Ư[�^�m��L�Co�g��q�E����7��v�����C��Q�uE��D��.���mu��ڇ�AM�5�򦂓�v;�4q�M�'���r��Ծ��ψW����#�hg�����%���\��C�U����	ڒM���.��/�_��߶U�\�+�z�l��+A��Չx�����qX����\p?Wb���TwU�X�q��d�'§�f5F���
��?����)}�H"�~ɴ�#�q�d dw�#3�$+~�d����+ȴ�*���ıտ��K�P��

�`�ry]~/1�Kq 1�S��lM\E�I��D�23�߳��1�.P��k����]���$�� �S��Z�����[��!��K�VRgHwS��34�Z��&�� 2��#�0��MrS�}���R�1~t7�J2�S#0Iʲ{���,�^�f�y���[9�8i�Y)m�#F8<Z�y��l��5������!���q�K�6%�G��M�H�xr���XV���������|�ZD��i$��y7�<�C>'��$��	hM�s�-�{Z���Wd�E�M���:+���-�q�;���Vt{��x{�`:�d��Hb�}���v^$�Ž�_[gb�2Ͷǈ����Hj�WeX˨��`8�������1�-l�E�U��l��H�p�wY�*WySAb����8x�hmٟ}��b9����$�
��N���b��#�1�C�&�h5C�*��n"-��ߴ�`���x d׫�^�%w+��i
�V�̳o�t���q�)B��qiݕ,��y���~/���pنSF~�#��|`U��x�oZdٖ:|_�X��qT��E������b<���YQ\��vy^�U��tYr3�IQ�4�p�&�6��ApLa�M��%���d5ar���?~�-͍~��S��''4�I�ğm�����eho�}�@��"r��7��G��YTx��a#�I�"ܨ쓓��>�v��bB���4f�c��8�'N�ʢ��	)(�fH�o�8�E�n�Ka¢��kQ�H_��B�53O¬�j��($���p�Q�����ڵ	��:D���t���|�ʇ�v���sO��+˚�Z=�B���g��~}��r��~a��2�wZ��XM���lF\=?��=tlM�
�3kq]�-��
�����.hZ�A��)U�՞�с:7H9��u�j G�h{�\��OnPv�}��@�t��Xr��
�n"��X�[O�];̢�&c��ܩ#��F2�aY� Z%[�8�\Ec.�����N��R�k�����-t����z( ��'��M�� k�'�#�����6�j�f��1�O��Od�ol�Maݪp΄c�ː��P4)"���^�/:�sP����1~���S���R
J�j��\q�`mfd��Z	9P 	�E���S�b��lZO��Ǖ1���0i#�g3}K~vd��?{�x�8E�1�9�3�/����`O�����H�L�c�1�"�Z��J��~�I��.}-S*�jf��,;�}T)2!V����zJ���a��m%��	�K�pKۺ�%As�\����Z��:|���]^ε̝f@LCS�i,`?��W�q�ho���UsJx�?�c#o��
r�Rmt��a�?2�w�*T���__m���qb�]G?�u�/��'b��[������O��H7u�&��P��2/��G�T�"H@����8��N�`�Z��w���X�^L��{h�GJg�i=4ͬ�*O�^c�qz�u�4�)��N�F?mY,��b�}����7p���d�Z�n,6L��o�Bk���d���=�"hϧ[��ي�?xB��\Ǩ�o8�� �,�Gl6�^	�J�)�ܜd_�G�Z�"�ܘmJ��k�G^Z�j.�[&zS�ƽ
�����0��+7 D�n�szG������'���r�2�?�:䒟b�L����o�|��c��q�L
��7�ʁ��$3y���;�nr�ӵ����6Ǉ�D�,Xs����c�|����U�l�e	1���k������z0�D�F�S�	��r�vN�1�b(]lM�{楴�	��	8�1$3X���ԉv�z�!�(��'�?����4
�=������0BV��{��7�x�j�ȀF��Y\1���g('�Ek��ˮ���� �����Z��P�N"��������#���랗�j7��w6raS@�7ٱZ�^=��a1��0
��,g�]�$��.`�ˡ��]/���p�6B�yr*�Vg[��J'��O���O�JⒶ'��y,`���MH��(-�����~H��i��U�xL��֔e�w�W
I�[�������L��%}�9]Y���6�2~L��1��:�)�ឞ���s���R��^�I`A�Kxe�{3Gp�ў_�bC���X�8���A�r2��R�a��%�Ì63���Z�4�����������k{�8�B�mŚ�6YQ�jB۽_L/ui���r����n?
(t�~�e�)C�nsO���&X����PR���卮^]:?��]h������.T
Nц�c�ע����O.r����/S��$>��7��$S&�����,��Y��c��'��>t�{}�^,���JSA5C]��������"i�r��-����'OB����Q���Q@�*�}O��<�x����{��ԝN�{P{^�7��<'Zj9H�8���_�i�1v��ykFr�LL��4��D�Xry�{)A�3�s
��y�	ZO��?ލkBY�)�&Yo;��'	3���
\���|�"��<>��15�
�n�Jc/eOä��}�F�cLs�y�nuD��L`�O�3|��c�	լr؄�.|��A��F.�J����W�.�e�f\z�`��aG�|7��eT"ȗV��,��Y9&����D���ʓQ��ub�!e!�Ѥ�E0F���������8�عT0~�#Y?�"[���%E�P�cG(g�h�#U��")R`Wkw-Qm�}����9|��qC�xl�_��y��߅�d��
����1�.\�f ��o�p�Ŷ��2�b�ԟb�l�,��sF5�ai�|<|�����k�o�g��u�e�Q���2B�8�O���ܒ�_y�8Az �B�;%^�A]�����l�W�9��Og�eM�۸���o2�}�8�oB����hڽ��9����'^S�Q��~y^pW�:�>�IV�7գ�Sh��R�o�E��Mwm���:��s�L�A��l��P����F��f���Lv���E��V9~Ȧ�ᙩV8���y�<���3�ئ��p�L�����e�����`����]a�O��]�_��ڿ��
���\�gvO�����@��IzI�ːY��2ast*�h)In�z��X�.6V�zD�� jy͎�H����ޔ�L TF�� ���%��-Ya�\?���Xz�\�(W��~����%��/}ȊM< ����B6L��rv���͹�j��Jjl��H�f��m�ʌ�<�X�b<}�`I��8A�йO(]*r�Yl���/�U1��I�$C��4~0S��B�Yvc�c�ZI=��ZY�ؽ�:�J��4@\_Q�mxɋ��C�2��j�|�}�g ���C�mc�y��C�@�M�E�ecqޅ�o��ӴB--ЈQ��b��N/�zy�5���6��A��G�!�R|]k[Q�����0��a'
��i�vo�s��A��� �3u�}ЍW��a���t`��ګ�UC������BI��^�÷+�nc�eS~8N�ɠw�12DTK�X/(���*��vtx��m���Mm]Ji�u���=rԟr/S��mTU��ӏ��#V�Α���l���>�8�;�??_'�OM�[�tH��c�j֚χ���0M�}�E��X�e�S_���u�"�}����(L����`�Uwo ϗ�|�
�dD{�E�3�y\�WVc�4�!woDq /	��͙��Yuu�)�������e�G�&�����qq)�5���EV��ǘ���ԋ�?�6����2`�Rj��R0�B>�_<n����`��c��)�#�qfa:��Vp��)$�8�6O�/MfS-S I�3�[��78c۰�G
��7�Z��n�8:2HLyx�<����O��䘣W"���$��$b�۔�DF9���rz������;1�3~�̣���?�ƱS�Hsf�[te�r/��w���V�P%�$�j�9�T��gqm�y��M��D�P�$ ��Y2����+�X}�
׋4��,�ד0�h���1O�LA�x�_�u����\����-'gGNn"�4�Cه�Z�ά�KU��0�:5,Y��ϰS���-e���r2��4O$M�v�A�W��\�@�1۰ʬ�[Ƽ���_�4���z6��A�\� \+x�܅��4���u[IG���d��63űJ"�؍����ʓ�*��j9��w��i}J}N��vd��aI1��ao�������
�Y�����C=b�`��*�n,]�L�%�@�M߮b�{f��検t��D����'!g��n�����"�죜_��:4<�d�3�U8p���#6��y��G��_m�y(Х��$]�F���5t
`�y���B?�2U��p�jb9��?��on������7�6���5驼D�O�n��B1�yۑ���6c��$�M�Q�D��$���� V��k"}�&s��?L!�U�I��3n�V���r�,���X2E� ��@�c�s� qm�
1��!��$M��u��N�����k��S�j~E�Z��P��;������ x���c}(����W�&��L�6�5��݅ǭ0�����x�����|�je���՟�2H��>�E }��[ �Ɋ���}��������o�©D��/����NV�g���� ��,�nd�t�0�nJ�J�*�?��I�LJ1�Y�$x��H��BvW�k�}6���^�&Û��0��L�6�Ov
u����P�eßQ��]�U�a��=:'=��2}�k	fМ�_D<��^+��G�N�ձzEa��~�-W�y`,���������u$uW[atx
ӷ+[�c����W� �a0�{]��5�a{��<�u�y}�9���2:�@ s57CN�(&���Uڇ���e���$:f3�f�R�!O���=B�gN��t�`��S��"/\㙟��h9���Ou4+۞m�+������@�<�u�a�}7=y��2�$�(X?ݏ,X3��'U�`��Q�W�_$��42�K�M���O�"}��*D�� Q�l�K�k��7�5����o6��02���6Ё}y����T�3�i�������*���"̎B5����ى8w4���3A/oլ�_G$�F���oB��4;&ė��lz��(�vl��J�P�#;�v�b��̯@��E�(��e��ë�g��\�\9����N�g�E��tf�m
,e_��ő��y��� �44N��n瑏]���5�;xX�}�*P�J��y9!��#��x|�ՎV,��g�F��684ݴ�8I2٭��n�y���A�:=4_*(�s�CvK���������Q�6��mr�I�D��c�����M)����V]C!|$�i|H�$1�����U_���2�������
�l�v�2T,��1ti�ߡM*(�خ�����B93��O�[F�6[]Y�1{Y���N<��u�Q�t�0wA~	Րi|}���SJ�w�K��[D:����7��22�GO��27r'#�_��O���/e�հ�ODՐZ���lg1���gs���q�����Oɩ`籟��.鲑�tL��p�QD�W���Қ�C@���Z��;�~O�Yn�J�z>�~pqH6:����Y�qq3&�7�qz�B�1�������Xu8h�0I�Y�� CWC�&���A�K��jr�	�2��o*		1��$���7�|��[L��7����l�l�j0�l��.�b3� ��.K���5}�Y)>l���n {�SA���_P*�v�[�Wj�	�����x3}��e�����V�ܧ�a��*X��d�W����d?�����p+�.�����R��؛*ePlF�Q�&��N�P�
|,FX�ɻ{��81�<�sAb��4�{K���i��_�<� ��n�� aO
�Ðs���S�|�ʌ�c�AB8�@��Sf�fIς*����|3:�e�{��T*�O;�Enr2&���=���|������F���f� 2щ�)~�9q�/n�:%�t��it�p�#�{�#| ,6���Z�#��n��C��0���ΐ��o���b+���J�9���%�;ڍ@``�5��'ׄƓE*��@�����t�����ܦS���������R�����=5��b�1����D�yb��>)=�����C��Ѓ�ZT%��&}ط��: �t7!KۋC}���	&*E=p24gs]9/v83 ��h̉<���b�� ##��G��U��0r���,�sӯ@�g����dEZ�e�5&!��{I��	y ��N��o?��u�0��]Cx�[���FFH7Ж,qr�RI*(Xa]w��N��.��n������%]T1 dp��u-��M���R��|26����_T�.�!�0��*/�>�@�lx`��g�S1���v�so�<'������5j�xö�YJfT������)�TW��tUS�����5tDCtC�.�h�Ԝ�o�z25������-a?_��C����Ň����Rݸc�&/A���M����Z���l�aO �ȧ@qZ�f��x{�g/�.���,��F��V�)�:���.n�rW�[�:�M��ӎM?'2�Rw����#��RSŕx'#��[(�h�k��Ꮪ��� ���Qx�T	[�*�nȨ�ƻq�'�۔;��?�[U��+?>����w5�Raj�@`$ʖA[N�P�1�(������ k$րw}�_�1OYɘC�o$�p4�o��U�Ek���HV *%�����x4�t��WP<�g��g��#�s� J
�WR�V��-�Dy/ʹ}M!Ù�T�K�r���d���ͺ�t{���򡬅��o�Uε�h��D0<���oA̖%�ME�-B������@��,c��=�>^��.P���5�lۧ3�U�G9�F�K��t�@N�U1�q���
��c {����h��!��(_�I{�=��?�qf�mg����c��1?�?U8LJ�q�q�#PE��T��uLr|���Dn�r�ۺ�Qp$iF�}�N%m��.��8Jְ�+�e[�����^�?���������DF���5�@۬�F�W%S�K�&3�nT�D��ʼ�_����d���/�ؒO��T7��Q�P|T��w�"�����di��yV$����mV^�s5��d{:}ӛ	\��Bً��M�nceI ��z������"��0|fk)�p����W�{S�!y肢���
�4�U��g��v�����3'�)�Hu��$��2����9Ȣwm,��'���� 瑪�Y{�go��0��U���ɑ���N�C�4��f�z������
[PTٲ%��W>��(���{�~��3A0�+f�Z>�OF�hr@�N��_�ozVs�#T[�6���Y�����{~��k\��G�MT�������y?@��gإ���7H�X����P�,K`�$'��9�E�-�� /���%�P~ކ+jzZ{p�[55��M`sU:za�Ư�Uwn�[���LY�U/� ����1bhBP8��_s&
�NQ\��ӢϠhiǈV�k�?���?*�#�:�h ̈92F�����'9� y5=,���'5n'%q	�� 6�c'�(�r�C|�w��m;�9�;���ĺ\3�{5s�n	.�l�y�����sx"� ҖQO�0:&���#=^�T�ᢑk��g�W�a�����˽�BJ�ġ6���/ș �,#־#T���s4Q�4�\c��4�Q$�H�Л�0i�	B8��70�,��{�72����I:J��D��A��_E�a���t*�fʊ�:S��)Hj�2��pD��8[��\��~�n���L
�+��F %'J��DP�@q�9���`[Q?��-���F�LX���'�Z�#��C�{���L<�)F�KL���c^);�ڐnH�Ib���e�?&�a����MBn'
vE�\Y�B �;���� )lh����6��m�8WE-�hsv�]%�t0I0�qŠ�ҧ�o�E�-U�����7
��|�p��c#�}YBu��^�1�[�E�FV������F����ְ�Qn��]�	Ǥ�0�$�lG/�%��9�CiI��RS��z��?���Z�y"E剣B��ڠ���}1��ߎM��	�Jb$�W+w_'�kf����$v���b�!R�UM�yf*~�O_��w#�u��R�zT�t�+�:Z�8���I�	��]�_�}~}��NX�=�`=���S'r_$U��D�J�'ʰ�i�k]�
�l�X7�m0U
	󂻅���oU�����j�M��E�e"��P[^ձāM��ઈL�D�*���� HA}5?���!�g5����ҝ.�͏���L���b�SJ�2����xxō��W�+=P�G�tיNQ�{?� �'n����x��:?C�8)Fv���]��|�9�M�Z�j�c�/T������H�ȆŰ[�xW[j��B��MD���"��F���T��L�'�v���X�fT�l�Om;|��dh5?B�xD��)���b�}=�Yb�����b._��{u�Ƒ�ㅛ�o�*��W_�R��7��`Ϝ��b��u�x��+Nx#׽I(3>}�61��1v׺��ё�ǌ��S�|3Er�oϹ���$��1�fq��Ƽ�;Ng���N���K���MKn�f�9_$����9��$j@$�q뇶�Z�L�[��,����R��7ֿ��Il"��ގ�t�U)�8!��u�*��'6
X�m���׏� �<��G��s�^Ѡe,�>V��i'�M&�	:�����]Oq���M7���㪗t����Q������srHB2#0���S5:/��;�=�Nl����c(����	�P�=)�ɉ�������eL�OFȍX���ۭx����g!qt���1����I�e4��.RWU/А��f�
`�%��,T�a��l~A���H77wy���6S�Ϩ��whџ,�5�e��F�Q���� �/�T
��>���c�PV�4��K�OK~�ՠ����V�|v.���rZa�* �5H�:����
&�f,)�#ndv`&�&�Q�55{\C���1���6)����G���G�=0���tx��_�\F��r�4+3�q{N~��A�|L5�~�ǐ �{�Pc�$v��𬐫>�D!�4.rI����;�p� E^Hs�_V��r[�8�QV�'TK�9zC��_�k�PD��n���RUX�E��C�y��B�"����u�$�4�(�$lߺ�H���Z.���'~�񀭯���ܶc�D�4���%����ʭ���=?�E�n��߲ܨ��]����M,���Jv@;g"-�ڝ
�PQb��_�� �������-��6�<.��IB�2�a� �^�W�X�=�����̑z�Lԉ�ς�;�U>���� �8wѳ:����Q0ϔV����;��l����7M���l�͇���QY�@����I�%����&S,�Yfw���V�գ�>8�vc]��M��UA�&�O�3�G �wr^7v
 ���G��O�PG�~��� �@ߕX��D���?Q�00Y�Y��()���P�Ϗa�"3��e�w��t`��S���/:�VÔF�����/�!�]��7��#@�"�����f �?��.U���/:��v��Ԁ/��\h۪
�� 8I_�����@�,�E�N\^��U�tUAy�8���\n�U��g�uػ4-�S�J�+ॳ��N���xFn�e�Rƪ�n4;d4{��AN���G�o���)�aa,�s{w�Z��Z�
oQ���[�2p�l`�:t�0���	�������j.����~��v�����)���l/���j�ɭ�� �-�r�}@�\��3�F��¹�?
>�h`�)&�tZ0׫�X�ßq��m}�G0���Y�q
�^Ș���?�֩�˞`�ܙ+�>㷘��)X����,ř9&�(u���LAá>�9j����d��MyI�yu���cB��g�������v����\d)�&{w��]=h�ic���O�ڴ?���F�~t<>4fgb[���_~̩W�A���K1S�R�%�.�}��rvay���p�5������8Sۧ����\w���֘�}�Gܾ��
�ȳ*���[���vjcd~��I�z�}�N�.~��<��y�o�.l8B��II�s�$Lo��׳U�o���ԃoB�+3�bn�]W���&15'?�!A��l��Ǜ�U���T�a�y��{�dCSO��
Q��tn���Z��e����7�j+n:�I��e���[~�{���P���~��~/�j?M�|>�@�T��=T���t
h%49�����C4˼���G��<�-TV��R� n��D���4�ܯ��Z�{�N��/�l�����7z�fdv�r>G[�}����\�V�����lU�.N4�j.Sy�Q�ޕ1*�U�lF�|D�trƇ1���G��T�S9�������-qϬ��I9R$�����9]ķ�V���FWR��RR����W=��<�_kg��ˆ�v2���@T�>�]�w� A����E��(���>Z?=�C��s8�[F0�I��%،��{�����<�q�?/��=0	ǟS^h��ٍT 9�;�E�$W�_�E26t�m~�����j�V_����^�/o���m��=�ᦨ@�
f�>���U6.���f��"�ӭ�{yh#�6c��]Qڑ�'�����/f 9�u%�����65A���t��v��yk8���X�[���Msс X%5<�O:��dJ�y��Ȥq�D�O�}�	5FC�����I�$���K�S����N=Z��[*ya�<Pٍ���jڧю��UI7Y%^�������$h�=@$�i^�
)���U������7�����f���݋S��ȃʢ v�tN:�`7�Ns��S��*����) C�`��x�V�3��^Y8r6����A��M�����,O�l��9�j��S�/1�.�����A��qd�9F���j>G�az=�,��ɕ�ݕ��+O^|�v����=���{Q�`��Rx�e�Qz�t.+fs�x�ʨ��R�\щ��+�
��k�$�;��uS��e�m�:��4(�Z�5�36N�Wh��(��~����2�L�{�E!�Ђ�*V�R��VW�h �����¥��OZ�_Q��O�H�D)5�ܱ��4v�J����HC��u{%$�!5�G���{�\��P��\0������Nd��A�k#�H���0���\.�6�YC�����r��Fh@�>V�=��z��=�5 
#����ױ�ش��D�r���_�mR��t�����!g�����KR��F7� 1♅3�s�9��F�EVJ�CP3���o	�ml;\�el�C��u-j����|=��|��`j��[���!�wA'���Xd�I�H�E�5�P����ĐX�߾�ð������B�� ry���ǉ0[t��d�ņ磣ܣ+aaE!'��� (�Zz��Z���}����*q�0:���վ�"lly�P���7��ϟ���Ԙ��|	���Ⱦ�H� ���x|�'N�H9�ɉ��S�f!!�n�������h$˶zEb�zC;�%��m92����s��W�p�A��s�N8�n��Ȩ���x�c� ����v��JNɥ�FBy'飪\�5�	,4,^�
�|�`��+���Cu�Ɔف�f�C�L����f"�#X+�d��:Z�~����ק\}/��_!Q�g�4w�9+{���7���}�X�WfO��>-�!B_�����������%zz3�ؗ�������$
j��B��C�-d���u�QZ4��ʬ�b�"��>:���/Dd�h��+'��'�)=��0Sy�H��=��T���4�55�@�e�r�)���[M��?^�vF�u�C��1��&�-
���)��RX!;R�=Gi���N #HEwN���H-��N�{��9�����QV.gH��bj��U^Ke-�`�k5��<r�.9��x��#�}#�KG�Sݡw��N�ٹ�D�׶��Y����/�bTޣh��o{LT�\aO�_4[rAP�f�x-�-Ď�,>��W	��&p�2�IR�jҍ��1��5�'M�9�ϒyr�R��v��K�m8�b�C�j�M�FC�1�_̣O�O�v�c��@ۨ��q�?o�T�c��6//oB�M�t0��S�8��q���~�A����#-��g�1�Ho�+3s�H��%d�ֱm�4O��p��3
����X돗��@4�՞h:�c7��3#��2����c#ġ��{?�v��K���rk����ّ��n���gq4��L٤���;a��֞$�/Hz��d ;���B�U����@���$�u��"]G�m�ߖ�Hw{[�?���,"O��[i����xp^���O�F�ޜ ׍=(���gu�
���	�V�&�QH��3��NT���h���]���g}W��j%�޶ް�"��3����\��8�����e��E1��<�1�A'���6�����vɦ^��#Nx�f�;(r�#���ꥉ�6�-uP�ZK�7.ĽJ�E�1]���0N�Ҷȷ/�Ɲ�������$�Q�i뵣53+;ՙTJ�4$�U��'SK?�,O��B�Ӆ�&�nwUnGDXX��m#ܾ�|��Jlb �](ʃc���('�	,�xl3߼�$��P���:.y�d* �����~�^g���QM�oIUb&T�~�3��tV,�| ,�Ha]�ż8��P(�o�~G)9���W;�>�7Wr�<��zG��r���M��S����D0��!�����C�x욗4�Ѝ�d:���!!�G�^�$��L�Tᶮ-�Q��L=�&ҫ�����	�Y|����������c��&Z��2Oj��*	�ez
ڦj�4&�N4em�M�"��
�ۜ�/�nn��Id����q��{e,�6%O���#��t��r�n	�]�ߍ�)�A�������i�2Ai�?�Z�O:����X�ߓKL�d���m��.\0Q]يߕՑ�{�:�`	8|�	�/��|�%�h�����mI�80g�Y��ѳw;K����M�
����}�X��IqGqȳ�30��k�D�\���-BHQȿ�d��>���0���\�^{�U�c��ߺ��}w����e��Sd*���9r������ؤ� ���ą9�t���u