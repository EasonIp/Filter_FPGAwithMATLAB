��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$���G�S*J�Ш��jk�bF�����\��!G�%V���4�<�S��n��X��"8�u����erB�,��o1�K�4t�.|IV7���E-�bOTu?��~}�e ?���.����u�� �������O���E$^!j�����J���A�&��o�q�6�D���O�e#)�O���PC!n�}[�)h��Y���R�P��e�hh���^J2�W��༭
������C�@�zq]������u�Y�n�S�A/g#}���߁8쥝�O���$jo�:�)��Ng`J�+
3�R�X>�M�R�`���W����n�+ηZn��!�e����5�\��e����!(�j�0���$�2��p�� Z>K�����Ӳ�4�����0R�kV��AO����7Lu��4�S��������_��T��zV<@ 2�R��Y�P �[?2�+{H���#T�x���¤
���^�oR�և�r�k�cUmWݼcb1J��͒������v(�BFw~��
?�~ֵ4}�#��f!\�)�lW �`����e,s'������	�'ʘ�-��(Kxzv�dI����1�^�S���)ӣ2�_r�iWK�(]s�l
nP���m�{�r��F��仁�Ļ�Qj��j��#����i�xBL��?g�Z��6�Y1����~Y�G��H�J?E v%�:X1Da��j/僭�.����W���'M-�Ю"���Bk6��79�i�*�jZ�2[�X����T*��%8�ay1��w,��\�<A��	�1\�����E�~�3s�l7�[��r�}���L�����8�UK�{��t���A�T�����\��5�F������Z6�j�o\���-��1�g�%.��N_��7�L���j��6Emp�,�k8w�10¿�
fܩ�æ �;���P�RG�K�h!�W8p"���$���Lr�&���q�[��P���]�Ї�>T�D_E�i��F�m�C�!R��D������ͭ��F�" S�ݼ��0�X��I�)�S��W�����)<��)��$ @�6�F_[j�5�uqT���R����8w<kn���Xq8D�u�t�͛�#� H$�7ik�gs�f��uL��Qς�+�BQ�|�����K�C���/6��,��{��z=��Q���6>��NmF��-(3�??]?��c�r�jP�d�Z�S��{�}���Ong�q�X��;,T��)C�Ԍ��>=Z�N*M����1d��-d7���".[2�z�.S"����^�KN��T^�v��/]=�79+l	.���