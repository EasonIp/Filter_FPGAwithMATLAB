��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$��x?M1u���Uu�'H�9}��J]t_+����n"�$}H��5�E?i�*_��%��\�ulqÜ�>�bH˯��猇A-�x��L��7X��.���U��dB_����Y�WLD�i�{���n��l�"f�6q�y�o�g���T�6*}/�+��tݿ&�c�֤��*-Eg(-4�����2�⳼2����,v��E��"鎎�����w{����%�C���_	67.�;r����>��^�{�NS�u�_.�Wp�ʟXCQ���/�:,f��E{ �	��F3�y��g�R��w͑T���=O���0�_)/?HB��4�.�0�,z���Gṯ�ZUՍ���!�Tcq��	;O.���sg�R�W8�a�W:eEP-�sr�x[��E���c1x�O�n���c�|§%(<�5�?��T� A���e�ǔ��%�Uz�4g�}�� ˉ`f$ko����L�_S�X{������f̬�7��Hǖ��x�T\�B����Ɣ�lNKΥ^0w����H���Zb���>&��d��y�,�iP�b�H�S�ј��̃�������F*$��H�E�y>�ѡ��8��i*r�3Ɖ�j��#������n�j��f�eL���!
��&U��,�ױ��t�?��ږ�#�+���h���ltr]��ā��O�$�����y"2�z<���I
3@�TC��JS�dBԣb!K��Ѿ�K���d�)ߓ�_ґ�5�  tcb���Z��%�jy@�
���Y�o����j��d�K�9��M����	�3w[�	#d�E�v��MTԢ@�࿝�XW&��<HF�|N_s(�"�����>�<����2nq��ep��*2ш.^I\<#�S�I֋�hx[�Z� #dշ�������m�~~@����I����ՉU��ΐ��`b�4Fe2=t�0���F 0(���V����~��G��D�R���������2���g��P:\�Js������:�����
:�s`/�2��������w:�B
�)�l�|V�V�P���^q��	>,��9-<��7��C�� �b�厰5��qE�씋�kK)),	\���V���A��@q��^�G_�ޗ8)1А���4���]L���ڪ�)�!|HQK�Y�S��a�`o��?N ��3��'��EƸ���b����D���9d���ǣ�>b�%�{�}3W�aR��C��i;�qz�ʟF�TE�l�%�߬�V�_�d(rwi��6�m�5�+8<�T�� ��_0�r����g{x�u�.z�?��LJ0\�i���ז0��4أo9��Bl5ɦR�����p;�Δ��h���m��}7�A����Y�U��B&��Cr�e����
��{J�����:�,�P�+���:��������v�:x;�0��pt��<��V���+FA�~��F�>�[�������O�::����k���=�hTH.&��NDO�� J����qk����u�
��$AM�����G,�9��	]�ʑv#5���:�z����U���%AF����}��(��9J��3��?*|���;Hs�GM�'��	B�^L��ª�5\j\����B��g*F���!�;����uvͽ=��SW�PI�����"��F�?�98H�Oi$�_�^���Q����T�ľA�
��8�)T��7螳pr�F���CER8P5ٳl�Z�Ҏ`����]j/ǲ�"�� �����j�#�«B~ǆ�a�p^���5��y�o�~~u:�:eX��.8xvMK�N+T�ݖv��)MC�n�UQZ��ءP����D^��]I,W�hy�C/<��5������WJ
�`q�m? ���f� ����Q��\K=����0����D�K?ʑ��&كw87�\eA��O��e�|�DЀ�c��E���-��wYs����WP|z������*��`�-�]���X	�v$ћI�fレ�=�p�?xoao|�q���3����!U g�<7�l�� �2un}���Dd�xa./-+�2�e�Ҏ
��Z.Z`�}��Y�	�������>;���{�_�$��L�_>'�	���^F#=�u<l1u�PA��D���t˰9��L邟�P6������ҭ���aU&h�����+ڥR��33I]<����,,악~�m$���	b��ZI+z�ȆT���eu�]��β�X5�a��n�XC�c0شx�X���J̡�j���Gft@�&��p�=�;M����@����Ό��l��yH��Kh�H+�(�I����#�K�% t��:�ߚwF,���qc7Os饺�6�2��������U���%|. SZ���¼A�=i:蝮F�L�ȺK�|�;�1�ǵA�Q����k�q���B�1q�@7w��j|e7�>"Kr{��]�|$���8�j홶��{R��a�=O��f�8*�$�Mc�[���Vr%��^ʿ�x�6������D3�3��-J�2��Hּ|�y��:A�;�|ň��U)4�6�B袙V��I5�9A���`�_�Xp!f��}:��{o/�An���ML�`����a�<\�,M�$�i受�(K�ᶚ�/2|�)xo��?�Q�;��M^i[��m�q�^m�(T��WVk�D��.��Ԉӄ�8�%���������(Xx�k���A��1o�����dbm9��1]��)��䩞��e�9���4��+A��AB�мd��O��y�`�������~y���0�w����pnW,vwu{tBy�To�Se��t�ߚ���:���U)?�tx�h>��A���(���`ߖ�ArM4��E�M_F���.��I>p���Ϯ���C�>��Ϳ��xGi���]�!4�	f�}�H�������(�ꦁ�?��y��c��r#'��L�U.���%�N�!��U�L2�Y(N��P����2#���i%A�:�N�s�d(��]3�dIiT��!!�MjBzlH��H�u����:*�M d0>M/r�e���6sԙ��S�س�IΖ�5Y���(�a{al�u�0w۬����哸��%;����q֠�t����bNp�|�?�n�_���N�4Vz�xW� #m��?F5�-�.h::])��~1y��}��5��M� �,�9�A]����>��&C���&�`5 �cf����J�.d�B�E'B3S�y㤨���$8(|b;�W���~o��-�z$>*�\��v��!ю\��,��9h�f��߇F/&ܫ��%���7S#!�9����"JƯ	����M���<g�����B�r���2���<<%1���t0?,�Z�%�-��6n彠���DG����`m6s�=F����V����U��ݸu�?�H�Ц��{�9Qb�[oʔ�T�L}D�
�Q���L���"_Q�T����5�I࣯���x-=,F``�����_�Zi�l������P���V�
(��ܘ�3�:.�5�Q�%A���ڸqB>h*�3õG{01��𐯦(Y�q���<w�gQb���*F��V;AU䷁e�yT�RRP��{��d����|�K�fA`�Y]��\!�!u+'�2����It3�{��Q^��1�1�HR���[?ozJ�1.�<�6.߃'rM>-,�-*�F��q�Y]x�y�����_޳9�3}͌�8�S-M7}7�R�dyT���� /���[ ���O��7BPpua��!�"8�"M�2G�d�[0{(����OO�:�l<������t�k����[��|��a&8��:��.�.��WY���8)��g��x��qH�&��������$?���%����*�����N���ioJ�!�����&jF�(`BI�ޢ�p���ae[ۓ����,o�/��h��	����0㼵�<fqꂖ��p�j�pW�����$���ZL��Tf�(*�@�Q;��gݗ55gH]����$}%bs%�Vm���^x���Ni�k�4L��"U���,�R��d�]���3� �/�>4J}�ͅ�B�E���]�Z��6���K.�4v�X*^��@UC�ABf�͙�a�fT�E����-3|�a��;���ٴ�+j��'�g�H-d��E��/���V;�6Y�Ճ��#�˭���Da�A>l�9���(�.���"�s�H*i��u�-�H�JRs�u��f��V`P�f�3�Μ� �DDke��3��H�t�5�<s�&��UZGU��谀�C�k3ۮ��/��km�j�_�5�Ѥ��[t$�e��� ����@8MI�.��r�S���H�q�N����ެ={��N*$�Ç�>m�K�򯚙X�g�RS�c!�AX{J����ɱ6�t�&Ĥz��<���B�*��3�+J2�O�n'�@:sB^������~�"�fn�h��Q�T"���������$FS&��_�Z��a��-���~�bjj�E.hi��'� ���s��lGޖ�S���pg����)�{ 4������u��FI��$\>�7�nz�)C�����B�D7k/j�#K�,e{)�(�hk#)\���,Ju���,��	�:#;ɴ��(7�J��m3uYa`��<�n�)���0g�>/��X��j]t {�m
7u=�����R�k�ϝ������e��m�չ֒�_��i_���҃u�.�rxH���cIi�
�]�b�#�L>i�p{�A���m�a!],���_�,JHf�!Z�8��56������$��7~���/@t1�+�ڮN�5�.<N̷h������NS2F�+�D�&.��-Ӌ8�ڎ�:��Ƹ�W&q��J���@����M��X�bC�
k%�#�z1��<\�I��-��h�=$q����ng^�d�?��hm��̒�Z�Y�����3;���R\��e�6�7٧�� ��"#�()�g�����EQ�*y�i�����.�j=��
�O |��M;>7�>]W��U��[�¦��LR�;�&ث�>l��� 漁a��h�ܹ��")I��nD|G�u�q�ϖ�q��o%��G�������He��d���#�����՝9�1�c08��\�B���Z�>�`;�g��l�B����[����w
7V([��f��-Y�[,�ܐ���9י��7�qw�a�E�)��g�\�hg��Z;�U�7uxÁ+�Q�3���m1a����I_껻4�PZ
tq�~G��5]�($�9�m�h�H�����I��,��k�k�<d�|~&z;��p��e	i%Ko�}���|s�*�����K�C�$�<v�\>�-Q½�����dWb�Iw�2-� ځ��rfm��*杷1>��jL�W%p4:p�(_���RZ��Θ�(XS9r���np3"5o׻���m�B��n�?���
�}Sk�s����"�ySɤ��$����S�:a�>�Q�Ow+��A.T�}	����(��c�$�S|a%�Z��T�;mjh(؜?:��:�|�����6�Jͻ9�N�s�%�UTue�I�y(І��Zn�����W��.^�_�D��۸A��b5E�4.ٺ.�J�z����Z�o����٢�}^h8K7���j�_-�I����l.���<$�~�２�7B���n�)�w�E�g-�fc51���U�֎����e�]c}��rTA�f�b�S�Rñ�֑"]�� �^	N/H�H&4�i��l��j�	��\�r�ʨ��5>���͈�	"�U��>�]���1�7w�۩�.-�]u9�)�th�#�C��.O�aA£ ��,aMf�D�P��Mg�( 1m���c(/�� �0��7��l�\�m�a@��nz�7��`1[���=R#��X�E����1�<��bA���苋���c.���)���7\��8������]����ǩ�<]Z��ЗC�;pZ5=�?_��;��55��EhV�	���>��!9�)���ɞ1A��lG�Q_�Ub%tb�ՀƇ��
M�ݣ�R=��G�)��TE�sv�y��Ȝ�B�x�3� ��o�����!E1SvF����h�A��.�9�1��j�<��[��TD�;L�v2�����$�}�8�+�IM��ey���:�
�B��2"}�S��^���QƒD���ôS+n��,�.t��'���hr�����8b$��,
ެ��z���D޲�M��L�ʰP*���U���_����P�at����e��_H���T���>C�3H�d�M�K7�	����!�V�//,4��g,������sy�0oV9/�.���P+���/pYK?ű{XZ��w�z.?�C6$�vϧE����)�U�f�|��1P�>�R�{�xm�.<?�G$�$�����/X�K���×��H���`0����S@9v�|��W���n�y�Wd��ͣ�Q�7u0b���D?N� �K­#�*Q/ӣyG�<�z�0���AVҥ�:+��G%��z���8����̀����4?�(�ZF�����.:��_=�¼W2ܖ�S��=��4�_w���=��5q2գ�̻���S�8�C����D�N�]�؆�A�a���y�;ӄ�oCDSg�1���xRW�S��_~�5��Q�"��8&�d�Ѥ i�HPwo�>��S���2M020֥�'|rk6���Ǽ}�M(�j����ct�̏5,%���Z�_]v.�w�x_��ig�+�FY�
��6���^9D�{�Ѯ��Q��?6�iOK����yg� �x!p���QL���k�(��y�#�bxWw{qA~ʬ��t(6����}e� ��v�IntO�ڝц�b���$� [h�tBm�����қK�J����#�w\\h껧�Mgɛ���4�K-L����-�X������g���)씁hy>���:����;��N������9�d^zFv��6�#d�z�r
����5�m�r4��'� �������d�D�b�DW�m��-c��N~�9��Y_�]��i���gv�c `F�H7ǿ�-��w�_9]��o&o78XA�� ����ol�@m5����x&���;�jۤ�����l��M�~��a�����P_e2t�ˬRpﻕ_��g��k��A.t򔏷̐�W=��<�.��}F�_Fd��5��.��J#a�aQ��2J#�'�<A�e�q�Vd�WQ��i�S$��U�g��ljP�n��@� _x�wB��=�SN&_eqێ_�V<|r�q�p�]	�[>��B��H�%��PeP�[󭂲r�BG�XSvC4왾xM-͖��E��_��M0� ����ӄ���#F�d/��H/��ݭ��J�{�
����f���^�P���y�����+@��L-�I��B��3IL]�3���Bg�a�ڎ^���~XI�7+j7J�x���C4���
gB*�9uzT,m�z�Ԇ»�a>�>4D��?G��� �T�D�g�@0�U}-�ݹ=�[X�{�&S�o��-��gt�׹�}�<Q�~�ם#M����Hv�Tyh�K��Y��Oey�-���J(��ż��_��������>�F����`�j��|�V�����Fۛ��##������I?���-gߧ+w�Xʉ��>Xv�Y�ion�x������Q��n䙲�.��ؐ�+�7I/�\Pl7Ë�@�=D F�,D�r����Rp����7M��o��KAQ��#�2���Z��,��¨*�Z3���сK��~�Z���8@��/=MA�9C5V|"��NZm~��ռK�EY�gm@~N�
�`w�=R�(p�u'��u֧�2�5Q�`�ٟ����\�v)�\�?��}h��Gã<�E�nsJ������]��ݐĚ�� 132��d�r�d���V+g���� �S��ʦ�W����b�5�2��F-RfA�t�m?�G�q-򃨻0����O���I�b��[�����b�cU
����H]{���Km��O7��!�M�/E'{�.n?���5�&_�Ϫ(�`�;8�
�I��Q���V (\+��QG���6��?��MݳҡS�`�cß��
1&�!v���3˓�j!�:3ge�ƚ<�P�)]�f�{�J�G�/�<��-�Kp��(�Q�e����#��@�Oi- �����d��U!���� ���O����_o��q��E^��G�:J>i-��B<�>w�B�kD�8�c~'�|i� ^�JY�SUK
��
�:�h������#����4�X��A�Ω)ai�YϚ ��'�Qn��~V�Q�<ʞ�O�I �geY6'^l�7���$f���K_/�T�O�bJ���ާ��M�כ�0H�o�Y��>s=�0����N�<����Fa��j-6Q�2.�u�)ǀH$�l�AAܜ��[w��u�?��]?,������=��Ǎ�Tj	=������!�,t���6��J�止�CZ�d�,��k�V��y����P�3B��2D���ԝF���b-���KJRߔ�����FGX�͘�r�.���a#��p������q��Kl�FxS���9'��`�G� �^�PǸ,a>`��� ��ȿ���3���T/k�Lh�n���F���`1-�V��{����UF��WB��ݻ�����s�ڈЬ<#_~o3}�}��,Ȧm������qB�����\�:�$	E�^ڇ�pO����-nR���΄Ľ��8���6�qX^F%c]�j�*0;�v�b�J��6�*��)�ެ�0��T����Q{f-�=�����Ƌa����Vs��XR'-�ӓ�VFX�;[�]���D��z�se�
�`���|g�>H�������9��X��X�)�w���q��`)���q9Ly%ņ�)����%H�T2���i?P7,���%��6# �첮�̸�p�/!�:\(>�ߙbJ*�I�+Ơ~T��xc�e@'�e �q%�,1� hn��.T+�F'��!�s���^��*|��'ړ?�d��򽉆`p�)��[�i^�{�g�-�g��]��SYR {�v���Ft�\�|+��T��3���%�jkA	�8��!Yd=_{�ڒ�8XkPV_�C�]]u�Ԁ 6RQk�`DԯD���Dm[zy��(]���pÉf����$�`˒4��N��<����mQ�]ҕ�	�8�����Ltr�fQ�}�{׏�x���������]#�?��P�H�W��/Z�m�M�yNJ�Ƕ>Pu�_g�g�d[���q�	�z=Yqc��]w0Z��"���r鳒.Q����a�n <�D�X�J����
��ŷo{�;2ѓb��DM.��⮺aV�߭&�o`���<b�eD���0-�S~�/�������)���@�O6�<�,��.��,�eb�P��c��Z��q��"Z7�J �^(X��5a���TiWY7�H�H^�HʚM�g���W�6��(�Ba�Wſ6�9���%�V}]��2�q����	������B!�Yϭ�g�F��H RWH�<}�O&��JZ��f�h��Ρ�À��$�,��1�[�@!17��o �	h�}���Tq�UJ,�r��%A������6ǻv�����x7v�ꋍ���<�N�x��D�����u��"���J�H"�����!��|��w<�.B�O�c�=:�CI�:2���Ɉ!B�ߜ��n1��I��_�7A1ܩ���0��?vR1VX��f.X��7R�=X��e��^�eƱ�p8|�6��K�$F�A�.n�8�T�$�sk֕v������Ԙ��>�0�������rƼ����A
�����I���w������ɉ���i���2b��]��J>�cݰήf�Êw@F:)�r�.��&���L&�4+}�K�i�3=q�_�fd��/�%(}���7��$��չ�^��w�4c;]�ds	�N^[�wbAZ�U���D�$"�q����[��S��]�B�3��eضS���2'��$����-����+�^�`����|��[fc�ysb�韉\�tkӞ^�@ng�:��̆#M8��^\��!Mԟ���[��a��)[�D����$[AhI�W�P��L"���e��>�����E�1]	.�rg(�w;h+���p�0�����",�b�,ZK]�g�%���ś�,(�*���]�h��������� �;���uv���K�w��X�5�%���i��*�#8��iR{����c��P��,\����ER�-�bd�Oe!�뺅]9�l܉��m�˴?O��ga�;�c;��(�U��d�^�U�D��!��~��3O�������z1�`go]��,�(2�%U
�-�T�I(J�\�v�[���wR�(ħ�X���åKs��`S�,�o�`; ���_Pu��tWS������F�0u�' �`c��M!��s�F�o9#��������r��#�C���1�/7�+>{~@o%����K�}�r�� Z�{��'1�|��*�9���B�|E�����>a*��J�&z	i΍�J��G����B�-$J ��tGc�x�	��q ��~�� �D�be�{ABnR�d�e��^���$Jl���X�sZ*��LiW-}�B_bQy?W�U�Z�HgZ7w8�	��t ͽ����T�w��7Q	92�W��m?p���a5����q�f�O�o�Ʌ��z��(���7�
3�2�cP����b��`���!��^��y ��OK�4�w��4kN�Ϋ�3�����#u�eg��l�'�/�X}f[Q���M�O���������_2��ҴP�@��=��)=;܎����\5�8���7�i����
���zL�-!Q�BIS�U]:ç�����)7�0>��:���F4��v��]�׭Fj v��0���܃a%���7fo�u���)Dm�)��7�=�8�?=���;`<m`lĵ��g�X7��O��u�9i_b���D�5>W��DEU���9��L�k��}.C�ok$����<q�C$|�e����%��z�l�@[�=��R�X���IӠ��[ �:���7ޚ����R�4�-�:�K��y��Ţ�P"�7����`�L����?ܶ<WZ�bV�9���� ����R�F~��,��+ͧ�4�z�ƻL/'���kk_�cb��vi�g������}��{��U��b�4|.�͠���{3�ڢ=���\�Ĩp]G�������!%ݘ _	�)j�(�ښ���̓]l7��u�76�����CE�e:1,��mݽO:����m��n�.T>+��,���]��S�)�w��b�����U��Zb�m��Xjq�}ZAUaЀJ��zX���i�HgV۩�\�����#��ziZ"	t���u�36͞�ԡw��)������4e��"�c��<Yj���C���DյiVq�*�A�W���N� J���?�����ŀ��g�if�Nv{ސa����u@=�������ᚧ}!ik�˿��I��D�<�d�:�=�StV~%&=;�'��Pk+��9a��<K��^Ð��#h�9�F?����J�@���Apq4���c��a�q��N�S���|N2ga��wSB,�Ȍ@qWV���HU�M�ĭ�;�%��w2�rD�����mO�[/Uy�m@>��	8�J���!�l��K��/:i��뾋?����x�8��ٴ�S��-SV^"���.����v���T�{-��5��@io������f���J7V�?o����J�V�u�܀j�^��E����Ep���>��<���b}V��Ð�,�a�Q�~�S��ph�\VG?VC��*�-��Mq�<�/��<G�$�xp���T?�!��%�Q}�Gw8��(Z��Nw�?��lg�z@��ӝ@y����Ų�Ͷ(	�v�6�����9;�N�CS��>�؉�M(Hn�iȰ�bQ�*g�r˰K�`X|�P.�j9��jz�D;��L�_^!��R��#�Į��x������p��� �j��U������b�՘��ҕ�ΰL��	�X����MO�skZ�5� 6�	t�(C�O��6��&[�����u��K�.�9�E� =A�����c����Z�Lf]
�C @d�΁ܞ�����`�e�6�*4"L�<����K<�%K1d��@�K�U�b=I�����91��C>���@"W�*{�.��
�%�����($~�r�����l@������Z��9�I�f�q�Hm㥋đ�����E���ģ���e��ߊ��dr�(�Ry}��f�ϒ��&�"}���SHs$B���"���	$xa�l��L�]���8��}�r}�N��%12��B�w�UM"��څ2	9��V�G��a4��V�6m�aҘӮ����e-�0Ͳd�Q�{+#�!̢r�ؿp�4."�����`g5�jc���7o�z�N�ISixK���ޜ���+J}(Iƹp�Rƛ�L1�A)�ʴG�f$ÿ�/Z����8we5��y�8�r�6&�z@I�x�ŷ�ج��4���K�V�\C� �E���hE�ľ<j�S�d_�U}bK�M�2��?ɜC���zpԬh(���t�P��dF�"�x߻�'�Cc)ʍ.����⭶&�N��Jϧ�"�,���9�o�P��r*˕���	_�vjj9_�D��Q��d�Ty���6�\|��|a������p���]h��~
(</��.���Nq)�d�-�8�[��IkLD��::V�-83n-0�`XHq;ţ j6�Z�_=�Cȃr�gv�Ờ�;�{��hf!����W���$0˒�+}d,�>�L�?�W��1�v��干c���Ra�����"�6���G�&t�?�M���(�*[y�u-�*� ���.w���'ʶ$���5�s@��@���,؞���qˎPЍ� �g
��I�`����t�FAT=񸻓9F���Qz�U!O�����ӿ�Y}�F�yQ���Ư������[j��3�\���f)��`�8�/V����LԖ8o�l*v{�1���+�>+ľ�:�ȷ� �A���KF���V�r�7�r�ġZ?�8�kP�d�ـm\�yo���6g{
��'�^q�dJ�ִ'p�+���N+�U�+Ɔz`GS�s�C��T!>Nպ9���T�����Az�k��C�9�]�W7�N*�ʀ�A�T��&���5����7��><���T����=C�,�����m�����9{�>�yW��mb���C�#J1컴�у�! }up���zŬK�d�8��^��~���;�ڇ�!<�7�wSx�jx��%\��~G�y�A�s�<��'��`G�^�*�i96w���⚤��[3�����j+\
���%ߥ��<9@��::��r<�v�?}�w���@���Ẃ����MGTp�FS��(7��E|L�f7������������L����������?�;4[�aE�,���nf�an���`���p��#�q�u��+	����׹��q�{5����!f�>�f%`�����G���ή�&7i�y߀Fvf���"��iW������j$��ɮ/�L?z?|�ci�E嚳��i���=�L�I��\)�<xYh������FfJ#�\�ϣ���U�)�W��R�wʖ70g��q�mݮu�a����v.Dn6��]D���v���n.O!�1��L�"�����>&�C�))�r��U�$���w�Gw����Kh��~�p-��G IIak�2�u����m<g��V��I6ׄH�	�AF��x��y�ёΓJ�Ȯ��s�$L��h�Ь�.��}���|a�2/���X��)��i1����4*�b��k.���!����(m�������~9_�=d����<�X.���l��sߕ����M�,
'w�� ^�7��uYW�92��vM�csmJUIj��5�6�7�pU0���ն>|9���wO�$}4�����A��V��Uq�]x�@��ё�-COT��
����jE�$�<���)�5�t��*�/��TA��ȶ-Y6�g�Ր��phU�`��p�WF���4%��?O(��UFSo �'��V�}��-�	{����Bɪ/E��r8̳��%�7�٣����BL%DHQ*�0����Aί���n�}�l��݄�K3ז6��� �VG!r=2� ��r��3�*��II�&5)� n��@�q�?���ӗ@������^ad���	�@R8x�����k�8�xS�V�'|@�B�^
O�K���{��+� �Tc?,����'�%	�>��5�V'満�w��Ѻ$��Q�3
��ę(a��oJM7j�<�=�!Y��B�v�Y�&��X9 ��5�is�dgQ9^��Z�d�آg�VM��/�._�:������M�)광'�%vl,d��B��*�ņ�$I/��-`3TFB�+�K/��q��c��_�]����=�> BG(J��=�Z�s��ui6� Q�ǆ�o8-ֻt��v���4+�3��K�O���Y��?�"���~aUYF��B#gM:%]��������AY�=ڠZ�U6ɝ4v��tٴ5�ݳ�M52Z�~��`(�\O�q�����*��FmV8k��7-V+;�;h��s���e��
B[~09��2�2/{!���p�'���w��)��mR���S�*�uo~�c���G��}@�P7ز�����9��k������y4/�T�1_xo�V�����-;��ѥ�y͍�jׅO������8��o�"S��!��>G�����o�б�t�S�y�g~����5�'#0:���<Ȥ��r��w�E��̹����̡��Ú3t�y��F��;n��0)�ɡx�4��nzF�aB�-�H��pڷ؆�Z��X�f	�S�_h.ROIy��?�A�S�h���F�T���x|�Q�07�*b�#��[�{��u�k葌��Cm�]���u�� KSP��x��G��ZeЇ�psX��c������@�~�+w�&��
]����E��
g�f�_�v���k�|�F�l���h�ͦ��8�?r�{�Ż1ZQ�f'+��O;�E�Z�D�3vD����
����l�������f)��8p�2�L/u�0��$�o
�Q헪ݧ�@��8t]9��ќZ�"o���#nz[&CW���Fa�h�Z�1ԍ�$���!I^�f����
QO7*d�4�����"�N�z�0�0��""&�I��mm��c��r6�Cpi��2�i�]�܃-���a�{s;�u�[r��er9��kha�PO@�F<bP��^R�������Oհ�w=WX�׆���6��\#ɯ��!9���ɬP>�J����~ݖ�6����Q�����J�q��nX��c�~p�f؀���*����+3���{���v����󠬚0P�#�p�=J_#�-��^�ĸ��cҟ�*�>��q���[0��q"U b)��ч3��W
I⡥y�>��	���5�p�,�|#�L���}ab4�kO���:�� 9G��:G�&��5�saY8�h�����A�1���L�W����z�,7�4�\b����S��I�$�xtz�o(��xL�jE+�~![�0u�!s%�ZS)�t�q���&/��$.�����N�!��"�>_�����E=r��!�0ד-�W� �pMIjyQ닽@/���_F��"�`�2VN_v -��-yZ��|�B��-�����wȑ��Y/�lK��&:rV��YC7��S���PcU���a,oMs�L���ᖬn���ۣ�p��K"^�R,#@�"8�E��H�S�����MBQT� �$m����<O��&�����sv�@�rYFN6�㙵�v��"�BGCSL�Ahiom?&g���r�i�i��AN��m�|��U���V�Vm�剗~��!��^N�-c�J󤩪5�)�~]���m��ke8�@��R��
��"ʀ�W9Z9���@�����J+L0��u����������Al�������"�ɝ���4��5D|�D^CH/hȨ,e�/"ܳv�!S�������9��Y���w��3`����%�i�<�~=f"�H�#д��*�~��[Z��Xa�%l�ȶ[�����])�'����dY��O9�{1z?��B!�!�9	��F� ^�VI��nl��4d�S�-�'��n�4���8aQ��Q��(P�&ѥ15��pa�e��8�~�&�ǖ=� �������Ÿ�17.��l��=�α�g.�Ih#b�|"�9mr/��S�&EE]�G^f��w:c�8���+7u������x����;ۺTb]�7��C��\	� ���j�����>�����#������"۰���^��3N���^��#�B޵v�.��ӂW<�VNr���h��-���!�Ƽ�乣��p BӔ�S���ɉs2}*H��v�����3]zˣ�8�є��;l/�;��6u�����l����8 �jr�wGo�l��|�J�a_��� �k�\{��Y6�������z�����`�e|�%ˑ�]R�͐j�6`��.h�Jph��?#%*nz�	t��S�
��ޜ���9Ќ�z�L�RO��H�'�����}Ѡ\�:�$�f����}J{�+��ݫ':�7�w���n��I�K��u`�R���㗺��g��i�>���l�aٽK��MF�]��1e^b7O��9��d��k���v'�ey����h��y+"6�@����l�2n���Vx3͍c�ޑ^�]4��e�d�4R�WP�A�% :���:�բ�r	�\o�'���u��3���-^�S���8ĿBh���`��%?t��{��QRy�ت���dĘb�*�M� �T[��UÎ�x����[���N��m����X����#�b����J��<�� ���[(��(�SrNon%!�������B�KN�Y�}�GKW`�Ҽ�E���(�6l�{
���PvB�o:���`|������1
a0���Ty���A��X:�x�IĦ/��E��
��@4�[��)5���e���b%��[H��ou%&a����RK�I^v�c�(t��R����c*fwl���>+v�wH�	�K����d����gV׏�y�^9��a�|&\�EV�?�LH{����]-�4�tpQ�-��|���H�w� -� <��zqV30���P���uO`�90w7c�;�mXX�c�C彙��l�v�G�R�AJ����Y�����&)q}��&����O�/�#f�]�QcB<�"=}Zf�Q���l
Z��{��}�zW�m��������$�-�i֔�p�Ԩ�O�-t��e:�C��+m1ڼ��=<�5[^8ws�-��u/,k�c��O�4�x��d^,���ɺj�H	0����G!�Q�Jy�L��k��<�^6Ԧ��Q�@�>.g�q��H�����Zϵo��E�)���NPT�&��GMI�����~\>��vm����p$ N��[�x6O��k���9Ȕ�9 EhM5��>qH��EZg�*~S�c�(e5�	!�0;�C1ȥcg�=�g���R�b�[��7/7�#�h��m|Zk���+bI�=s�l�$�H�㕨���f�1���V���b����*À-z�����X��o�9��
C*y��2<��Hxm��*� NI�f^�	��^6E��|�[��駫=�"�͹GK�ikoA�k{��/	D��.��%�UT��B�f^z-��2��Z�$�v�p�%�!��7��CZH}�'���c}�AET�F�Q[��{E������5w����kc��Y��pJf;�Dq;
�m�p�+/��ƿTD�qښ��gzU+	��ʤ4b&�-�a����	�%�֝s�
P��M�=����U����[o�R�"���0�,�[i��Gf���D{Eej{�<�^2<�EJ�c�n@
�\��̥ː��$�a6C�j��皐��=�Qs<�_|�B��,�+,#���3���_�W۪�_o��CZw�7n��ioف%b�	������_ta=u箠."}L�uvU���Ă�&��M-{<�4�tif�P(u�H66��}\HQ���r�u���U�Sv\�#��B7�!�2
4K(XotױG4��(^' v��,�1�y��9]8I�ѯa��_!C�_�� q/-u�Փq��������x�]��x��IM�\N�p�\�>����0�s�T�a<#S���� 1�g1�D'�韱�4�(Vo�ςa���)[Ǳ��E���m<��B.���>�����Բ�����ow�Δ��`>���LW�����zD�*о�8^�F