��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>Q�y�`�}н龓I�����>g������w�O�������x�d,p�ܞVt�}�񺮻�G���-)?������"�c���x��B���_"2$[��m�8��H���`�/&���
{�90n��2@�Ԑ4B\���EB(�(K2�O�#�c%֩�q; �;��&�eb0 R�Q�H�ec⪫xd�Q<�>U�w���G��`�"�m}�qC�y)�巍�XD��òs�ه� �Z�$��6�T	�0�&��etoH�ׂ 1��ˎ�)3����fڸ���82hI\}�[cF��bQ��C�}���K�w�X��y8B�������+j�q�A��k|���_[z�꛿P���W��mv�(�E��� �WU������-g�g"ʱ��f�Rm�Pj�v	���b6�*+���B�FEy0v���.���	���	�N��ay��É~1p,C�}I��@�JzW4{��g0�}t��F� һ���O�� �!W��*ٽ�I��z��m��F����N��wS��/gV�G)5�p6ߨ����L�ҜL�U��[�Y*%���R?��KE�'w�`O<��$Ƭ�H����v��_&l������Ұ��=O����A���(�����Cs��G���Hn���-#��OY��I)^Qz�Ǩq��.qr�Q��:iOq���oW�{*!=���3�ǫ%�(>�&�a'���h(6�&��q��Y�����E���nM��<Pd�vի�-%���g����Lz��R+��i�7*���NzK���H�+��_ <\X�`�>�j 05Q���iT*��c�.s�ֹN��5���i	�Sǜa���W/�G �D�r����ӌV~�����\��l��������\T~x�Zf��?�Wӗ���� ʆ���|m���}�V4����u�W��Ռ�H<w6zq4	��^�wJ�"w���]� ������pN�Y�	����C��E]���q��q�������>>�A�� ��\������Ku��H���5�қ�:����u�KW�Ni����m4��YW�S�P��w�㓇~I���Ja{|�H�\*u�P�r0K������X���Z�_-J�3�@I���I|��f6�F�L8	�y�>5��f�>�-�Uy߼�S��;QԳ|ų��5��q��^�C�r�LFc���P�L�kC����	���<^<h����AK�O"Fc
�` n���ǜD�џ[�D�pD�|�"���g��#�c(פ�&bn�`qKO4s8�u?>㌕]���m���=ɸ��CX������}8���Iݡ�6A��ooG(�/�i�[���
���J��z�g6�%�s���3��pZ|�o�ֻʢ�w��T$t:gDP��i⽜����F�3��mwr,/�p-_G��_w>>L��s�� ���?�?��
 �xA��5�����؋w��b1)�2.c ��y�����
o�#@�����S��!P�/��_h�@트(t�%x���$�"�#��{�y��<�Ԃ�`u�+�T�ז�!nEU=�S,��qX��l��\���׉:Ї�������y*����d��o�5;�M��Mԝ^��{t_�qA/Ǵ�Ɩ�عkT�y���	��!�9)�+s����C��*�l$�.t��I����l�K�r�ֵh8]�	E��+�T<��]B��}�1/2���`�Bq� Q�w[vU���S�ր��"��Viɶ��+)�U{����Omx�PzPu��~m{��W[[]�t�1�>��!6�R�č|�4�ltQ���'�@"�׍���Q�Q@�E\��~0���G�6�%���gT�⏭�<8*&��ҁ�`��rZ�A���#���t����opd�Y������"��p%lO0���}vN&�B��A���5/4:ĭ��������0��*��������<C\��Bes(�Bm�Z\ҟ�q� �E��p�(XM��K���B.D>����n�B�n���@�K��̋�2Q\֩'�b�+s ��.���2XV���3�w�������ӫ3��
x���X6���f>#תE�cp�)9���Y��S�VwUja���B������)�M�W4�*�lOVV��=��<\�H�*��}�r����s������ޅ�&q�Wfq	�\0F!ϤS�e��ߕ�>��Ԭhw�k�e��w&h/V��ù�U���D�7�Jb���@�Zq �9����b��K����[�I��o���{XʧBy�f�)������,�:#cBw�w�k��˧��:�c�#�h�K\Ro���鞵6�)�6K���no�3��15��_�\W����P(S1fxq�\�Ry%�������@3�����<�{po��O�p��_Kƈ'�����[2���>2tηO~_�Џe��U���%�����������@ ��`�b6��%< �P=~?�^�v���NH)X]wU8��CCS�n��.
���ۿ��2Ach7
�w:����b0�e�.�n���'�%*R:��oy�L���k^I��.Ѡ�@�ژʪ`�|�Z�E��zm}#��az�y�y~,O���<�m�%��0v"M�ړ�],�0y�w�n=!"��ާ�b�vEz��Y�ep���#��XJ��/BC�%Z	z�aD����O�<�*kC�r��t�.�r1S������/�p�K�|�j��?�jJ`ÄQϐ�nr0�Kr�	�x~�с p�􀾇ۙ�h�ߵMxR�B;��&����j����A� �Y`�	�\��ѧ�>��,���� 3pfD>����^זWL��CB�n��I�a8b�������|�	�<�z���aVI�n%,�w�:ۖ~y,o��ݶ�<�޺�����C�,e*�d��"\>��"qU;�$�Z!f���6�\�]�����r���Pk�U���r}Ȅ=�v�⸂��j�1��Jd���ɠ�sD�δprm���<M�">1�c�E�hi���Si[��<�-�%�L^G�h���$V�� �����m�,LX�] ��<o�4jcч�N�2c�v��o�9�!��$�a/�۲��#�(Ijȋ3���p%����H�]~'y5�sZ>�s%A��r#��W�#�� ��=`RWC>t1���C���?�w��a��0�(�Đ�q1����NY���P� XȜ.T_���p|�NwW�Ke`�����A�
{Z\X�&6�FK���2�Ž��k`�Iϯ�}�I-d�	�dʩg֜����˺�2�o�Oa2��Hc����ߊi۷��s)��wq��d��KA�ӹ������6\��d�Lÿ�{�@e������%54O�q��z/W@ p��"䓞\���w^df��]"���w�Q�WԴ�Б��Rq]y3#����.x�93����?V��}�2�Z��#�(����~۞��㉹g#�}��������;<(ߠ��dQ��n"�D:�9�#�]`d�)�^T �{��D]��o%c\�Ò�����߿��`F�Î�L�)�	��tF�}H��%�y^�����՟
����x�M����~� ���ƈ'U$X�cEƒN�]7�e��@�U�ڶiR���ثI��Ȝ9�U�7����fQ�6�N��S+�P��N���j+�5����cs�������%>��4x�fs�*�v���9��h#D=��aq�L��W|�ͨ�^��NϬ��T�W��K$B֤J�w�<Ψ@�C� �Js���ж�X3��ݰ%?[���ަ�5� �ѱ��n�4�WJ�v�]�����o����
�o)�BuS��Æ�~tg��t�F<�C��9�O?�x8I$,��,�{{��[-u�Ҽ�����	��w�1JyF�gx������j�=S���͟frDvۢo��4�y4tK�W����r�)��lW�k<Z.��:^?��]1���*�'A?��|���,����U J?�Cև�L�::�E�C�x��V7������i���}{�Y��2�{/J~H��suhy�,d��&jO�i�6
��Q��+�M��-��:��aC٥�R!�8M�s
�(����0�vH[�N�Bl����6�������<��6�j���݁�gS���n�!`O�����D�e�P�3����.C�O ~�6�ă�,:�wv�I�Z[,i)Vb����.��}{DC@���"
N��{<�΂����Q�*�ɏv_Ov��/������c�������~�A�=h@O�|�dg8@�ߡ���"h���^��X	�����L�͕�b�6��xT�T�*��9�����߿L�9�d��@ߢe$��Vq�~{��Ay�_L�=��$Gh��,_iC �^�Y#��I>;�G׭��\mT���o�g�+Z�ǁn.�p\��7H��|��Y��P�G�a��>�F��Gx��Niq���5���,��Lx�M����BO#͐����_e^m��g��;>��s�mp�ʘN�{����l27�K=�1������3͛����$���"�4�^��nF�-�M���v;��͵�b�ќ�pu���V�ĩP,��ƾ�ω�Oǌ�"J��g�oD���uf��@b��:�P��N0�Ñ�Mic���#=��ҖƲ�-��fH���-��Ϥ|��u�2�z����-_�%�؈2��O�7#_���@#w8�|dc��`�,�d��.���tCD�+=�Z[��E�G8O���Sjj��UZ3�"�{��L�kz>C2-e��|<��������N�Ci��H�%����>��!��n�W���1u	'"T��"�L���N�N�3������ӏ��e��V[��k��s��^bk�����>:4�v�S�z�h>?��I�� �KK g��M`<��sO��7��o����z���@@[��L}[p��?�T(ț���Hrn��VG���W��ǒ�Ԧ�
�Ê��`*Gy����?9�da��n�Yu��d�s��IJ
a�ò�K\����m���F�����!r�#9�PG/-�a#�DX���L�}U�g�i�`k�9��70��=�ރ ���oER̫�F��`my{Ϭ���فc��������-��1����/Թ��%������o�:"�v�������b�69G��.,�!�{qNnq���|T68~��A�^X&l��ƕ;/���Y7��1m�R�(7ڀ����r���YjJ���%ƛ#�jF��X�\T�@9Stzs:�U'�`qt�d4C��e2#1�F"�|w`�V��p���w ��y~� ��L��Ww%r��#�$R��m�ܪ�`M����b���)[�����.6d���0�6�� ��x,$0Dp���Wވ�S���	��L� �Z� ���
۽Q3��Z�W{$V�r,
��-܈Nw�h	W����%s0��AO6=f(Nݰ��c�#1V�UV�4kq�Й����V�̈�e"�9(��J�ߕ�����k�,=�E�ABdߦ�Kǐ��C��:4ˤ��	���mb��3�2w8�H�aQ2�U��4�Kw)��`'���٘ǳ�g�n�c���2�|֨����F��7>�"l0�]P�he%ݓE�G���P�g�V@KC7A#�����|m�ȱ^,
����U��.p��u�7�+~�Tz�ʵ64��<^�C)\d^Ek�,��n��wIk����~�Matm�r�R#����(�'Z;4Z���;��L���v �K1�l�1a ��Y!@�|tփ����w[�ha�uD�eZ�d2��\���]���M��W)׭{�?��6���d�?��?�XkK�t��f;��
���� �B弄��Y�А�����!Q>$P�T(�_~�s��W��z,T�,nR�%�J.&}�� t'��>��w�a5ԋ:u�<���*'ǃ<�H��
k�|��h�>��:�*�vҭ���4lb�٩x���<������u�wc�ͤ�{����{E9�q~{��}^��*�o��l��j�S`*�3b�w�Q!U�V�{aGCU�$�;w�����Ó8�ܳ�ķ�mr��������"ķ.w:��Î8��/p\��rm�e�)jrs��**�c���~e��״v�7oU�<�|W��(�+]���Ì���A+��.H׆�܍C`�u!q8Xv����)�^�f�������T�8��t�a�O�"x�bDe�0D�us�5S��ܕ}��K\�ȟwQ���a���a�ѡ�2`M$�_$��
�mWe��������-5}�<�JQ�=�n^׬��M'͒y����~���3%����hj ,&���R҉���h��ʬ=����y�����,�#,�9����'nc�HJd�Մ�j��ox��Y��y�� ��>��|q9\��G �2�,�ǣ}��H@�~�A\�!��J�l�!�q���CCq�Tp���P܏X�����o�y���#$⎲�e���v�[�l.�y�jǼM/�����70}���Xƹ3�|ƛ��Ck�b1����Q[H�TDH7���#h�"��1��C�x���u5�7�F�Q���a3�'P�*ꍻޘ��gu=&���� >�z��Bi�w��~3��Q����i���l��Ǟ�b��B)W��`�ޓ�;A/9���u�s��z����$�"&Eb������,�d��c�c�
������qpŇ�$љ D��m݊	s���dמ�$/vJ��F������@E�B}v5��Z	Ҟ
���GM�p��(�����Π$b��(>"���T$ܪq2,����ڤ[:�?n�����7�Ж�lQ?0KR�i�S������Y/��ة,3{6�,�� ׹��ś�KgD��H�Z�2��.��4-Ԑai���
A�F��� $o�)��H��
���b��}����#�Q3]��\�K<4����E��	I��\�dPF8>WOׄ�[�	K���g��x,�����7���H�mp��'��G�2����s�Kc[b���g��5��������TCLJwu�<�$�%�m �r��\�N�"� �[>���S��]�e��yң-5ԥ��,nʺaCa5�@1��w̓��+���n���rn��^�;v��.���o�N�t�$�7ۑ�o����>.�ؑ�z9Ř*`Ŭ%�qGm�R�.�6��6JP�&|p��J�	w<��ڄa⃵6["m>�B���l�D��l>!��Ъ�)]O����!Lh��	I��+TLoTEЋ�j�h{l�='�Og�����xP�M<��w����s��D1h|����M5�H����Q�u�r�;�������^�è�ք�Žb�>��M1�md�PMdg�u�֚˖��� ��o�\`h��t���.*�����"�s��X���1���h��Ǘ���1V�;�!�:_��GU�'?���BРtPM8S��?&����}��/;|3���7B�D��X�]��R]|��`�횪軺���ݡ~Jk���n��͞�>����\ǜ�1����=e�龘.�(pl��R��;oh1<����^N*]�d� ?pf0f:��M�(D�vA%c�?�(��Ig���E\˚m%�m6@R��I��_���(Uz�L=0���޽y��� �pB>1s���e�(�'� .�����	�+2
�r2,��qv�-1���; ��U �領՝���}�j�T+D
*6 �k��E˷�<Cu�v���A��H'C�m_Do/�;%��S��FO �;Zm�Li`����H�?t>��g��+�u6L̈́R��7�'}�'����D�7L�?< ʸAP���P�\�3�27u�����������8�VS��uO[��~����!yl(p��'���PP�L|Ɔ�X�!Ap����!�����u��}�����I�Ѱ�r�܃i�v-���t4�<��' ��\��cp^���RLѝ�w�+�BiZ��\BZ��h�	��P��f5�5�\�U�Bc�}$uN���p�<ւ�Y��fN�'���Ϊi>�	r��o�k)X�\�m�õN'/���⾳n���:M�ׂ��z����R4��F��8���t�;��uo5�D����,p�&�:֫��7�ܟ� 
� ��A�ƶL����N�9,N�Ԭ��yE6��6��F�a���Q9�#�g�B�:�)�Xr��R���7E��֋h��0S+�qċ�Z�����a��Tm���\���ߧ�E���q���ve1DD����!�1[���e�&�
A���n#��/�bO['�]��P	=���k�x{'B�" &� �$"�6�ޒY3wiia�����.Q�R���J�Z8��s8SYf�>�,4x���0�Q!��^w�} EL8V�#ǔ�=����ڱ������ӛ/g8¯�=S�߈�?�G)0��q�j9 �)P�-"p��ӷ�G�$������s֑�I�"�+DT�;>�.4wR�mL*w����L���b0�;h�O��#>Yx��?�7x�\�Dg�ZA�J���Nvlx]`[
I\�n���x
�{�B��%�g�n��͘��I������v���i�����Ο�4�S~���G�)x��m�5�1��nn`}f�F���JXC���Y\����S`�R?2�n͛F�{{�z��l65��x��h��B��TUT��Ȫ��uV�@X�՝~0��'���[3�5�g�A�ʮ�f5T��A�����$�&�CP���ӏ����q1G�>֒��%��Ì<��G����0�g�}8bMk�X����+�S�۲GiC���)��lUɼe�!RL�#��,�@�Je_�!^���_�wjz©�`��>A�����Gk�t���b�3���b��#��UQ*gA#�QW	L�҈F�����CE���^�E�"m��{�@:����e6�+&��ȩ�����˷8���ϭ�3�)i�Xy|�O��E9}R�K�XQ̭׮�B��Q���LwD��,^+�H�'R���e��e�E(�Y�4*�0<.�p������ ��n
�0ԯ�F����>���e�h�$~�I�lnG}.'��>
c9����JXJ��i��Ҽ�«2,)ya��\K��t���N1It����и�i�Jr?��<���-�lA<��H�����@gq��L�R�5+>o$�|۶�yr �k�����j�3��9}�X�#3�%'N�:�ߧ �Hi����B��t���]a�ёj�=����͂��p�D�Z��3Ċޡ,l$�Ȫ�̎]����u��W��h�M��d;��Jzw��L��n��-��J��ah�����?��K@��G���_bmвS����x�ʈv�]9�(����ּ�?��(t�¨�T��MЉ���[�6�ٵ��}�h����&7R����\�,�xBH�r1�ֱXlB� M"�-Ů$k�m�-�nٔ�c�0���NAo���)���a��D�M1Y�6�2}�}j�B{^�sT�f &�]��.�s�ra0L+��8^X��l������cj9���q���F��e��BpmA��Z���X�w�LNsg?�
`?f&���J��+T�����$����'$%B����*������	��X�_�5��O��lv�,���c~mOS�l`Օ��o�������Cd��ڏ �3���|��2 x�����������pÑ��S-i*�T@ǣ��D��u�v>�Da��Bj���Ri_���8���@̶ϟ���h��%�����Vh���]�^(왩��~}�%���_��F�v�#��g�ӂ�*�Ddd�#ր�y ��u��Y�n�I#v�/�]�B��������d�X���/$���M$����-�\;� ��r�?�M��Zb?��TG�Xs�/��ƃ�������":~$��s�c���al�f Z��ẞy&�����UnKMg��#?���	Ew��4��5G�����w](�Z$�FM7�F�Viqb��.����ɝx������9)r�ˋE��R�E��e��\7G؆�;c��C ��D�JʑM����ܧNM���R����Eֺ���]N��I9{ݴ�}���ٻ�ʖ�+'1��2�QÐ�;��]�X�����6���f)/�
!}˥`�ӇSZXOľe����T3a�k�,�
�Z�y�z�ڕ�>�߷������V�D����G�4�9�w
�K{̣[T�$b)_&Z��ܰ�,�s�_�&?�V|e�"I[��� Ք� 	G³9�>����yL�#�P�ǵd3+��:�L!vS����)�P=��������hj�.�Pq�5�e�3�+ 4T�)40�w����}϶���ũ����BBr�F6_� �ݚ��)�A*҄�L�2�����̜C�ԇ�6:�2@JI�&��&��f	���;Fw����T�;T��'X�N��K̞��v��nt<ׯ	�E�5�9�O��|Ѻb���vT���жE9��℧ƑB!�Q��y4���6xtꑑ�wx5�-��
���7b%����]���Cyx���,�*�X�0a�hڽ���*pl�p��m&���o�s�sjo>����;����EJ��8�Q!'=d�f���IL؂����mu"�Ts$��-�;,�~�RU �_&�#b�<+�����||�wo]#��u*5�U�; ;]������OK�~!7�9�w�M��HU��R'�������0s���]���;6tgT&B��v$�\#�DF�@Aw6�q�/7�WB�x"%��3��i�p|���4�!ݳ{��������9YJ������F��y<�A36ت�	����ǓI��a{^����پ�%��#�4Z:�������lL��PyG�/_]�X��>��=�`41�J$�E(�`B�F�#p��rه�������]���9���X��J�Z~�}����G�v!g�����W��ݸ�������aA���G}0��ħ�.n���a��rh̆�SY�g)0�=pO�M;�ߊc�;N��>�+�'Y��8sw�E1��	(��Bdi