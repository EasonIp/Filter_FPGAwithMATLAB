��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�tڐ�!��Q�����xZ�H������
��(��B_K;bA|���.-ƍ�B)�wr�q�h1�oDu�j`�3|�?l�d�U�J��%��{�.Q~Ѻ:��E�)�֪�3��g��UvT���F���ћ�2�&�7}C{ ��e�9�W���Z0bnf��*�TS�n�2%�"��=E`T��3}o�ξd�ـk%xUl
��'V��\uJܪ���$��g���� l�.�!Y�|p�������]�N)b�l���rɛ;�6׏���bEK.�Xx"O��Ӛ�#Q����H<^�Q[J��������]�����j��u�ѕ����6�U�*��k���ɩ�so"���d/�������M�s-0N�x�c�Vj^P�����K،)�ql���~9T�\b	�TXPC{+�*'�H���O��I\]��R�O	]��_�Ȏc�����È�9��S���)�q�u�)t~&�rG�W=��\{�Zo#�{D�.۵�u�&-���ߟ�����4^���T��(�U؟v��'��~�L"�k:�T�~^1�l�[晲:�Ä��F�]�����9(���C+fV�Č'�=%�U�x����B�)@ћ�;��±��?���B�7,���1D���0d+�!A5��nB�4�䕇�L@�s1�ãKFU_���#�	k�I�	
����M5t)ǥåxm��It�����q���`y�u��Λ�_���Iy�^"����~Z����~FU�����ڠk�1t[�}��I�����@	)z�<Y&�q?٘w(�SU�����B�X+~��Ч�l�s�5'����,>�	/���;�"]�	Ma��O�����7�LH:�f�dKS4	�B�\%�Р-u���6�k��z�>��=B[� ���J��]P�/��$�����*�Y�[3���[x4�p���c�kZ�W}F���&7��m�ԭ�M���n�5��Ӱ��^��
s�׶l�ЬR������ɫ�HW6R
g�_t�� !��Y��kT�K�>?v��'{�&7�c����<��>Fҿ&W�v�P���S�w1�:/������mj�u���$����zp�8��w>3^�<��]��S��4wP�'@~陱�1�l,4
�T#\���>�j�vc�E�_�-�ö���$e����O`B 6J�<��{�'�����<M��N�a,n���L^/�J�N�W1���c?�:n#`��ܡ�K���y
���?�Σ��N���S�8\��� p���C��q> B7-�{�u��m�b�"$	��i��Ȋ.�(5i0��$��=�a���{�����<�$GVCS��@��=H�*��;�ﱯ�*n|5�]��w�\��1S��$�Ԓ�mgT�A�E&��Akc��hօw5�y�Оj�ne.��ᙦԪk�(�*����B�P����%����Wy��Ur����CS�3{F���,��p��mW�X���/�v����]�LGR��X����A)_�-T� h�-�O�U$�����"���hER��B�e��[r�߂3���<d�G�k�g�s����52!�x�m���iB7� ]���,Q��*�ȍ@ٶ���4s�tg�Zp�o�Ҭ^��û�ȑ�ǚ(m� ]��A}K�{C�0,��G���z�<{`�!��OZ�@A����-��7����X#ư�i8��Z��2�'����W�z�*�M4cH�< Ľ�ό`���M��6�"��
'n�7�1��e-&z\m�T.� !{ƈ�%��߫�&&��#y�(�%\o�&��ڄp%�O
���᳔5А3����CO@��d�/
ug�S��1c̠)NY_ڙ�$^A	Z���C����U*�ERp������^+�H���Ef�} 2.�����/'���Z� ;[	�&�#�u��Y ��i&������/F:JB���te�+�[k��}|桷u;�|�~��N�H\<�9Q�||�p�C�I�D& �I��ʫ�:DO�<̥�j+4+�!�n���(�Z���$�x�G։Rd����"��rmZ�0�J���o�/4������������n��^\��L�0��yO���N|��~1(�5�\�߬�h�94�}�qK
Z�W�[_��/�J�+W�:����e�[�