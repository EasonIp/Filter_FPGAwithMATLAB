��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�rQ��7%gN���i��v1��(���:m�>���D'Ͷ���tur)���!^���p�NW���^��I<:�E����Gd ��L�y�V�����`�N�_-#�ì9y��^�+e�I�Xɐ�b�oѯ&ioY,��z���ͺe8��l_H3ud����C �V�����5q������Jv�Zr}��pj��5X_����a��H��|���6+��g��T_p:��X��I�o��C��pz?�*��)# ��TMq�҇ �~�-�(�Ͻ��3W���n��-ҀW�J7�j�����@��:�s�6�%~��X��%�'a�CQ>���I��W�C8�E~�Xnϑ��;�6�f�����4na}�|�y���A��F�ʒ�3i�'�H��7@0�x���t�5x��b���S?���v@#B�'`��M�R���/�
C�������T!\�<�0��#(:��	�>��x��H86�騵7�������n�݅��������Z6�����7o5�Zrѐ��m�X3�����2�z֐[�AC��ܜ:U��O��1��Lwl2��`8�����Z ���B�`��˗����kƦw�v�-�iɑc��d��-�d�[�[G�����!|���M.��Ñj��E��-�e���r�����|�_7��9.��yo��hY�˂ݥ��Y����_�b\�d؏Жm>�X�����5kO�h2�P�`��~S��� -D�tB�̠0;D��I��
�Yg����ߌ�I���� m��δ/1�6����Qĝ���m�W������o�{zw�n��4��A��jQ��:G	�,؉+h��f�1mC�ɓ���eeuSo?���ٜ�-��U�d]��A)1��p��XV��r:J�#�����Б�:�{�M��=�����鉪ʵ��h?sy��J�8穳/��hC-W�!i���PË�u�T�O#i�M�S�ՐV	*�~hK�qR�˦�9\�5��#%���y�Բ��8�"��M�6�+����|(�'INB�6��ߵ2|�l	��0T��s�!�~BL,Ԫ<�F,D,kH�������uN�<�0�.y�L�"$q{������E"S�[�]�1��S"~�ixrF��d 7�X��r����P�ɧM��c~��"FU��|��F!�%'0*P� ���]| �E D�oY5��~[,D�y�lb�J���N�r�L���Y��i��o1�Q��T'^�0���3�'P�|Bw=bc}�m��w\���ʱ@���3�0�w���x1fEdv?T�~\��_�w�@�1�Y$FQ1m�-���"!;*gO��<ep�ט�4�
S�f~�%��n����o��,�9�rʾ>2�'D��η�hǜ��(���<����wi�sN��c��z���t�6G.��Oƹ8��z$�d���l1"�A�#¿�ހ<�a�v�#a.U0�dm����x��"jO�)3�����&�\@��j������OD��_�D��eEBz�bQ_�yt��-3_�4�k:6ߊJ�9�S<���.���{���J��
v����������S��u�`W��h�M�>C�Jb�^��]3�!���D鉈{���0݀��vI/�����q�|9�l�+���шqH���b0������ټG�I �򀹅.����i�L���_������H��c�ɾ@�GJY|��.ٗ��j'��!n�puQ���!�)�'va�+p�a� ~'H,z9a�i)��ˎ�ؗ����n۩�+��k��~W9F}��V�@��E$��i�m*�����jL��ZZ4wfԜ�1�g�e�۾hT�v�釒��%ۋ�v/��lPqZj���?3�I_�ߜ`��^���wΤai2���|�rc]$QM!@ܴ����9��[wkw�i�i#?����?�3�]GNsB�E6�dyD\Q� �`g�˱ji�+N&�NOm��p���%t��+��w�Y����$��@��2��m�y�1�����,�f��#��r2��z�o
�����.~'T�Mī��,��ք��߅j��p�M�y�~+��N��Z=Z��u�	DdpÛq�]���*�EG{O���u2@9���~tX�N���[j���ʿ��М��Xe��]��^e'HN��0y��c:5�s��޵q�>(��������Hk�:w\(��t�*���t�������$�$�<}Y�5��u�p"�y�q�5�o���d���o~IS��U�3EM.�3Sg�5
��d�|���T��<��� &���g#7_̻'�%J�L����M��	�s��G�%�	�� ���|rk`����t�إLo�<��qz�q���m����u���u��b'=�{`���%'�ZJ����EK���@)����/8� �V��4J/���!﹜�0�7� ��4�-Z��ƷH�ŀ���i0�L�+��mX�,|Ku�̩�5��Ǯ���K7���$�����.!�
� �y�UX��r�'	s啵�mT'	'cƫ]㜭��@��4�I�W�2�����y`u��i�`�yu��6�ˎh8养�2�K�=:3�m�T�aJF��� ��6�'��G&�gx!�uup6ۮ��>�C����S-س��PE�e����@�H��XI�;;W�,�xPI˟n����ή��e[�Wh2�Mu�:�s=
��d�k�d]@A/�%ט'�떫�^�
SDSo�[�@"�f���~\��S��1���e��縙�C0��8�� :Dr�%�jG�� ��2��SA {��H����OY�*��Y�B
�����«�:��3C~��^�?�������ı5��w/�RDZ��p6˕+⟑�!��;Js�ɨq3��.�B�}ɗ53$Q���V�~�U��6vϼ�t��?����7Ռ������fJ�o�k3z�K���[c�`,v��|Ig+�-n�ژ�fS�-|S��!c����L�l*�
��Ȫq�t��	9��&�~m.T��c��)�F��W�_�����Y�HGԼ�yŐ��bQwG�/M�hr��J�s9��ц���[?A����7�{�^A�ܱ�1=_�6_�,[��pXB,�h�߆j��sbu>Ep� rb'ʪ ����}
^i��j � ���9�Uާ2=?���4�ۜI
�A�ʇ���	��7���d\�����v�P
�I�Q'��=�&�bK�V���N���u?F�V�m���P�4�4Ô�{�j<����'���L�OoN8�[�?�:�c�,J���{�|�a-˘]VG��pEW2��s�3v����M%�7���HG����X�11��dF�{r��I����q�o���tB����^���p!�
���δ<�0���o�ki�!�Y��������/F�<�BK�M�´h	AǘT������Kf�4]c��ɰ�{�*��j,_D�u]c�Jk"�9a��ط����]��Vy�80�y�o����R9��+_��C��<o�g�yd� ·2<ݭB�chB���R��;��U�~W�ؚn?�C�0A��d�7�T��fc1���l�W�\	U��^|��� �B�w�� uz����ߣ;g��p�53Ф�@�L_f�TЇ �xixHba�����~�P���Ok��x��H�q�l7[3*�M�G��� �yV�VP<��}h�FOα��g8ۙÞ���LB���s���������B�uO G�����)-�?i�\K[ޥ��E7d�Ih7,��A�0�,�W;
�Ǆc��`	NG��ѯ�s1d�Ũ��� �w4��y�GŅ���`9<O<�c3���=fRL�\�C�z�U���凭Һ`�a�Ɩ<-�^L�4
�,����xV�IJ�
���!���{���j��rm_��<�'b�z��]�S��Ѽ�_�K��|���6~+I�͋�_�/����>^�(�f�ܮ�0�nb����1_��r�̆�J<I̚�^hYBn"_H8�V�|&��;��RRvH[^�AL���08{A��gC�����%��v#$'Nx�Mw:f&؄� �>��6h1hM�iF���Ē�:G-Az��D��u�TS^ŗ6p�!r�v:�z��w������̏Ͼ\��Pq�QX�H��_M�Vs�"R��?߿meǚ�}��;I�FcR6�2�s*�śun>v���W���l  )���:��l�ive��f.<�G�r0��wU9���&�;�9�r�C�E�C�m�+!�+�-6 t��8�lpϨ���)�}4h��M��V|��J�P�U���.7��*u΃����W4@ҞD���̶8+_�ň��'����ϐ���,��c�t�h��3��>��@�a�V:Z��<�?����~S���45ֆ'�������xi�Tw��A"�md��i&��m^�U�w
��h��	��ك���L�f�Z�X#ɻ�oN�N�����y��%�R�\Z0D0����������0H�/�ӥ��8��0 �K���-4de2�An%�)��Mj��v����I�S*U�ES)�����/m��C
�i|0�4��Ϡ	�%��C_��T�S^��NF��*NBЊ�dGǨ�1���mV�Ɖ�S�S�b
��?�����n���3�j�9
LNJX�6t��̀�Jj����}1ũ��h���+)Jc���zEh�`D"߫�f:0�ix˜�v��l��?���W�f�"O�����N�"�sC^�q�QH9[�_�f0T�hzM��H/�W�Մys�g�*�\"����LE[�Y��{������i{�[%N	'ƞK�Ƹ
x�㞼 ����a�H���^ל�Ĥ`���	$-c��"��p�u��j{y)��eTNW��y�r��~2)H�����R`Z{J�-]�4��-Vˈ��4�
z�re�lS.�KT	w���lK!9G���1��Fͺ@68�5{6���~'��+;FV�$���S�9.S�w�{�/4Ԧ�p c���U����횡$�(A-rgS��n�8s��D����e,�Ev%m��k���Z{����2�`�{DkM��D�7�Z���J$���Ĉ�b����O�e���@q�=#�Ey�PeS-�����y��4oD��f*�,�������^��3<��L�Ȱ��b��Q�恂����zI�kF�jVg°_��:E5����s���d���5�J�lu���T�M�z��i�Ih�c����L�.g��oTFmg�h�I�	Ø�(��p���ϴ��wc��]^�4���z�n#��]�v	���{��o��bU1*�0ߞN/?E�ƺ�J�a��9v�L`����"�؃1����s5�q�n���޲f��9���"��C���#�:	�sPMO�~Q����9�=���
)�5���3���]%j4��Nƪ�K�V�.�����E���{�(F@m�G_�&��7��n���4	�+��e]�*�{�Wua��<��UAwi�3�$n�z��((p�(7�5oe龒�$����@�B�.�嘙 ��5��O�V��O `��Q��Z0���LV��4�=ؽغ���*T�%����L��e�!]N�FS9p�����K�p<_3f}�ؘ��y٨�4j�9�N5��JC�WP;��h$��)�գ�C���(�x4�嗆d�E��E���!���ri��L����)��;���~{}� `��j��w���#�6�g���4�i�W��o)" 	iU&�vX����1Xz�nV6o?�狾��/6������ǩ���}�eicte)�J��zJ�M C�Ț����3k�/X�!��!�{א֮gA�R�1���{�ӹ��q`=��
��>����{�Z�pw b؎'�}��>���/@��dݮ����kKG�����s��*��8^��!���Q*MA�cí��!Mݗmp��3DE���hl���,��P��X�.L^v�F��\(�Af���\�W�䃩܇����ckf\�X"]���������|�)���&w@%����/qQ�^�:�'LC�G��Cd|"�[�aSOjIF���X"�^���.�������G#��p3%qΖ��1�Ҳ�u e{�>��iH���I%���0�W��e����Rgwl:���a��s�����6P�]}Wq�^\'�]s��z
�є��&k(��uM�h�r�AL(?r�&~��Ȃ��>��\�u����h��ڻ��L~�o��^!��w���~vλ�>+n��5�z��]Rhs��ǦVq��BɃ�Y����<��y6��ؕM.����G-g���	������)�e�c����7��(!���l�eS�E��1��o�V��#�6π`���x��X�0��}U!��s����U�u��?�J�u������w��ڮ 'uy����C_R�"KS�ӣ����ɕ=� �r���ps�!� ���X�|�����
\��2�c��#�Y�GQ���P�[�Рヹl 	D��p�=A�V3�c����Bk���I���F��r�GJ��'���\��۟tjy5wEE�(ޒ�a;]�D���F3��(x�����ɼ��⫈��Gs��4h&�� 3t)r�fQ�W�o��c��OI�z����?�7n@N�s*�;���|W˯�M�XD�hէ���� ��ɍ�����K�<��aL��I�o���!����ˌ���ڞk��¬��Ⓩ\2�D��	��o���*���'/O&Q�~�����=�%�Hu�4'��Yv�ˆ�R�<6�M�	��<gs�|�}�ݯ��X|1l�����q/H9YX��\�.��g ۢXBC'�,:�UH������l��6�$S�e8fN�����D��x&�`���E�n�ٞ�Jl��ڸ�`o��l���Z��|<�x;��Uu%��ѷT�y����>�fQ�VgėE��Z
+lTd��FY�G)OH!X��4�kHo��1���F�]�K��!hu9�dT��]�C�<�nC��4����WQ0����	���\� �
�ۉg3&�	��bm�7W���xQ��F�ʧWY3k�嚧���}K�~�G����;���(rʂ@���u�t���^�Xk�v�D� 3����Z}t7�;v<�B�6'�I�V��+�)�NB�D�n��WtM�xo8���ƴ\��l���j�,}U��Q�TB;]����Ҵ+�9�묅�"l�@�n�ب ����Ezk���&+��왡vx�֚�/�����]=p�*�n�^�/�!74i��
���gn� c�Z>T,�m�"��.⦀(��W�ى����	��hy*�xC�\�W��Kݝd"�Ka���Z��T��1�L�z4�ؐ��+ݺR�؁m��*!�����W��;��^9�7Ŗ����=�6�����-3e���E5��J~�����Ú�Ծ�6ӹm渑��I5~>S�|,���K@�o��C�I�Z�3a���]F�ĿGA�Ɔ���WXe?7#//E�aZ�0��SE����ɣ
�w�E=h���<"Gg�p���B(7�����j��*����o^�s/o��^�C\��(l���wz�����#�p�1�R�dG_OQ��� �&��M�㕛�5�D�lϻVBZ��X�Ƕ���T��k�),�'J$IL]!~"��n��-�K�:�X�t�FW���m����|�n_�J�,&w؃�8.�����F��n -w�?�#��ȭ<;�i��/m0�<^��ɿ*��>	���N��c̆
���N�-.��'���3��ѩ9/A�E�\<!:�D~��\]i���<T��("܄��̐������L�4Tm?�Cp�F^�L����S"���~�goZ�0������Vd"C����8�����|9����(Z�qd���iPe����2+����pj-,�MG2�$�T�lNYD�o&��C����^}ȿ��������C�����P>����l�6 �St���ˉ#��Mf彡����C�H��3�s��υ�lbK)(�hB��������Y�Ӂ������^���X��JK�s�+�L��J�-�p����8���9v�s������r��G��d),d�����++�d��1��_@�Gut�spچ����bcQ�����qz�N������S2Q/�>��u��ҸD��v}�$<~,��]
�[� ��n�X���D��[S�t+&��}跏]R��i(sE�,��'��W1@��>3�w�/�BĴf�
������Z.	�G�"�\K/�B���5�.��u2<�D*�HC�h��K��s4	�c	��r����͋60��-�A�UL!�MJ#)���P���Jqc�ͧ��p>8�[J�i=4�n�Z�|6����<�,/����&m��QE�(ڕB��8Q\b�*~۰��y6hU �;�>8���o�Y.��ֽ;�#l|�6,�cALD�kv �����n���_� $���}YE`��A�I���߃���̓�.$.@���UF~9���W߃��Vd��P  }��n(i&��/U�=oj "��r;a.XZh�:��G<��)����U�;b;F+8;�gY��+���.>c4�N�'o)����^���-�0At�L�J�h4����u�&X<&9cfx-��z����c�'SpD�.�C��Ͽ��yG|Ic��_���
<�Ԧ��w��Ŗ��?j-��)�&b�� ��X�A�~&�I� .sP�,ly<^CcN#漜q�.3�G\_$���}R(�X�b{��	��p`E����r��g杉V���'\7�s��G�>.��ٶWᷕZ:7�H
�D��'L����3JIȔ𨒬$�_�8�|Dk6�W�~����A箬�,��J�O���`�P{:�P1A�C��sF�^�ӝ�b��}ͺ���|]�]������!q�Й��"�ڭ�aV��%�F,X�;O��o���> ��H�%��=�BV�t2�5��s-�E���^��Eϲd%�#QB���D��beK�X�u3������&,�Fb�����(j.�/$���=O��b,��E�i�����j|D��̺��܊o���A��w�I\*�Q�#>�2��l�A����xd��P�7bj�`�x��A}����t,�E��E�Ϸw�9�ڙ�:ُ7J���Ȃ�2����#%J��S���k����ׇ5a(��jm�M��M���,.?GS�p�w�D���8�QvO��G��{����՟��/2̿�©�n�گ!T��l�i�ͦ��"��_��>��Re�Gn}i�O\��)e��o�`�2`����PZ�����SO����PbZH��w��S����+��,p*���&e�k��אp�ź�ɒ�Jʾg�^!lJ,�J��