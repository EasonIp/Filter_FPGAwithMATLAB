��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>�m��`K����٥J��5ƨ"���Ur�
x����.6P��E¡���Y��ا�o�j�T����� 7%�gE�V�}�eZB@�'��ӹ`��˟���aO�EѸ��^��PMR$�?�QH{�o���KW.��0n2	BE�\5�J��K�8В����N����?�-��zs|,����զlP�ʆ��t�^)�T�%��~l�{5�M5��<]�=�-�8��;p�����E||���G��o�s��>�ďw�oÒ�$ ?�A�(�k>d���Cp_�}G��6�c�ȰA�ٔ-�nO0�)�.oss�� ��#[��1i�Ա�0�q���Ic��K�W����g���tމ��#��ܡ�C+1���:�VWG���ͳ郔�GE�pT�
�d�׎9ld�!�Se#P�ψ�i�Do�54/B0�R����b;Q�*e�R��ˍ���q��Y�A��,���n�I1ڤ��:�2�����j��z(	��Y�_z�	���1o��.���Hg�x;��� �-&�������)7�7���I�/} �!� g/��C+�ܩ	y���|{ `��(��+CP6�C7�D�39�{�����B@s�a�ӏ^��k$�ƚɋi(/�秆��y�L���M�>�@�%��u����|���	��E�� �N�P��~�-gt$Y����Ɲb�����Z�$/m���v��b>EP�S*�.�{���鏔��Z����
kZiWm4��Ʋ����"�I-C�g��-�C�{&���!��|G��8�P��G�)���1 �ɯH����|7K�"�|�����y�ك��o�~��j
�_ȡ��C�ك<�٘�-
էY�B0\YY@B[��⾡O�Aˣ��B}=5+�X�{p]E4g%Y�%u�U@HJ��9��Ռ�����iEo�)�S�\o(ug7L�0���ؐˣ��\��. ����r(�`H���R�~�F���B�A�HA��<���==7���[��iwf��@� `.z{U�5R�P�[^/1>JԱ�S�N�Z���j��4�}͈Ly�X-���W�H��c��י���C�6$�����b����A�-���u��u���D�$q�rn�Z�d��r�|������l��~�i�ˬ�����:	�e+Oc�t	�zJ���ĆR����V�eͳȁv˷��asB{��;LS�����Vk��i�)�D�ĉ;I�B���nP�G�j� ~1)���o�EhIã�!�͒ʍn6D��{������ӡ��KL�kmگ*��L\� Ȯi��$�a,���&7��7Kcn���K|v����F�W�� އ���<c�J)=�A#z���ڛ��2s: �|�:.��X��b����Ӣȭ�y�%�Ec�RO��P$�o{�� GQ����$�T�T�qs�`��|�v�^�gA�U�]��o�������8{�(�⛆�e�3w�//a��텝8�]�x����i�h
4����C�>� �.��i�뉖	Q ��T����)�5�R�z��-'����Ѫu�y����@W`��-(W) %�l�/�'閼�s�(���{5�=���A2C��1�M���#1>&����A���l)\��b��"=��d���o=lu��m�l^ިiX�ӲҿP�v���&浍~�5��æԐqɭ��%�6�y�i�wS�z��F���zc��=�*�����������h�����D�%�֑P~���6F��a�R���Dn��Y��|nh�K���n?h����t����WX4Z�_q�A��$�O6���5�9�TВ�e���#�i,��D�+�E�(����N�v6?���(��y���T�g5@D=/Q��P$_U���Φ�&�z�̈0�	�b�|�MW��d�\-��-�djl���V�@7VO�~4���67�ۘ��O�2tֆ��yM��UQ�7������St��O,��q} ~7]%u��/WM�3�	I`[� �Z,F�}�$�EFB�H�P�8wA��n�_[D��\�/�'��Z&2�ݴ�"w���[^��^~�X+.�*k�go�t�,,/u%��1�ʌU�Q��UB��c��&��H)�Fv�{Λ��It��]���ЇpC�_�vN|���^�7{-̎R�-_sՊRSn!����Ib�7�[jJ����ך���i�<p��'�����m�!�
o�Qx�Α5͇2��bm��
��mx3������*.��u�M�-j�Ak���M�wp =�����ЬB�|�y+���k.vS1D?��=�	����%J�xz\#�b��,i�b���茿�A�F҈ /y�(����Ȫk�ɋO���uQJ�4Ԧ"	�5fߨT
�5������%�xw���^_�<ޑi	$o/�X�ї�wѪ����$�h��4�\޽E )�[ڰ��Ñ ��Fx��,�)�ȇ�hs8����%Ӑ	$)�?�)������W�����<Y������G=�X��L�o	e5u*|�,��8_�T �ϧU�H�V��*G��n+��s����$�ِ��#>�'ɹ��S���*iajY�JM���)�A$N|h�Q�%�؄��x��@5()�;��Y�6N�9�E��4qZ���q�*��0�}�K(�fi��:	�D��K�=�ck���r&�·��9���>���k��g�� N�x2B���{��P�c���� )�����/O���G��x�F%1z'��Ǝ�/�Ŷ�����Ep�ёތ�FR/\���Ĝ^�k;��ݪ�jfm�����ߪ��קɔ������ 7H����^��8�͡�Rb9���,�I�`	�	�ah��O��%f_,-���@�jnjĩG�����{����T�bu�eٜ�iT�J�-�^���9�nb���$?���G�3�U�,�!]��~���&�ʀ��s��m�#BwL?��t�ZĪ�j�ڀYP��DL+ �h��Y���c^%7�,�;C@��~��ߔD�K8V��j����Н�*��9�P�vh�:(9�գ}r��d���
C��(�ޫ�2�*Sҷ�<~�	X�-'����L��as6 q6ׇ���d_u�}�+�k�`��0O��~�%,Օ(=h/^���UVjP���[[���ynj*C�i��Y':>n���U�ܛmlY(�����C���^M!:���C@]1����w��v���l���BT̤ڰ�_��#URȂ9]�,)��iY]`�p�Pp�������D��n$+�x�W�W�-��%}y%;� �i���J��(�~�q����>�ߤf��=��l�	 s����2Kd�l|�ڌ��k�Z��D�F�fS,�\|s�輷Ҳ�/��w��˭F�Z�p�<߰�(H觻�\}/�6S�+�