��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��V�^�Zð5-{=�8p؍� �]I$�/L=���|�+'B�����c�*wZ}z:m��G�WJW�0cYb(+i��{�3%Dp�$=灆#����3�E���5/,�.��F�� �A�u�@�/5OA�E�o7skeEp`��1��a��4�\���_f��|��w��2�3瀨�ul�)Bc�ۣ�.8�a�V���/Fm�(l��b�u�֙�s���u۔���N>�0yD���
���}Iw*6�׽���r���glD��{�v4��q?�K7��-uq�N�Q�t�C+%:���Q[����,Ds�e����ocG���_�5��� �X7@9v����?L�$1�F�0n:d�5�]�5Ӓ*ڻ3�Ӷ��)������w[[�ᬑ"�
���W�������j�ie����8��������j��O?���8���Ҳ��s�򜗩�?E�n���:fm��^����_��`�B|(eԍ`�V)P����<0�[��/��&�Q�Bx Րfb�M[�:i\�C#�ƍ4���k$)���E:�P\N� ��{��6�Rw�����<ג��/��Px.�g\�+�	ΈĖ�cY��y^NM/(�l�~DЏB���NJ>ߑZoNV��<���!���)�< �Zԗ�"� A��kσTZ���O�p|+K�݂��M[c��LE6{���H�L�.ǺqoQM�~�[K~6+D>=y��I�(���'�����(x�DD��S����/�8���\����^ZYf�u�����۸�E�NjM4�x��h� ;�`@-*� �Ɇv��G�H����q$��q�a9W�L����v��4����?T��f�]�,S��G~L����)�?Ml��?�,`��m ����.�m�������ɨ��w�����BB��~��P�/�*t�	�[=�qr�+�+r��uQZ�l$li>k.�{7a�EM��r���	�M�z5#��n����f�H2����@k�@��ŗ�ø�T��S�\=h�wMZu�����m��я�����b��wQ�7����)�TI`. ��v���k@��'�Ɇ_�n�4�%��	��YV[M��&&S����!�n;��:��8&Y�����>���'CQSC��zO��zi{�B��A�i�A���uܢ���X��aʠ��\��`���#'ŲN#/�<�3�s�s��o#�[��s���y~,���H4�Ni�%����gf�t��D��w.5[۬�!ёw�n�,��g����Z���q�XN���Sq����Rm�x���������1*2��3I�7�������*u��٘x^�O}�`T���g�u�26gTƢ3��~1�L�	á��&�u#j����p�.:ފ>
 `����j�c�@��L[��{��b]��QUI��m8(g+��.%}���[g��p3��^��h$��6x'NZ��K��m=f�2r�@s�A��T�g��e��Z�k!��1z��	
c7n6cV�?�~*���BUo�2(S~��{��%�����AyǄ 5#��|�"ؓ���e��ͪ�2MƧ��gx�x�������J;,;.��N��ni�����l��G���gI��񋘎kz�8+�Ѓ����<��v�!F�&�����(Y+��4�2��t������X�#X�g85��""���{��ǆ]�W��O���I�Z^�3Nڀ��w��-�X}���������ML�
l���� ��?�}_����_�U'���$�����-�*-����S)�lI0A�A.�� ���ؠ1|�b��ã��x������U��bֺ��rN�g�4������J?��#�a���Z{�{R��T�US��!�
�V��[|��6K�U�.O�""v���^��>�̎���+F�e={�F�Ҳ������Dw�M�(M�����x�HUP�K�sF�r�����]2��$�{-�x	w`sN�ֳAɕC#^��&�ʨ� ���i�m���9�Cy!�V�����aM"2��g��LO���(�����h
I#|p��s���@�d�9���/�l(�D�1f�a�;D�xNlFm������Yd�\9Ų�*P9ƁVZ�:e���TXP^��<�̤
���	
��B$�ˇ�����2 �̀Eq���W\�o��^5��b%�:�{1���a���7��5���+ȼ�;��8����$rm~jݶ�?�g!�
N�`,��L�e&.\�@f��y
�/=��g�VŤah�U�Eev-V�j�1"\�)��I��
��Y�����G�
��.�%�>�0x�r m~�T�d��:iR.lIt'���y_��\��
���yV�5�5/�&���x�_�6L����q��/T&��3�bG�B{_���)\��ƛf݈��B��4�3�(��j��bh�ل�"���V���Dl�4ި.��y��f?�C���dbusݣ�yN��{�?�!i"hv^�H*�9��z©�,��%3o���;�B��)��#)��%�F��]�N%c*���@(��Hci�2�dn��J�e%Bj��u6����;B[�(�W��$I�3�\$�1g �>wr�L�N�N��w(��]�[�>6b���s[�/�i��-��g.jT�<@�K@ &�	�h�j%�*@�'ﱚ��N��*��^��$=�R�~������F�CBB�h�㒚<c(eԲ�U��E"�x:<�3���C�����Q3�=R�\%s�����^�@�a4�*_��"_;Ga�]C�OԚ��̴JHSg@I�=�D6X+;�4V��x���t�3��t�k�ol��jl%X0\�G6��H��$���|"�ݻ�۪�ֺ�,��������Z�hB&�M����9�r���+�:'Ի:M�;S��G���v�s����U���ݺ
�����J��/��gm!VEnP�$
�-�;*������:�[���,�����S)\�7[�{��N��ªz���=`����G��[�.ZXP+�����\-TW2��RS����n�/�:���a�3���Y��zn0������d~�vܶ�^&U��������T4V� E���ݝ��c�dkd���ݳl&��}����^��S�)F�I~��
�1��!(��.<��b��̄�2Ŵ4X㋫�V$�ʚ[@��&΍?�K��>ʛ�e����6ރYW<%M$�Z�<Î;��bjmi�c�A�Ѐ&[� ��]T-9N�(]�W$��;��T���(67H�|W�Wb���|����7�W�R�~[�O�/�E��pk��T��ޑX��b
��iKlF\@�~�B=�}U=����W2]���%`�^2��k��o:�� �hCآ��oc��h%!#h~5�� Jr��#�AZ3˴����\��!�!�.�׬�ƴ��Q"IL��(�W����({�>�0�O:k��xywPi��Gp���N�z�%0��i�'��D���ˀ�Y�������S?�M�3��
��	nא����j \*���$�~��8�.@��Sx;@���G�w/P`R+�����Ź:p��|�	$^B�˿Iie9HS8��� �����is�}��>t�TgiT�
#���i]���H�����nYX��y�[��a.����!݌//
7 �w��̂r^g��=�fO@_0˼�^�oe��E�$��~�Q�f���{5�/��<�Q�|Љ�(�[���@��`jmT�|q�0͵�&g��Y#�"���$	�ȏ�'�Q'�U�:4�,��V!�/�w�킈T�5�@�G�|�����.�F*L'�;���{K�永n���Sմ?	`y����p6�	���}��-�����y[�Hp�P3Z������X�1�=y��0�^����"\���ĩ^�����A�E��M�pbi��<�Cy��қ�T҉��ih�K_��͸��Ņoa'�����:�q;�%>�80�	9ٖ�d����Q�=��eL�(ٹ��}9�tG�&P����Z��� (n��\)'�����[��� ��+��S�v�)}n���n�hm\�0KI��Yq:.��!L镧����ˬ��c�X�.�U�e����x�t�3��4�c�z�?��i�:�]}��[��FTX���������h��鼗�7�f]������Q�4V�K��&Q%���;W1fn��w��J�ҙ�#ɪ�@<����n���U�8����<6FJ�Z��Z�h�`n!�T_&i����8q4Ϋ���"*mv����b�?���G:|�NpC�������q<�j���JGa�$6�&Ja�J
����Y�t�i5��*|\ނ�ۖ"#�Ev�����w�q�~q7����_��z�L2Iz��K�e�V^[U��0f��aD<*�'���H�mS2H�l��4̹�BD��iΆ�2qSEs�f�}�o�*�����%����,���;q9�"��0�VL�q�V�Y�����\���c`���o6QۇI {q���#���dL/Y�$�E:�C���������-�C[��vj�x�#���<����U�Cހ_+���2�9i�f�K蜡5��y/g�\�%b0�X�)S.�#N�>�k:!�뺇h\�l�
n���K-1UR=NY�;�jr1DM\�gw��Z�����L�w�^�����m^k��]{���G	Q�����3�?o8���Z�uҮb�D��5�M~�ԯ�����>*�2R �R<�|�B�v=�pw $~�I��xl7���X�� l�7���j]�1�.��ǀ'E:[^ѮU�Otatu�9| ~p��e�堚�׿�~ג�#�:P����uVX�I�G�
d�z�c��o�{e�x�8��ޫL��Rk5��`E���+�jh�!BV�R>]���.���6C]��,�4|�"�����ڽ~v�,���+�(�W�
�S��}���3�*83�>�+e��"|�+$@��C����������43n��*�W�Cח�W�ޣT)��?�����HBjQ�V��07��7	�ќ4��w��ܱ�v�?�g�C��g:$z����8R٘�	�Q��6Y�!
�`��@s� �RA�t�7�oV���O�,o�: ��2�W3��4��/�� �E$+��I{6>����.܃�I������Ȑy�9X�&AB8 8���̟�����p�\�y����2�@�1�p��P�<v4X"��ǝd��H 6VM3����8�������b�;b6�>�/���N[C:�� ֺ,2L��ղAN忯�?4�.��F�t�?�$��f��Ie����e����Q����ѹy��Sk	OD`I���/�CSI��dIS�L^�c�ݬ̋[�+��[Ņ��b|gDǽ2��!ۧ�׀yKo�N�ן�
��q
�ŵ���	�U� |L>q!��_ǻ�
h��$�?;�}��U�����>�0�C����5c�s,$�m�}o[�S�v���[WG��U@��s�e���܄�<�(�q��0���i	��H�4WV�sˁg)�||�[���	����=kP�C��mo�ZC��v�Q�*~)������]�J3/��s�ZP����B{r�Hlb��uU�U1�y�3eW�����B��I��B�;=G�5��C��l:���S��fp��_}�*�b��������'�J�a@��k:_�Kk�֋�|�ܻ���
{C��G�Z����N��N Z���Wő@x5_J�G��Q7/��-���m,-���H��-��NGľߒ�;�%����l��/�V�C�+}O�&�C��ݹx�uW��=�>ZV7 ��H${p2*L������t���w D�L�@�7�H5��}�BԪ�H���4��!+���	�`��}eNݥWF凯�ძM�uHj�̓��F�@Ϻ�9d�im�~�.9�ۖ�\���o��P~�㌶��/��fNV�W��%��
��(�m�ު����-���Q��y��N�ˠL>;ecr��Q�T��堇s�]N���8
F�+�S��kX&��R�?�����?�Az��B0v�u����z�N��`���d7#~x+�gG�T�ں���}���0�A`��ԙLN����`���"��S��l��96��@�(~�orB��!�.��r�%�㏚>u�V�[8ZPS�;	HM����6eҴ I1�Oz�G�E��n���g�c���7v�4.Cz3lk:i���R�JG�����W���o��h0P\:�;$� � �	>���էL��P���2�ʯ�-H�����c �������)3�/
q�6�#�-�B6N���G����.�����ʢ�������&t�z�mW�H�˝[�E�v�?���� 'j>������L�����X�|��ú&�C�vQR��@;mԞ�0��P�� ��s�hl#�"~f��/tĖ(��#����z+X���pi�<��X�-8�TZz���H�$A��6�znv���H�u��Pm}ԟ�oډ��<	���׫��{3.��t�K�!$j��o�Ol:��V�H:��
���Pk���J�Nb'}���S���.,��M��Ք23A)�1]}�-2��DH�ax6��tRn��ٵ�Q!/��n�u���X:zxQVMJ��d�M�_������/���S��97����yzM.�#?j��y���r��[�u&�d��fK�^\h�n"�ݫ���VEZ<����Μ��}���)�x����t�y����m�^,��7�"w�o����B�%$Q����*��4~$�o��,�%9�03k�W����Z^ 1q�< к�OCT4�\S�X��y<?LSC��_�z��߀��`��
K�Z�}>pQ�g�nNsk�ٱ"I�Ը�P	U�?�F�_9��)���]J�D�;5�x�Es/*�&P#`-%(����]��{�M�i���_<�ȥ�S�6]��1��� � ��V�^��hy����|�K��4�=o�R��U����4�n�z�{X59p˩�#�
z�e|��NpO;`�Պ;�&�l�	��ہc�������Ɩ侕!�䨹K��l�L$S��o\�G�RÄ����n1��P%Z��C8��#<9E����ŠX�G3�������Cv0���-S�	��?���{n
�#~�|��A�L�L�r�9| ^��e� u�0֒��(�Ҏ�����=��'���X�b��0�X��
+����S��ya%>�������-6�q�(E�I��aΠ������(� �E�խNg�w���Jk�7\O�tH����2]|�^|5�n)�(h.��
��7�4���«��+�-�w㒨' �Z�8o
��b;W�8��.$<:�,�8�6�:6��ﾲ����f���`+uѱn�W�:< Q�H����]��c@�B��03Y��X���H��(��3�r!�&Q��J����6�R�z��'��^ȯ�.�g�g�p�m�p`���gg�ӵB�k��rN��/5�(�:�������ž*�@4��S��=����N0x�O�Yb�f�}+ЀH�hԗ)*�En�{]|$kFL��k�ѫa�B��b��4E~l�v���/��	�Y���q��\�U�8�s$hl{�Ts'��	�ǀ�$�~0%S,����