��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L���"WYj����i� �N�7A!�@<e�]ң�;��5DXL�%�����f�"|���\y�]d4�V���(h��_Ϣqn���RL�/� 8�OK���a�Z����IL܅T?5
�Nx0��Ϳ�7͋)]��2�� ���S-��<�&42OƱ�%�N�H�s��)}��Lo,����;��?��'[\�W_ ���������=��hm@W�)�c[~+�!?�;7�w� �٦d|}���6�
�{��b%Cq�SM�f؉3��
���{�R�mbQ�U���j��l_No�w�0�9�t����d:"�O��;|`�c.^9C��
�6��=6�i��|m�~���sK�r�i���%���ݸ�iD�L/=zT1�V����Qf�A�����;H��Qh?p��3k�ԩ���os�k�����cG�|j�
W%�%6�Z�퓔���鏹��1z\h)(M<s&c�v;��=�*�1�6DiX�H��QM�;���=d�$�������n�3�e(%��+�ʾ�'�P�s{��G]+���.��Xr|�����B��Q	e��$hN���-���ߴoĭeD�\_k_���y����l���A�Nm��@+�c��J*��ׂ����`�>�]�H�Y������BB=A5���ω��C��@6����'�@\:`�{�7���:�5��@� �C��1�Q��&�s�O�[���of� mVڨ�q[����K�̗�>"v-�J!���!{�����I�[C˕��5�ɍ�Ӈ�0Ձ�S^˓�;y&HCȠ� m�{-lV��� �b����ru)������"���>KL]�C�EmЩ) N#e���p,���O�Y�g`���/-�r�^Ǳ�f��N��n�@e����,�;]~ڡ Z����bU�^F;'
 RhE���G&�];��%�8/P^�!�/���Crބ�XH��a��bԘ� "��JT�4�\V�;�D�ǪϤ���Q+.��#�p��!���Hܝ;��6����ʜ��_����1w?�s���D�[�Pmoʮ�_a=�^K#����X��>�i��H4�I��q8G�D�)]�uxj��������9B:�΅�8A���fp$��/I��n�Nh��4UΗ����x.թ����m�7^�;�cW�s]�)�-5D��k��$2��;�� ��?���p��o��i���[��|���I��t�C������(ʃI�n:����߳^�c\$�X���,4��A� ���Ʀ��:;�5��)���1<�1V9MH�L
q�{S���WT�@�d��_]����J��Ĝ�tYd˛-���2 }lnޜn\^�W��d>;�j^b�z蔧Yg���2r��&�0]�t�s��5�����8�b*�R���AM
��8��/CJ��*b[�[�)x��rT]9��lr���GD��)�Kl	;[ѷ�~�Y&uo.l�kQ�%�=�+j���#i~�#NYMti�
	�IІ�+q�r�k��qcω}����,_l)�����jz�]<͙�և�K���4��1�[�7���B�Ϫ���;(���%�ۖ�`��w�旑$Ƚ}c�0�h��]��(|Z�t��Yc������?���Ϟ��m���9�RP`*��H-�����\�RO��#XI��,�]KG���Q�@�l�� a����H�u{�gg��D��P�s�u!ms�I�r�yrs�0[Ӹq�Zﵱe�H�[��?�t����� v��c�K�[��L�N��E��{Y3�h����#lEnc�ı8$�}�r><�xc��_Q����Gy��Gg�J��%�#����`򴿔�֔y���Z���a�[�h��|B�0�J�B��HL�U�%�L��2��\.=Pڰp��ȓ�J����z����R�X%/�l��%���ܴs�_�jT@A�ʌ��a����κ.����/��D/*���}��E�����)�Q��u�\�׉���������L��I`���G� 8�N/��5�|d�;N�m���#�o(o�RA��}g����۱l�B?�p�/�G;���2q�v����]�$��l�!4�C���6� �[%�D�VX]h2z�ˀ�<��o��Ą!� v
s:k���T?�m��Y�I$��G�*�6�U\a_FG�$�Tj�u&63�qPd�%D�w�B���Ǖ,��S|��s4�o�v��r�E@��_�4����ӟ�#>�$�^�c_�iź�|��������#Yu�O�`�������>�l���Ii����Kg[�/���)��^Zz�r�dPN;W�q�v����9�����3P��ád ��h2e��}԰�մ�H�j��R׷L��E�S�|Z����~M�9R��J�Y��u%3
��2đ�4V����_���4�>�.�&KZw�7��΂��<��֌���G3s3޶���h����Q}ӥXu?� Z��s?�d�j��p�Bs�i�E�Cx��R���9_Bn�<�Y�Q�_S�^]��N�a�DZ�sv����l����c]����b�����[	����`��z���b%��W��f��Y�=c����ۇ���" \��t��GCQ�ߖj���Q �������j�����Z����7t����G�*|�B�ޛfv�7�!���0�j���ߦ$-���?.�,bn�9��^������Ǿ+dE1�֤i ��b���� �E��}�gX�CM�9���}�&��&=�L��b�Z!_ُ�&D�ʸ������#%b���䏐߾	����������H$���^�xY]�nA!w=<_W-�%Ut}4#������l���6��	�0��}��`'$�{���7aԩ�}���.F��]t�UCV�*�@�6�:8F�1ؔ�6Jz��B�7\0��{��q��D�����K��|5����yJ ��W{�P�5Ka`�a�.gV��]S� V�ԩ��lH�CQxhD���2t,v�a��ͽ],�w�A��5��"y;��Ua}��!�@��g\�o�L�ϡ��GO'�}Ux�Hp�W�O�sd��@讝�vބ���Ce��o��jyB�w�=��	?��8������"L�:�Dҗ����(?)�Z�w��~��^������zG<�]H��kԁ�Fڀ(�QĬ���1�K��>d���;�n�~��RG@�*�:��F��z��Å�I��7��Z#��=H�� s���g���1�n���j�����ȣ!�6�k����1d_�E�_n@v��Գ&�ZI�$u[�U��ۄ4���w����U�wLȠF��}j~	F��Z��=��'�������'�j.��<���$�o�U!� �"�x�=הٛY��c��2�͡���jv_��[����3��$�.�٦+*����|M��l��8"~�!�l��h:���&��t�� `U�]\��f"����>s4_����d�=��uO���o��.N��Q���-��7e4��֪�á�F���c]U����-�W\�x̱]��o�s6�3nm��$[ ڕ�;7�1�:�Z[��J|gV�g+n�*�A%fHg'Aiv�F��U��w��i��v!��ș�7B:*�����8�I%�."L~[XN�}���[��C�����Y4�ĦL�� ^�SU�~�
�5��=�܎�o�#�N��1MRװ��o�L��q�}�X�.{Y���'~��>Kw�NU�{�ս�߅�1����y�� 	���-�� ���g��g �?��>�|���H�j�g�GzL�VD��=�g�`�m:G:&g��Z�9��P�䰩�-�W�F��d�´!.u����)$R&���u�*M��>�!�̹<b�'W�D�����:�.��00?��.^\A�������E/>�wv;<��!�y;D2�e��t�:�1�ݧ�����QǷ!m"2%�6c��

�7E��n�$ziTN�|��a��m�?�#����c#�M� ����p۫y�-B'��Џ7�ϐ�Q�F�N��O��j�c���p��{��ձ�_2��:��;���a@<��Kk-�dc�
_�z_��S.D��)~���wDC���C�ݘ��W�C0�?�2�	ƻ��^@=���&�}��2�����u}ͩ