��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������"0F��}�h'��8��<���9���-�j����,W�_/�H: 2���x���CH�^�g߹+�F��0�tw:�j��{�)�0��H.�'�[��'0���ck�D����L�Lq�&��IzV�G;]V0~ݭQ�����)�47�gP�ILO�"���tAf�?V��-8�/b������$�9~�
�l])V�"q��&=��b]��[��rL<�\��+��1:����Q_��!>5
9�͖RT���/��Ől��W�f,���th��sC|�o�lԾ���3I�*�)���l�넢�}�����'�x�nM�Y
8SE0����K�!��I�C3m�G]�3�����v���:���fT�~��g�.��\��܉�?+���{�]b�Т��2�`~�U�mԞ���n���7��x�^�p�}���5Ss4�PCCv�˼a�A/�}χѢo`�����	
���6*���9�����7q��|s�I)�����cj�+�ٖ��Xt��4�Ef��v[�`������\���	��K����t�(�!��u���Z�k8QS�aF��L9�g_a�l0c�_N����;��Sԭ��+�����?Ջ|�u�,��C+ަ�&99���\K���&q� ��L���Å
�u�#џ�
�M�U�6v0ǎ�N <�ʒZ�HI^*�KF �h�[mA`/�vk5M[�o�L�0��&<����w��~3���7�<��p}Cjy���<��ą��*s0��"u�Ū�ߨt!	�w��j.`��.ǀNe�HB�rnc���W�=^���hŢ ǁ��ɩ��h�w�� ȶ�gB�,iu�S��;��N!���{�~����[�C����&��x����p����|�6jw�;�ৠ;Ω��h�Ǌ�;����Y=�������;���8b��4q*S���.��OZȒ.ͣ3�)���Clh\�,�껸y���a��R�i�Q{Z�N�6G��w"i�����n��yϮ�!aq��2,���l��;]a3%�VI�W�JS�����3��m[�V�Ȗ�G^+3��!ӿ��	�1��V��!X��a��q�&�z�üOh���Jl߹H��s:O�v����B��d��SVI�q��XO�#�5�|L��=�m~Y�ė];)2w�hM���������	\)�l,��n�<�������pի{�GO�s�Q�'#���)�b�m lC���Y1C��X�RT�w��"��D;�ܡ�� � ?���Բ#�q5� M�����7�0�kM�]��?.{��ӂ�bIଓs�ɴ��
R� $���Ҿ��[Ա���]�0�v7w���뷷C��E��00����KZ�I�F�	���y�ۭ�m�7��R~���5�Vݭ
��ːEa�$7qꂬ�9�,�F��?bJ�t�y�$r�i�M��V�֘;����]e��.Mj���jX���$;�L�z- %�ز*��M����P�+�k�J�2Dq�S]�o�����3^3�J4�%P��BO׫�.׍T���9�W�Cu]j��~��z���O��K�M"\�8�9];(.,I�M0v���U��"�]�$��3{�dhL��#�/������d'�<!A��B�/�K����!nk�|<�X�o$�x��|bM����ȸ�*��f�7��\�wBH_2cO��gX5��
�>$�Rk���������g0C�C�N�i-�WIt��aQg8����K���?hqs7��W+V�60��3���8<� 2<7���̙�LMەy\���0V��0����g,��C���n7�L�?]���,T$�&�֩L��R�ÎE�Z`\��IW�o�����e
�
��q�y���IĶ˂Y*����!9��H4�9�\�CuqAj���:B3����q�R����u�--]b+���"揍�]�O^HA=7����J�n�6�c��~� 'd�:���$���F�ɾ���:m����S	v�Hpvj�!+1��4�a+=��6%5[f�JAR%iH�/Q���+EQ�<�ɍ�K�� ��������l�����[R:��c�n��\7"Sޔ�X���d�?<`�b߯t3�$�_X�G�Sp�M|R�3�O'��\).�|8OJ̽��a�o���vOٿ�T{����~��8X���=��>����F�Օ��o`��~��8��j��5�َ�?�w[iMy=�Ё{ �Ң��nÞ�dT�<P^ �C)�t��A>�E���K�z����7c�'�Z��P��LB����/�Z$_�T���ۡ�J>��P:~�����u�In����`��N�o� ���}jrG�+�?�ق߶L�N��	=��ǭl�Կ�X��6y6+T�(a�x�=ۙ���9� eԃ�bK��%� 6�\����{�D]�A�}�_��f�\�"�I_p�0�%ͮ>��u�|�),���V�~�窘�u�4%�`A�� �V�s1�T��"O0R�4��**{�|4�E!YM�X����ӏ�ޒ�p��tQ7Y����h�ʞ.�Fږ=<��p{e�~pl�oT!�R �����Eb�h�q�5s��r�pj���)��"t+��v9�ބg�Ϥ�*����_�@�В��NgV�S��~}_�W&�y�htJO�mH(ߜ鈷	9�`��z/{'�S��m!z��&'�J�Gn'�f�ؽݪ[D�c^k���=�--:�oo�-�[��z?clK!��t��V��,��I��M܎h�k;,I�F�Q���O��J�.s�8i[�&��\>@��DuT)��Gy�K���ǟD�f���l_�QժjH�����ea'���j��Կ���Gƪ�Z�b�/'GB�<���VK���_�~uP��ү�6}ެm��|o+�=\P�]j±��^Y�����(�x�Ns�����LJhO��Ӓ _����O��dClcm���<Z�>3��uwՃ䟳sK���j	KF�a������m�X5��#\��n0�Br�is�EM��:��B�1�彐gï۰�!��� #��N��OLD��cNvaoCYՎγ$+>�#,�D_��%s�P��i����ڤ�	��d0�`�v9̎1@Թw|�;b�:N�A��RF^�5e�d�8��:�
����L4Ƥ��d�����*fE� A����.�6;e�V&HҌ����ϩ�Wl��F��\-7�P8�O�d�/�v�5VG�-�ns�~���j�.�m��)����@N�SF5��/��~yc�&��a�Kjl<H`*���`Y �ը�(+V��ʴk7:��to}B�|IȨsj�tS�A�Áj����mj�H��x=�3��g#��	�����6��%�A�i?E�K���2-蝹��U�a�is}p�VBM��I\>d��cǙ�W����P��1�62*����3�ؗ��;I����G.'�)�N�	�t�Q'�/�}՘��%q�Z���K�n�,��~��G"Id$b��G�Q���)�Na����̄j]i-�S,t�J�K ����?�M����lC8��N*�?��r����"B?�X8W0�F��YQ��hE&V{ߑR+44bN�CN' ��I ��LF�aO_�̤�6��)�D���`0�"('۪\DL��:i��{�l�
x��Rho�|�����Q�'�������SVt�-1�u�H��FlGK�&�4h�\\*n����w�C�~zJ�5]"J��C!G-3aX�K����#����-�M�չ�TV;��lN��6"���[.�S)A��qr�W��gKk��J�y/�����;'T��H�]���D���P�n�P��*ֈ�ׂ��x��Q�J����0�s��t��Rq��#���������˕�5:�+J���Ѷ����}c]#j�_
Tgߝ�7�q�HdV�f\ V�|��d��<��Y�D
8��j�e��<�(!�eA�β�I����j�ݥL�fB����N���/ʓUs���wiKj,:n�
���3���apsy���ZZ��ֵ��U�� nR�c����[�k��a脳t�Mkxcx�L���"^���)�����z��A�&q�G]���A]��
"�}�V�<���Gw�:{U�6���"�(��]|7'fw����S�̖f ^�'�|�տ~�^�S�oP��$JJEL@ϯ5��C�]�ԏn�٧����T��R.��M/���*���BK@�ڢHN��c��nW�:���@B,׮\�w�Y���Í-&�to���>��⮻�VR���	U����Z�;`�� a����so��U�^EUQ���I�];��}(+����	N�x���-}��'"�0m��]�~u�S�e��|���Oɰ��}�3/w�_h�������]��l�����a��#OV�?����}a\�|nݕ�����Fބ0n�0�$+U���7����%Kk�X
o0�����-g����QN�ނl�ڠ5���I-�Պ�o�-��8<R��%�4�Nگx���g�C�0�k��c�a&�~X���W�dwV5ͦ��Й���޸_g =�t\ݑ���Ԡ2-`���L����0��m�r�)��néd��hO��1t�oafB5=p�(�s^6)���tpe?:u
��&xT��j��Y������u|���y �����]E�m@@_��]�@���m�1Hs�R4���y$ڳ1��["dz�Ch��;I��]u���g����4}�e=����%��
� ձ�oAH���x >d��m���~ys�iK9g5;�u8���4q�E��e��F�k�n���:���rk��94CF肵���{z����B�i��a<T+�[N�וU��G���.#TV�I�Dv:�]����F�Bs�����C ��e�H��dAd�y���#���[���Mc1T�B�kr�q�9ˀ��*�ʼ�4�Fܓ�5�C 08�M|�!�b)�\gn�����It��V� �z�����3���2g�`���g����k>1�ߪ;4ȿf*���
eN�t�Nu�f����$�j��(�x��ֆ��z@����O�r���w���M�u~�cO2YP빓�|�8N��17FpV���u����Q�.�E�:+%tY�m@�}��5Wl�	#���f7 GB��$_�f��-^��1>���ٔ
�^�bÝ��HՍ�2w�3۹z�����X�|m�Z(��0��Ż$�P���Ksb�ùO¾��5�K�ͥPm��Z��3/����9 ^��ƗC8̝$��I��k���T}�����h>W~1�&��n�;(á�@t��=��_�D	j�.p[�8�PV:H���MZ��Ӊ��m{��2=>��_sټ��&���#ȓm��T��G��ɪ<ǈ�O�2���:Bw:'Uy�v="�}�S��C�����u"\�Q��I�Z�-˔H����>p-���z�9)q�+�1t���_h��Z�"/2�{�>���c6��� ��R#1.�&\�<��&>��|ҘM�>WK�M%{)MApg�΀��w��ֲ������/O�0֝���'������������(s���g��sY��0KG�,+���
�lX!D~I�j˞��:��d\���,S&�����{yc�	^`�KX$ع�@_�x���Nq���A�>{�I�f���4�Be�3�a����	?�"f�������gq�#Y�~8��)�3���u��)�@�U��ٌCCk�=5Դ��s�4� k�3S�A�m�
4'~l����jw�.k���4c����z�7���**[Ot�ɳ��Ϡ��>HxG��\�����ov6w��q�:���b�@UcrM�tx���Rm�G��N�ұ2~��3;=}S+��5�U�mJ|�ϭ��( ��8;�;�|����65�g`$,5����[wt8d������o+�S���&x.��d	(�QT>[.9>�הB�~�Ǯ��<��$���wIfQ����pv�I�H�R.��z�]ą���!!���J}�E��+b6��o�$��7&t'ǭ7��7���X|����
f��)�o�����h��Y�Kɛ��I�ȶ�3	˂�v���E�L	%C1fN�{࠿�oaY�Q���d��4����9��t�(�r|\��_�p��逞��?P��՞^+�7��̼T�ӻ�{G�mr7�}��@�4x�u�������d��s��'mŒD������5c������nӐ���=iX?g,�x]X���^�H��b� f�����/����u�d�qi�(�1���fMm��a���㐨�A���-;�8V.�/3Hh�$&w��BS.�)������k��� ,�O���|['�K�}pV�;'e�Fu�4eJB��C��@�{+����39� ��X0�K�T&]i8�A�����+ª��^a�⍜uH}#��;���'q�����-���bX $j�� ���b��ɼM=�����x��<��L�t��}@�	�h��%�v[o�����`Jpk�'v/>n�c���AA���S?����KIC�(h5��wN�t����q�O����*���1��'��e�T�<yqlܵ�eȑ/Y�,M'�(��k��a�yk�'��AҶ�4M�ҧ;NF�.���ݮnEC_M�(;�$�if���Ѝ��/A4",CK�֘O������-m[�{���Z����] AQ�u8�k]�-�)F��!1��ȼ��V�ic�M��4h2�/l���7���
����i��#R�eĻ� P�����x��O��slm�u4X�'��)DE����~T�~6K�g/��.�j��xhT� ���CDx��6KȔ��u+�E§�I����R��A�]��E����k��P{�6�J����;��.��+�N��?V�Nq]��s͓:�oEw��N��aݰ�N�G��fZo��3��_�i�>["-� .���@jv���r�wQ�e^��ǝ͔�a���N��E���H�,�:��Ehވ:=H{سɘ�dk���U�d�l���ds�ऍV��~��3�Tʻ1�E��y�of�LI\�5*kG_��~�󾅛� �_��Zin��Fq>�8�T�g��x�˂��,노��<�5+O���m���u(Fo���y0�G�׊���_A{p#1���	,n�|<	ϖ�5���B��'J����
}#��������&mp��;�f��Ak�������؝4!�)������G:��<5���7�������G�]EI����a9J���Ս#7� ���n�<��D�$���6��{\gٯ{�lJ�hpj(A.9b�B��pR��%�{;M`-�R���9��=-�
e���P�gD�@��t@�る_�{�'��Q[���M��C����J��Z���#ߖmi�m�$��{y�qD�����ԡH9��K<zZ�f2��&]��׭�[D_p|�i�.�?T���٣�M�SH{�� c:ftp���1*zXZ�� �kf����������	u8Xy%��x&d��UE�=A�H�:�L�:~SEd$yw�A4���NU�1��pE0��c�^��m'�N����&αK{�i�X�
1������;J%]�o΁�}OsЫu%D���Y�D���&<�6He�/�n����FP��p�Ig/)�ѡ>�X��֢9(UЮ����+�]V��6����-�}(�+y��AAI�u�#�I��1��i�ށ��t���!�j:]�G@�D�?EQ��7�7�A�z�<"~����$3|гn��`{����)@[��ej�Cc��l<Yv�?�����ಃw�{���>�֑�V������X�R�|��0�nݢ���Bx���נ��&d���~v��Ϫ�q�:��xH�.U9��d��Ix,�#�I-{\Mo+hbg���f����.g�|Q�/�ݺ��r��؈���sAGT�sP���s���Ϸ)x\{������_�Go�E�� %L�3~��y�(׭vķ��e���.6�"�B�ԇ@��9<
�QC���si����k"����p�u����8�O�/��������$�e~�o����M�P�+�tN�p{~��)
�N��+�� �5�C�U�
�꒙��Qv�12K����HV�������h{i��a�f�L�jL�<Ńɾ\ko��q�+�=o�Gצf�̩�eDw�9���oE�9��:����]E�Q��~��iEW�>�*(�D#;�C`�[z��տ����9�gh��&B:�}���9��"�WEU�غO�&��U���W���60����AF������hHE���3����-8f�t��Q`h��X=?:*?�M��<mK�	i�sn�!�S�N�&?��5�p(�����U�l=%�`���Z�pE%x����󐖁r�j<��-߹�@�����꿴�g�`��/aWv�aTa3 �!"L��NM�(2�9K��{���˻X0�n�tY�G�t�޷1Q���F�������[4+���l	z��F�U���j�����k�{�A��S��$Y<"s�\�깞�@c�A�S/�V=:�� �y�%k�N4��V-�-��Wgk֟s�eB�	�"�#����9uu\|E�}���������}�7.-�o�/�e[v��?���O���=���rB߷Vj�UÃ��:m�&Y���9e$�Ϥ`iITdV�@�*�5�Z��8��g5Q��N����՗�l�pG�C�=�٢�Yn��Z�pC,RO��j��_���rT"*>SQ�W�T�F�	$��r���QY����oZh�[p6&I��;{y�R��Z���QIvP?��w��	�����~XU��]��/��5��Q.ʗ�s����H�����5�lou���,9;��|&]����f�y�����ɕ�hTl�|u����o��
K\�z+����k�vgJ_�	�dA��JW}w�zX�}�wӰ{-v��yt�	�����*d�=�\ʌHꧦ*:�E����%�����
UgQ��w��	J�PY����8���s��;��	M�~��1�$���f�gJuw�9��O~��υ��f�5q��!��f���/�	/����N�Q����@e/N/B�j]7⨰G�� Ӑ~�.�ƻ[�(H�.�E��dM_�����D3/h�\N�^~������t�W8��,�B<���?�
�c�A��ƹ� �f��_���6�r�jm��p�����<��Ypv�P��jU0;#��R���:��	+���=�+q�ϻ�һB�$@�>��VI]qǃ�Nf��r��y���#F��G����fkoہ�<]��P���/w�vW_�o�dG$�����{�Ӫ�II�o2ۑ��F ��R4�����ո�A~R"���<K�\#2<DFS�ζ�Z��~k�Qo�]���*dQ7f��.ge���X����v2�R�ö�gr0�镔*���1xZ6Q
F��.����ۄb%��WK�l��5*�m�j�gk�\�K)�" �:�m�h���!����%.czF�n/�07�$���۠�Iup/�6��$~�$���1��_�iЭ��v��c��@�L�4��+�Z�p�aಞRk�#잀�].��f(M�0t7���>�.%'��1����~�������xQOo���g$�j���{{<]�*����E#_F}�$�][{Ԫª�I�-d�v��֒W����p9w�cؿ���ȷ�{�g��/�3�!K��hV����"u0h�Z�ѯe�(� #F�B=Pk�J�/��+s<�4gYМ[{�D̯���Ad�G];nn
�]=ױ^Rڕ�b�H�8d�-�������2�_7�j,�C�{FsǪݜ}^g��
>����u���~�'��	��"�Q_�inHQ�
��R���T��D���6�F�~�+�����I�7-ǃ�v��x-��1�CK�� >B���'¦�r���;8CB}H�Z	�e8x�F�w�y��y�^g�� N$Ws�=���-�.+���7\���O�����$��e<�\z�	�`�@���g�5c���a<� 9�MB�/�[�My��uqi��)}�K�Ez�K�����_S
�ՂG��+�e>s�a#t��	�J�gp]x̋t��O#󉣋	�Y�%3 4����^ݲ�U�9�����Z���uC޺R��$�4�$��'�$rH�t|o<�+*	A���t5f�a�%��r�洲(Ц�py���\(hHD2��P�GlZ^K렛5��$�6*i��_a�n�ߒJ���X��elh'g��:_behN��� [C��	�L���-�̣}��%ǌs'��lQ)NAGM.�E=Ʋ���TW���T<Y���	�!ք2;n��2����U;�;!3��ȚJR�;f���.��{�m�Kc�v�~D��4G=��K?mt\��:?%��5t�/h���2~��)�p�l�:�D��_���YCP������jaH��)�˗�t>򃵗��W�OT����[�\�OD�a�ʀ�M1�Li�|�#V�^i8�2R.}]A�C�)�e�*�\�k�q����	�)��\g�h�j�����,^-�.T�d(���㏽�Ӆ�U���Gx����C�' ��c�K�{&.;�����=BeT"걭jR������܆[ߡ������ap	x:x�ېWؠ�4�������~����z&N�'V���e��NBd�e�`}�K�5`�����wؒ�Ն/-w�8M��+�?��f�;�	,U��i��b�X���`4�	�^/O��׾Md�ك+�.��� o,��Rab����$r���+I.ev�v��͹��mr�4;�*ǚ�Q�.s��1g�*]}l"����
G ��]� 5�: ���`s�U@�*�:گC��˔�Kӯ���9���*�p�r1sܲ�/q[��B��p�NF���3η��_�e-�!S�w��T���/0i7X[�Q/��sn$\(������&�
�}J^��w�2L�6�ZS�g �{X��uy<U���{ݝBpqkC�7�< �7�6B� ~��2��
K
�HЈסoeF�,�Hl�RLv17�x�x�Ç��w�_L��Aq�Guhv�l�=J/�i=8%=���k�D^z�����=!�uo��S�s,R��vM8�G7��ks�Y���t�Db��*g�;-�J w�P�Q�l���K�in��Jˊ��6�ⲵ��{�ߐ8�Z����9�ޙ��F���
!�����/������G���2�׊V�Ö[���..ܱ-�Z1�GD���C�YSV�$�x�J�_�:_X��&Ŧ^��E��?q�)�����pw�;e�V�l�0�p������Js_
4g��/��5�Y,�ѐ�
8����r�`��ð�H���|�����:���6��0�)���ݽ��Oa�OP��3d��m_���Ҭ"��O�0K�r�*
�*��y��ơ���;�����Uy,E�(����&�ܻ=�5��\�Δ߼�[J�	R�
�dk5Uu#�n��Gn<]�xc~I���g+�(�Z_I�N�vR��󘡄�+����"#(���R����%��0:	U93-چ�VX���=mpw���w8���*Tv]�q����/D-���ar���)�}�t��cz�Ymook���� ?T����Mc_�u��'~b�;i��t'<`-z[L^�T��V2�N!-�,���/V�&�cR%�8�|i7Mv��+��˯�J�9����Br���ÊqT�������h��D��VZ9�l�"ޛLq��]��xv�k�(�)�O��\��h|��Z ����1����W�-u���e��k������.dj��ԉ`��C>�k�P��@���ÎV��E�V���E��m"�=��uq�is�l:���z�Cq�+���P<fO�s�Vy{��݃���ҥ��.���C��dX����U�i))����/�kU�0j��pR��	