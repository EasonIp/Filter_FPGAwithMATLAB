��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��We�����9�b�vI�2�ȏ�����
G�Ӱ���L�`/���谙W���?�U3M��,w,a�*= <kG�m@(�I���б�OTc�]A�\�C�/h�>�����\a�1x��M�%��ʼ7���+i�N�.�q���;��m���/\��_2oV<��y彊��\��0e��5�}|�/��uKN��$Ҏ5���ZK��9���A���@��T��K,5�ZK�A�t�w9�Xi��z����!����-�Х���� �R��Ik(����}�����!���l�=���0���i4d��xJ��y�y��+�A��'��"����V�Y�`�<�n�����
�A�5��
���1v�j��?�̊v�)q�_'�n�S�#ݩ��]�蹛b^�U�� �8SZ��M\b��6-|T��x���_��ڴ�a8�$1K��+VSėpc�^o���f���롲�}�J7���FW}�Z��b	�C���z�;v��c�<S�$�V���WV����O�%�?E�]A�4ڣ�̾�Hl�؁��ׅt�5��H��&(�O��;
4V���8&���;�oN�%u��'�ڰ����[�� ��z1���l�$_��>qw�s[-HE3WT?`�|w1�lfi2�Z���1�W��FANPJU��f
��yG��oj��=�M���G���- ��kST� d�D��ԓ��}y�� ^)f�LHuW�����қ,�!�@�yv8+v�)Ez����a�:b{�8U9��	!RY�4jbS��k�+ׇ�����Ď"T��)�����L5��������yd��5�U���~۬���M�Me;�*�LW}��-{ Z&��ǡ�FRa��QT� �I�#5��R"$#���'㻺�� ^�y���Xw��~���jM��Q�Ǘb=P�������(�i��\ؔ���f`�C�ۭ�ͯ�͈�����ب���e�
;��ƪ����|���5SْЇ4�W4uvj�)�J俤��S�7��RЪg���8*��E�3��,_4����O ;z;�\�3<�{�90e��4u�l����[N'�E�C;6��rkm��.����y����Sȫ5̾�!������/5��OOc�]l��~f�m���C�u�}�n;D�TZ�����p>��HW�-L��P~ЩU�B�q%��[]Γ��j��x�s���5��,L��d�����8Qg_���9�Z}��'�g�ҔYj�؟U8g���H��A�y�w��Z�;R���N�ߑ�"�i��&y}��G$��O�vl�XWo9$��< ����6�r_��c�[�}P<�_�N���s:R����K����������_���ir� �sM�؎��X!�/Yt>ץ�o�w���qH{���f�w�~�մx�X�ݒϞ�6�w���S�bQvo"P�6f:X����A�\�B~.`�'�>�o�e5LS^�N���`�ٚ�����>�.$��H��ƍM>�B2] �5 1l�y锃g���W��vM���Kvb��k�j�5]�j��!�k�BU�^��(�~Az����`S���X>����c�x""z�Oq>n��%[��̚9`�I���MG8tgc.�Ds����#*�O��i��ԗ�vr�z��CԈ��h�'�{Y�+Y�|m���A�욉gm��d�r�W��#����\ ��l�u�̡�fg�q�Kv���`dm��;!�^��P���mR��=���H|+�tcQab��}����Z��F�]�s���@Z;�h���a=�8�͏���eze��4ݛ1�-����3��FB�Ȭ�u����P����Y��b`��&�bǹ�m�{��~�3,��_����T�]szXM��1f��#�������=�L�@%ݤu�D ���M����h-[��e�_x�n���% ��&aLq+c�wd�.��圴���+q86cx����2\t�k�vIj�����@�ʏd����9�������J�p5�!����ݐ��h�16tFI�צi9늭��%qb�h%��O��� fP�A^�po�=�Q�?��(d�o]i�jaQ����!�Dw��i�Z��<E���H��r�$�N�0:q3xC�v����[&Vĵ�k����*3V�˟B�ܡb��h��Z�Hi��Y{i�T}�3~Է�M;��2�ќ�X��:I[Vu�3>��}z���H*�C�����E^8\Q�[���>��\L�Q�̯�	@��,��;�.�Js���F>��+���Q
 V��&UJ��!s߈�B�W��<�=9)���4m=-�KL�i�Q{M`�66�#�����tA�������nx���,��T���S�BdG�LS�uH��u�{d � ���B��N���
>�O����&ڋ��2=�Xp+�eg��v�O&��U! j�Vę��Ҏ6�Kp�by�x�ߗ���e���v�>jl@rN
V�ZG2����}��P#����m�uѳ�w�љ�G����#B���Cכ�"&~�RA��Ĉ��{,]��26'D�,Ft�dj�Bd7:Dy�O��H7'x��^(�v�R��K"i�_��5c΄(�`��|��6Cb��»N��|�	�;�2P�V�(*3+�p)�Xs��"��$h��}�j|8>X�H���=�x@V�������xn����\�j���_6'�Q�r�E���[�=�J�b����y�Jd&���>���ap�)�هjB*l��x�֬����>�9R9��'� �k��UC3H:���t	�C�ַ�a�E;����A��Rz=��@`����0o?�D��q���Ee� ���C1��s� ��IE�O��6�����ʋ��qj�z���Yx�w���'�KU7��q��i)ң����~���خœ�%�T^xSVW1*��I���N�_�����X�.��ũa�0��q���"_yJJj�H��v��sKte�:g�@��=T�#*k
�U|x ݇�J(�]��%��'�|��R�1c��N�y ��Fui-�]�--I⣴St�-��q����x�*�G���&��޽,`ݶ��<и�U-֎x�p��\�ZՓ;�7����(����2��$�]���_̳�QdR;�������s!��呭��}�=�K�Gǩg�����3tf�*#pY�^����g
D`�������봨�r��Ǹ�u������$mm�˙NŘ��:A��8f.c/���z�x����'Q�SC�4���=���*Ι�lB�A)مI_%�#gG���@�6�7w��R�;Rϊ~�㤻�ٯ��l����'ቩ^Y�h�������-�l�#���#���x]��ȗ������
O�zf�-w��G�3� jW������W*�N���X�)��"�bB,@�L�����ˏ4pMQX� ����_���J?k��<P4�ga#C�	S��$	���j���^q4�G� sp����o��'�d�5�kTT��`�PN���*H���Y��p$Lu7���:��H��ߩ�F�8�2��E�����^:G�d������eMZ� n#\f�?|�ŉ�v�Zu� 5!>v7yϋ�DRX�� �XP���da��,�x� K���%���T5��r��(|���,���c:z7iG�Q^�wy�A3�6����d5�~�Ɗ�:�1����r�6�Pm�T�߶��4��ʥ�o�[b������$ �E�xs�7��~
")����蓑[Vf��o��dz
lxOj�q:��`\����c�J��s8��az�y%�����? ń#�Q�\�\Qb2k)RV/��3a�h���5�������(�kx��&�!�$ŷa�n�[�W2�d���� ��"#��O\��։y [�7wT<q%��a
�Z����Ƈ�_N���_1Fu��D�ܶ�����qBj�Dړāl�B	�j�H%��*���z6\SЫ��vK��@��3�(�33��n�����~�0�|��*G�N��<]�!�M�6�,X.��|x��R ��(yJ�uJ�Z�9м���2v��.7�9��- *�<����_���lg�~ڑ�E�����"-`$��_P�	I>yU:��G�)�v���� �Ia����4;� `o���۰�r|� +I㤀=�yE�C��<1
D�oJ�Ԧ$|�@�����{\��o�9s���t*�k��Ů��L΄W~俔û$��1�����U��ˤsc�v�-��.��IV�]w!_`�S��F�ҁ0�H�{i�9�䓇�_d�m�n�<����A+L��YՌ\��q����A=�F�������y�J˹z�jJ���0#2�ңy�9�08�z}�z��<T�<!�Z��b��}��)�$�Z����}��r񖭸Q���r� 8���d�ٵe�nT��� [���=ʺ��/�[��`�����Y�\^����1��G�Ep�T�$>
��Ʀ�;�-C`>ڦ`����� �\�/\w��j::J�����~������u�����^����Y�����l�JSnD�rl��v�� �u�'�k~SO�!��#�/]�~'*a���Nwɠ^w��t�ra�����QA$��BK�Q��v˛�;�1.�U�#�ʹv_/�IE(���ȵ�T޴����[* S�Z���r6��\�A:�<��䄷r8�d�!����y���	-C�j=EҞb��Y,8�^�> �E���h��@�[x�N�k��Ռ�hD]&�:�W���\������mD�F�P��zB>d�
��̐8E�jCN����J

$Y�w�+�j����?��Gu#��0QstC���vڎ�%�c�yD<�� �z@c��2;�<]����+vlҀ�&�bR��[r7e�����>z��ٷ���B���r��ǝi	+��5�4�S=D1G�>�b�q�u�Fq�A\���aSz,Q_�,��r-�f��P6m�����؅&��Xf�Rmr�M<[v;��z���g�?G
(U
�<H�`ץ�5�]�����[��
���]����48?x��`��"�b���
\���W>�ū����wn���er���&�?�u!q:w�dz�1���*�0�Xǎkm�"w'?R;���4�4��^ސZ�Cw 9�b_�~�2^�a0x���M�ɂ1P�B�!�R�FE�~?��g�H�KO�Z,f�)��g�pF�]f)�8s;���8�>����(��d�r4n^�0w�B��r$��P�
�%�t����!<r����w�ͅ���s���&��=sn+w�Ωy�#"ݠ܋�5@����O��.��LcYT`��ʈ%b�.3W,�r$�p�Q�ƶ�$����6�9��b�A��Uhv?��wD���~��g�D>�U�-�1�����5��y^�e4_�bT-��#���b�������_��M8�h��W���('U쩏��Y���=���@  ��u��p:XL2�mT��,�w���`�
��Y���okp�J�xD���:��vOõ���^(rt�F�,���~	��r��G [��&���#�>cq�R��贅��� �<B��2���^�t�'c!�2ws�Ϝ��S�]oY�X4%�����.<k�i�8�0��.S�c�� ;F69��D�w���F�{|1�=->��Jp���^b�s|.�r��):]�.>��a�B�3O��1�l}؈�;Թ��n���*��Ʃe���랤QP�.ֹ�ǝ��[��-�aS�N��!�հ�K�b�4H%� ��4�tf��"�C�ŭiau�����(���H)U��ňC� !\�� �K�p���y���,y��L�$.��q6&����!�2Ѱ8;��J��[P�
���t��D���������&�g�1�'Q2�B��S�8�\�p`�{���q�||�*^M����Y�ℙh�*�b�ZĔ��
Ǿ� Uh�C���V<��h۱�$w�����b�)B��&2ZI	XM��G�Ȕ�H+C��fs����۸���������BE�J�/%� �/Dܳ&G���#i��M����v����{d��-��%5�^!m��h�i�1'����i���_�M1zmk�(���>�̤��W�[Uf�p��HY����$ܜ�^�~�)NY�b�Ҵ";��_8�P��Dv�C7���|���n�$6�9�mfaۢF��H#�.��;a�]�J�Zb��g ^iH�4ubl��u%X��8�5��M��1����u��{$�U��5�[��ǂa��Oq)�U�U����ء9���{�y5�Sq�<����~�ڏ8/��5�C��rgl$Y�����DFBś�`�{����y�1�
��G�6x�}t���H�s���J�0���ig�!8�1R:��Q� ��n���a���G/:8�����.����G��gt�Lk��S�����*�+��f�̪�4����H������ç�2l�b��p,%]���a��YsK[���lC���:�n�<�V����l?�^��e�	H�䰓5-�� �_�i@b����ب����<�wW�Bl�#Cb> �!�R�W<�/�`0^R"Ay$w�E���s��ѩ����'�ٛ��?5Gz��o�Y���-�"p��A�\�,��g��f�d�:0�4���,6���}��/ϼ���e�՚^��Mֻ����g�F�`��r�ʃ��r6>Nx�ۡ�+�Cōe�h�1��5��̇O�E�BN��>�2�vpZBN෉�������|a�CLz���/����gc�R�����ύ�e�>4�mڦPʄ�6�o3�����ԧ7����l���Zz��=���C~1w��h��S���gӦ\̹�_�<X�Uo����;F�p�[��:
on�EK���/=��$u;�hD����H8=*���?|`�I���#xy���ό��3�~&���֪��̩��lpTq�'W�9u~7���k� -���YK�O@e��VI��՛g.���|����켒�b�i6R��gމL?֯|R{�H?���^����Q�ݻ��A�w8�bD����y<�{��d��j��T��n)�n���c��Zf�F�gGYV}T���MR�>�Qm8UNr���GJ�\|H�P�ِ�Lyq=�S� �/�����`8��9#��Lفܨ.���c��-y1^���-1��={w�ӳIZ�ʣA��q�G0z�d4XtA�-g�b�5^��1�S���C��S$	x���ʷ�Q���<����
�����ܺ�G"�9���S��������v���*��*C�zo9 ${^s��?���v�붭?����#/|jFK;hA!�q��	��la��"t[�76|�+���z�����D��d�k"��\��4ĳ�����ݪ}����V9��OtDE��<�����ʷ�핅=�&��ؒ� }W�d$խ��Dk_���CYЛj���^��|.��v��ED��߬�s`�9�5�k�n[���N�'"ʋ��Y��݂�G�J���\�]��&l����|/n���b\��^��MH�-F�{�?�F�Iܡ�Ar�zkٴ�|���m�)�&	��1��A���B��� <C�7���t�鰥G���I��exUk��z&wk�A�Qb�n����~�g�1���~؃sqw����������%s'����<$Gh���q9���&��(-�$�"��E���0t�2]=Y�I�t���GKg�D�!��X}Z��c�1�3�J1��Q�7���&CQ��_2z)`Q6P�%S2F��H��kX�X�?�?�\;��E���{?�^���<[Â4[\/荠u�+A<��49��k�X�m�6p�� �+)_#-��c����h��ݞ���t��0�8'�¦"=p�m��_��!���:����C�?c��aN��ut���!!�"
jV���9�Y���N�����|w��a�K����]O[aN�5�#� ��YӞ���q�c���LV���q�P��ʕfv�\��/���՟�}��B�K0wG���{�����P`^X���&(��ti}j�ւ��"����*�[8��O�QOAޭW阔�=��H_���]�G��nSk��!�o&� QA��cdo,t
w�_нᗣ�� .�����N�B��xa��ٶ8�h�!�[Q�r����˹�ݧ���@�"��7�7m(���J�������JhJ*T��j��\�5������n�B�݅�1>��\i����I��$S�ĸ�к-k�u�K��Y�OW������J�k��O;���),�{p�yTݵ��r �p�Y(���-܃��ua�F�C�Zd,k�������]wWB���4��)��k�Yƻ����o���M��qBm*͵۷j'�2E/,�y�n�f`�p���'��z�D����u�g�5����3a���D@p�''�'��#w�;Lҁ?�N�G��q��Yy
�-���\,�#�g>~Q�lKz!�����?:��ڢ���|]c���&�'�������f���G�w� ��/
���2�XX��(ذ|4�M02����/�l'��)d��^64�͛�����F\��<$bmp=��w��i,V�=6B��иې;��	���X{�UV�!��ĞBs`^��-ֹP�g"��\�E�6c�4NGl��������dpg&@�˿�B��_h?F�ۀ��<����b��e���j���e�������r��ۙ��.���y.�u�NQ)��K���V��}�u�U��8t<^�L�E J�r�m��#U�T�Y�i��H�՗&��'i�FI�39q'��û�c�ۘ��@p���1�^�%Eb���(�u��� ΄r?�� ����/�F�?f�"�J^)�S�Ұ�E4m��wǖ�O!@�@���U���p���.T^o����eutF����4_u���=�2l`��J&/���)�	�lZ�#!�����x˽	�ا�=#���<���s�|��EI�-B:/�u�F�� ���:hA`A�j*��A�C'�n�d�ˍ�R�^&��7-��':c_����{��R��sIRki�}��@A.2.XԂ���DT�l�H��$�EY^��#N*9�� έy�_��ɵ�&E+�Xvfv7�j��+�Z�������/��pz)/�-yu�w9@�H��C�YjB������^R���>�uF-ʥ�E��]M�`s��d !��A�uBg��,:�y���Ѣ\�Ъ�r��P��蝉b��#�ٲ�W�ܡ\�<?j�)�yN:���l1��4�"����
�E�eZo�<�,r�HI$	�}
!���"s7���8�Flt��w@~7F��3	Q��<.j�L�<�����r�&)\��~�!���=�|�M��`<�;�ON��k+<m�ʸ�Y/+�������ho�Yz����(1\v ���o�ŘI5�e�Jn�[�c�m���%�}�z�ӯ��1��U�c�E���9
���N
~1ƥ���M�B���E��=ϰ(���ѱ���C��O�6~�	�Tzw�cM�B�~{�Բ����Bl��ň��c��O�h
wa|�\�Z����l��y��+����r�d�V3S��.>�8�;�T|���\N�C>��ɍ��奞cV�'`�6�K�7��z#R�;
$Զ�G�g�~'�r�ARy�{l[�1)2i���.�Q�3{p� ���y��L�ʧ�g���uG���
G8��ƶD�մaPY��m
i7J�k��0B�y�P�C�0�oDB�Oۄ��
��P����҂�S��(ɸ&+ �DG����}�M�ZR��p����r�Æ�hJ������@����uv���׶�m/y�w(�?��h��CW{�%��b�Y�ta(�y��Ytw�H���W�]^���%��#!j�G"uTRv�s�K�d�L�T��|�ؒ�h���yf-A��O�J�UTL��=���w�?*t,���`���09?�Na�L��,�ڝ܄���^��V���"�E�_�н)Ƌ��?g?S�Ћ�=��_k�J��3�T��o
-L����,�$��T�'������q�F�#Ne�.���ޅݦ654�\g�H�$1�BԯLkL'�
d���V�h7z�A_�J~œ6��8>/*�� ��r��q��Sb�&�I���[�rO&�v��	IA���	�J=����b�%��Fr'�C�oj�/o�X���8&��cw����~����t[���T�|S�f�&`��ﺮ������z�z9�Vy.����Ģ@�kFM��+���R�F�������������67ې�8{S.����h�cx�s���A�w������ǖ�Cµ�� �Hfc*7Y�`>�Lb�4i��v����Ed=`��l4FY�P���B�m�?��[�z}r�=u�Q&���En��Bs0؏��0�����X��NqC���rW�z�>���ъJ`O�r���z����,Iև������\@��&)�4��#�i�$
�CcҾ����@2r��16y�Y�4� ��U�ʓ~+|���Z����Vo���e���L��O�����������|��?�]� ��b��0�(��6���ǹ<[�?��i�;�����Z�'5ܒT��(��/4�n���Y/�G����2�3�q����,'�>��go��[0�s[gy����uP���/{f��[m���D*a�i*����66J�E&�������GB_�ǹԪ5*��ץ�������~h���A����l�>�AsB�;8��.J�a�
r��cɎ�"�.ذ͹�Q����.�	�A�/���5C,�` A�F]e0�:Z��Ja��k����C�������O�(.�-��8���ʭ��Ƥ�����>�BN޻�.�10�Ũ*Y/�����b��҉��y�|��&�}-K��u�MD �=�Q�F�����N�����/��W��ŁT�1�;�APW�9.�+����L g8@K�B�{�[.�H(  ���I��(���,b