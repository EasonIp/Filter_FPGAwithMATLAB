��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ۧ[���v=k��J.�b�ԓ���y���Y �g栦O^e��8�����W��}C�͞u�!ēB���sy�,��7�ޡ�nѽ3��.��HI
�8���b
�S ^��y���"E����ڜ�e,ɓ@h�=Kn��+��$�O�&^(?�� f�I���ĝ�+z�CM�г_��A	@��by� =���K��.��Ee/����$�J�bU�i��\�v5�Q,T�TҳW]G������mU�H�gKDV<9.���Mi���.	�uv��ͥk�������|eA��Z�����q�o�=��w2�64�O�<S�g��ޗ�}��A (���/��+�Ҧ�?�b�7��蹳A+~�,Aq0/��0
q�
�5��<��|�Z���B�?ozBA���1Πc�:�lA`���\i_��n�=cm�z	��1���� ����ʸ��ķ1�,bYC)J-[BOA�~��iCu_=}#�� چ��gw&�F�OAO	��=z��<{|���^r+�$�#�*g��aҵ\�O}�{~.?��1��m�7���)Ɂ���WPE�@^����|[��������kG�=d���v��~0u�֫+��H��4|/��Q\]k����@�0P3��`�6;�!�H�c��bz��%���{�V�%�~2¬��M!�(kl��#P�M�y�@���~�]G��z��M!(#�:�kZ!�x��l�l�BVש��`����A�[�(F_��m��"���^�ruUS��#>.�lj�>�J�$@�u�:�qq��%�B��eI��5@w68�и���Lz6���)�>ȩq5��[~�V��9�TK�3A����F�=�5��<bP�T0�|�$>߾�\����ڹ�h�|��]���y�ȝ�Z�j�y~���¸� ͸��.kb�&�9p���4���� ��(��$G^��Rh�S��_���	����q��0��V�-��O�c����60s�p0جF�$�6ѷ�Q��Z"*���"As�OS�����H��v;>����qU�Zp��n�/J@j�����&_�x�:W�א�do��#�������(���V�+qidv��3��·Z��0��� 2Uż��[�^�����m$|��#�}Dm8[aJG_�K~��Ǚ��Q�F���VV�6My
(�����<����h��}��b�\?�sٹO�ނ����T�y������������:W>��-dJ�G��H�ۯ-�8���
!�P(X~L�	��ׂ7�L��/����@
�T0����:�9iN��scT&N�#�m�ț�>�q(���"r�N�}��/�ʛC��4�Smw���u����։Ԑ�UTx�ww͔�9�����6u��sg�[b@�1
f{��Z��M\'R�S��)�ƜL��hvx ���.��Y�c��ԣ���w�z ��(�sT,�p�"ȷ?,��t� ��O3}����d|�G}J�V�4y��:lI�m��9@�t��85�&<y��*WIl��(<bϣl����m�} C@Ԃ���nHϓw�G��?��+ČZ_�M(��Gn��l���֡J����W�M�5��!��un��c�Z�΍�(/�.ª'� �<��Bw��Z��`1���)��S\g�l�!��v� 0�/b��x�Qȭ1��D�cm��%`CD��t&w��|�1�n�nR�Z��\�gH�V����'h����A�3�B)�y�Aj�zf�#��k$��BBv�Pr7܍K��@o�I�Zw��#@�nw�}��3g��M��베,��a��̓�oYe��	��JH�IP;�܉M�$���e"\�V��4�������鋋�A�����Ö㸈���r?U�O�齃��y_�Ē�*�-�{>��g�ZǠ��Q��bI�e%�=���ٌw�{n�r�XQ�Aڀu&+�=/�.��Q�\ȹ������u���1-�"�;D��z%�UgjhBY���!.��D�8�%r��pVM �����x�p�ͻ��o_�
��Z�3��TA���5:�m�7#z�-��d�$��Va~��4q���v*a3��+��ANX�<�ǼU @�����c�;.��e�zF6xf��GC��]/�VZ[��kz��-dvĲ̍�}�nB�4[��Mm���^Ё�LD�Ą���,Q}��L4a� ȱ�tg	~K)�'����n�d@K)ud3O��1�^�J+p,gO�����h����T�]�V�pY!̈́MyX�6
���Ȕ����;u|�MJ�91�Y��n�|����B%1���e�n�M�r���Yu�B�1g�G9�!��C�s&D�l\)��@�>�����. 󆱾۫x;�Z��x)E�y����faC�~>һ�B�B�)��g����������zSL��7��M��nR���Q��kc�o���a�Ry<i��`��̞�L�ee�?�J:�-�����/��f�C!<55��g{��E/��ڶ{m\n�V�/�II��>��G	υ%�jּw���,؋۵Am�[�>�Ȍ9P�X��0I:��]H�b�% �I��v)b`ȝħ��Xʵ1��Mw���N*��1zPg2#��u���ժKR��p�^�ݤDc?��B��6��\��u}zDȔ��2J am�2�li��2QS�5�EH�.^����$B�Aq� �M�&Q��;t)��OaH�p��F��Ū@�4��=�����*'	2n������e�ݦ�{�^�j�/z�}��.�"�2=� �@�t7Hm�Җ�a!q��Ye��1�Ȳ���0��8j��y�3���sD�'4��)0W�lA{l���*3!XM;�"o����iP{�xow@S�M��x�$V�'�|}�{#����'&� �cE���Ra� ��R�En��8N�5/�Rޅ�o,�Y�M����ZM� ����v�ύ<N�"�!ۍ
�)C5~۾�D�rN0�����}������/�Vg38�)[�5L����N����fA4�Md�^�}��
,>o*,Ǔ������3r.�k�0���z�nO8s�I���&N�a��*c�iT����YLlc������h�5�6��Gd�;��k��=\���Z�6�$D���д����u9(�P���'�%
�,�V��mb%	�=�~E9�٧��h]��h�����rK`��J!����5��ۗ�*
��p�K�.8K���2�����;]���"[��͞�%�l�����Hk�FY)���_���OL��I"��ƞ�_c;	H3%)���ɒ�$G�*�-o�9�g(G�h,�S3��I�V?;�&��߾pfW��Ե�v�9Hi"�1{���/r�X��^��/'�(�<���'��7*	J�����3�k���h1���n�W��lQh��(;jb�q`�)R�d95����ŤК�X�Je�#�n����U�]dn���"�V�Yrz&C��/����4��;�q�0� L+��[��2�]��ٚ��R��ud���0�tRz^�~q�Z�x	��ɛ���*�֧��S�<��M��U�uxc�~'E:�����������-bZ ��}�^�O��x�?n�x�DS!-�zz�WB&����o�T�s/��uЂ�3�D�M K���k��
=a���3��}���1���E	=f�B��igQ�y�
+|���В%��/]���Ơou��5��� ��Z���uB�
����%�~����TҸ�2.8YU�#��	��\�Ȑ��c� �F�����A;��h<���e�Y25I�������x��<�,�\tN�Z5���^ߺ8(�q�!=��|�p)B��Qv���7��6������H'��
Aک�{`M����A�gzL������@��.u�"g��a�4�:Ѫ�l�=>��=�#Vk��nf3K��a�9�Ǧ?^�D��X�x�Y��Kf�i�P�8-t|��:�]�ӻ��W�x~r�50��W�fv�9���ྒྷ����<���D��'�-�%�IVM8��D�x��6�(A��A�S���W��`�?�V*P>���|z�!g��)��#�LRے�\)'(EGgE��ڽ%E�D�U$nܴ�SB;���Bk���lr�����T����U�m�d�Q��,�_"}J2b���/��)��mJ]l�t�ZRG��S:v噩2�#�}�Q,EO__dR1�H9�E�fG}�s��Mv�p	&
�C�I�\(����[�]�Mp����
��K\�>�ɊK�����߯c|�|~�@��C�fA/y{�(J��C�ps�e���;�;�=`������he�?�q<�M�mF�F0N��#�~Fᐸ�_y�mc����0�S���N�2����"�D�D���"0��׸��_�0��+�.���a?J�)�W�[
^
�h硧?!,��Dw���C��g�V�kV�|���O[���L�-����X�:.f�|#�h��j�]S��P�זë0��z'�f�OJB��V�n2U�dw�'Bd��9ц�%Y�:�.�3��r�n��	Q���ׄTs;GMޘ�����*�B؆�����qt�t}�h_�r�UUa�$�2%5Ⱥ��N��0�r�M��664=K�3K��a�ݥH&[���%<�-��K��`+5���n����oP�F���LZn�7$�ӆ4՝�B�}�#q�	ɜ
pU+Lb�z�Je/�⍂���g���")��c�o{��O �����Nͱ��Ӣ�:�
�U���g��F�w������<-GFxRr�^���[�roj ۢ�8M����.;��u�����v��	���O�������x �Q_2�ws^�a|�װ%b�KQ����%7�13�k%�%+m�R���,�0�~��A(v�l�'��ޖ���?	e�g��K��h�+5C<|6���ވ�	a�n�4�����*�j����6cD�t:�k뱵ͽ��F:���F���π������c�'>�r�eM��{��B洬��`ۇ�����1n_���Pk���I8Ho�5~1�j|�=��j7��bf���Q;��h*&�p�!Hh7w�]�Zu,#��s�d4��~v�l�'�� ��n��R"G�U9/a����ikOvq\�_� ���"�δV���H�.�І��{�����I���M�&k��A��FE�ve>p��,Z��v�#��l4��Ĕ���M�B_?��֡����0@�q�p��ɑm1V�%�!����/���5%�����?KH'� �G��f�rh�5�S����l���2p�����i~Ձ�i��{��C���(˫��Ĳ�fE��v����N�� ]��+��+�'�q
(ͩG���3hC��Oec��%��؊����x������?Ơ�L�>����	:(��J$#]:č�'��jU�x��ז2�+Sr���gK�� M��H\��ѳ̊���!�X��f�GȞ���������4꣍O�)@���"�N����W��)�޼#�A�OG�Ѵ�!���˓���QA*j������Ä�@I�!���Z���M����5�L�=늁Lu���>hF1XB�QNg�Z	��G�c�0`��0���m?�o�N��5�.�%Ei�T���_�J(�;�a����`O���@Fꐀ���X]������o��!��M���B�,[S������2/�)t���l���KY��������մ�G� e�ՓK�r�!&n�at�QkQ�u����P�ZU��� $�3ۗmV{)c!vm| ����Ԃ�8S�v�j}{N%~cF�Gf�+��I4;�q�+ JR�c`���ʿ>�{֋��ǨK�0��C8���QB�;
�DS��������`5qӱu��p:��(0�� �״��i^0 ��n���Rk�i��1��1���0�L�͗��q����+*�E� .�Y"p��:�<Vs�cT�}y�l���$6��%��e/������H���*�y( �w�s����+�.�:�!=���C�ܟ��>�*�'*pd��9����������P:�N�5�ǇN���nT�ho�@\a��1#��gy�6��|Z`���1�gy�m�'�?�4��{\{G�<���ǋ��V�I68���4Z�� 
�n�9�>�1�Y	�kë��c4�5��2�tŏ\'*��j[�M{K�O�pN����|�1H9��)�o�(@�j$!�f*f�h�ྲྀm4�-%/-����3���jw�`���:��ĺz4��@����!��|}�BN�n�B
�Kv���gqa7���~)ȋ�@�e��TI��Q`���0�	C������bB�������D�tiE��B��F���NH��㡖R�dv��!DH��%��f�s����X���BI74�򻪄�n�2��o�C�RD�e;LC�j�X�3�5��$� ���"��(V̔{�ST5�����*_����g7L��mc<�,A�65Pa]\,z�nTpp}�(ֺXGU���7<�xr1���>R����<.�8�x��)�M������\,w���j�� �$��<��Je���� *����_?z[b��}!����+}	�����E(\�3�`�W�<��A�g��
ֿ��P�1���O�k;��і����=�N�=SP��@4�J�E���$�&�ο�qU��ck��*�j #Ѹ�b2tak_q��䑵R��C^���uz��Y���޺�,�NI�]1���8��g�#��Z��X�J��\*:�^-�xU�a����瀱�F���>͕����O���0r��W�=U����� �^�f���d%z+(4t�9��-�6=�R����}����Y�����!%w��t�e�!���uʆG=��e=}�fCH�"�sY438��S�꧙�i'�+�$��W������
���$^�����.r���kP��CA�8����Oa���P֭���B�����r�?�~�}�C��m-ZH�*�h�PF	.��ݫ��IJ%.c���a�:di��&�b2ג��x�OJ�bZ�p#1��w:���;"0��6J�o�@�L綟��
DÚ�@�~Zo7�)u�/�
��p_jS������^47u�;{���:!�b*x^MXajƬ�����r�
Dw��������μ��� G��e?eo�<kn��.��K�+���U��z���ݥg�ƺ`�Nw�R����@�	~ߨڍzјv�u�tѻjQs�,��,�G�5����cA!Ys#�D��2�dU�pk��C����ݚ���2���9[����g2�Ӫ�<w)��R'˃�#��	 ϿVCF��wv��b�"��B���:�q�:�,��{����/%�����~}:@�s��`�̗M
x{���2��t�ΐ�nPE��r*�J>��ۖ;P�3�ÿ�GlP~�kaE�s"Xw7&+��f�Ny�x�1��~�sݙ�p>�������TK��Hw�I�嶱h�Ɍ&�R��˒�4���z(v%�B:�ׁ3b�ٜ��r �z�g'�1�o����CK! |i���!��U��m>\�?��D�n�w)��>���x�"���Ev�=�߼���?4�*Lֻ��B�U_O��R*��2�$����������\���g��G�e�_�k�y�x��ʆ�(mg���s��{7V��5g�ul���F�V��K��:'�,�ͧ.cƪmb�w�桽au"�z�v����pM����с$t�sOq��;�0����w�������7�x�?'������t�̙f�%��5�2��e�Y.�n:ޓ�i����#hƷu�"QE�y7lv��s
����H�N5��*zq�o�&�%�`��62��Ε��r�4���@ή>������A $5f%�j�[>b��!�̚-�������;�$e�UXFڇFf"��9���XZcd��xhq��>�^��c|tN��,܏N�C����h��w�y%��l��h��0bh� �
ɜku\^�W�}R3ńB'�(Jr%�P}���گ�6���*Rq��~K꺟(s�4Rr�ejm��#�G�%���
��\�_�(�n1Zd������6Q�u�S~g%!�*�R�&8���Ͼf�qA���G'��	���u8D�3l����������9/b�AP����y��I�FP��M',i�1��4�&� �[��i�5p���/�o˿��4�N�5���y�0��MuC���1&��fR]zظ��Μ�.�`W�qB�H��%�q���WI2�5sw�� �K��Q\�v��h�!���'���e	���0�B'�YZ���A�Mi���ݡ�WCF��]+RHz�o�t��'���-3�t�A쏐�1��j�B�=�e�Ɲ3�7v�l��t?z
�W�z��C�2;*Bx� z7�Ҵb��4pwhU��{�0cBM��DsK�M��y��j�SG��_K��[�`�ׯq���}����0F��Xs+��vRle��p*�����v�!�	�T���1dZƏT�B[���e%�rӃ/6V��F-(B��\��R[j�0�6�٦�����r�Y&#��,tjH�b(��t�����.�۔��Ԁ��T�y�q�*�6ٰ`�mY��.L�f�Kq\�/o,kX�/Tm�0�fx�NR}��<x^4�����/�m&%�vKE�C_5_׻��s�E���+Jw��.(|���ab��Ϲ�;��n�I�D=BkhL�%�|v.�|,��1�M�v��C�����!����&�R�QQ<�S�!�F��Z�X��B�u�6�}O��{�y�x�2����ėB��>��vbl\F��� �����|�-/5�]m;�q0�4(6�,�)��BD?�1F�㍂�X9��<.�R][���ٛUn��f�� �pt�u�U/c��c��E�B$`��EL���J4n��Za�W|�&���1[x!�0��򱙇{�	+E��؝��A P�2����)�ct)o'�Υ��{�1f�U�S�d�aa��'/�슭A?3֭�,�r�N���$
�Bjg!2ΊV�V�Wt��y�5�/��~Ws�^}ҩ��/e�����Yv�5D${�k�x{��fUXE�����5��1�i�
`6�ĶQl[yJ�w�Z$��j����g���A Nq.����K��y��H. Qyy�e�-�5HK@�%X�	�
N⬎\F�&�21x`��U!צdP!�J��-է�_�4Cz=[b8�_��^xV����}M�.?�[�����`~�=� ����U�"��YS8n>˗i�Ru=��o�
��Ia��	\���7j��M�j�Fb��@�.����6s�s�8�Ԣ�ES�	7��j�Gm\�(a����)f0{@��Gh[�aH� ����5��9�~��C�-�	��=5Tqz�|�p"��5d�X�͉ꚢ�@����yG�Z�����c|A����c���is]
�!5����Jx���@O�5(�y�@�J�SM6a�$8���F)�������V��;'R�udL�kr�꣄���L9�u������Z[�k@mn�1e"�~6Y�o�!D3�ErsB�A9���hA��	��a`���Mυ�"w�rؒ�F�i����M�I�����d����z����s���W��}�7�s�#�oh��{IY&O��mO�ߥ����,;7+�$$��g2�������w�x2j�1E��Xs��u��Է6���s�Ex,�W�?ymH?%^��AN�0�}�\����}.�2F�j�/��^S���T��J#���Y�pb�s��zvOs�"U�g<�z��O)25j�\y��ۈ���WΪ�D�r��#i-����g`��y��>d��GX�Mw���2E���TB
:��C/߉@��;���8$eє�⷏q ��;1�����v�&� ���J����-�H����J�Œ�MN,���kA)Ⱥ��V��>fB�ft�F,8������e�.���MELއ���%o{�gv�"�F��pR��M��������ss�:�	��������g��H�(>�~��Ejh����;M��Ū��l�F}���ql�y>N2|O�\%{H��)�5�Xq++s���"�)nqM�վƴ:���f2�O]�k,�L�!V�Dvӭ��>B@���� �	�
�V��}�M%��^�>��Z�ۍ�9&����~�y_���
��4���R��D��.]��M�s�זvaA�Ȇ��`��H��g Πnk�'���.���P���~��Z�=�;�52�嬙�|�͆��`��i�o�l]E��	�Jq�O"O��������6-��`�e�S�S4:�a�i��Tl��.�����	��`�b�x2�U5��?�:�.\f3#�v�}&�_Z�=��ꌷ0�T�%%�~'s	4k�lN��],�u��C��w�@>������֒W���v�h!�����]m�!z�3Su5��=]�(Z��+��}e��_+,�QՋ^��Q&N<��t16�Xo���SJӡ�P�����@dK"���:Tnx�����Fo����������rX=L]���%�-�6EnQ	�g�}p�O�i�17V���;8�.�Jjb��a��N�!�zLV8��a�~u�����#:��K&�<�g"H���.�V����g�ۢ����Dq�~�P鿃m�N>Ax���tz���ܥ���=�P����:��ꪉ�4����ѡ�<H���r׫9?0 ?��/�]��[���v@����9�r��^|��f~$��6v&�oF�I*�����~�>1���s�t>0���Ԃ5��d��^*F7Z��\Ģ��G�9�5��H�+����V����%@���x6�r}�.R G`����ڹk�N-��2�t9)?Jz���p3C6�:����21��j��)0��ZV���%&X�p`J���d�M\��^x�����h|M([���Ʈ��
o_�l�q�m���3؊��ye�e��̪�U���3'�F��.Veg!��>KX�.�7���R��!�g��g�L�P�{�6��}ԝ�F��;=���F�F���{|�>)�3����禾��a��U��}��P���5�v��~�G�{:Q.7�h������H�f�W�zF�DR�	7J��C�׏�l-C?�ò{�������`�P��K����6�=��L�n!JNg�lox��O�ݰ�B�dD������aph�!8A�KM\@z���7w����V1w��L��;��Ys�����"O2Y��a?�eR �g�h�I��9���/�ɠ��퐰�����?4��v��0~��/Ȅ���KBn��>��`��/,�h�Ɨ�'�!G�{�A�����S�:�<ÚD�_��}�����`t��p[�:s)����	�]������?��wP+�R _9���Bm�	��=<�-����`: �Co��\��/J����V���6�Cn��R�#�%#o4����i�����Ա�{�I�����꽖�M�� ;���2�Fi�K&�=`�9���	7��桝pG��A�^`-�*I(kb~�P��REd;D���`���V%����m��d��z���#�?����~Id0��$ mZ>��e�j�>��|��C��<���|��R��V3����T�1����'�u<1�y(��;OMnɪ-�#/0 �j�]��I�,�U�����A���g�)�1N�p��}k�c��H�<¥�͡�g"	��4�H�5�s���Q��W�@^5�3���GA���A�f���Wz�$i��3�|�|�a���Da��6{��烒L�?]5��C2s�&4�ׁl������k�ty���zb�W{�OE�h��h�d��Ey�R�#qm�k�S~���f͇�$]��w�
E|��9������6t�g�7���>���W� �5J'MgHH�7��Y��B�����6��I��F�3G��<����_��*��5��!�Yȓ��?aC�XkV�`�0Ӷ*���/��m��5���LA&^Lg589k����^�UH	�9[�$���o���>4K
�)W�"TGy�7�:M	�).	'����?��h'/��ڒt��mb����(lQh�s�< ~�J��������7�'e�1��\���O�s��%0C�j4{������>ws����oxb���Eg�p�L�3E��?�^4��y�K�V�����K!����pX�t���놔ȸG��2i�G�C��bQ�ҷ�:L!}S�sG��б�ɩ���Q��˓�ߑ`i�;�O_:���2Ə7����E���	�s6}�S7�J�#+=Zl;1ǿ�:3��I��5�0qSj2
|�l4VO��k`C��L\�i��Ls��hQ�O��J��Y��a��"1���H<<� ��~����&��0k��4�{BH���,J=�
t��|�3	��q77�L;޳g����3��"�:E�#����HMIٰ��;W�wB�0�s ����sD���/7Q�`ò���Ԥ����0����Ah�3��������zW5�T>�J��y5|�w)��# ��=�=ڂ}=��3��+&�)�þJC�� 2:�E���z�p�E����+����h�6�d�U��|��7��� �g�],��'r�x�@�_}� �/D����K�g<9Q��!,�X�,�u%�:>��=�'cB$B�Z@�;�*�����y�BhK.�J���_�� �0��`o�1Q�[�GMq+�>\]��Ah4��d0"�F�ͥg�� D�I�d8��6��x�x'����`��]����p�g���B"��W��U �O<jh�9��S���
��ay7�a#𠪔�s}�,�?��_�.�z��g��l�j�9&�/�E��$��&>I����a4���S�c�w���L��<���)lC������A]g
3e׻R���uF��K"1�������L �}��z9�>*5��+�p����qm�,���-ٓ���*�U��$.�W���b9��5�k5KS2M�"�Z�`������o��Ug��H��:>�*����r�-h}�f��x�I�\Γ����2p����_ �Oj�o,Q�1�R�(�·�|�:�M���y��.2T��MM�}$�n�Z��d1���7��3!���CP/��cf>�n g/��2�+IC�)Ԝ8׃�-H�.`���L4J����gqL���a0ػ��~
��kq��(���Q���,�������pl7�����hE�Րƍ�Cj�?���iM1��wCv�uAĥ��.b	77EС�szM��ܽi��Ą��ߐRX����R(r����7-R
�V�,F -����#G�%7"�oz�o?9��(?-���|k�j�����!īW5��c�M=E���EK�J�ʔ����H�t��<#-���kDi��_�O��5�W2v��*�`Å �H��!T����.�#䬇[�}æYo��p��~����{6����M� @�;�$�3��� TE��?�;�iz������1��<�I ��a���HP|���
�@^�:&��#hAb#P��2��<
Q��q�H�*;%@�] �kN
"�F��Thf�6)ޕ6���8%ad�U��g;����T���Eq=��f��/��k�P8�p$k4:���B��b�a�2e�!���S!W"ľ4ѳ�c)���8� C^[dF?�˞���8�^�駑��r:9Q5ց�.�J�}�i�7p���Q�7�J3Ĭ�G�o(��}�(3g?�Eİϱ�wt����Ax�{�Bj�2m�i�ÒV8}�M1e^)(D[�ugt��3_�AG]�a�rԩR�Ru�s q����[�Q���aO��y�`�r�GJ���ĘA�o�wt�����������yzR�^s����������n$�55���/_{_�k��zڍeQp�l�_�P'e��=@�K劣+����
ww 
��8w����ͷ����{�=�"]�^=L�'q�W�� �o��G4d��V��Y���U
aX�c�?��@m>����A���'ޝ�a�Q-��X���rɔH2�r�������ɑo���K�:թ�H]�h����OXm���yήX�s�s:�?�!*�y�����e���;���q��=����v�:b�%p���-�Y_z6�[E,��XwE�:��k��)�n���h���1G�b���B�n�G�_	y��) �8
�w4o��� ���Ÿ�0	^�j!\F:ǳ������Y�{d=i���[��ٷ��Dܡ����^7$�N@�O=`7zӨ���{���V+����(�!$�r��W�|:���s<�U�&n���Vϗb\B�'"t1n,�����:�����L�;16�Ɇֲ�Z���܏F6S?ȫ�&(6���kw�'��k�(�矄�g���*�>�J��Ŝ�&@e�4^�u�,�,�>l��"��h��xK��'�T�Ip�J�z./�0�����*�T����l/�寽"*��S@��+�\냫Փ}q�{%�s����M����P
����1q)�!L4�[����HC
@���ڣᝧ/��ӆ���}$nq�$�԰hlu*�@����&�1�G?t��O�//�5֗��7��F��a����hU��C
'Gt�xQ��Rƚ�y�E/̄'j�~��U�ks�o6 �8�Z���g�d�'�3}P��HXv��o�߾��O�h��2��d�W�G�oH��#�M�S��\"�Ծ�QJ� �٠�DD�"cY+��� �r>�Kˏ��`��*'���6���i;y#O'�#��A]�>��(S���n�л���kũ5р��+�$�]�����٢�PI����&������N��3�~ٶ.����,t�h1�gT��ʃ��'�Da\��f�δ:;�)���ť+k3��+��"�BtO-�hT�\z���M;����l;�E�"z;�u�|Q>Ds	���p�%�k
�����ߴ�z�}�j��.h�3��v�Z�g�
�A�?:���P�&����By�9q�> l� �S%T.��C$�t�������N؉��F���}vj�%����E,����PaJ�X�aG,e�	�"'�O��n]���E���;-����h��'����N� `�	�a���ͤu���tJ[4���������;�Q��Km@���Q�EČb�m-�Z&��ڨ�~���Oi��]��C�F	-P|�NUA�#C�s(
�L��$)c��P������E��&"��>yc��O~U�
\[��b����'C�'��A�D<��a�e2��`$���6X>�S������ kXݪ������Ě��A,��v���k������*Y �[w�OV#��S����oz�t��
�`��(Y���7ی�f��KؾOI���7�eO����2��r��R���n�� � <sôܧLt�@-F\b���!�]R��4�|/�ՠoS�Ω��&�.m@�%]ᛕAƗ0��S�jB�ע(�0Q{�Pp�$3�<)W}ɋ��>*����������g럦��>�Њ�h�--��٩[��*��.���n�E�i�����(���Q�d�{ik���M�Hp2\�����*��q-��;E�N:(�.���{Rx�����<w:Z�\���Q1��z�P��㍞hW����<��٭��(wa�{ט>�������}��BrX�S�l�q>ߝ?�/)ӟ�>uy]�D������C۱�#�d���EʌM�hP�^}���E�hI�д��P��W�sX��/W��H���ò��yZڵ�&N	�������eD�[QI�NcD�ɐXC	����o��\���Ft���5MD��猛�eB/Ctw�B�a��.$x��qHX��:Ė�,T"����A?ĽD���������E��~\ؾ"+�4����]t��U��YafH0Q}T���p���J�������qo3 �>����	��WC��w�Y5[���x�u�>2�Vw���=��6,Ϻ)��Ƨ��a0O�9p��0d[h���u�~��M��/X��-�:���Z�vR�d&Pz�j�}���M;�8쥷,�Y���w�[�"�E�i�|�x�ѓ�>0'g���U.�At���)�r�����
_�f1>���|�f8�B�&�h1k�%���a2��'�Fh������
Ps�bl�h��Md�Fƈ���	 ���g8�M�� `�ڱ9��v�ޑ8�'��n���Yc8z>؇}�s���J!G���B%�D���gVnV��-�����o��2�<r�XtTivHޱ]8��[=E���:�@�<{G+�T�o��^;���!��S�������c�/OǾ9��	 z%A�9�X��.��̍���y��ѫF���s#Ξ8�[����(�����8w����ig�r8�9}��I-{�}�V)=���t�pd�ڋ�WmZ����F	�	�G����_�"�|�C��-�JB�V�x�w#��/��^�����S���C��T��b	��x�X��Y��,��c�/��̢�'5��ŠXy��Y�_ޕ���w�2�%��%KǱ���B>
ۈKK��1����M�I��� ���=��Ї�2��(�,��W���L�[j������w�Li5 DcF�Q2ڶ^���b''�g�d�I������F��?R��<�ăj�I��d�x�
h�	�41X��W��~\ȑv.I���gLZX�;��1!�#�S���`�.��W{��+�Z�g���M�F�ʼ��F����&�d����&C����?f��� �/��-g���5٦�Dʶl�j����vA�y�c(�����|$��7������r i�t�'�o�!u��G �r�`y|����(�-{�W k�g�tߕ����=�C�m�ffA-+�߱ժ�E��<iϧ���R���.nU��ܑt�V@����H
���7��q��,n�d��p���#us3s
� �_�tn��?[}����NG���s�N����p7�fC~�6�qB>�04�5.lG	�?�
����D��~Ay�)f�!)�~v��q��� �i�5��|� b},$?q����+Q�+ضN1��r-Q>��Ib�rř5[%��Rt���xi�ikȶS��,[)uES-&Y��y���p�t8k��E24����B�u��C<��@e��W�~nF����=��$��ml)��L�'c򚚗�GO���`E ��웥f�'HBt`A�|�ݝ����T�A%\�����0j�F�<��L�PBr���t�	�p�ؼ����>�/v:��}�0�#�]g�������9B!x�g������&�_#h���l�������s���g><Jl���x����q*��V«1�~�ذ{DdveF�,�'O,����sye՘m�WJ��1�.�� ���=` }� ]�z�c�vGm�'�Y�xn u2m-4�P�%�3#E��֖2y������L���V��ld�YT�w]B�[�֝d�M��j�n�8���g)���`p]HYMP��:�]2�HчhdW�N o|�D򋴽�fǖz�]�D`�WPYh��ڠ�̋Xp�qfp��n��
H�@4D�ȧL��(^��޼��ԝ���{�@���).��m�����a�`�b�(ǩ!~�%{Jl��G7����4=-�4R�֨�\��?2�Lx� `֜�9�a#9�r8����
�]�Hb�Y^ĖdP2�k2-,��E�E�K��w���X�te�MC�RV��}���ᑒv��a��w�s���$�nց���U����Yx{�o)�7X��)%�����2���f���(˓���/:Q�$�͑ݚ$��P��M)�G���!�"p��^�TeLӑ����hC��j��`�D�����{�W�
�Cg*#�!�5-�.M�`��%a(��̖�b�	M�-�h��09��V��9�Ǡ�E��v�Q�/��K�Ks$�v�%>�[*���7��L߄�wwaϸv��r+�70�\G4�frϟ�����,+��fp(���!����r�`DZ���}Jb/��7�|`�w�>w���BML�;��Z,W
$��{�)JK枪�iHa�S��.8�����o��9������F1�&������"�t��Q�+��ɚ��y
�v�O��[�hS���Y�dV�ul�����ѣ��>|DMFR�x����?�y�˖�?N�.�^���Hj���Nln��,L$����e/��:����2����s�F��̇�l�
�
�����*ʪK�&�8��'Ij�c!P"HJ���FѬf��/�����!�OC,^���$�$�BJ {����W	��:�7:�M;:Ѷ c��̪bp�K����Z��{�X���ɴ�gMv ��}�5_�gO� �Ӟ�k%$u ��9��P`&�F��4�X&V���j.�����s?�_OnO���@�y"��~U��6)K)!��������R��pF(w/��:�R�s�/Ţ��xB�U���S�(K�}�P�Vj^�_%���ƲWz�C��دe���;���k�Cw�V(����A�Kڝa���|,o8��K�� ���^ x�E�V֮�i�'���#Ҹ�"�|O pTnfEN=� �����>ݧ9-#���3̎/�z.�S���B�8�
tp�b� �r�ߦ���ʵMi�!2���sE�n'��.{�eA�ޗ��M�p�쇋��
Xee��.�(�+�k<tn��˅�T��+�K�>i�8쪒J�:�U �3wD�U[aNc��&d���n��5]e������I���.��l t��I*��z�L��{��>rj��ޢ����>=���,�Ԗ.(�5�ez��M=�;��h#�/r�aQ��'�p#.DF������8�1��Vvi�fNt��Z��Jm��҄pR�q�oU'K�����J��C�Li�$I��.�L�b�Q�c��ij�祘w���EoP��j��Ѱ�S�G����lV��v�f�W(v�_�W�h�W�l(7����|,?ȭQ�P4��+(U��"m��U_�����6�	����+��wZ�u�0=gL�ث�X�[+���I��8 dXD����Tc��760�2�O5�!sf��0�P�w�BO�a���H������v�䕘�\vPk|��wl����r���{�K*��84p9�5;���FjUi�u��� �!%�]��-�����p��}"i*��R̙:�[Q����j�I��׆��f?��
��*�@����k_3��$�
���=H7��)��k�PDkD�-H��q�������S..��Ę+Q$�q���c��)�O;�5xU6~����Ã���͈G/��t)t;Y�A�m@��� �����f��w�D���̷C�M� ��7o�c2�`ᡂ��9��!c��RR||(4����u,������Yd�OCJ�+�]�"�=�}d��68��}�sP��o�O����k�Z�_���XH���O��Ivg����C�����]=p�1��"�䵼6�%^q��D��0� 92&��En�{s��K���R�7
���gσ��#gP�Zw��;=��Y��+���yEAB��8��CWڊe��T¸�|�i�]6u��%�`�9$�E�̯7۶G���x*�>�l?�����G��'��xJ�6�ߊ�L���E{
�%���D��&��ɑ���ÜKL`f�+��g�+�W:F��z�n�u�����^�&����}e���h�5'V)̱$����X<�KG�Q� g�8;��$����#	T�
&+B�БxH��y�HlMJA���P����G^�7�GG:tд�q0�27��8�����pA)����)��*}����'w��{���]� ��Zh��_m��:�q�x�0SQ�~����r^���	���}8('�D�l^W������n�Y`\
f���bnzQ�A��e�q/�P�a�V&]�I&�߰��7?��h"�c-���kj�������<ēj<I�@�v
�j�����o1�Z6Xy��0W�N�3o׮n�?y�{�e���>ܫ�W/�I�0|�aٲ.D&0k��S������8y=�>Ϧ��E�=Y��>���Oّkm>�S5�D��;�L��M��҉#M
�&�|=�o��Ү(��7bn�m�8�Er6;�����ع&��Z��ބ��h/:ɛ�֦����_�!��+J���2��x �n�<�K��aZ	` �8
9�mb�%��`�|�	'a֧�WL�%n�� Vi�!��L��MЎ��S��P�`;�&�/N�F�ê��:�hH�Yp^v�dt��� /e^���qg�mA�H�	@i4���|���^��Δ���`����5�B��{Pz�Z.��K\�_ǒ�6Z�L��>�N|̾QP��Y�m�h��'���^�	H����H$��{+�6�B��<E4&��k��؈�u���,��H�J����I�!ژl�KR��#~J�,�9_��z�j���=F��9�]3o�u��Ey�a�i�A~��Dp݁$r�3�^��^qd�ԇ+���ƕ��r�y�����cL��Փ���4>)O�p9�Ѧ["�?�ل?�~OUǺ &j��H>�_��x�t�rx,5�a�Z}:�J��A����%���s��_/�"|�:c-0$|�y�Nc#}ߍ�:^��!���`��Ϝ�8�3�{_2D?j��6l��.�� �T���O�%͍���`�ĉ�F<��p���ᯈ�P�[/'�nג�b���X�N\�[�?���N��t�J:W��(���t׶���z�UrSģ�� ���1��o<��K�B��&�q3��Y�(������1Hk�_-��Y�?��0�8���PnR�C�	�kwC�>duLqF�i
!��t����r�C��a`��Z�����:B�K�1d��~�㷷b��b�]���[f��9	�+I�tT0e�3�����<�� �:aϚ�S��z��$�W�c�YDP<�޸�͘`m�[��j�u�rA��4�yK��ơ��J�7�ِ���5�����\?7�9���Ht�d1�BNſ�Ŏ���e��,F=pt
�ugKw��6�V����c-wOVX�<4�� Yv��\��E�(f5���{�6��6|Ј㵦���ൽ��w}�[|��5�Ȼ꧇b�_\�sKo�#Wlm�Y�&�X9�}t�+(��wh*�t�:$(۪�)��ېUlG�ubD�,�xl9����t'�u����Pz�T��*y.w�
�,-H�Ô]79�*�9:k�%�
��%�ɳ�Y��?Нu���[!��(�U�౴��{P�?޻����o�ǀcC�֕������I:��g��z���)׻�:��hxmǜ��.�Ğ�-9Y�)xN ���t��g��u��7�B.�^5I������k��f�@$��}��+�4&���ψĲ0�O�U*1��|%e���"!0{����CcO��K]�,���'L��p��rī}<X����}x�j	�pẻ�(=h ��8q�W::�q7ȳv�q����C���"���r�@ �pc<�E�.	��7F�z���h�9rk^�Cͼ��ؖ[�v��� �Y%w���vj�_�+&L4��vfX��Ҡ&	9TE\S�)׍.��Q"
-�t�;l�P3�ek&a)���_+���jy�R������w���+ڟ��\Z�j$N~CէE����y=Ȟ��b�Ð)u����7�u�<5z'��O��_��K,�.�N��Y��Zy�5����hN�r6OF�2Q`�Y8(�)�azo-~�`B��QCH�ACj�B���k��fY��喱��ޝ�d�b��vLB@��ꊒm=$���L}��8]�xo�}���=���B�7�y�8Ql5D�m�U��U_��E������9��6>�N@=�[�(�19�?��w��*z�e/�tM����`�Z��+%�3~���4A����^�s���t��B%��Q��J`�T���E.�P�r�6&�b�Yz:[}P�ԏv J�����r�d�����M!D�����Y�	�S\�XR%
(Ai)~�BxB�t^�Z��m�7R���|���+kR�r�:O�&V^��w��\,C<�q��^���$���	�	HeDi�p��xk�
�A�a*�V
�3���6t���5S�b>�27}�o�P.�ۦV���K}�&Z2	�k1�xA"�`��nI���?����$��ٲ�c�����Y�T���[���\Թ}����H����⶗����x�z���
7�$gH��o+�B����+h�Y+��Z[u�D	��r:̝*x}��!�^�\.k[0�`\�J�yTR�z�!#��,-��B��?;�%Sy��"y���v�L<����u� S�7<V�({��*k�q�BŮ6P��=t�I��D��U��uH��z)�������ztw#M�㩵��	"�ɲ��U��$W� ?�;�WOAU�;V���
�3Х0�p��0�"�"��m�gY���f��^�L�kk�W
댆��(�6���H���B���5q��T��-hǘ���D4=�h��8M��p�w,��\��Z�t�x�#�ݰ1f����ʆ��#G���t�݊�k���y6`"ط�\����4�`�O�-a��K̽dC��>��d���e��Kxa�����QRi>|�����!�H')(����:���w�{�� �N^��N�������NJ�i�goNN�i!�-8�:���`��>Q7����,3�Y*�@K0���~��WQMŜ��U�|{خ�n���x{>�d��H[_v��R��r&��[Y@�}M��3F/QJ<��熌���x�o���*�Ʌ��Ro���=�E�N3De/�π;�w9g��?��VFN�y1�J@۹lVk���-��G�F��%�Y�ל�Ҡ�$�8DRL ���s��� �-�Y�;1�HX�5�-�V�e��<ǻ���6?����'.�M���S?�9�O97�v��Z�`�֙���5��:H�t|>)X�x�u?�dl�A��V[RIo6exPv(^�1c�Wr	����s+c/ս���1r9e"��=cr���]��]���rFL��{�z����d�lg��b��/6~�䜰<��V��&�k˰2"��ˀ� ��݋K���6~jqz�$_� s�,Orб�/��c�FO|�m�3��LsN+�m�MG�EMK�hq��(�?lm:K�w�	yJ<�{.V��z��SOY���&����l���U��/eф�	N��=��dK&�2ViL����m�bE�!U��s��g�d���k��o]�4�s�զ���u<�������GX������k�L���5���^�"ۦڏ�w���wb�E����ɝC�9Qg{E-���s1��K��Bl��U���:9��S�~�$��%�г���n��]
B�-�A�F-/7�m&�x��ؚ�n*d�Z�	�����6�\&�e�3����K�f(�ʊݻ�eL��@���^2�ؘ� �ll�2ĥ���]���_/4�-�fɘ�A��6�,P�^g�E�Rg: �	��ґ�F�2��ܸKKp��U���D�Ē�r�?���N�����ՁCTMc�sk>D�#a����JO�9h7�UM| K��OG��@��A���7�j)�c_��Z|	M��c)'2=;�����7�������g?�ZO��o�3E�\9���*�*ג�.�U�kaE��J?xdI��S3	����"5�o�@-(7V�DS^� T�J�ȢNЁ$���O{A�N$�-8��Y��֝!	���C�~h�h�����l�xS������+�_��t��}y�]$'����Ov�Qϙc�VN��|Y��
^Bn���'��F�؍D���MX ���Y�	2��m��\#��ܥ���p�Jf�e���|�^IZ��\Vc���]�d�u��5���h�v�=���I8��ֵ&���\e/�%��ׯYSt�B�d���"�}hɴ�r���fU#�I��Z��D'!���. ��kk�eX��'^�9��q�3����jz�Ӆ�lf�G� FCY��T'�b�&!S��5�C$}���n����&}�n��bu~���W��&�2��a��ƺ����׳��L�S���Dx��͆;�#6b����q�9N�o�dA�l�;h�`����~A�p���AV2�ORk�2���^��|�6�Qt��IwFa�8N���s�I�:����:o��Y��t뼁}�!��bYarqc9�lZ�c��8E�c��Z�oO�%��*+-(仩�Ҕ�i�I} ;	xvIW�߅ɽ�$�{ـ�ѱ����)1�M��q�g�|h�y��� QB8v2��J^.,���K��Vr�\CS�:M���y
��1*Hz��V>�;��G���:��������h�\�?0]�ع�$�e>��l͵�?�_��<N=�\C)����ǫ������_&��?��6:�2o�PKZ���3S��f{����.�#!D!��*��Y�l`���\��y�EVxaX�˻�os$d���"0�����B0�3�w�݂��H��蕞����I��� ��JYN��~�~�m�*�r�k��t��@��F�z�]�� ��Ӵ�lJ��R?�c�T��/�x�nTѳ[��� w�:����&��'~/�����O�����q�M��]?��?���-��qt�Z�A�CX��G�Rc�6a�E{��K92����ݏ� ���Iɭ�]��k
�w�Ne�����4Y�f�k�#��˖�����A:z�|����XS�+v���oہ���n7�Hp����>�d4��x��ֱ�Q�<�VD�̧M�fUV�^uC�$x=�,wPBF|���\U�k7-եͅ����	�]�@@�w����]@~�/h�:��PԽ�{a�^𻍯�����%)�S�o�3���� a��d�+OfyW*�shó��1�hQ�V\�h����t0!&�u��H�VD�x�|�vMb��zO�,����(?����W�&�0�2�^C��K�[\K*��)�Uv�-�k�/ЅM��X���A����Qy���u�,{�+ӅÑ� ���'D}\�;N�$�wYAlf�#,��߆��&����r�C3�]��G!���=�4��`�4I�Ȓ�1��Sa�u�+<�U H�L�H%��c�t����C򥫃����0^6@ �TЇ2a��!�:^����&~s�.���9���H�Ɗ��7|g��d���:���9+��5..������Q'�)�[����ųLce7�2�}���@����z����d�~֎�?͔�j*2MDMe9�}��E�������l������<�副
�_����N�@��x�J���b��^"�,��dA�Ez�U�o��b��/vV��<`���&>*o��\�(~�r���7J���=Z3��r;����DR2`J�z�������\ܶ�_jj%�f���|��U��6�2�p<�0�y��u�J|v�K�_>�i����R9���l�c� �V㱁�{i���>kC�����o��Q�[�!������]҅u�h�|qu��Rg}h���H��:�:���N�1�Ol�^Ĩ��&���,=3ʦ��t�3��5�&�כ��O�k �o�W6�.�.(4�U,.Q����we��5[�)��b6_�I��	���&82�{�t������fQ{�*^,����#��W��{���.R��I����;Z�^�jg�	9��=�߻�<PHrx����>N�ٕ�����m!Ւh�!�tU����@8�7���2��,�D4Y��a��[�Dr�k�` 5���7.P����Ӄ >tyb�յ���488�g�I5�)�`a��5��"�
��]�9y� ֲ���Y^#]�Ge�SS"���`kNљ�SZ�x��#J��Q���P'�� ^�LQ��E�	�Bp|��CVò �����!��n��*L.,�>T�/�5 �nr^��4c|SB�Z�)S�#��Ղ���������&�4t_G�(h�GI|-O����~K�v�VgV%�gΊq�0��00SMI�Z;D2u� ��z��*�V�uQ4n�c���i����t���G'�~�]�su�rS�}��Qq$���"U����G<�i;20K��'�K|m�ݟ��5b��$o�{	V��F1H_6o���'_�WG���^��w(��!�����J$6�X��m"�/c���%0�Q�(�d�n�.�<��#y�T�DRl�}�r�d
��������-�HDK�`�`�7����,�!\â�<�3RO�N���uIMKU�+�=���!���.���a������*F�:X�hȄ��i<U�6�Gr̈J9��B��mC6�j���1��O����!<����3���]��(��Q8�{
�:a~P?���4bG����3=A�����N;a�q�i��\��v&���`�`c�;%�0ƭ[U=+���X]�7�"s7�-GJ?�"}���w��xa��E�p�$���3#w�y��q�+[D�,*oP�����ҁ(`�;Ѽ7�L���u����'4��ئ��x���^K��9����*Q��ΰȊ�JF8�r�*��A�Xt���"�(�A:�N�T���B���xTe2���J���O��~	 ��<�~��m�f0�j�#�9��Z�3�c�����i��Nr���"�.��˕��A���QJ �-����0�R������ٟ��M;�<��¯�ő�9�Q�֖����6�®�e�@���]��}�G��2�'꘮�4r�f�]JR�����B{\�Fk�lzE�!�78}fvU�pcã��jك���ӼeJ�<Z��wvh˾�u�����%�d 9��쨟<�fbG��������ݓX�v�9KH�a�y��Y?���IwvY�s~��]��l]Q�M�/W�?��������HG3#w��rZ�C��G �����="2�r��U�����?����Wp
8	�����EDz�J3�n�寂�<�u�{l,�N��.͊|ڎNb!���Jf�0$����W+��#:<`٥L��Q1,��<;�: �P�/>w� �|�`Y�����wr1h��#�wGI� �CY�X�Bs<�s��no��qCO����x�XO'H��}�m�6�;�֋qeg���QGP�P ��Q�� /�td?L�S��x=o�/R��a�Z�¤�*�[M����oSs�X��)q,��S��YOT��`����m�$�A��_���q���9m7�]��'�Eg��~(/��S��seE?k��f��pz���Fj]X�{�
��e}!�é�M��m@2�r�+��4n�䙝M���E� ���a�=|����]*'v��<���!&���9
�<����{�6 ��@������VR�������+~���u�)��sO4�KV��{�3�
�xDg7��el���*�k���:�����B\hS,�V�/���uq����;�����c�R$�;U��D�@Ǜ�sb8���]@�X ��V	�_7)6���(�m�5ďh���@���c�@h�O�����@R9W���`�[�}�� пV�a�'��b%D�x��2Y�OR�oB�{ٺ5�3r]��A��y���3(PC��]�"r}��g�+��!��$��}x�j�«�z?��
!��ǫ.T���g�e�3Dב%۪6K�4��-��� 1H�f��No�L!�+��io�5vm�����||��{�ðM{jީD�<�Bc2&k�	j���"|��Eڝ`<Ď�Ⱔ�!2Q>�kdo
�� D�6׭�����R�!gHP#��.,��������b~��ZZ��j��'pH���l<��䍊;Fϣ���Ԧ�w9�ש"�V�ׇ�ID"M��f�L�����:�[
݇��`�)E�������7v݌bf*d��Z�b�a~}Y�^��T���W�?��"8�4h�J(���+����HݹuD�tč�!����g�@)�y%��a���%��2�oZz���JH������H��1 ���>��DC���[Σ��@,�{"������2�8s�����q��!-��>%ɞm���ߩdՉ�ߣ�y��������`SIU��UA[S���D��o{j���@��Jx�o��Փ�����0�i��VND�WS��|�s�E�t�p���+����#�5���$7�5��	fKˮ>{�W	��hd���U�h���<�q�,�j�CB�<�����n��d����Vg��y����h��%^LДd�Ѿ��t�S��vB(���ZU/�K�{�Vq�Ǝ�Jۃ�Ul�f�i�&W�EK�W��8���(�Ȧ�"݉��z��R&�u�� A#��ֶ^���i7MQd(�p� �.�lQ?��7�ͬ@�� ���@an�.	�}����f���7ؼ����WM��Z�x�,X7���Q ���8)����
����+,9�7{�w�C߯ �HS����ҳ�V�3?Ȅ\Bε����їKGqDs�+r�ۼ������ O>�(A?��	M%*]�7��cJo��]X���&�d���K��೶�n�D��P����F�-��R��s�%̚���b��*�x����~��V���=�z��M R	�Hy�|p?����T٥r�Q'�m/=�+�A����wR֎ȑ���6�[]�lj��<���Ҹ����_L�=�Z@�v���1U)M��]��kV<-���Qݘ�J�}��zZ:=$�����i���D�Yo�:ʯ�Jsx�w\��l)�³�^���Ҵ�$�-� ةѱ�8V�|������� ���7�Z�m+ʵx�2P\Y��,y@h���Q��m�F+}_���������O�o�b��R2�|N2�g��1ӂ�1�j���	���[�#����)�Յ3�\��M���Z8����O��M��?v>����*rŊ�ɭG(ݾ�w��}l�B9����m������L�qg��0�M��_�)�I����	&:���&��܅�P�` ���j�]�������{��Z8+��J�)�ce�4lx����t�M?w�0���/+�+��������Q�4)�ϛ� �;MD1;_jE�HV�9��>�H�����vDVl*+��*y�)�$y�8,d�L�`G;���ҏy���P�)\������Y�LW���-۩�hl��u��$�ք_o�ԗ_���6���P��d�;7�e�M�<80�U���G�h����^|	�ә)L�"ߏ+�Ng4�0��n�AҸ�B��(��b���lt�8�����BZ
�{�=KC�9���׀�F;,���Ru�H���\)F����%�5"͂`�`i32�a4���<k��wnd/S�#���Np�͂�Y�xqy
5�F7�
7G2`�D;9=��Gb�#��
c�4�e�j
����{��@	ʷ0��\(���e��	f	i��Dl��4�3�+W��?�����Z�𝼫��ٿ��)s���i�M)#~��?�9,yF� (�5(�����\�LI
�1��Q1��٫�m��o�c~h��D�cg�6�e�ȂV���-F�B�A��� ��[RP�մ� %?`��ąW?Q(�ϥ�	/X��Ju�ۙD^^%-D��Z8���'��<��naO�Z�ے,�:G���:�P�QՏ�J�s��.�~�i���U�y�Vd�\���@��wh���Ry ��>�-�>��O)
q�ڐ���E�z�n6]�TWޢ�XCG�(����b�\���x������C>͡17�SH��:4V#Ōp�f�RV��w[8��g� r�-c�B��5z!�O�r����c��/�V�N	{e��G�dvx�����z�=��kXC�x� ,�Z�m��ɣ�5i_��՝���`�g��Z��]RYp4�
�e8�Q�j���'>�0U|m�0_]R�TYMI���@j,�# Q`Aȯ�ȂzFR�U��N�\�F���n�6~�lb�ߟ罒�=A���o�j��O_�"G�rӋT�G~����a��Y
䣅��o�;�����M^��/f���cKގـ/���ogN����R^�OgY�;��M���Q[
[�g��L�D�HI��m�b�bV�0�	�DP�s�~&�vl>�y��$O�1B�y�܁	�Ҡ�vJ��r�z�^[C6�!�d%��*�Z-m��n�/���x:��������S�x�N���+H�6��N���t����-�����|��ց����"��Xs��7�����VQz�T�U/�F���J[Q���2A�/��FLO~q�?�H�D&�����}�-������OO����?�^=����K�����L0�t$�ziszc!UG
�Z�	�f��I!r1��=A����#�!�	�~_H�@�3�!��耴���'�y��+vj��H��R-�`��-����[�yCO����xf��-�Ɠ{��Iri��K��AD�u����';^�j��9#��=��8�*��t*�qؠl^�	��:��~%����"W���rRx]��.Q��h��}ˆ�D���2p����k���4y<N-�	P����N�x_;hg~���{�K\���BTi&	�[��&��he�q�(/4
���[��7�i5�}��D�\�M氉�J���#�钐vjY��>����Ls���o-� �����yC�9_tM�,{i�0��߫C�^�/��yS����L)��-L�AZB^-UKh�WM�^}�u$jR7�s���wF6�$L���aW����A(������Bh�!*4�m8b�:��KA��A�����w�sE;1>e�؜y�IĎ-ܢ���{�����gx�v���G�OW\����C����O��3�B���1j�"�Լ��"�M5�t��돹�>tUX�+��>ɶz;Eu[���K�;�zm�̣-���y��#���\����)�H0
��O�l�>*u�e#WZm��C웘2��@[�������<i��eyA�	,mh\[�HAI QJhUq�M�ܸ|��T#����ƸT���꺂��W ;�ER�A���d$��)�n��1x�-�T�#9p	lX"?�JE�KF�6���D��� �aR�:	�zo �4��l��"-������������tuN�&8�O�/e�.��lG��?\7aB�<"�.�}O�[�[~���l8@���r���!�v��2�5;�F)����`��;�?��~C��ֻՕU�U��}�^�n�-(����hZt���H�� �Ԡ��*���DXO9�ZҊ��IR�m.����m2��9����o�����Y��|��>Y��(��R�R�Z����Ύ����F��q�p[�?�%�$w�h��rd8�ط���+wm�<A/[ZZ8��yN�b�m* =D�X@����1@�ςevgqQ��(�L*�c���4�t��0�Kj����j{�$G�â��F�Ӝ�8�D{�'E��Q�ו.��Z�sB̖BT�_���&͹��p�.|�J	8X�"��D�f�y��_c�8���o�����O70v�V�az���������
������*��.>���Կ^�7�g)�2U��
=1������L���%⩔����/�)�	թϜ�F�>�x�)�!��8|�/eAۙL�W���t��!�K��طY��vuEyR�.�tf.7���.t�{��F
�����>�/���nnh9���!�]��|�v`�F�d���]k��V����\�!���}��:����$=����911�A��+��_$X�9\�ʔ�+�͏���Mx��BE�0�J�5�w�@��K��$�:`�x���dd��ը��%DPP����":g�] n�éߴp� ��N~("�����DJ�3+{V�.�%SZ�Y
�Y�tC��A�����e׋e{k�R�G1�oQ8+/(:j q���o�;H�=�6��}vG�j�ǹpuPk���!�i�I�����N�&`1=�����Z-�j��O�/f8	e�:Dй�f�(lxj����X:�/��f���c�Z��>��k[��m�p�]c�y��=Ǯ�̵`�بy+^#�8$�[�r`�WX�F��V6�J��P��g�F�mI���~Ou�z���� ��#�a] :ej���rs�Lm�� ŷ����'�	�f�%=���e6�48��}�'9�wQY��<Ni������%�$��˔B�3�6=�Hj���^��	���_Z��7^Bh�2d-�%>�|1�5aK�5���N� 	l�ƃU�:o�Q����&��� 8t�.�:�/ꚳAm���z$y ���פT�����@�P���_2�X��>�\���<���f�ӂn�z=�2��D���Pbp�u����"�"k��	�3�a�i�^L-�H|(v�F�� ��-�`j�����C���0�5�IL{�1r$����0�Î����1��:<I:�(���u:�c�{W��y���߮/���}���4�IL�7񯑜���ʰ����C�s�K�\i_a#c:.#:�����nL��P����G� ��Bf���Zg�y{-o)��%���tET�]/?uJ���J���J�o�2V�=�n��PÍ�\Ҫ�[_��]>|>jv��*gsN`D��ʤ`?͆�i�] �2��}B���,��}�Mk����6g�n!V޳R��SByb9�v�����3v
4iI�xh��L~S?�57��:R�����_�i�_ ��W[%[m �Y�N�P!�e'8�.�p\�Lz�����yWLE�?�>R����-����DY͕aL���-��qז�P���U���Xwu���e���Rf����E�Aq��~1W�Xf�4�gT������������ԃ׻㴰1c�����H�:S'�����+��^N�lw��(���Be�u>���B��ʽ�.�jS��[>���K�I*����(��ݾD�F�?f��_p
E{����?
�k 2Z@W��]x���8�.������|�rKC�77-8�\[��KZ�4�`��0�,b)�r7�@��%�I�,���քMn/�֧H���Dۗ���p)�|+bi�0�������A&����imHB	��;��&o'���R��}V��r�*L�y��)�a~��!'ʹ��4P-=+�+�,�a�;�ܣ�'P�R�d(�����C8�r���z�,��W�����85AZr��R���m0vc��Z�鴪~�J0,Bw��*�.�.�K����'��� 0`>���i1j�+���2�fc���ٮ��'�7Gȩ����Iƽ�c��r]U�`-z�� 3���γ���*��	ݓ��V����$���,_$␎�n%>��E�}���Z�oW�3f��� �z���җ��/�.���~�����I��P�g���~/���ί-'�!.VOkV��<\���;ɞ�_���+�y����6���/��,�D������`��u�J?��!������*lk
��|���q��L����K���)8�9ڂ����S��:d�߱��޾�Hy*������i]��z0�H��C�y�:
��6nd���ﮕXm��-��i���qC��oS�v����r�I)��A��؝[�O��y��1وC)9rP��a��� 6�>��@���ў5+�g���>wN�DJ�6��ǐ2��h���|R�]VT=  ��p|xmA,JFS�۹4s��=��|�4Y�+�e�w*_jMH=�E��o1���h�!�u.e�S��!���6�x&�Ԭ�*`?�r��)�,����}�뿲?t(�V���µ�y��w��;��?�~�zEDR�W�L�_����ݷ���bp�MS�u�C�4����'�K,{�al~E$�ޜ��2Fw��^Z��(Tז���3^.D�'ƩX$�٣OP��v�Cy��HBT��Gv�X���T�i�H|&mOI�ש+}�m� qģ��LO�7G���`z�i��ϧT��4#w�"0�<$�,:Q=rɚ���)���:���[��\�	�<����0�-"������z�q�����r�y��Tbr<0Lshjޔ5��*���{>ѻ�߈Aj>�濶�Ӏn7��C��������K�)��]�TM}�K��%v�k�/�E��4��Bj���Nа���7��20�¸hQZS����wvGA�f��wv$;T���� 0���8�Y˫!s�e'�EH����$b�Đ�H�=�g���;�]�5�I�ǒ�?^&�_�|@>��N�h�%��q{L�n�m,�T���Ga�g����@���&�ܐrV�߸�c���Kԣl����젬�ω�������;r�!N��H�_��i��	ª}1M�^����N�H�p���BU�K/i^d���vt�]�2�س���)N�����A��8.�����<��(}i�G���j��"^i<���|��[%:��i۸����'����Vl@nN��{�hٯ��G��њ�q�w��x�����^-�p�̖��j�aʪ۬\^�mR�&c֧�r�a�1x�޾d��g;�.\����ޏ�i^��d���)͂;R�S�㘫F��@�Lfu���f�'��Ӿi6*k]�W��n�Cx�2����<;�Ց�&t{&�� N��$
��?�i������Q�a<�$�+�1�a������R:j�Td�^�����@�ģ4"`�i�	��O���C�qK�L�q�~T��2���6.Xd�UÏ,�ϵa_�Pq���H��PzI�����{��n�pq�>���@���XsN�s��y,��B�����J���B�)ZVCC*?��BO��f���j�`P`7\����'v�j;��d�x���;��=-����$;*��6]���p(̞h��q�'��%�ι�겊Ѹ���N�κvF:Y�l�F�00:*5���䶇���}A��]Uߖ�P��}�xR�"%�N���U�qbbF�_h�����p�-�^��>���O=���<�3��O��5zr��̈́f��,�_M%����E�ڔ8>/~�BC�	c��\���K���=�j�v�V��	jקV[(j���)%��6�X�7����)��V���[W�I�����b�.U��'�!���a�М2F�Ձ���N0�TR�Sp�Γ�۪��/S�$�E�Rdbcu��M��f;|ICT�.�>�>j���&#������G\0����(_�����~
m��Ih����oy��!���s7�
Y^��9�)�hq��yw�s�������
�?aa���?��VXo� �.9HG����B�`���D�7��8�t�²��ʏ��_�u��7N/�q�^���xjY��xИ��1~}�+=�;�Yi����-9S�)��ʸ��֌5�vksc��^m�-�`�� @Sr�ݱ&�����X�
��c���qc�f�җ�1g����cLN���u�+�S�P�q3��;��`_ �jf�1e�k�A��J8BAc�V�ރ#@Ku��\p4R����Vf��n��7\�����5h�{O�nC���"�	�X :�OT���K�w 3�п�D�ըq:��0�����?ff���\[�����
9uG��Y��-.ǭl�L-m� ���r�k�ԙ��	���uw�7<�������;\��K������])�W�W���pާQw�$���A%�T�E�L���D/k��C�w6�>T>B	����'@�ꩰ� �J�I�ݒ���!�3�=��(���V;�W�rv�5�¯ʄw��[{�]��'��y�ĸȕ��F/��!	�h2��]N��x9Wŵ2)���^���2���{�����b��>%���m��%�����&�����0��.^��f@�C��; ]����X�J`(�_�C�����a/|Sm)&��%^��O��(�����6d���z���^>-�&��ĺ$�0�q�1�����w�|��5ޅ羒����>�����ex�-�WMz{�^)!Yj�F����H}K�E��b-`��"E��OS�dqg��n �i ����+!��f�a�Fۣ</W�ؐ^x�O��^I�R�[�~���H��z}y}��n��ʗ���('��=�D�I��-5#lf#��V�q��В,��5�,@s�ˑ��/�Q�5Z0��ֺ�;�Tm�Y����I%/8��|�zL���;��Z�X�쁤��sj��9����5���RJ��:�;$f�ӭxɔ�F-RO�����5������i�H!(�P x��??�*HI���K�
�0��1Ꞙ�]�qF
0hjs��~=�K����5�W+2i���`sK����N�>~9C��m�?Q�����e֭wW
��{n�t8��p�4l��隁��wUTu���VEk�e��0��/V��I�`��|��P����������9ÌN{�@�ǥ$u�KU�q!%�1���#P�9Yt������{��*�B(@���_U���E��ŅH�&7!��OH����tٯ�:f�>M��t�oǬoh<L\��>l��@Ѱ��$gZ2��k|���A����'F�?ci;Q�ud���R�$v�,�K���/�q��Q!��Ԧ�����n-�.�-�����E�&�O��m+�L�֮�
�`��a��"p�t���m7�%5�\^t�t���7]&m��j�$�aA�X��-l�$�Ƃ��]��0�{�8��׻O�3�
#���Z^�w�q�$,�c;��ܚ2F
]���Ў�)	a���y*�]�4����>��C�=05n�������[��egS�� R���U��Yj}�2� �tRX]N�,��_s6O�8Y��o��(� ��'�WTv����)+K�E�l�H�����$�Tf����DA��]:�����Iގ£J���`��V�~#Ǥ�jAe7WQk�y{�ؖ�g8.M����8ѧ��*-R�����M����ri,&yW��I�a߈ ��E2O*}2��EA ����D������-����q�5�6:��jA��o�K����I�vl� �>7���� �#a�P��6g�E$h�.���4\ZҜ�u� ��_�q}{��ʓ/w�tPն������6d�T�h)L�(�[x�b��"����ɟ了�f*t�����Ԝ.&=�B��.�BI$�;���A(p��Q��2 ��OUR��* Y5�׷����N�j:q�9�6�s��$�9��e�#Unn۬GE6[�2?[����-Z��������CD(ޭ#�~���AŚ����:��G���
ޛ��|�U� �(Vd8�O!7��Jp��ZF,%��s0^dj2��8a/����b�����4�Uu�zc�����"8��d^�����z��Y�"�Q~�	��xV�A�f��1.��9&Z����s�f�Ո�l�<�>uYD���wHS�=���!`�uV����j����2�n,�M��#��
��($��
�O����9v��L�Q�}��;��p>�
A.B�p;Q����`�@;ʙB	�Co~L��v���^(@��_"7L�;��'%�V3�%��P%�~Dݝ=��/�i\��J�Q�O<.s/���Eb������i�,	,���n��A<�x&�]�U�Ct�$7%˞�6�GV$q���D�p��Ս�
yf����D���'����9l���tp���׋��,'�D�}�4�����X�����1 \;yeLi�Iv4��V�Aҵ��E�M��hȈ�Rd��9�P&���d~�,�`���Ɵ�~�w=���t�7�s���B�`&��k�>D;_=L�>�zB��Պ�i>�(u��y�%�P������%'����W����Dʲ����i���g^nА㛅�f�'�zdG��m�0i���3b"�{���DT�rvuӃ��GG� ������ r �c�gD�d����+�2Y���n����D݁审R�_>�r2�t����Gѷ���T*"�Z�E@�1�E�l��F/5�(�p�#f�ِū�}�7?����?o�V�I�\#PH�������6.?���1���6�*5��-�*�-�9T*w�}�y��*�h�t�P�.}AN�Z���M�n�r����	^.�*���gYz1�	������6O����v�G�R���*T���-5��|3n���F��E	9K�b�Fc[��S�s�s疞Y�q8(���C
��Z��nC}c�h�ou~��t] �/�t5�1Q am%3-�R���C�~���ʢ��VΕc\4�p�1��1�0����R? �d�IagR#�u��PI��Б\-v}]�'I�&���Ii���I��(�HM�Dt� �~#NC��cD��v���@���X&f<YRq'L��`��OPiG�Kdd��QY��|�՝���9$�F�5=8�2�OLZ8$P�:_�/��9C*����4��B'y�8���ͮ��Z�-46�V;�Iy)A��B���MQ��6S�w.V5i|`;�:���vԵ��Ԅ8�[�H�ύ�q,���n�c�W�e��0u�YM�D� ��b��2\ՔW���HO�Y̆���xȋ�+ &q�c��fQ%�����dYo$r7��zx�S���(^7�4�/b��f�}`���`r��Px:�Ei���n�R����x�OnU�c4�X\�ޯ�q������rb������3jj,c,s�/E�az�n� Y\?8�Uj)�� �,��s�O��M���<�
Zj[���� p�{*?�N�U�����B����թ��F[�.���C�Ex���GG�I�L��˥�W��}~�tQ&$T���̩A��##��~h��ן��ށd�V!��tx�n�v
r��M��p�R�	݋�o�d>p9#vڇL���q�>B.0��:��ie�Bi��Q<�`f�ȕ� j���5qq����|�6�]7�h�h�*֗`Z3�TxXU�st�Ha~�y�i�ؚ�St���`����#0���(�����X1?�t֋rt��2n�_��|KFhm�W�x0M�%��`_!MMw�?�0z��X6�S]��A��y47P��� ����hYв�)O#-|���ܒ�22FB�z��_����d�4��gg�w�%�N+v�X�U�$���@�e�b�C`��Ք��;t��-?��঻�Wj9��1�i��dD]�Ӏ���(gg)=�t���#<�e6}��No��-c�����k��ضP�O7�u}+lz}1�e�Ma���+� ��������{�[>}��M'C�m�lð�*�ِЗ%uW�i���5��rVM`��g`�Iƅ�[GP��J&)>�9̈́�J1#
2�2ȫ1/��3&>�L��#$W�-*\J��gy ��^�39ݷq��ok���F=��@Fq���S�
o��ʀ�xR ��tj IY���	`��|S �!c��e=����#*�j@t�뗢>��O�x���[����3�;�!W���	�Q�i��B�j�$-�[8Չ�G�i8A_#g*_�a�_��4�VQK!H��狠L����������XQ x��]ʬෛ1����Db�Z��O]Ii�h��C7�iF�0%��%�K��"��׶�$��cs��8�����4����-;���A<L�C���%ο�ۚ	w����?����Nk��
Q��#�uj����LD�_ ��c����������c�̐)��ZrP�}Ɋ8Z �<z�0[|g�u�����Tj���y���<���{D~l�����$li�s�,�e����$�����gi�2n	���H�4Y��6!D��8' �|���詟-֋�Z	�S���A�R�<�h5� ��0�����p@�/�ݷ���1y��j�|��B���d@�Hk��W:YT\�4�v�\e�1Gk+�x��S1�ƹ�Fɘ���k�?�#��/�)��}Q&w4�H�  =���Q�s|ΟxdM�S�2�ܬ��b�k���ӺE��V��֩<�����8\e-�>%��5���;�6$-��gq�m҈��J���o�WRW����ۢ�f�3*�Lc��*�Ҁ��2=��;a�щ��*v�Sc��/��s����������A9��T�Y%Q��]���<��\�)z>���C����&�UB���*��p]`<�t�A����\]0iMVP�u�p,�[��ݩsO����>�7g	�Tn��~��P�u)ѣIU%�	:������~ji}�KM�m�*����u�0���-�+=��^@�l�z6RʄT��zn@�}��f����]�	�c/D����a�;�#��@�<) |ubu�b�!}�ˤ0 �|�����4H�E��.(��2�0(���� 
	?nT���u'���V8���g��j�:E�e �[�qe�������_�v.B���PD�O�ї�(+�iU��P:�V�D-���I�W���cP��eg��}�H0MtV��� L��2\�`ux��33����$��EP����)�a�3JR�*fĲ���g�"��g�I	P��(X=ًhP3����l<i�_+�7�S���L�B"��uB�9C�n˃��J@�:庚�L����r)x���A�� �c�����A��|��~���~=9$)�8ags6�PO�����?���ӠKKǨc����A�Ӳ�g���3� �1Ll@e�Z�R"g�@�v��Z�H�Dq�C%�}i��!�*�R��$t@*�I�k�TL��v�*XP�w���WH5��$�ᗎ�W�Pc�����}4,z��ѷ%��-��h3�}\�g��v}��{�hdͶ"�x`4�t��E6b�a�͛�W��,jz�>�FGm�>� �v�Q�0w�~����O�,
��+�:z�@QX����
��%]ϗ���¿�FE�\\=��
҉P�v�3������h�;��a�"}�q����ѮV��x̓m��mOw�牆�~٬�0/�L���%̩"� (�O�w���/�����|�8W�g/"��L�׮��x6|�/I_��V�z�Xa��wH9��]���6�qj�z��/3��7��Ö4��48t�&��8Ր�UQ�ي�������ai��}�e�j��Ѱ|�9�	1�	�Ѐ�o����#?;��B���H�e���ٷ���@�`.e:��W�M�z�	��l>HMDV����\W�=�U"�^-o�#L��Q3x+�}�c7Z�xĝ�TЬ���Y}���?�~p�va�t�/����0�ˎ!�~��H�WO�g��{�w�qB�pU�f�|ۭ� �v�7��^ĊrQ�A����bȏ�Zjcn녣�H�z���W�v�mMk��y�Z�um�xb*�@�A����pA�����N9Z9aj&^�raE��MY��٣�M�9-���e��G��U���y�#��^Kb�nFo/z��BVhb1

�
�����*���;�b�����I��@d�� ��t�����F+=K[���ݿ��N�-�ҙ�&v���ԐD؃���_M��NȞ�5�*�+b�
�Czq�m�Hr+X(���̆EQ��h�'�5-���mN^����ܦ�tQd�`�q�e��l9���6�am����;�g������lb�w���L���T�:�gԻ8�&x�1�����V�JN���e�װVe����%��3�ty�����(��XƩe�����<�^�{z�u���P~��<o��L�{#�k)`�����9ˆ��y;ٳx��C�2�X�v`Y�E�B�=ީy� ���#���:�h;��aU�lo�5�����t"@Zϊ��G�,�i�d0_�`���ҟ�b�Q��|�-As	�b�X$?w�a2zt2������Y�G�O'q��|�>���(#s���dW��8{�*Qu����@�f�.���W>��b_��a8��JC,_Ǿ������!.�'�4pɕ�I%ʇ^+J�s�-��$�q:����a���-��������A1�ǉ<������r��G^[��Z/Lt�/�(�N�Ŕ���������-A#a-��K]��R@qo���|����T�ђ�ԕ�T�S�����"T�	|�H�祮Os�^��"&�BOyP?/�"Z��N��}�QW���
5}�s�м>�k>.,akU[w��M,(�[0xs�n?V��П-&A�54
�{�-ڳ)�����0_�\��7*QH=��:FM�h�Q���g��;�/��U�1�Ⱦ��lq���S���1�E�Pe��4C,�.j<�9A�+�ȉ*4��@w]u���5N���|aC��Bx��K�DB�F	9��}l�$�l����d���H��= �ذ��'=���MȔ�i)t̋�<����T���t��#W���b����b��V^V�!p��B�Jԡ�@m����كѢ�VMBƨcFzb5�� ���.�H w�.�h��y�`n;�gڏ-Z�?�z�66�n�˵���D�u~�T��Z�:g�i�!�tb@�;6ӷ�^L��aa5Q�o�:����8Q/������'z�"�Mؑ)��f�e����!0/)D��
�,��#fp��qVÛB���}/g&��ཱུ@-���M�Sh�i �,P���POU�)�[�(S����8F�B�F �`�!�m/I+Mi�D���s���ǜI��Q�Pj��W�g&
� �}�edY�rO�O:�T�n�[�6���ܴ�� V�a"�b�:Y�2���@8<�V2�RWiya��n+E|^�߹y���I�r�[CHZ� �a���@�����	�g��ֽ�nFp�����d�y6��b;�г�3dp�<oCe�y���~� �Z�s���@�\���J%�?��?��r��AQ�m����h�����8f3[HD��]~{U��;� 7	t���Z����){��(�/���;/^b�u|$��w�������9z���V�m�����磇��v�}}����|�vWa����ѹ����U�N�T[�]
���s@���щ�Gj�?`Y���B�r3R3����+8>_*�:��x��E���a�Ь��%y�� {zm��n~�2A�'����t��i�fp ���*�u�@|0������cl���a3�SWo1�N}��Z�nA�@@^��d��*��Xz<�	Y=��o��E?3	�����9ك{yh��a���+�`vv�*#S��ЎA��q���ZS�~%O}�z��<B�W�@��N̰�Vx�yw�-����`� �xT�Ǧ8�yݍ���	��<�XA)�k��X�~����kN*�T7�!q�)�KK��4�H�l��y���|�7�H�߇L`"������M�p�p�����\&�)�|F7�Ո�	uD�~:����0L.Z���������vV��H�,n���G	�c�}�|*;�KZ�m�)��
l7�ȋ�)��n0�n4�4�f�T���H#��~�$��5ַ�����x�K�
��𛜇Gt��"&���[H�)��t3$2����x���W�?,�� ��E�b;�5�X�$��?v�OnU�7K�ƪL0?��^���x:Dr@��E%���{����b�g����y�r�))s���gk��)���\W{��3�8�ئU�Qc
�%ͧa�1fn����+�J�G��:|�Џŏ㱿�HT�l�J�S�4��F������G���^�闍R�pg��΅�#�yv��_+Tr�P�QS�+�]�i���)G��l<�:�0��>��oynI
�\*�T��nevQP&��i����:=O�&��Ba/_�K&�R	{���)�6�J��v�9S3���4r�a��J��Ϻ��QZ��оy��5k�uP]�G=ɧk6��R�R���t�9%u-��-�u0����3��m�7-���I����yR���n�o-��i��=��.�71xjM��V���đ�P��$'k���i�a���b���א�\���Gۂpm���ѴaԊSZ���ML�%�.17=f��O�z��`$�<���u�`,�C��'Q�A@p��w����î�&��1+�ݵ���?�i�)��/	�G����`��w�O��?�$�Ԥ�.(eu�}U@�t\K��q��5a�<�n��#r�7�?�>�P�ˀ���z�|^�%��j����1BQzi<�y��օ�105��v@�EZ&z�m��2k���&��t5Okό�8YZ=3�a39^W)&�<� {�|��,֓�O�,**����9�S`���Q�G�	�~�4�,I
�@��Eili��#�1�N�lïf�`n���k�<�~Z�?A�B�����ŮA�%2�?�ڰsJ-�U��T����nf�TU�Zm��� _;���?�r�=W;��e��8��1�����R��)��:�ݠ���i=���+�R�b��0����2-K��(/[1����$�l��<7���a^��[����[�n`��_�l��h�|��FK��O
��Ie�]0@�'�gl���*{�2�m�y���!�����* �K�f�G�n}R����(��8��?K�<N���� �5Y)�
�0ڪR�k���5�9 �'T�m9�O���C>�����J���0�2�/�=vڒ�ɂJ
�fTI��N�V��b�aT��Y��P��G�FF�	�4��Mj��5����4L�ƻiBV�O�����i�6zz�#N嵱��L���6Ψ�c��������}��v�־�E��h$[��бJ�LnK�]��A I�i]G*�;xl�+r�\+���7�±�~Eg��XxxU�B��P�������h� �s��v+��<��khJ�����S\7��[j�ܽ<���J���.�4ֵV"k�����+�l"�w�ߖH^�$�̷E_��<�T�Q� 6�O@�v_�J�Z���+�ktO�
�(�F���/���<�"�}\]ס6�g�4j�����(�>`A�ƪgr9S�<c(���T�}�/��/L�u�T��B�f<O��ڏR� !��m �^D���f�� v��fI.u��*�h��q��|Qǉ�������~�5Í����1�3W����5�|�#@z2m�x�[���⢚�]�M�t���_=��y>�`_��8Y��\�+��oa��sd�Tn���Op(4��s5�򴲘Z����)���~�!Y������f���;#g�����Ϫ���v#�H�"V��6���� �]���lCf\K���ə�R5�Ȧ`��2~�|f�P�H+��(���Y#��|Y;$�lIW�Z#����I���0n��2���
X]�fC�4"��He�a���$4E���$_��eѾ�4���a �/��Z�@���P鬨c��Y;���j~�̳�q
�i�-�lf�����	�Q�S����c�s1R{O�ر�������	��'7�f+��UHӞ��һGR!��s`'B%i���}������L�{D
E��zV[:������NW���|�^kHR{�Y�Q[Ď�$L�!>~��{�D���
z�	��U�,d-ض��ڰ<O��_�~��P+Ƽ��읆���h`����s��T��ڿ�����D�/���X�*|oH�L&� 7	��G����+�Ə�i�H;�H*>e��q����8/��!�"�t�+���]���=5����1����u��w��qU��@ ſ����'���p>9�P$�b/>�ms�@S�0EDhO";�p6A3}k��wW:����ih��O�:Ċz��~i�q�i�r-`�ޱB	]��MA|E�s�a�(h�zԯ	:�54g�G���w�T�h��!��h6�:a��V:]�[^��V�q�O�_+]Bӫd�ޗk�%:�@"G�=�����*���P˸�j��j�ar�����"�jf�q��C��7��<��h����;����ˎ3gk�)�*���I<LI���ވU;1����@�Z��K=#�C�����M2��j��!��N���?���Km�C8��^�u�5��'�a��7��BԨlX��>�0}�k.�~�E=ZbxDA�3``�Z���,��6�+�p�k/"$�cKd�b�
�s��#IP1�o�Щ�B`\f�k�N�t��� ��~ �ء=f7��"2�]"��l��>����&��T{�T���s��႔L
�x6����6���!A�C�F#R�+�
d# �]oP�"����3�D�����ly��en7.�Zr����V��˕�/��8����J\�Cy�#8�V��"p��.|1YO�_�n�!b��1;�v��A,���K�Ԃ6���by4�ɏ�����HT���e��и�_�lζ&�����c���|�O��>E�b��3���Gsɹ�b���]ǐ��@o8��M1�.����c9|��;�̸�dE�Ĺ�ᙍG|������H'i���U�{^���Cw�V���]{5���B����	iVP���Zw˧@���Ug���ψH�g�ۇ��	ԭ\H��X�8���~�%t.�yZ�n�1��DZP�ŗ�ë�P*����2��c�[v��GN�V�5��U��O�Lݧ)��)��"�w4�nx�����1�X�7���GLR����&1��Y�����I���T'6�!�EĽ�(k�7�F�@����� Y�]0�\p�p��$4�ۙg�� 3�+�+����]a��8�;M��Qq�%s����$)s���
g��  vH�oʃ�3��$�@�fj�����e�r�`�[Z�_g�1�z���`�3�0� W�%k�pCg�ը*��s&��(�� l����q�r���F�,��#�YX�ټ1�}�_��4}}Xb�O���Ӫ*�ĵb�f�y�Z'�� ���Ic��s~��e_=�B��"���'�T�\2tC���F#?2s���iM~�9��%c�bWh�+:�s3t�ݐh�� ��d<�������"u\T�hu���SɎ�n��Ch�8�bro�R��z���yt�7�����܌� �A�n�N���m�~�^ +����Ϯ� �[�T�����M��d��hh�)I*�=6��ABbk��~y��c���5FnMЌ�
⏙tRK#,��N� �-D�vi��^�Db~ׅ�U����W=��B���X�֒��F۞���VT~2��f����\�O�;�v���/�Q[d�e�s�A���"_���یlG��}���e��ۅ�4q23&�!���)�/��И��>���v��bL�ћ���þ����iٸ����M�	��suM��4�D�=�E����,�N�3y)s�u'��v�d}��|ҵ�E������V�����4����F���?�9_Ō�ѕ�t���܁[�>���  &T�CH�\�*�D���6�r�\
b�0ܾwf5�א�w�b�櫎��l�H���>�|�K��8��m-�g����դB�¥PػL#��<A
�ė��]7Pܶ/ٷ@1��
I�z#/���,���U��_�$������jÜ}��Oz��q6R���@�C6�z�L.�d�z{�3J�����x��!*�)�WL�B3xȑ���Ҥ�g��x�E"C���с�J�"��&�$H���+�v:��0�d�۱���?�[(�ޢ�-joK��.(�W��]�)�M�5I�
za��qM^��t����],����!P���6z8k�\��;�D�Po�?/�x�#�_ �w-���TV�nM�\�k�Hu�n9&��%���h�
�H����e��[G�-e��"�:R=��4�k�)�aL��K݄\�]%��Nļ�Wb]A�f�p��m:�%�����pf�Z�n+��w�2�꿥�x�M�p�:�??�$�ʘ�	�{�3�l�}z�DM .��~Z+����!���IL֡.i�A^�O�:�����q۱���3�:0�C�0��C2���&�c���u+/	�E��-� `�A�P8���ʹ�Lɴ�R��!}�p�c��i;�	X΂"���/���W�+6])���H��:ji�,d-�
Z�����%�>6�@M�u�$��גǐ+͈�w���-�8�ǞP�ttjI��-�=��Ϧ<���t�k�[I!��P��ޏFZ#������s�dRx�+l�'3J��	�rW��qg�΄�U����T�^�?�23#�[y.wW�r�?��`��0��"R�� �=M��8��	�W��'�j���J��˒����zH_vc֌�iT6�ϓ���e��,V�>���7�I�M[jx?���1&~ݣ�	���fvw��ǎa�վ�Pp�[��ٸ mޭPϛh�経Y�a���E-��k�𷍺qLE:C�52����ƛ!���5S�����:i����T|�a3:S��e��\<Ҕ.��qNu���Ã^���c��̒��n�êG|6�Jg�n1���pd��V#]w]�LP�Bk�9���1B�H�S�`^��;���,�㭧8���QXi�:�So4]M��la�*�A�X�z���u��������5��vx��Z=]� �Q�߾f"u}p���v6v�n��7G�^)a*�!qu���P���lEݚI��ACO�ny��ќ9@	-�w��З���AFѯ.�pf�Ȋ#Q<���q��=`i�ץu�m���"�tTʻ�������wR��"�G���	{j$��c&�=v�B��F�J�U�\Ʃڛ���m���9��V)KROTO�G栂��o'�Ƶ��!	�Nl��k�`|WK"L����i g��h}�?��ֵ�v��RY�Ȑz8����%q��Qld�����&ؓK,��~��~C��ė[�Ee�j��*��W�pʺ-#�P����o��15�wJ`S@[+�ʽ^`�F}a~Nƒ'�{����Ae�% �Z���h�n��O|�Ad��v����h`�����A��b�oh���av 4��47.���I���v�,����COS�k"��-��S� ����$��&AS%��'��6���.H�_0��T��Wq�39��Bs���7�<�)3X��8�g��i����(G��F���ꆖ��qQ:2lK͊�%H�d�e7G��s�I�Ito�ݨD�6����@d��r�*����|yZi��4Z&�|2nHѓKfm���$��; �2eS�4��Ĳ@\��N���t6Q-�)�Xg'��6\Q�V�hz7~�u�^[T��*�3�K���ڱ�c	��qҼ���4z��1�I|��i��ӈ�����X�����d���d����S�~�W���s=�#�9Xg(~DI�Ir`��DN���:4���AE�<U2Q|8�����n���wGD�t��u3Z.E��"����Ӽ�f!���$���_��N�@��9 ���*]�<���� ����&�2�og�Ձ�Y�T��v5�_���ft�lE�A�Og�z�� ��2�|�OU-�XDs�X�H�P
iE�v��{�i
�2�k�?j����a GΌr53 �OE1/��!"Cp�	�g`>��*#sewb�0xpǛ�7S�E����,Z�����E5ЉC�
;,�<M��f���k��*?�G�ȯ�2W�&�u�\�w_��?�z%�L�b�<qǒX^WYf�ކ�G5�tفO�jG����m7��Xѕ�ݷwx��{,���6����X~��,m��? ��-��Nd�a��� 7�?3 }��}&�a���L9�e)��τ�H7����_���'�����4U��╳��!�\��]��wA�,��1=D6p�I�|v���)�OI\���z^_R���O�r�
`)z�%�j�*hL#�.+�������$Kk�2yMY~L��3��C�m�)ĀNH�(��ڸ��v:)-�ˇA\n��m����2����(��U�vl�ȿ緹�&����Z�.^�v<�b������-���i��Kk&�6��=�_ԝ	�F�v�[�ӥ8�æ#�|ɧ��"�W6Ч��W@��G?0�XP]�J6�_V.e�aju����gap9���3�����F�xO��ɨ��3]�k��?�+�c��
��������=�ƾ�)D$~�W���+1H��mSsއ���,���h�HC�h.X&g�|=����)����>�n�vڲB�!�L1,&2�/˾�h���řp!M$=ԧ�V�X&���C�g?]r c߅ކ��r�U�;S�f����}�AI}46�D����s�n]��3ᣳ��sWYĊ	��vƺ�����g���5�����0�Z���;�`9:��rbƱ����̃�֜�s�O�a b����N＜o�,����)z �7$���{?׫����)S�����y�+��f��,#N	�[{�Kpe+L�����b(>VdVr��7Q��p� �t��|�W��3`�F�+õ�G�m�x����l�z	��`����`�p���*hW��@�<|�M�����	�x�CHI��ܓF|W̍��8������=�\I�Y���=����{~�����+�U����Y�u.α�,��uma,�1;�&�*hS�����AZAf{���r2u
��=D�ғuE4UoM��85�{]�N�_������H�W{C^�˦�2s8��ʹ�P,�(87�TL |gJ{����~�gUF�1�F�C�1�J�hJ��z����y���g�	�e�#���������ņ-�	Z��X~�:3��L���xƓ(���=z[�T�������ȕ�}O�<�S˕4�T*Ю�/��\0Ս���$ Kkf�n��|�gS�x�9�uS��DdK.7�k�n� ��"`nj���$�H8��!IN
aace뱔��#�����жes&c�xR,�ʁ�[���C(~ =J�n���E<ӟ8�Dೊ��9D���qm�z�⩸�����!�� i��U�!�J8$M�-��RSsQ6���\2Ɵ�-�ͅ(��qa�Q����$�-c���9^aQ�}��{���s�Aԣe�1kEA�.����U��@+�8�<���5��v�/���%����4E��bm�� ��%#��Br�%��Md<�r��&:_����_�DH����U�C%�*����=Z���٦7�T�����H3�����3�Ԁ�
\P�{rVl�WE�D���0�&?u��?>��؟5�_����zE"+OZ���/����j�����d�K�b��/c/[�-y�
�)o��{����~�v�C.bG���u�0U�N�`�\��a�G������\��jB#3Ԍ;�pK��*�\ۢ9˪Y����z�@�'5Ô%}J{����7ct�D��n��[uf$)��7��t�英�S�� ��:\��:�x�C�w	�.h�gj/10eZį 	_�M1H�)@Y���lCҁ8�/���!�铯�|�T�<H�8�YQ`r�U�ٖ�`x�M_���������}�M�vT�*:,y̧lݙ��ϥiS����**�
g	������PZ͊�r�mMT ?�N�)"D�M���
d�?o���*<+^$up��E|��B߾G]��I<�!t�Ub�f¨�y`�o|,�}[�T��=�9���;Xq�)��]QNT��I>�F���N+�D��yp)����!��G�A�lD�<�'��w����ZH��:����Rp!�J���2%o�0���A8����!�C3�*����$RQ8�TK,ٰD�zt&�E�m��$�dJ�Xs��Å�ГUi���!�S0��u� �T�oW{���m�&��~WR�o�,��@�z��U�>4e�Ɏh�<���ٞD���c�����n)��30�^h��Xm��(�(|�CcfFs��L*�;��<e��W�c{�+���6���4��F*��ǒ�u$�x;IU�AD
O9�V�`M��Hǔx�������;piK�u�zKaT}�:�V�m��T������9�Z���H6�$ky�w��(��u���İЉh*ͩ_N��+��@��P�j���I5�(z����H����S�K�s؀q�~fK��*&uV%?O�����L���=�Ux���|ĉ-��`�C{nx�乹"
)���a��o����T�7�3�0�؞L&�)�Z�����ܐ�3QGr,n��}YxL��oˡa�dq��)�6�(B��7݇}[+.c��{�@L}����-o$ң�����I痷�3-Z������^,��ٖ��.;���}��*+uu�/�+S�tԵ0��m-=F~"GFZ!�o�w%�!�]|JM��'��J�_:�8��'���q��)�� ��K�+\����:mV�����I����&�r��(�-D�"#�'Ͳ�hȗ�J�z�w�3�+wΠ6}O:���}$�G�yb��I���	�/n�o����̛vSڅX��?��|#H�yXN��=ơ&�'�	0�}:X�ZS�pV�N�c�%�5ls{!�H��.���0��4��۟�)��Z�D^w�����X�GV��Ό%8�c��w��s�9��3���Gs���D�u��v�t'W����-1�z���I� �q��6d4[?[!Q�}����E��іg�8�.��Ii�5�>B���@�dVc�{/q~���oMr
��y�p���g���j[�-e�!�9��ؠu9GѺ�
o�;y��ni�B̂l9��k�`ѝ%g���6�h>)�.t6Y/c���p?U���E�f�w��f-U��� RRN`z��F�b/ə�҃�:�v4�%(� ��4g'�i��KJI���}	�Yl��̤�[�BJ�A\l9p5�P�5gń������F;u��V�
Ü�a<���)`�����C�.�t�̼V5�1ɣ_[?>�&�ٶ�n�Rn8�Ick3�շN��*�n�$��	�o���3
e�VOG��̇B�!���I�x��	�ڲG���Cn{";3����Y�b__��g\퉰KR�$��b�@c�Ϯ+~D��9s��~}��}i��2>�h�\�wUo�տO�8�<`��|��5(�ȋ5!8	��mK �ǟb'��A8�$�v�,�f�ڭ���[�Vk�|my�8��?9�T��$:!F��hp|Ry�YtP>�B�mi~7P٩	��6��a��&��b�+@��NOvgV�����rA4��4�CL�_��%8�W�2Y��I�ޗ���:s�������gQ���Мw�sE���D�T8��>�֔�&R$
Bů�D�_N^�͞�f뛫���S�Ŧ���|�3��P�������#I�Q�a&9�����K�XH!O�����1���`70����D�4^�5[���Ӵ��q�Q�|��a�����UmꟐ�q�tvmEl�y�3��u;+~�0�z��Є�yFZS��IQ�����5{��l{@bR��������W���X�b�B�Ԅ��J��tK J>���+w�2P|u�L�΅"|6�r{7�#3�&K2M<����	�׵K�8a:�c�\�!��z�=K�)���dP)g�
�j�I�Y֡�&��� �SH�K�jl��#�$�jW�Dε�;ȼ	|�[��@�I��_��@n1�/<�d�����QVBn�:�D���e�88�^�����c=܋�I��7R�W�s����Q�S����=z3�:pB^�R6���Ŕ���&�T� �lV��Sݚ8m
r�=���zQ����@���J^ՌB���'Ɔ��8�a�11�>;m"]�˪��|���W�!��M�eqh5�z3PJ�u�����߼�5{�j�|�!W.=�@J������X������z���f�B0��'�і�����6��4�S�7^笪w�p	m�0y��_��1K�#��V�_�;E��'*em=�����^/��u����m�3���Y�<X#����1�dϦ.�a��-�A��ث��m�n�m�y+S߅ʨk��Q��G����{�`ݣS�,nDq?��Ռ5��<���QC0���Het�R�zu�;#��d��.��S>֒�Jן�� �,&��S���{_0�թ}��P��[�g��q��Q�x��x��q"��Q3FΊ�DF��5����9eb�5p�3+UWI��C��(����X}�����$x݆� pK�X?P?$T����"'�C�j�r�-d��P�%�\"sX�+b@����1r�?�ĕ?��3k��/:N�ON*0L���h"
/��bd�y�V�u��W�.����zu#��T�Z�_�<�b��5��%g%�������6�#���r6j�cMu,
��C���"���T �}Yo�ͫ�ε�lq�Ƹ�I��DKªy�^�y�G�O,�o�õ�=e���\�L��}q�I�-��݅ǡO�⧗����x���4��^������]%gHd6�����P� c.��fd�L���~Ǵ��U[�}�覒5���Jn�a?�؊7�L?��5���H? H��zDhZXZ0��Q���7��p�o6/������W_职2���^xmD�¾�*G�d�?����E*�ͷy��|:�0�\,j"��·��|�Y���~��0��	v�ƞ�����P��u;�:��N��֯�&��#�>  >`xLE�8[�8���a����@kb��I�)��n��ِ!]���2ȹ�?��˗����Q@�o�C�)�4�aY,QIa�$��G�y�&x��-R~*�Ƣ�w�I{m hf�@��
��	�'��ݨ��,��˨#�����ye)����V�L����5�]�8t�C8��r$)1aWy�#�26�䐆U8���� �_i���ĸ���/uI�*~#T(�CL��"3���X}�&���l	N��щZ�i�����@�����Ǚz�����s@�5�<«R�z�i�+��+�Ul>C���ڧpv���(H�lMu�׮i&�A�K}}��`�^0�ԡ��v'w�4J0oɳ3]�%�B0];F�x}t�m�3��%�(bv�J�|�1_�d�a����|�#,�[~h�8��������T�6y�L�e�!k 
��f��0��� �YZu��gs���Ɓt�-9Aӥ��&/3�O�	{i��FA��W��I@��˞B�%�s,������h>|Q����<�łj�j��ʟ�qF�$Y������w��ܠv����Qiֹ��T½v����;\/�'Y�ܝ�a@�ϸRJa �����u�50m"�A���~�֝�/C�v3��wbٌ~PT�x9��g#�CSyQ�h !�ˏ@-O�8���7wˏ0z��%��m��o]t6<iL��@��!B
%iָzf:�����FDݏו5t0�tzߔ�.C�����M��eK�v���>�aM��:E�KS�5d�SK��$�@~$Fs��������(q�fIU���̔ݴf�uc�����o�y��(0�F��,����0��#@;h?|bn�Śi����� ��=��>_�ͧ��s�Z�����Pa�z2���۷�ĳ�y�`<�ȤF��޿-�7"���e�ED��D$�盧_��um���U?=9b�Qaգ�~�vv-Tb�B�x��<5���)`��)�b��_�.�����ߤ���H#-�ҋ�?7P׮g$�]D�ST��<$l�c�d������.k��y@I�n�9}����}��5�����Gm6gƩ��m3�;���*	#Z�@��i+r���z�;��prЀQ���4Pi��s�3&^R8-��`5h��V��jK�3Hг
g�zԌWi!nWu%K,R�g�s�H(�7�2Cш��G�G�IP����C���Id�0m�^�<W�� :`^���p|>��<�QT�W��̾�4��B� �X|~�Y���Yy�2�"��4:i/:�����x�,r�� N�*�2�I�
�=e�G�H�BvZ��������
��n�hP|���F'.���J4ч��'��Z�W�#ˏ�^�Ӣ삟p��n��P�����?e����s��kg�T[PO��A�X�9��*$Bo�Ϣq�(VI�b��?UA��r��i}dn�5a�w�<�
�ˁ��Gj���+�����	 9���G�T�-�ņ�뭭6��!���&�n�T�Ҁ�#������4AL7.�*�_|h��Bͣ:�!��aOW��LF��ˏ�z�����zU�й�F�?�~�S�T���D*�p7���A�.8�u�݌%׶�4l��N2w�N?R��c,��R�D�S�L��@T�+u6�]�Z>i)�	����Գr��߻�v�Jq*��s>#��8o���@�ؖX�s@C�F4�nF�:�sDe]��ۮR��`�>��2!�3���T�dE�`���&*��j�t���f�}頢����r�š��s�f��QU�~�� ��B��3��������ߏ�M�8�>�]X�k`D�͚���2��b^�SOr��;-'�17?�,�+1(��ΰ��Rd�Ptrq��2���b9'-)�f�L��*v�y��L��ҫ�F���"�����u9 ��d��w���V 
p���$�I ���Eρ��r�c?:�G���F�'�kMSﮂ2��;�EW
�/y��i[�L�;L������Ŵ?�5��sew�&��ϗU�vl�8�M+f����l�2Ŗ}��Ⱥ��� �3i�qwiق�u�Mz-�_����C�a�$/}/�q/� ��dds������Ė��ӫ���l��~�U�{(���@�t*x���k5����&ƃ���X�x�'�"Z�l�o�?� �)�^׌����0Gz@c<���g�H ��5�YX��D���)h㒔ϱ�5�(�r�h �t�-��Ӊ�ɷ:w�Q��;���¸�]���g�6��ict�.]y7`��5��ͧ�VI��_�����`����Sl�����;G�ue�^A�B"p�7��� Ý�5�P��w��9����po�i�R�z���ԙr��t�ҫދ�OL���8o����	���=����#�'�YO!�)��s�H�j�@Y�bʓZ"�d�EL��n;�t��m�y ޘ�lm�ʇ:��
D�=��n	�5��5����a�f�%Ho�6���
�0+�4eشm#�I���oY�}�d[��4c� )�:��@�6�����1u�U%I�#����&�K/��G�#�\@X�ac��~Fe�`��"��*� ��C�A*��Q�0͆�^�|���o�JN����W�p>)� .m%֊	x��ϯ��D�[��6����1��mA�O^O0N"�j�C���$���7�ז]���p�S���
�69jOO��Ί�2<��S�oa�5�	�(�&�hO�_������f���=����C}K��7��q����E=�W�u����/���Ds��a��r��9��?�[X.�ު��5�h���G�[���^�G�1\���[������"B�n�����1��=8B3�X�!�V��)%�@ޙm���0=U�-�#�qH?�G�e����G\��x3�^�Yᘐ�Lyf0�(�u�x��P�Ґ/[�M11�ހ����L����̑�Rs���L�����*	��>kk@)
n��c�v�e��J~O��^4�*���,���[wY�;�ED���ZS�8��5fl���V��I6_���M�$���EL?*�_���M5V���&=��3�;T�h���ޥ�b\<GvX���3@I~�+��#)����E�d�W(�M,�w�9GjǶ���� M���Db$tY`#�}�]n$Б������#~��r�6�+��I�@a�Rӄ<	g��c��g�6�)�ӦS�L*|�-��%��y���A�����ܝ�>(p���;o����o�K̼�~��9Psj ��j;EY�&3�M�VƝ��f4P�E���Ď�_�L֩�@l9���g	�]Շ�EdI�蒴��:��p��MI
РV�Z��o��N�=s`$�����V	� ��� t�l'���
f"����AVO"�N����g¸�9eA��2�S[�<�"�;�2��t��OY����{��}vHUшߔ�g�z(z}��9%���ťn�hj��._*������b.Yg$zXV��Y�urF�G�s�_���3c &�<x9�cܠȶ�&��&c��ܿψ'�ġ��4�F�_?����-f�q�:�cD��e�g�����!�hNa&4x�5F��q�u&�jtRX>�?��M��,#^������(�tz����I�7����G;���h�
S �2�|�7jĠ�u�p�O��3T��6=��s���1"6�ρ"��3�09WR��,7WEP�=� ������"/�N���&�ǰ��Ȫ����#a�����@��覾�[6��v�5K@4��؈�l�C�آf-�\	Jn��w���q|����y�j$9�e�׷>O~2�AJ�4V%WQ�݋<GT�؂�.2Ȇ�K��נ���~�������9eG���?�V�f��N���_���ڏ��r�W`W�o:3C���L�ܷC�B+|�����3T8��|�1���!���|�ߙ��&ȹ>�:/�J<�Ғ����n�rA��`����N2{Z�"CK<&b\��=l���RCDrQ����2��F�4���'���W��x� ��nv�3Wڙ��vRw0�Ia3��"�b�ۜ�i&�-t�"��	�:�ehl��֣��>7M��,Bu[��2 jYh��Ј+���t%�R�G�"+%����!އ�f^�/�W��D�S0T��S�ז��t���")��Z6	�*fE���R܍�<`T� p]q�%�)-[_�;���^��˧E������z��_=�_�Շ����\��[�n�\�sUMe�O��Q���G�Z7g�����'a��"Yp,�3f��;��9J��f����=��/�=ߗ�z&� �<���=2�$~Rq7� �s�Y�jSuUR����j�A PU���jJ|�&�l�܃�NWS�Be��F�����#��WE�1,fՔ���WjƤ���Y�=����G~	�f�n|�N/�>���-4�5�e�7��n!�p~����~K�`9�Β"f@q�~b�3�Asd5� o�N F�U��|�U�� 3$�TT��G��pux����!�fȧ�R�+@�BX�<,]�+�B��S�7R@�ˢi�Y;�s{ӳ��qZ��t�V-�b9�w�|@��`�,"&XV�=�d���M���w�Q��.���2�����_F
c�b֟����;3n�:!��@&� �.s�2�q�k_�C��x��H�{
���d�K�./�@Qܺ�CH�U��#&����2_`��+�bRC��ͧ(�q�t[��M;��'5��Pб�?���=�.U�o��(O�-8H�hpm��B�5��8���J��ԗ�%z�v�)��k���+3�l@{��~�` @1�o�tc��Q�$�m���pz����h�>��ᔺ[�>��g��,d~&!��R��FG�b{�(ϝ �JB�B# d�}Pl�x�l��`e�,0�'��Ӕ4~�> �<�b��y�UB��)G��i�H/m�Z�)w�x�A�k]5C�q՞H���>���>l��@|����i���qoN���L��25 ����y;��no���.�]��l�18^I�|�.}V:/��Ũ��Uͪ�cH�֦Ʈvhjq)@�{<R:A���p�{y%T������=�_���@�w܏��W�E�l��O�.�\t��s�M�'$�j�9r8����w�"UL�����SX߫��$�_b4���V�So0O�N7%?�Ȟ`����V���������2��YK�Ii��(�|Jo6���S��ӟL7��\0�<F ���N	��&Rñ��L��u���� �O(�ig���J���y��lC"�3�>A�fP|?�AB8�Al�IB��N��o��ە�Nm!�'{@��g��_)�Ye�Z����z��
-��F�>CyI��ᶾp���;����mlJaO*�;��*~�cOl8k'$�ւ(Y����K�!c��Kw�Et�uZ�a`�� z�@�� �}n��ڕ�C�x��R�sR�񝒡H ���k*�eɧ�I|�^�p�L~�˛l�\,��h<��쇹[<ٿc�k�^i�w\՜�A,88��j�ɯ	4о�ʷ���_�i��w�o�o���/�R�-����G�^������#N
P��)��c������
NE�D���u��b�Ɍ�����Oz57=@�������.cz���x5 5��0����.��D�k��<�.W���
%Lf=��8��q�ю#�G�ͦ=��E
�q�|磊<��}�j�i*���������:�?ñj���g0w[I����U��k` �C��Z C���	�ʰ~��/��D{gQ/t[ a�E�Ñ����b⒌vWsc�N!�`��7�����fe�I�Q^m�Z뵞}����p�=���ů_�dcNүƸY������O��^���պ��6<��k#�Ҟ,w�h��ha'���BbX	-^(�v��m���äЊ�%�X81���+1���J�o���V��U;I��`ƫ&���`JV�,��2�8���^PoS���OӢ��WT.M�'>��}�4�K�k���U��b���m��I��g���b��e8f��ݸi��|�n G��S{Sa�+�F��n����$v8u붆���m>��PlsO�@kD�S.m�a��s���Q."Z��f5��(ŧ� ����,PP��%���nL~Z���C�����	}N��g�).!�q���h�Y!�>��k�~�8��6{/����t=�j���'}���r��d��E�"<.�#Q��L��wm~�. V&��_#�S�d4�x��� F@��V���.O�0��C���`�����Ʃ�����|�B��Lƙ����� O��8��ء���u���> �a\�X�a�o^�z��vx� |a��DS��/����+�/���H��Iit�%~&��'�ZJ.x��,�y��9"\g�z�Ὄ���a��."�-������w�,P��؉���L�}�4��y�'/�
�J!͵�U�0_�~ʄܤ$����Z[A�=�/�9�ߊ�l�M:���#�ɯ8	JN�y����
�q��2k(r�����$���c���=1y��Mҥ�r�Ī����(�� W*�徭I�u\��'0�[�QJ��?�b8>m�q^�[d�3�2�/���N��c��o�>4�_����m]�og���!~WsZf=/�
w����0o*,[I�U����_�y����Vt׭��۵�FZ?��ǧ�ȶ���]R	XCv�c��^7������A��>1�Y,����wS�����1`ɖ�z��;}M�Ū*���8��\j�R�z����R5	K�ēd�Ŭ�|������Im�Tؠ�A��3[/�[�%�zyh}�=S�&�C���۰�M����@{���P�\�i�-W��������E9-h63�����H� �L���f�M�s��"�Ȍ�v���'�ʯт;�ܜ�2)0� �?V���_5 �b��\JP��"�F��n�C%u��yzF	�� @��J,����7��u+�9����/)�`@�]���U�{�[��d�7h�����e�4/������AicD��h�/�h�e��}u���Q241���JG `CRk�1�Cn��F+�>�X�pY��0$����� �����i��O�Qޢ��a��F�	�P/b�OZ�T�?�Z3�g'J��9t~�d\�FY��c�1Ӂ�^WY���$i��_L-<`�t�	2C`D��9���<�ʐ�?�uE7U��d'������Q���9�|�-�͈f�>`�!O)��Grg9n�
 Z'`	h�
��.%��<?W���\k�2g@ᾱF����gY��4l9U����΢߾����cT�N2�x)+�o~~儿�:�Su{ڼ��i��B�%:E'Z܁iU����>2g�E�~<��y�<����A1��1JW�[��yH�J�Q�=s��@'��i=bg���܎}}�<v�0�L|Q�W��ᙼ�,�,��r��&����Zٽ��ҷ�?�D|�m@�sN�!�ۢc� ����a���*�.9�R/Ui�\пq�ۢ�J{�W���\«%��RX���Q|���1��S;-7�靰�P# �E�xGU��f�>v\n���Li�F�}W-�+��ɾB���q�� ��8���|Q<��f�m��u���[�@����oع�KW�#�̪1�8��;[w�t���B6r9����~)�!T�.�x�I�rt;}7�:��m�у�p`��܂�KO��`"gX��;XUOX�l���4��ɽMB�,�p�Y��8��)���c�Mq��w�������M;�:Qe��ˁ��J��o��0R~���CX.٭`�@�{2 �3p�f�=2tK����t�����c��#xttk�����2y�}�bXQą��`R�=x9 ��bJ����i'��~�H��XD-j����4��]��llP�E؏;�������XQǼ��������- ���C�&�jj�ps�L�W �N�`|i�(���w6��a�9�#lx��$�X��n��N�C�ϰ��?��O�G�4����g�̝7�S�*n!�7	X�!��?sۢ����<���W ��E�?����̕A�i�`tqO�Mcxj4,�6L{ch�s\�|�4־@�௯x�wߓ�3rc��MQV�	�Y��.�2�����M�UH������-�]V\a��As���N��PX��XM�~<�S�QC��)Y�u�V��1����W
>����6S	�����6`�NF�ҹb8r�Б&�1S�*lhH�l�Z�]��͸�Q�8�E.�U��wZFać��՗�6�nS�£��4��7؋�޹-�c9դbd]�L�XD9x�{�^�����5���L��$�N�ml��Ҹx����_������x��:��׆�����Qr[X��mH����n���v�ok�f��hxLI��85fo&�f�>���(j��-�r�A%������~�D�WYM�VH�s��?՜�K��@VȦ���z�G�� W�3a[B�M��eʵ��P�,~����M�Bw����ɓ��\�ڔ�g<��U�_�,����/��?��ӿ@��U�g��`n����!���S]���]�C���1')5q[$�x�K�G��a���c��p䲶8ݴ�R�v�ƽ?����~���:YQ�ӆ$J�����ty�R�'�+vs}0�d�-�:sO7�F�&��d_���-�	A�w���9�s�/�u�(Ym�c�Q�6�9��p�����"�Ƚ$�*t^��L)��utɓ�rM�Xw�HgH1�P��A!'�p�L�k��t�^"�~��Q�H����@"�2�#�k�������0���M�������.��I�˱J�WSG�b��[�� ��Z�l�~��W@�1�o�ȟ�i�l��#l���Wz�_F{�U�8t��@L�+P.��Ö�1|t0@o�����W�]�T!�L`5\3��>-�V�>��%aD�8��F1C]}�NR5��3�^���C&�i�c)��`�/�t�RE�