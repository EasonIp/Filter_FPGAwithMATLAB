��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>� 0�ʪ�c�}@�+W���#��Uj��mrϐםv�����%�͂�c���&��iUd]�)Ve��,� ��$�aWg%��4�J5�W�y��(�>	_�3��_��HV�x�Y�κ͑ԧ���.��1..PeZ�9�X��W�w��K�d���Χ�f m�ԾT�T��M�[/?� �H��������+��j|�\�έng����~������J!)ej��gl�*')�K�N+�$�L�U�/͈x}�nk�U���i�xÅ
e�.�Vq.P�}ڦߟtt�M�;���s���1������ �4�.����[�5=��c����u9��J��$�._�B�fi|�.�Y-m�k�8� _$�������MT�>�nhϺo(�뜊�ۃ�I.�^���1w�%����K�/�Y�7��Xm��kN� %�6�����a���vQ��9�rb�N�U�_|�E�;U�9L��x���)�Q������T{�&�`�\�w�����AU?m9#'��UQR8��,�"s��9�6��n��'�lY��/��7Ѵ�������wv�K/��\s��g'v[��k�y�D��3��i �fO3�N��Ȫ�:��s@��"���m1=�"�e`NY*����|]╓�-$�y��\� 	Q>.-DG!{�W-T����'"Y�?�+d����m��X�: �3#��4���y�0����"����.�란266>����b�p��7T���B+������~"L���đ7B�C��g�Q��'�C�z�~��ʘ�Roi?�#���W>�ь��hɵ��L#ń�w��L�܊���XB>zg�U���\+:��4h��g�3�+(B�B����S�J�~����������|�ӶB�j{���t��RXܹ���i6޻A���:�Ma��%�����h��5� ZAw֨��hT���$m`��~�E�/?+7Y�߅a��a^B���"�y��Ɨ��z�ѐLR�-;s*�X!�-1%�.�T�ǈvA9b�"-D�L1V��4�d! 4b&�e���{�ߐy�.ᕾ֜�^�ԑT����V��ٔ�e���&=�J�!�]j��|�84��L�\�P�t�}�[���X�4�}kY��4B�a�WG�FR�e��e�� <~A���AS�����>E���<��]������c�*Y^z��S��1d[�]�$7K�%�m$��t͒�7�t��d��py��:�����{�=����g���-�*-d�D�"�2��d�#@��ܖ�Lɲ�X3'3ږ_�vb�����LUWv�6�;���A��SF�ꦌ�%��ߤ��g������ՙ��	��^�}&��W��=���~9��51�A�{��I�N���j#2� �����~����[$�_u�*��iq`��RHL��=�?����l&H��j�l���,G�8?u�Y�N��������AiS���DBh�k;���?zk���gf��܁0gv���u�U�C:�w���oW?Q{b7�a�d��јoV\�6�s]��L2M�C���]��k/H@���S��	���G���导��"��k�"}���q��*���ߩgq}��j�-��/B��߹q�����s�K�E��J���'^��.�j:&amfq5�#N]��o�+��Y��D�uT���q־��W�� �=gN"��X���M������:?�Й 7�݀�^���6�(�L��*[�j�ŉ���`T�J���ȇU!�G>�&����?�i��K�-�y0hΌl�xn�@*��¢�K��:�Pw��E��� �W���B�$��j�Y@ł2�hwLBm�;�^���Jǔ�K���Q���l+4ímӖk�R�?le 7ب���O��K�̬�2ʃ��+�ɴ:n"�=Êv��a _G<�Q����i<b)�--T����[�~��铀���W����~k	�j�s���A}e)���qo�ђ&��j>8�Ey���|��Z`.2\T�f-�}�ړz��ȯH'|�V��������P�MX��Q�\�搾�V���|��ȀTe�O$bƟ9�ĔR�b���v�Td�zŹ�"�3�{ҏ�d���:���u֑3��[�ܙ�ȱ_���eA�v`yf�\�+���U�����B��dK���]��>7���p+޼ց�¹a���w.����a0��~G;�$jar���|����^w�D���ecp�\%yQ�}SM�Y�y(�r��A��x	Y��T1t��&����Z&{�]��cIgHu5�i��.���;����`���7Z-sR�8*����5==���M�K���Ӈ-�-B~�-��|��.� �hק� �Z�`p}S�OZ�}�_�5�T����y{f�~s�'��� �e�����G�?O;M{�c��䋘���\�j��c�g�\r��h�*������g��*��Q�m��~X�?oh[n�=ej��$�^�ҿ"jXZF6�����=F�c�.���������R��	/�J59�g��;������m~�ff�L��B�	��dex���ŎZ�3�E���&_�|uj3i�Ǉ�"K̫��ۺ�̑W\N��m�+�o�a|�}Q"FM��#(<���t��*�Z��Fѥ����x:�b��@�/�% �"8�
�No4�7)�#�h9rNs�n#k�XyR�ˑ��i��?w�T���uR��Q6"e>�NH`2��.�!E������x;]��Fc�
w߄]�u0�1|G�}��S�U�����H� O�+y���y<OmC��ԉ� /%?%�$ܛ�n���Qnn�W�9��?>���:~���$/�Q�_	lkg���!5�����+*��Gs�6��z-W7X��0�^�"JQ�b5N�I͜�z{TP{�8���xY{�>(�4�e�	��=�-���C[�I�I�j���ga"�+ M-4v�9w�����
�G����"w����{�9�_�H��F�yHl@���B5s��AqY������O5
q�+��W�-�;y�3!J�Gi��Eh�/�U�%���G蒅V��,��,�$8�~*�g7��7mE:��ߗ�.�/笴kh��s�&X�o�=�j��"���O�5�pu=�3��^�ߧ5���b5���n�,��T�Î���āi���m�]��Y//�C�"�D���!�2}�$D�y�I)���i���5�?0`�7��>�G�Z��lu��R.(�����v�����NnUm����Ȟ�f�;�!z&�-��d�e�h���Gu�Ӥ��C�e�}t+n).�ʦ�e����<BȽ�E�:s ��3����L�@� �vW��:\�6I���f�0��d��ͭ�`M��W�h �;}a�3