��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�J��"4�=�7(�T�JѺ�ő��,\��s���ӣ�F�؏���5�u�%U��6F���[�?����
"<U)�O���а�˾cm�4{����E\�k�����֘������vOG�R
�Xp%�n���z�?^���X9�U���_ׯ�6�v�U���i�ݥ�'S/�I����(���;��<uC�o,�e�+��;��y��N�1#]me<���c�#|
a1��ɐP�F�����z�{�OW�/d�A�gޕ��\}�Y�I�e�Ԑ��`�P�ΚB ��#��	���_��qU]y��Z4A�U���'��5�Z_��R�����d|�E)*�l�� ����湴��y,Xv��j[$�h�����)�8�L��߻��`��g�M����#�� �y�@�8���(����o=�>������#�&_���y�u'qM�^5�6!���D~�{^N������}�Ф.ot�@�ؒ+c'w�.��@|�r:\����5ҙ�l�O}}������D�=Yf�u����.�,v֮J[�*G:���ݗrfh�󁹱7[����	����+ߊ�]�-խ���0�@���}�$`m��k�z�R(�E[�w�
ƿM�Lɼ0��gufBx<�z���۽�圝�t��&�bk��W����d�a���j*SW�?`�P�����竹�p�r�$s^��2�s���З�D9r�\���3*İ��Z�FN�ۄ��sĹQ��J��!]q�/��!�〴�i�F^T�;6 I���Y�����Ov����L�a2&�:[hSȺ���/ܖ�!"�oC�o��m������(�%g���G�|,�LH߹yQQ�ҧ�8o%��1��Iٷ�pT����k��8�ܠrz&f�}��7����T��*Я�v�J�8!����E��)��|d�F��8�$�>O�+tT~��i���ޫ������RP�����c)	$�z*�ZIϴ)�fa��t��<T�>��Q�_F-W���W�fV� �]M9�U~��Mx�����Ywy$�&A$E6�V���E��2���#L����Ē�| �$�?�V@=�9-9
]&Z���d��7V�+�ju�sPm[r�z�f�-���F��?��#����6'���K��8�n������8KľtC� ��i�	�H�5X̞��Ց���wWC�>�9�\��'�D��Bs����B��F�����p�_��|����Dkr����쥟h,��p%���=�_��_��3��̀��đ�j�o-��Q��3����6�O!����O�,0�9�4� y��N�:�]�Qj~���B��[��W�����G+����9ɸB�*��(�#�"S��`^'m(Ҷ��)�Y@r�T�2������Y
fg��r��j�y�vr�HB�Bա�[�"��Ir
G�
����L�t1�L��ƒ�z��ٺ�ܧ?<�~�1=�]����9l�4-10�� ��	[l�t7i��q$����j�����ƭSd�`��7���DFX�}F���U�Ӌ9��e�uN�)��Lݖ�*J�xENK+��
���Yl˄Ҭ�j��%�� >؞Dc�*�M��a�Qޡ�l^����͆�O��d�Lߞ�8ʩ]Q�=~>�BN���C�� ��L��XՌ/�T';�~�H���x*C(��� 7�7��iSb���/sS��޳M�@R _���>��d���y����z�����L�фu6/ �7�K%���T�M���@�f�;��nK�==sV��M�4�'��Jhߊ��EAF#���%���=�(������mN�#�|��`ֆS]����m���|�����e�#Q�+T�#<V���f�?���Yf�D
,��׉]�6֗@��t)�˟���>"ɡ�s=~�G���N9|k���jGW=���fR�ϵe7��z��C�0�(��Djե+'���a��g��+��� E���p��CI��8��M� �)�:A��^I9n�7��i���\�x߻��N6aǂ&e	vO�k|���Ӱ��8�.�)�F�e�Q�4m�kA�ҝ�n&�}��i�D���xC���@ZS��;����'��U�+���\Xe�=#����G���u�&�S�ufpP|�{ޫ���y��0&�"��N�'������,@���Pt?�����'ǽ.�ae@��ܦ�H�,�ժ�gA�>Q�5�:���s��6�
��RT�5�8���)����r񙍭�)��At�˼�ϓ����������i1,�f���?�w���:�ٲ���6BϺ�SB4����ھ�!���M�0N2����9i�o�B2p��X�ޡgX�5V`~R�Qv*XEP�}� i춥�E5�TRO_�.%e�?RZu�_Wg�H�LX2nLl*���qO�}Kh�����t9�7�F�"�ћq��z<���ā�d�H0��O��~�?]h�ױ�.
Kԋ3Ef�*�L�|z7K�'�+r	D'�
7|S�od��cdR�6��}�M7>� �4t%��nMr~7������w�ǌ!E����r����3�&Ȭ��5�
U�rj�9��������]i����(�j\�"j�J��h�9t�b�"ʡ`|Mw�	1���i73��~JJ/�\ $r��<X�P��s>��ّ��R&2r���(\���������
����Z�_�$�Ƨ�Y%M��Xܐ�~6��vϓ���0`K��| �='|�Wp%�=�S(xp�
��ԋ�U!m>��,i����C��?$`@�N��"/�g�.�
��c��U�a3~3 ����V~����qe�4�x#hQu2kY��F����l��z���m��4�TD7��ӭ�{�7�;�.�	G]'ȇ�-xNf)�۫ś�I�G*�?Lb>( !v
:��)evK.� y����7�g_[�-Xl���l;]���ı�=��*Lc����M��=w�S�?��� �g��P6*��bPTtN�?��w6QA��<�{�DJ�YŽ���_���7K �� �A4���)b~�֌��F�ۍ��!=1�|~F�R���.�J��l߶?6�g�[�,���g�cY�%��yk�*�?K�guK����ʹ��ࣸ��s��*��g��z˕솟�-&c��R;r\�J�� dl�r���$���rs���F�%$�'���Z�<�_���g��&��P�~U̍_~�Bj�PvY���E���̎���X19���R��jg������q�ʝU�v�k��A��o���n�{��h��)4��%z'��U��ɵ��&G��e;�?I�<f;=�ݹZ�0k*s����� �!U�X�8�0gum�Q�����D�z�����c�̖h-@�1e, ^J�����uId�
3�S�5?�)Z������xާ��`M%����d�-�/¨����3�D=�5��3�׌ۃ=�X�rw�.hcp�V���������Dh�v�kc���,������W��W�x5�;�x~.�n�~��ul��d��%	ײ�)��s��z�CJ�ss0`E���O�E���d��`
�����0��v�?_� �3�E���6D��*|��i 2kXZ*��j��>7����b"1���q�\u�#ϗ匓�Σ�>QҺ��ܢMv��S+�A<���+W�O8�:B�>Ս+�����fڗ�����V�ƥ���ِ�/|h[����� =��Ә���$s�稨���s6v��wT�?t� ���sC,��q�Ov�����琀R��hU�';���<�F����J��ڙ�EM���y�ka�!IXf�|�����j�s�r]�R��ì��J!!d ��N:m�c~7��Y�����&�:���X-^���Y�w[ig��vq��|U H����(��)��T��bp�:��v�l�V,7�ND�|c�;;.��7j�+�b7)�*y�:�N	:t*F7Oԣ�`����Gj(�ՖA5/3w,���x�$*�KMЊ^���ju�84��8��6��M|<j\��su1K�f �<��y��]��@��&�R�@��(hC5�e;��23�7���Ϩ���t���6>��ݛ�ĐG�g,:P�h�@*YԈ'|��h� �	L��ZqV���u����耀�r\��
��XжÒh�Р(:g��e�#)?��5P��}W]s>1�x��|�жn�;I��\igT��q��IG��d�Jw���C��-�0��zغ����A�f����*��=�H����}����.�uq'�Gؠz��u4������5��tK�.�|������&G ],��wm���d��k���b/R�tϷ�NWl5L����y ��o����u�/$>�I%�GM7)[��!�屇][�M��ݘ��Z�[jB;�"��B��\v�h)�Rf:h���u�����3c��b�C�Bp��w�N�[ ��Hײ���� �b�M�c�y�2�D*%/�^!�+��	�1�(��	�6ۧPU��v������}~�Y[�y""�!���w����W��{(�^�fU�g�mv{cr�(uZU0����n�d"up�V�� N]�ͨ^��%�2 ^s�Pǅ#��KB��T�N䙣Z@E#y�$����A8(DC��h��rq�-��Miw2Kr�%T0b����	��qu��9�>۳�.V�P�=/?�U0&g;�ܭ��+��}0Y������(�BR
��D�֟��l k�<���o�5��Bv����3'�}2c櫵�!��)�EBEq�%��1{� �ul��g�wR�S�U��:f
* G�f�H/��U�kqV�IA�'��^Rfxj̨�����-�xK����t�B��Uߓ� �l���T��i�a�U���u��P5�Yϳ)�8	�	���9A�@��=�	wu���v��%�AxD����/����Ɓ;)|�'�1OsZ����������\W���W��\������&�A�f�wВ��;�J��s ��6[^H}��a�s1�;�+v7���[{\�x<ːP}@Lk���On��C���"�	M�2�n?O��sֺ��>�X%4��!d�\�$�¢���5� "`�`)C�`7���I#��� Ҵ�Ԇl�jx�e�7�yg�����
Eӝ��ѢV\��h(��x��fN�$���NO���llpth� Z��EjB��TH��M��b#b����l2�4��p}s��Cx;���O�w?6��]�v���t_xC�l�B3'k)U�����Ud}ap�O����L������4;����FYl-V��:��	���X�l�c�N�5<�7��ftA5���us�j��� �oD���Rc���%Z���`�x~��(��ΨS1<��O
&.�N���Ցgy�kj/w�-hŚ�8_���FS�G]���Cn�o�,��͸xL� ��+��>,f �J�5�����Gw�;ǫ��<��pSXOe������o�t$􏞂̸����Eف��a��P�2

����{�Hm1�::p�
ʂƿv�.n�=:p�N:{&��u�D�z:����^byWS�C^������<����~}� پ7n1Mּ�l`�2`��������[��O�G%�>����r	ፅ���H�;A�Q���E���9G*�� w��r��c����~�6v���-!���9(v�jp�i����I��T���!DWJ���-�jd�xX����|狕��8��;HW��t6�!o�&�q���0޲K{�8j������w��*}��?�ej���
i�fb�����t=60-jliO�TE�Cy$x��[���ď]S;������
03*h���N��`MzN�yl�;�|�e����Zܯ�;�u�.!�c��F2;���#��7�����R�&�ϰ�Az�':�6�K�q_-��������x��V�vw!��O���Mm�ψ��R��H�)�h��_'oe�C������D�O�V>�d�/by�_�'뗗^c����%��bGȎẬ2�Dn^�}�̈�9V�w�9Fz�W˰�4<a~/L��Ԫ.�,]���J+(DĎNV&�B�l��;�A��u`6�VMP�,wRx��r��:���+(R�����~5��nB���c���&��&�,�����&�$��K�1x�3�i��K�
�����~�?�k��&Nlݍ��2mS��TN������ ����>����B�pCFB�r�ʡP��W�_6(Cy�6R6��Bq��l��e�U��7�l�!�\|�G�=T��q�X2�@05��)㗆�h!61�lT�����G ��r8u�#�ߘ^0����p\��߸t��1�8�����.hk�n��)8N<��ḡ�ᅐ�9��RK�>�#�D�7��JJ��&�� ¡��{�oL �U=zɴu �܏n��~J�3�`A�M�=��j��H�Cc�(Dd�0J�OaIb]M�����WN6u�g�)�.�z����r.$?ˆu�}o����~G7�{]5�h�Z`�Ÿ�^�TJa�hZ\�o��\�B=_��_�V�5�=�8|�d�X��q�r���e�	a)E���.]>���7.I�ǻ�ݲ��	�xUl��hl�o�Ш���kmڼ���Wv�n\�W���W�Ћ��*0���ƕ^�%�<5��U���5f��}r���@�ـ:{���2ۗ�h=�t�P5��F�J��H697Gg�f�;��#b�(tT�n����d�
 
�E%��W�|��A��J��V�Z�L��E)��s�>��4q�La_�ό4i���x&�TJZm�WF�>�㟕a��̓�o����"���~?|~���U�\g�a�����L' <y���9����m��a�VJR�^� ���Uu���R�kdd=0��y����~�<	]aN��}�A|-��󋝈�c���@zK�b��+�*fzӉ�,�z)�I~")s�tYq�^*r*��X����.��<�6*�\ �� 0XK�K�s�y%�1��j����"��fV�<J���-w_�%���S붪J�bt�fp|-
���4��q���<	�c99�ixȡ�_�´����$�R�U����Yx+�|�L-�X���Fjv&��,�MS�R\��#��_u1�2&7$,��;B�[�'9T5:|�b8�\�a�
r��Bʾ��q@�n�9�2�"��]��[#$3��ཉ ��{��0<_��B�\�GD1�ܐש��V�2a��ԕ]�9�I��(+;bs*�#�2z�x׌�Nl
2j���I���rFk�&�Ro���S�p)��� s(��9����|m�����z���U�����㵮�c�n�I��� �S�jWr�1������R6twn�P�������{l1���lQg�S"Nxk�!9�U5���d>=ok�̷��<o,"r��}~�"�Sh~��_��~�ٕ���P+�`t���Q�����Q���	A|�_n�>;�A��m�U�.j`]^����jw���\B����t;����;�,U9��N  ��=�X�"�䞭�0��ۚsul�V�t�������o�Zo�˂��z�aá�+'�=g���D�N^����*F��z�y��~\��m%r��y����o�Gq���[w�g�R_;�R:�D'�p�sB�:��g���M�(L��X-q��z�/�{��S������W�n`Vj�g4y�v�i��[y��:{�>>���� ��и.q4�4��]��Hkی=�Z�!9���<��Ղ��_`W�����!�8t֗���\�{
G,����1����R�b��脤�1�.ME���6n��GF�%�ۋ(�m��曧+&DE#$�v�+�J�"�T��O,�AoeTH�>ݎ���e��F��6������q�Ƚgl�K3#(=�w���Zo,���&��vB�BO/h��◦��|�x����Ҷ�X�]���G�G�6?b�_9{�aC�Uf� {�+�<��c��Ԣ�~��`�e�߇�ݪ��Y9� /��S�PF�!|��Bi0gHƪf
��n�ϥ��۬�㢊��*Y�]Z,դ��T��Od���E�*,��x���|cY��%�[�\K���h�a�2����w_�����j����H��֗��%~�{6^�B�,�Bֹ�4��ϣR����3�v�ql�N��Bx��Ծ\RX�?į6q��%+适C�ڏ�(��X~3��_�?��>�h��Q��w��\US`e�J������d\8�6��7�x�*�^�L��e�Y���w��/��w��`)�*�6����Ί��Cw������X.��j��t��}�U-K�`�dp��Z��w r��dY��������^�
~v�'�X+*nlۺU޳rk^�l�R�ї(Kf-�ԃZx�g-��B�a��a���%ԁ
�8����m	l�f���ܹ�4hǄ<%�O�� |���f+�a��t�����!.(��}KRt�K7�g珺s39��&?UD&$!��ҕ�Z(VjE�ۭ��==�s1z[���oRM�[�+Uy�zH�h�T���\�qh�����m�ɜ}��,����`�ô�Y���~��D
��D�B�ҧYqpbg���U#�]{��J���e@}��!��A���`�c	Y�9�%C3ᯯ������6�N�e��6!��H^a�C^�Λ*\#��d��$f���*�(����+���?q�<e<v���$��!n�:$�t���;S�/D���ڃ��l�E��r6)cl��R��$�U7�ο�j���
`\�t
��5��<�q/H�ɉ`G&[ۯ]_�5���8VW�Ëa�@�� ��Eg�K�8�� .n^)��m4�p߀}����U�_��Jc�=Nu�*��A�4�hd�k��S�I�6rx����G�����Y�^ e�ڽ����;�f����L�G�6y'�|kܧ� ����dfE�صZ��zlҵU�^��4WWi �����;�p5��T����J�,��tQ�KJ�,�,w�9Z/�������R&�r�T���� F�f�W
�3��g$�[���1���j���]iI��<��� �?虦t�|ߦM�/e������<�OVr'H�|�����$�d�a4��I �(�?�v_��J�7ҩ.�4O|��`���D>M��'��Ĺ�{ڷf�6���O�+X�ȥpp�T掐{���������a�����^�����[<X~*e�4_ �r�kk$����na�gĜ���1	��!��'���
���}��%�N
�V!w��I<�X�zt�
�xij�,0�a]I�6#+fVy	�.
��bɫ��-uP����E9-���!�xp�5�O�^�bXzl�"8j�PpR	������+��~r�k�K���U��I�D��#�C�6��3	��	���ߏ��ŦNs��F~�u�����@��搦�Ү�^Ĭ�k���/<1��y��u�&��?�Ƶ�7�<M^�,���&�ݶ��U�/>Q.�#f�)�^�W7�&L��3�+#�ywo��,�1ѷixn��f�6�esw���w�V�7R����,��vh�i5-^u�����fs��(�N�"2h���ȳe�e��6y�H��r��qUw����&�=�p6Ǽ�,Vl"��o+[���a6�n���2�Q��
fn�,����P~�pcuy�+�T�Y�.,�$�J��k雕p@�p�Dcd6̊�_��q�I�Ѣ�i}��)!q��S)��l+7we�~^ؒ���;r���w3"���6��W��E�Ffp�B* �(��0�S��>�/��o�W�W��Y��K�O|�3�
ym��qR#@lR�����K�����Z�9DL��	�%�W{C������=���cFk.�����K�|���\�jlK�v��8�|C���M!T�9b� :��c�fCmks�M5w�]��G�t0����i]1Y/0�R7i��ď���>\4���P.�L,��)�oh�4674uJA��Sc ��6������<~N�8���a8�D�֨�~�rUA�rMJv,[ͽ���ߗ8z����|2@�YBD����L;�_��s#�}��>t��p�8�����I�g�旆z̕���[OP���F��@;&b�,�Gg�����^��7� �pv�῀E>hᮐ�ܙPŕ ��8d���~�ct� ���wg�0;1��V/4�� ���z������g�jZX��L���1��V&O�>��q,�	*Ȝ����u�{�}��^B�V��j+���]�p�i]&'���r����L�O:�b_j�Y'�x��%K���1�نu�����\��VU��m�5谊�6�#��s����xlj	ڬ&4"xQj*�Ք��A:�(���2���V�uv�߆�oa�I)e�,������rZ5�(����K��h(EQ+�sA'�/���*���e�N�ڌ��ć��$n�<�o��;fu���/��.�mDc���^-X����2D�3���G��������^�������������3iD�_�����({<�=1�3A�_�J��%6G��Y����6h����̹�N�L2��eI]IΩ�R��B�s#J���SY�P�I^�W1�Б�k�͙��zu��~rg6����������IRhd�P9e��9�O^~�O�OJ5����[�B�%
�n�lB��A��s�M0ݨ�Zk����*CKC��]��)*M���66)�1��ี���r��J�k[6�H6	`�np�o7��<��p!�H������#���=�����+O ^��^�<$	��RHf�����-��H��ǀ'�{�r>�U���q�9��d��#k.��0���~��Ѝ�w&*��6������ŲHyk�N��o�����&��O|�!�,>6X\R��η�<���&w��X���mǴ��WL���"�fRq0�<S-]	����a���?�lu������k�b�cO�����;���d���7X��r:�\D^�@��h�����m�N�W�{�!�ǧ��q,장���<���s�"񞗝�,4�L^�z��c�~s���Ŭ��a�6��VK����5�Z2X4:��|��$��h����5���� 5E�3D�N��ּ��_��e��B,w�~��Ș�s�t;�2V���e�0���� �h��**����1�KQ�Y{#��V�������>kp!x`ij8 ����Z�O�`���H!��h���V��*���Rd�]�59�B���N	�h�0������m^;���t;�Q�
-t�E��n��=Cz��3?����Y��&���b��������сg�QW��0'u��;*����ɽ�[�v�^�z��׋����ԶE ,�3��-�a�V�����$i��@�I���8,���b6��odg��LC�ӑ�)d��f��9��Z:Ծ�m����شin25��ȑ�ІX�������&�f�lo�ғ���ť˸����8�OM;wK���۶�ݦ����b��Հ�9�[��OL �uK���42�+��0Ё�)A�WW^��Jrv��[4-W�i��{9��*���8�r���a�fn#xv�h�IV�D�#%@`�Zt���)y#<��T��ّe�u�b�#��J�cW�0��+��4���L9zd��묮(����rܳ��+Ba�ҋ��g�$����o�^�����/Lh���O����*�[��xC�`�\��c���^���?����NV�T�z��ָ�:_���h����E&�X]�2���+w��*�~�ˌxane���n=gr,/^�}���)�O��k0�P#��bG��×3����ʈ��>��`oF�4�ӳ�J)�'��uavza{��$����l>&t���rτJb�t˥��&/#"���H6L7d��$E���k�al��ā|�J�k_`*����#�-Z��#f�W���d5�����6�yyP���{
LJBВb�ܞќ��m��;Y�-Y_UZ��(�*	%4\9�q1�	fz*N��i�F�,@Q��[����T��i�AK9�#n�x$ o-_,W1��0��x���;Ma,��z@��a�'�~9a2WT�N8.[��v3����)�	��O 
\�_L��=�����G�Y�Tva=!
Y̾���Pp5�L����QE�h�8����v� #q�(�b�B#��f�����B*Ϡ&O��>\h\x�_��[�w�Mx����T��xѰd�O�&� I�-o�$�[��Z�P�v+��ٓٓA�ʫ1��r�9�����3L1�/�`!jܼ���E�F�[�(���O�ſڤ���[V�fQ;.4arr��ͩ3D�7�O��U���wUp�I����l�s���,Ն�`�W�ٵ��G淨�K�%�7q2�J0X��ͬ��=7��`��|���K��~"��زE:���ŀ�C�c�{��]"�Qhy�.�-�IV5�,誩��g����%�������iH� ̮���O�?���En'�����LBv6�[��[7P�mЀ���F�Ɣ^�������uV���T��|�R[� �B�h�[�܃;0q��M�H�&o�'w�ݼ��"��F���E��ۜ�DUU�4�VG�xf�����v[�^ѱ���W� %�_�Pڭ���I�������G���N��p�����5�o;�j*X��xe�P��R�^-���I��l55tti`�r��t>/0�~RPN]�)�DĘRW�7L��x��G����K={�w�� �Se�m_�[-��
=�oHp)?g���#1C��	�������H̦�
��]($��U8�IM�2e}r���'���Yy�*�[g2�%�1�6nb�H㩣Z@]�*]�+�u%EhZ:�-7�y�%�CBJ5�l��;�m$�%;fZ��w�G�B�b�ZC���:��:f� F$�N��Gk�j���u']�(���`��Z��L=d��|��v�����yV�5���1�Z����.&��Cs��ys	�������$�	�YT�I=��P@Ի��p�3��厌!�=*îW��-� JK���l��J��aT+k��&LY��P8���nx����!���\��j�:AQ���
p"�oJ���k�.��&~V�ȚG�#�\^ꓬ8�����s��=U�QI�R=�*jl���Q��d�h���H������x<��O"m�̛�62dh��п��R-��h��>Ku�a�Z��3<f\uBr��LF���֋� ���s�w�<ɚND)>��;}6gI��jS��!�W઺F,#9-��)�awJ�Y�˼}��|��ǀ�QA�����U���`�ւ�h���8�}gN	R��3}�!@'fԅW�w[���K�O�u*�([�$��-���b/+~�ݐ����ij"�?�?��/��l�Y5|D�P�ǲ7:�9Mt���R[qD�ݚlФJ�[��!�EI=�5u ��<)�_�tZN���k��7�M���͠��x
vϐ\4m=�nP�����y6_�~�n*#ˎҶ2�Hp8 �4�ތR��@��nWZ'G�轚���^j��s%��LPQoO�b�o�0{(��F���l��N&�p�B�����|V1�.�VqQ�Ĭ�V`~T�1���yW��4�zT�z��e��ܝ�;sHH��'s��n�w���a��0�F�&~�¤J���9����<�%y���}���[Ν��������Ƣ�~"�����^q�H\�}KP�iJqR���|������}9y�����	�Q:lT�i�,���1ծ\d<9E}u�7y/Z�2��a�E�W�����Ͻ�&��B[�R��Hz��)�K`���)**�N���/��[�����[kk��߾�M�)\{0O&��e�����`-�Y�H����l��P�n�\~��� 4���E;I�̨�2�1TȨ N�'c�0�2h�oInu)T��i�zQz��/��?o����^g�=����z�u��U�J�1��4>���L�9�6�{�n���֖���V}
��Cr�WqNQ����aG�'V��7��b+�Aĩ�����G�p�ā�����*�^Q�!&+����jC��f��Ƕ�w��'���f�c�1u���|O���̮�����Їw�Pk!�/�َ2���32�=��P���FJ�ơM�5wǅv�e���г-���'Q�L��n�]q���>��~ @�.�t��[�x�w�y���A��X��q,~��)���'���f't���Z��� )0t'<�U�G�wTp˓����كZª[�a�������kMH���S��X�y�̘��'�z�0��̌��o���=�JS�
h���R���r��R�?��#��)ÉW�z��;�����7�2�L5�06^*+�S�@Ql�o� _�6����
&��W��>!���^��='����S�1R>���+:͟CvN.�
Yd]��7`j�	Q����U�P�>�)���[[�C�s�j���I�{�鬸)�y?��A�0��Lֶ��>P/j��E�N�܁��&�	:�zJ�������ϰ[٨.f�Ԝ���\(��U��McV U��9��>����D��SJ�Nߞ/�t��7P��Bw V�?^@�uC�$�V���.����y���}��c�[��+���&�q�@8�r�j��㚵�c4�9����fTڰ��� �1Z����y�N:9�� �aU�W�H�d&��Ü����RTb/"bi���αX��d�E���ES}+��BHD9� �'|Ehp�����X�z��fl��u�gڿ����l�&̏�A���ge�ິC~EmW�0^�V�R�N�� Zku*/գ�;��ͭ4 S���̆������26��z�����rWi�YC'�l/�`Gc�?��z���t��(D����J ���}��*�"#�%���fX-fg���[	+�	]u����.����g�:j�ٶ3DnZ��7����h������%//ЭZ�
�=x�dͪ�n��������Y�i�.��ޒm�Z0�x�a�H�Z蟱�f���-�8�2�b�5h%g��#T�3^r�2g���)�[uиh'��Of������[7�z��8��z�TsF�-+ݪ�=G��~���V����\���m��~r��z�W�����3ң�sx���/"	Qm�;��0�J��*g�޾��g��`BN����:�}�ܭ�$:�;G�HlU���3h61�Z��ϸ0o(lN[y����о鏪�g�W��l������O�`�S&��Ź��w6,ه��������Pf��쀍r�J�=`�ʖ%-�o�U
��@ib:�sT1��֍�qi�7��gV�ar��swE~HD���~02X�f>��P�К�$�<�����PA����~�3�VM�qyor���F��BdcG��䳛��Z)]]�|�=.�<0�[�Ę�[�M�;�^J����I�4�{��U�CCə�^̼R�v9%�1�%�-x��C���H�B~���W����	����;���6"�=�Նb:�^2�FZ#�;#�NRi�S|4�5!�+�g�����B������n.r9�b� M�K��r͔b�f7��(��/^"����Mn;��^���B�V%b'���!K�8��H�꯷S�G�G<��:%�i�1��Lp}A<�J$ݸy莚/,�@��.���ڈ�f4�X�P�T����>2^:ֻ��>F���m!֦��9-ݣջ��$�#�%��J�(e=�D�>�$BiU��/4$�=#������&��xfEj�}��;���������٧�x_�Z'��3�l�C"���&�4�$r�ԯ�n'���>���6	+h�\E�$�����E�cn �d'U/<�N�",D��
>���睝���b*ē��/R@���b���OQ��cW� ?u�7�{,xAƈ<�Ayݗ�ojb�;��v�#$c���|u�F��F��%vJ���� �a������*ޫ�u�&2o�N��KN�1�_���⍳�9y�N�!�jy��U��̔R����Le�&�*��H�2A����6�?�,�d�œ�Hӡ��З��lJ��aby���ċ��wwÉt��P.��̇��=[#u ����V���9����_B͒�t����	�5�����V��P���x�o|bvq����	]/���N��}���:���;�/���|��cvm�$ *����8,=mj�{�;��*�޳��o�Q@��N�O�����Va��70/Ph��������Cڠ<�L��U����LU u��pD:L�%��!S���8b�$<���.:d[�=�������
�|��yAX��"�
��9h
V��}��z}_��1
d�����2Z�L�)�n��~�C*�F%��e�ZR����/�����y�4��h�>[������&Ntl!3Yә�[wo \��3�CGjL���AN��ZP�ҍ�w ��A�&<x�TCPAm�f�� �7�!+3��L �~��+�Z�#:�I���J&f�\�t�ɹ>9_�|�W�[����gRgI����N�D��$��EU�{Mh:�ח(�x��(I>���e�d5�A����eU{U?��T��Ϊ�~"�߮E���[!���B`��$����,V��}��ar�U���m�� ���X�f_�W�T��1�c2]�Wz���0��{yłl	��jT��*	J��W�l	���P��t�t���*�m��mT��� �'&�seJ��`���$�Uf��w���I��Uǃ
 ;�H�/��q����yH�<w��P3[z��(���Δ�R��|��E��X��G^�г��a�aK/n58gtt��t3��b���":s�vCx��#$�q������$m|Hv� }��� EH�Zm�3���Ue��s���h-�`�7 x������i���.{h�0���4i���SI	BA�Z���O�^�iwUH��A��H���;#'�be�wM^(�w,6Aha���.�Pz����iD����O��9ߓJ�Ҙ�E���R�<�9��1�=[-� ����ոcG�����װ��"r�a6�p�i��A�_ į:fjꟋ����K����́�:�LN��4����pT_��R�9��{pln�0Dl�0����"w_RO��5�B������dn
Z�A
�)Q|���:���(:�߯JF��%%�hyS	�Y�c�:?|� K:T:��O�dgb��w��<�h\V(�*��s�3���yz^C�X�$V�qb�Z?�g�O����"�>�b��e�{]jU*j����o��5�}�E�)��4}�F�=UR����`�<u>�/,������+i��P+u�"�x�)�p�T�.�I=�yV�>P@�k��[��ki_�\�8�#ugs�� c�*ϝ;��t������ ����Hz"[��U�Am{J@��@�d��]��N�M2�ڛh�Oެ��lq�&mc��N������?�i���H�|dG*��.S;�rg\Cdr���f�f�J7���w/FJ�NN�^u��.��"��,�0�Yb��{a���gi"��p�Y!B�cu��V%2!��/u:����c�S��񜦹�)m��,uW�4�	�ljWC�7"�6��#ι~�洜��Â������R~�\ahl����hP��)q
ғ&Yn�Z}�<<�^�y�7	}sS��Y�S���'�t��+]��~MG5��2�B�pG�����3}v��A�qɵ�@�Ks��j�fP�XX�7��ԥHS�����|��\9�^ N�XT�T�-φ%m����;�=�4����N�>p��6�.�o0��8�� g?mxa�d�dQi�6�x=�+�7:�Kx&�/���K�ve��[-�>�ڈ�nL��n���jD��q#�j&�G;�8������c~:�}�����Z,��a�i�f@�4��#`��͐��o�`������yKY/鸁���:_C�h��ƾw�P�3ҷ-l�����O�sT5�۞g#~�? 	n)=�-�2|a����Q����.Ek��L���v����[	0e�X��6k��|T�h:V�Ϲ�^wQ��M��V�L%f��]���$P��Ppi	�N(0ֿ'�<8Z�9�H�--�rl�y�����f���:����H������qg�<ڹ��<�Q��+{�̥����>I�/�*����(l������YPfYvԫp��ց�܁�.Y2qu��T����^��F�h�+G���>`y�������ŹNi٥`9��0��|�ް��������0�0��A�<Ef_0���� 
�+��y�8!ߠ��[x it�hW�=����P��M^�˖�lok<�P\�,�i�ի��k��7�
���������/� 4����C��8zTbp�rUPj����T
��hcxjך(��������aօ�w]��&�)X�����f�O��*D;k�'�fuy1G�,YO�s���I����b/��c7-�N� 7j��BT���I=��N�Лf��V�4��+g9}�M��P��s0}�	g0ċ2�]3H��ԯ����p�D�9�e�tl�V��k�V���I�l��F %j��h���Z��wT�$
�tW��}Fy�XcA�����		 �Hb�I������%��Sz���j�ŋ��Sl8��d�`vl1 ��^�{#���������p�ʌ �J�Z����κUv���q@�V�ϱ��c&��
��@����]x���Gl�!�l�d;Ãʼ�]�9PQ�x+�'&j�)HV�IO�p�:�Lz��	-�� ���G��"��9�#���4.�J]zb�.����M�{�p\杺�mɰ&ŧT˖�Zv��M~���{|�aI�l�����0E�1�1N&hUO���8�K+3��3>�@��	����pB�H�-IBG�"� N��% :�,��$��,�>��Ɖ]3�2��7�������P�	���^c�#�f�f�?���0�\�~�U���5G1⿿�t N����i�/@����Q�8`);׻7��K���-t���A�Ѳ��ά�n#K����d��껣H��T͉�l\`�iZn���/��p;J!,Ź�[����B79��^)	:rZ������l]�*��فܘ�96oA�;�K�:�O����^�`�9�+�le.V�c�iO꤬q��U&�54��������k� �����H��rX��F$�å�{Wy��O�5��4���wov|[ �	� ��/�pV���to�71�_yߍ�9
Cz��C��P1���k�q?AŊ���=���d��m0s>�3��3���Àt�?G�=�s�Xe���>��@�*@ZQ��l4��㶧Z�� ��� ��L9t����vO���yJ8V�A��>uc�M�-BU�[�lF���sbd�Zڸ���� LV`=TBS*u��t�#{�JP�b�wmÀ ���1=�p7�հ�z͆6|��N����X{������t�s-wX���T�#�x�f���Ei�񟏷e��a�)��G�V�f��vK��6��@���`�F�Ё�IΠ�}h�k}��B���꘹�B���] ���ftĲ����t)1�wz�4�!Plb8�����<���ra��K���'*_j���|��aoD '��xd�1��x+SD�����Ja�{�8�~��e��V2�-]�9H8H��KN����åSGOoS�0mJ1;[U76��ң��ͯɁ@��������moU �~b���L���J`�1+���:܇�+�;�|q3m�Ε�V�!~߮�8n���~��t�R����\�:@�E�������B��Nп���A�B���:w$��s����>n|���
���͡)v̡.xj�( ��E��UDnh��k����KT/����J�����0���^#�;A�#��ܔj���>�5�_
(���o����a�׷}���p��$�^-���vy�'���r������s Z�k:��K� �U(�bsUBƩ��#\4�r���J�Y΋�apv�嫛�-]�3����A!j�
i]=� �ߞ���a���x?Doz,��os���v^ $�^��ݩ�vN�|0�K��,�i���i��5D��C�Ie� �G��Y���kG-��`�L�@��2G�>qG�v����{�{&�X�Ƅ�}->c��	�5��5���EBp�2����ۢԀ��;d�,�����>�n�;j�j��ɐ����Il�r�%���J�wr��'e�BE���{4$��I��u�J'�ym�����"���Whޡ�s1��=�sЯ���i����o��ϒb�G?�b%<�c�c&Ɗo�ks�8��rg�yЗ�4���
�I���:<��uW͹I����r�&��|��F]7x�L�[��ũ�[�$Q���3�EOu�4����U��<4�����]�Ս�����_�+�5L��-�O�g�=�B�@�~���K`��_��l\B�;�q���/�Ƌ�
eʈ��hN��t@���dR]�<Ѓ��Rg��g�AR
 ���Ȑm��"Z�����{x�;?��?�ܳ�2n;[P�۫������>]�P'�i� ������>�����ȴ��_$�/]"��Lh��eGJn��bem,0$*c@��O޷� x#f��A��k��Gi��#�v愩k�E�	�0���\�Ñ��Z1��'�Q� ̖\Y��ٛ��&?|wV��x��M�4�w#k`����!��A��R�x�������y�6�{잣�dX�]XH-z��	L�mz~����ߊ>!N���#�AMFѰ����s$�j�+'���W�E�6]����0#0�M(*�\�=�������I�ϥ��A9l��ЅԿ^���魴f!���5�0O16����c�_��u&�'�o�d�h��ߵ�}L1����͇~�3����@�����.#އi��4�!���k�ztq��2�(}ꈮ�Y�CNͻW*�s���֢��7_�7��m���H�/6����&B�eW��[���$h���69��2�	�#���4*�1�-�M]�z�4����B��a_?�����p:P�B���u��_�D9o�ř{q�����)�ۢ@	���Ҳ}�#<�����!܂�]"�p1�]�.���Tp�Pv��[�u���+��RЧ�K�l�[���l�[���̶����݄��f�U���3�Y�ag
 M���mo=~�)�/�lӪ2�`+)JW@o��RcQ7�j�:=1��H!ˉ��I_7�����
 �?j<�v's�ٴY�}�x�p�8�'à��1cg���T�L�:�JQ�g/�@\�`�Лx�yT���FKg��$ݘ��t����R��N�\�(s�A���cFm��!�_��)�\�����Š��\�>8]�A�@9Y2h�u>4�V��D��KIt^E|�*q�7�t;�<���k6oJ��o3C�Ք��G�vI�����`EF��y#2�i��.��j*,D�i����B�XQW�.�y�
/A�[{ ��%�
�$�Y{�F;I?y#�R�#��\��u���aba~.{p�=�}M���&�b���y�)�	F3�� վ�T�}p姜b8�%��w#�-��B ���q�}���o[�d�Yԙ����I�IP����[������:(?g �8.�`�]��N��������ҝ��	�hG�ϔ)]6��`j����<�9%��Wp����!-��mÚ�s=�(B�fd������{����UF�9�:{#��ՂS|<DLy��w�{zx�բ�&M͠8�G�6�Dbh9/���5�:̳� �x�֣A�6�Q���u��^������=��&�(��C���t���D�sz�{��W�)c如MT����L[g�ɖ��\�F�>������K�������|V!�u/��!��JT���&_��})e��V�����}���2�]z�iN$���B��βd�z�n�j��%*CR�GR_���j���Ĥ�5�U@ȘK�5cD@����pc�t��ݮX�x�?�CM�h)����L���Qڒ�M�\�P*%̯[��`{%uI�1y��}���X�y��Ɂ����E�%G�=�%�G*
j�("��X�����P�DH���7��;�lt��Qe=�'��[{it#��ȑ�%��c�3�^�����-g.jj�(�	x���2qd:zLu߈��Х�v�V��?��7��ʋ�Ӵ$p&����E��03�!$
Lu/�_��W���0�>��%�wm�����GP��e
W��ߧ+�í�t��Q��d���הϷO�vP4jm�G�Gmi(��蚾���qԑ�ik@�ӪzS3��7<�m�1�R��g�{�D�����,�[1��"�Q�_r�>p�j���c�S�&k��Ap� �]��a0�t�4�{q)��2�>��⓳�ry��A�5�����]���27=�B���Z���?-4����\�Q�̔<������k+�k�G��C`z- ���y�\�]8�ueX|���JQ����_���QF��?Q$���* � %Q�Y��|o!�O�1��N۽�NِK�J#��v�z�)z��!�*E�~�]w�ћܒ����p.�QBORUF>j�$ ��tl~�(3��4k��P���3������Q�<J���GsMY�X.�����}&9P֯��P/ONN�plYA0G��:5���Uv-`b=I8|��������C�w�_�@'�	B<�F*�1��+]�CyTޕ^���s��UʭW����>�ˉ�h2_K[����C�;����h���T��s˅�g-9�9G? (�0B�;H��0�o�X��0c��*;	DJ����X��1]�y�8(3JL��b��0�<K_s�* @����g������s�����w��>6@-�;�d��v:����iz��VW'Js�iI���^�M���xICC�����!� Ԥe���$��jy;jH�)��Y[�.<&�d����0de�>OR�ȭ��!�!D.v�M +�/�g�-��uբR ������I�y�Գ~�R-jS1Ŷ��?�����%�G� x<랏c�s���<�W�AEX��q��;�!��
 �� �˛�Bd+�/�X4"2-I��2�����ˮz�(�"�7�Ӌh�P�����܎���$g#�B�Ahs"JWZ��$I�[2���1�k�if�!��X�A�i쾜�~�_��H?x�ɬ���5�<`�4|/�tb��&�mA�W���H|�O�����TmAG��sZ\g��h���H�p��>1���4%�j�9�w�VuX�(��P�RX��غ�ZwM��I����G�^?_'�^�g���о�QG.տ^R$<�$���^�;;��iq�-MlPeu��Z�k��߄����ɅNzf&[�\"ܒNx�|�Q8�����1SQ� �E���弬�i�fR�@�C��.�UDnn�̆h��}��{ą3nT�M"y�B��v��BNj��Jʊ��p������ʚ���W��o���EZ��*�5'�G	A�6�S�a���զ4���*r��Q�c�J�d��=���Z��~`ʱ:�اFn�XKU���-Y���}�@Vƍ�=��4��>R
��0zbd;t���iI��]sz�1ڍ�� [���[qY��
��4!j�ɔ��d�[�<6�g��H��SP�'d�[�T{�p�|�b�H��N>	��E8U
�ot���MD���V�x�+�^EĂӇ�,�n�F<%�|=#��$�q2�F�M1s=P���Do�ߢmN����a����j�)"'�k؞�jw��uw �Ƽ)��ʄ&uJ�'��{:8��̐��0fg饇�2���5��|�$���;�g���5�D$�`��,K���q��3���7U������"�L�?���O�5�KY6CA"�@c��mи���`<rK�=��X��a�����O.�����g��ʕgY(=���m�d�e#�uӱ}|�Y4�}�f��3;=>�ߖ.L"�-�ޯ�M�ԝ$�v�E :p=L[����?�%4���X"�%�Dz�*��bf���%�D����rQ#:K�VN��y)�P��"�3-]
&/ċ�\]�6��}|�CF��a�{�AB杬���}��B� �i��&����դs]��NNh?]�0�ԍ�"�z�ĭ�@s�A;���,���	����.+7~߻u���o'��^&��éY�������l �Ŀ��w���1c����VC�ܱ��x�L(nT��&6_�Vw|��q�3v�U�o�V�	Aa��l���ը?$�Ve9�L��0���YICD�G�U}$Ѵ	����8i�v����Y����i������c�� lF�P���1�}�UL`q�
!o���aO��]Ah-�xm=H���)3K^��J�=z�z���	�������c����X9�1��`�֞f�k�.���iS*�LuS�U+�~�-E��j�w#����z�"�H-�	1�P��,x�0���T̲m&J �r��ֈ�5h��NSp��<�אԡ�.x�X�c��]�8�-'���)�J�ShJF4� �B�W93���������a�v�C&�M�&�'E>��:-�c{?^b����Pa(��V���A�'�Qw,q~[�5���!�G��e-Q���"p<j�ٌ+@=Xw蒂<�f��vܻ|�B�ý0��3+(b �tǺ-�?��
~�ȭCp���c�b�"��m��;m��<��0s`G��?2�Iv"Mt��kD���1P�&&�N�2�>��Lc�k� jF�ZRx��x�@���"��ufA��^o��a��飰�F�7�!�C�#h�?��:�hwRi9WӈyB�7�_�@����#�h��fW�/��}��Q�ߞR��2^�"�Y��k�xI��`Q!���{����y:���e���O�-o�n�5���+'�jO�+]�L	+�T��Bx�ݽU pkR*}ϤM��ɱ�K�Х�6�9lǦe�41As������p���xMT��^F;��ph��c?A�8i�@<`#�)*m������YUހU�'&N��O��NE�Ek>2�ڐS�(0xp�gl须uvlWNh
V- �/�h?EX`����Կw�S 8$1�찷4/��Q����{�p�ET��q�[G��<�k�6�����ყ�Z96I"�:���k��Z=ҌlIi5���"���q�CB�p�,M~�L �Kwֹ���I3�{l�}�MJ%���#�W[I�^g�J��/c�y�# ������,`�_bH��k'-�/�@_j�����KT����ɻZxQh����N[�s�Ъ����!N�x�p
i����W���-���u��0��� �@��^�!~T��,�k.�M���r�>a�����<���Yޠz�
���:H$E��P3!n����tA��))W��ā[�~�����$�E0�M�@O�L0M˖��l\��9���4>eU��q��:���b	1�Tk#E����t$?�Oy�x]�!����s*���9ҋ@�/@��ê�30tU�Nv�o�9�l@�y�M��N�4%p��io�M�՘��1/�/(��*�Բ��1�l(�ه��h����j��������&�\��^�ȋ�un~Ja7Z]s�������3�sW-r�6��*�[�����*U1��s��h�s�e�bޣY�p��#/^�7q�R˛k�1y&��,.(�g�O;e�H���gPAS��z�yذk#ш/Ik'X��`�L��Q>Zp1LٛP��!ʖa7.Ia�H���Ĕ���'�IR�?T���+��I.��%��]k�_;0ݢ�U��ā��#�������P@��㔾��'��Zy+���Zj� !|��~'�Ӟ͏���Z���� ́��3��z����e�/�t�2gy3�l5�u�bCܧ�1�Z�ĥK��+�߲ćp)Р��%|����Hq(��b�O
�eF��.�-+����0�{ʶ�_Q%�F�)�t=�X��]��!��:���1��x�䂵�wQg�O�g�~���m�.�E5 �М	ƪ�q6�8�+��i���.�1���	����96�櫮�x��$GX�.��]�j����{@짦N9�t¶m������]L�8�)d�a&8�j3�b���3�|j-=�~98��3x�h������!��m�ԓ����� ����ߎ�j��M;�>>���!�$��<�}6���f��Ӕ���0�m��ږ7.��״�)�w
�q����RO?4��w����������)v���5<�I|�n!T��t�)�f:g��Q@{j$��.`�VN%T��UCBC�=����?%k��d�*VM��F�H��>���֞_瞦A=/�O&�Q7�I:�u�Aڄ�m�zH�!e/���LO���ѮJ�4��}:���:�b^�S�d���&���}J.�CvȰ
�\m;«녑_\o`
�K�y���$����k�|�k� ��Hg�ɅOf���1d���4.���{��Ʒi%��F ���W�\��vxq� hJ|[�2Ƿ��+G�`?o$k�|�ԧ|g�L��<��ifn1&*z���5��`m�;��qP����q��:��j2�:�kQ[,�R��?�Eq������f:��⏽Y���mz�J��$f�OD�'!�}A�!�{����~6��V����m�8ߟ�]��\L����;;�*&��<?Y�FxW���Kꨄhj�}B�sr��f��-r��{�Ծ�M��-��m�͡S�����{���{��]u��Zp�������Z��`�?&i��3y�쓥�.��iZv��m��U�d#SL���PO������iMw� �h�e�2��t���j̮ �9ls
śo��DVh!��)<Y#޺tT��������-A��e���݉�e_�,�k����N��#��;�u���;XW�������P;���<��_1��,8O�?�,H� W�K��3,z�7�n����E~��ᛒ�R���XC�U��@&�߱@9��DUf0,qK��vɻ�EH1�x]Y����~S�m��%��+�Q|�k$�L�	\�U�ct��˛ʽ,[�r�$Q斫z ���V6���n�2���-�ek�A�����ہ5��1���PO-G�D�0]}� �6��C����(8��3�cX�U�;��<�Y8����f&،0�؃a��}K&�/lsT��UX�������({��Ғ���'�),M��\3��T��eRq~9%����j��ikà�Ҋ�!��4�ȍ1�Y0{��P���B4� -��6"�c�n��~3�笄~_�%�lѢ�A��)�:a/.�h�=;���L�>Q�-j��G����Z��;�x�n�yoU�70�PtD�j��8�H"�7 ��'��+�Th�j��xZf���Ȧ"vJ�1��S�6	I�v�UN�O J�r����H��!>�Ԫ��z�Z~�o	Ʊ�-.[�Pr�y����@�o0y2����ʠ�5���q�b[~��9ۋ5D�!�^�����p������㙯ȯ����^n��f� q���c�,��5��f���F��L�H:��PY��^���3q�4n!x��kb���c���^/O6�����]��Nÿ�P]��`e͐^��2|�ұ�E*9$5{a�D�b3a�+�y&y�����>��5�+W�`�����A�6F������{�&_���vΐ�s�l�FC�; 4z��jHo(�:Z`��%B��Mn����/τ�:�L�̀����g��������%�	���.�.3G@u��s4!Wy���I�w5[���a�l��ʷa'�0t�g�?xfx�W;����Z`X���z�m����Ij��M�y(���f�<��i�кf����Ic{r`����K粓�3���s{ZD��7��[��<Z�q��k��q3q>W�A�Q�����Ԝ�hQ�PlW� -�z`ׄ`��{���ȞA4[�*_�#`��RpJɾ��4�者����.�vr���=�O`I̎�	���_�o�%�����S���<��
 �#oEJ���(J��^I8h �-�p;�3����)�BE"������0����\�	)~1
���)躭��g�W��c4�ѽ6�jɫ�[��Ֆ$������V̀�d�mP��%��Z�>���_�{���&팴D$������]46}����JR��p05�D�o���9t/VvxO�u�K_�d�4�ɏ����o�,Y %Zms�']��p�8a�Y�	�6U[���;�r�ʳ���J������?;�2�.DT�D��3�2�n�����4v*�i"�ˠ���Y#���"uLC�p����zz6�C�!Ka�C�C������E>#�]�
�{2�N|����&����g-�D֌N�oq�c�	
��['C$��M}O�`�-@I�������K#�.�>į'ǰU��pW �P��?_S��_7��g���Fx����iz����Ս[�Ö�2:�K�ϬWPc���	���CY�t8΋�[��̀�����;w�\���fX�#SIX���[8�@V- �N�%�\�3�R=��[�3R��v��h��iEg���
�N��޺_�ҳ��H%��xy����Z E=:�3�n��r�lq�
���OW;��S/�sO8��ލLʝ/� dpTNd}b=��^x!ϱ|�ڨY�f.�%t���*ib �:�����Ku����Ā�!�"��L���Y�ˆo�+n�����N����c�kª��z�u�"�\K虣G���0G�S���jz\�����8H�LT��Wx�K��i;�ϟ�?�qX(��آR@�� ��a� ��@S��i?��[���H���0h��d���tUV$���
���S�w?3�j6����A��`%�m��Z��o��ZW~��>ao�P�3V�j�l�2W����r�ǔL��u�_�^8Q��r>�Ts�bO�]�H�:\�/.o������7�/4�P�E�.v�"��Y�v2~(���Ȭ�p	W@�����_��=Q���d�^�
�޹�#F��,�M���b@]�,\�|z�A��!���e�)�1�+Uwi"�8��bܮz�3܍.�YyQhW��j��n��DbCܩ�w3-��(���S�C~
}"fcdO;����S�!5#*��",�L���7��J�w�����;i�@p��{Ο�/s���pe��o�9����wν��Xa�5F���f]Q~"t3G����^5Y"Kj�&��9��N��H<9#Y#��%i�)�xmۓU��gLz0��y�pųcRu#��	����O-s�G�m~Z`�h���� �Z��n�}�4B���ڧK�>F�7����$ƽ�VHg>�;k+B6qGxx~�z���q���ր��Gi�,-;:[W���m���K)0�����w�Ԗt^��K�Q%���f����q�N�	�T��Y-��@	*d�:�l�M�r�h��Y'Jܕ��S� ��։�K���yf����L�i.P�EP�/GӶ0^�^e7�M����$�����Au�TZ�`���r���	��
̶E3y`w��U��m:Kqb-��=̋��
yp>G��o�k	J^�?���S&��Mlh�$;�������2�� dL2��9��v>��.w�(���D-o��n4_`*�fwK�恗��Ɨ��#��r��8���gN����o(��Aw$ǥ�#���,��\l�y���Ղ�Na�,��>1�q8�Z!��ӽ��',��cY�Kw��VD �X ���3P�?>l����\FeE+߂���f9�����[X�>e���tN�V�6fk��o0�l{� �(�fM}}It�0���$n��L�&<���ZP!5���8��F455�m5��,T�хnZ\�u�WI ��j�ĝ/�,�i(��,�C�k��NB
o����'�����W�3��Cُ��-ـ|a�͘�uC|,�LV�e�c�21��U"L�����<����<����\8r|���LG��=�!8p��Ws+>̱�ĵ	L��`�WnJPa�b� ΢LK�j��aƱ���
��dA�a���B��:�5�;d��%�0�i�����:�F$8*�J��pC��od(�j��~���;��Hpi�pZ��V(	�ZO��E!b�cE��?�х�S�pP+<J+��d �i)�"t�D/���Y�x��x7[��6JQ�Fq�F̾dף`��(x{�/y`A�n���9��N�;���[��V\[Vj��p���)��w����wkO�Ewt��\n��ѯ9�\��{�}����"��
�Ԋ�R�B=�m��"�H�5,���ha�Ocb ԏZ�?��}f�Kzy��Kuo&�S*
U
o�Xl�e�u����#�ٹ�x��*��/QW_d��%�(t��/p�	���OL'�M�s���/��̛��"al�ZQ"�4!4(%�k�O�P8.#)��>��񉉊NX�{�60��C���;��f��_L�-�$:�<^�Ě�#.�iۄc� N: ڊ�����-���hU��@��><��n)ϕ�z��٭z����R�Y4Ձ�>B_�)Ӳ��J^w�݂3����<���>a�,O���Ў���ϳ}#�ȏtɷX�6�#F��&em�|���;�k���S��U%�g�h��po ��������3�.�u�=ܢ��\2Դ7ZMG	�<E)S�����/���*�>�������9L�����5e�(�eNXto�O5:���#_�fP����5<5�Dna�7�J��z���E��8�=f�{�k����k�@���ݵ-�e���- Wk/<���z��}�}�t�X��Ө�E�����V@�s���]*�jp����nt01I��V�&����D�5�`�R_D�2�����D��J'}n����hm�A�
�x{����ʙl�
ަI]g��d�8�vt2�JQag�2�R:�W��_�C�j���}h �t�Z*.9�^u���W�� �#n�Ce�CX.���s#c"w�Q��zY�N���WlC&���}X,���Z����M�
�{���\ǁC��5�p��X4{�G�M8��Þ��]GAH��JA+1_�fSј��F�xf�����q���eH��>pr��L�ьM��rt�n(D�CuRt}$���2�a�L���w��F���0�q�X.lkk3��ċ޵�V^M����<[���!��+�7�ʥ��Ph���2H�vu;*��ml�W�b�1�Ύò�;�;���A7ƅw�Z<�uN����KU*]pm������Ctk�ގ�!'�~��	VWú_���-�!&mD^�`j��<�m����f�خ�׀�o���w���\L�Oh�̺=@��;y�&{T|��N"�5�{�Ce��1��t����،��ra��FlrF��xbqb���ѱ�����z����. S�Wͻ};�A�{��i�c������3�[��e��h��-Щu�%���8v�w`�+�h!�=�;����c�������b�����8]��1�V�Xyv�h9v��m0�SlrtB�o��Y_>����/��R)��� �18���78�[UV�BT��.��0,��^�]���l��z��~i��t>�'RHs� ż?��	qy��6)+��G=�]��*m�ܿS�լÙ����/���+��_�������Vw�_ӱf���I�C�`¸�f6'5)�����OMI��p�`���`����+g�7�B��܌��w��Hq���6\hP�������;�YZ�E����X>���@~K6$����5����qI�,-�ۮ_�X�o�g:2�f�즘����=:t��HGuWw8�O�?E�/.Ԇ�Qae�J�C��'fmGa�e	�vv��QU����-��]	M	�׿ �O�xĠ 5A�̶�7О����Wy�$��&�h<�	�0(_y'������y̶E�5W�g�9����2�szf�nK�T��]\Gb>t�©%���N$Ȑ���+�l�rI�lB�̿��r��'*��D��̈�(�>�cQ���P�a2���Ez,Wo�M��c;�^̿<�'��w>��v��*$́�:3����G���Au��	�%�	���a)��?��A�-NX��X���'�Q�%#i'-�o<~Jb�-�y�\:�nmW��%ڻ��;l���@U���'@]U��_��@}����ǒ��F��6�c=䶓�G��Jc��t]���󠌉j4]mJ��l f����llR�?��f-���|��Pf1�s0��?�f���������)R���Օ=��"�q����,`D�vI#[��OdM�E�����I���Ft���P�]�5�6+p��h�&C�ׇ����Xtg|,]w��'��C��/j�{����D4f��z7v*���G�zJ	��7E�@A�;�Yz�4W��\5�W��%ٿ�-����ҭ�+뽃�@ֻ
���Xۖ&���J�_��-~�v\`�6O߃�;]�^�A	�G� �̔��~w/�e+�)��ǺI��?L��sM��گC��9TŐP�ثN�*�ET,o��^���A���X�Gg���9޾�8������EX���C��Pd|��E�q��`S|Tf���J���S��t� �q@mi�4�ABtx�/j�np���}���~jH�s�-�)�K6��K�Bu0��e��n�B�}i��P�ANn�C @�� w��V�bS{g�;=�?�V;�I��Q�KrG��Q$q�__�HlC��˱��^0���S���Omh|r��PӢ����>V9ujtY��f���"�����>��s{k�`Dr<��7�a*`K�|,00��b�̇�
"e]��/��p�;O�D�g������g��}lȠ���@ +Qx���k\xB�t�HË�T�$F�͎Iw>�s&n>�?�t�<���z�"q�OHB?1������J���M
���}9�]~U��M��ㆱ�,�H�S̾?|� D��zH���!?2݃��)fZ�&�-��s���A��x�g���C��̳��N4/�vJ�2�*i�t����F�[rm��A�\�~��6�6�P��Y�MC�b��eK��Ш/� /_�3��j�\zO.�GD���^Ήt�"ՔM��B\�\����>(�,���ߥ�Ѭ@�F����t�ּ
*S�xE)��Pq?� ��>�cmd��{q���D��x2vp��Y����j�/�^{���;@��[I�ɤ]�j¨�QKfcw�
��k%��>�T&������tgrb��!���[�4+�[��Gx���q�7vl������/L%m��$Y.$`�C�*&��V�`�2�e�߷o�nsm�Q���i�;E"�fS]�>�=�j3�J+���j�(&җ�X^-|��$��r5��ߩiJ��k��m���'+yЪ)�8w*��$������u�x�62�CN��{v��o��^�˜��?��e#�q�F������F�O'�TS�=9	���^�\�P�눯B��<[�1�L���B�o��홄:8��166>�_fP�E��P���!L�h�0�9�k~C�F�WUa�-�a�K|���L�yӰb+:E��mq	j�TK��M����v,����_���t��ͣ�Ry�`�wsu�����p�XMW��"'�1o�Bϓnݥ��Ft,͗-�ʬ��
*rx�'?r쯐�Đ��{S��7lu` t�+CHuA�D�E�M<�#s����8��<��QN�wRwV�����81ΒQkX'����f
�@xJP�r���ނK�T�^)בU3�����>��V>�^�,��R��s^;X�ܻ�am]��7pw���ۢ�SVr���L�����gbN�{�٫<�5��~��X��3)��
���>T��㊍�!p(���O|�\��1���?\�7����&���L8�o#���Ȗ��Ro$�����a���[�Mmwc�{�
ydP��q���+�4p-�	��^���o�־�Ϙf⟼D�I��B�H��F���<�,�=��4�Ba��Lmz�Ґ~�Qa��pOdp�}Bi��~��q���d��;���TF^��-,��*Y>��ު����2JT�x�)��=�T�����A #��)Khsypg�>n4.�c�J[qL�c7�9kue\�=,���8�0+�,t���Y���9�R-"N�mn���>�8�JY��])m���(s��f�;���oJ���*Eu�+��l���Е)�� �.����)!��T:.$L����y��Ej���?��+V�8)8��=?ANgq�|�0���U�i_i��~7��z}������ �;r\��%��}T ���&!����G���ɋWO��@W5G�r��I�wv�!��d|K�P�1�5ß��W��$]o
���oL�E���}#��S�p?2 ��V�
}"���v�0�K�u��v�h��U7��.���@�#���!��.�Z���/.�7JR�=H���$v{KʑA����Q� �*Ϥ�BU�����4KE�`r6��b����-����`�>W�%=��v����q�N^��1����/�_�M#K�vg�&��%���}�@��Ρ'��=�~��_�k=��r�Ƒ�ZBL�G�z��+�NR%���Ԗ��,O����i��/���ߖ�?���^Q��K��c���4�2���^��s�΄{J��)��_��k�pHqf"C�,.�}�(�ӂ|�f������*��L���V_s�PQdy�4	/�%?T�?���d�&�LB�V�{�Ut�����BVƦ�1ɪ��Fy��^�e���!j���?�+)����i�@��hh~IpU9�q&�I�or5Aqu�oR��M�]J?KCN��g�+0Ō�$Vz�
������U}k6h�i��5�\��	����Ħ���+�R�ޟ�᧏�6�ѭ�N�Ъ��w�ح��Ė�}(}3�m��N�:��_��m��:��H�{=ʗ�K�������a~?���x�WD���$ZH�_r3��h$S����G�Y�m�����r�yqv�:<'�_q����v��j�?g=��{$^�y)���ba�Z^"�~;�2b�=nTD�M�zl0[rv%|�W!R��p4�'�ǽI�0y�_�rj
�b_�[x�Oy�����`��%`t�R�㜭ATgw(���=Ƃv�ɔ��̹�c.�M�-�����8�����H4ڶ쁥l�]���	r˓��C�j[�%/P+O�����1K��|0����`c3�EL8riU�4+���+ŨG�q9��*�b�����/8�.�g���N�y	�8���m�b6�
.(� y^�h)VD�2�dMʎ �J<�uU\�`���X�s9�5Ϡ}/�j$��&>N�Mhl�oݣ5Y.!�1\���2�V�jvȹ�O��J������$�O ���W&XC�kC��l��#y	�E����k�?�F��U�����/��ZC�Fcグ�k$����Ӧ-C�S��#�M�?��4(r��5v�{�ʸ�RȰ�F�i~"�HA=��,�o�D:�W��*׽�Ʃ�e8�4�H��5!�Y����|(zõc�I,��r�iY�a�z��&��2�A���e ���&y�Α�	#������$A��WN��{�yȥ�u���h}ոb-'��~!ԥ@���.���T)i��O�P[^��݈�9�᠎�C*ᔩ�T�G-�j孈I�'�EG.�Ǣ��Ҩ?�|.�#~ݩ��5@�ʦF<�x�$����y������J�\(�� <M�u>Oe&�==�B��R���s%�`���J���	�Pٿ��o�Bn��G�^m�VI�Rc.�Q�!�؟rJ�e���L>h�G�jP�=Y"��m^B��X] I��f֚c��ER	�)��=���k��0�Uw�C�s�5��\Z�UO2����ڠ�*t�-�}Ĕ���$�|b�˝�6#����K��58���8a�8yfq*&�6�R��6���*�}���<xw���i���Q����P�O�Mi�P)\k�Ϥ�+��V�4�����u�Bb�l�tnAZc@0�֚t��{�5�,%o��F#P��eg�Xu�^Ub�����0��o{����5����w�g�0�ƕV�o��B�9��~G ]�����On���wmr˅��}lv���E���䫫�}���kSW�����WQ_��OA�Z,�OP�	4����c-[�	��:��&֊��8�.�T���)ȾV�ABH�|n��JaG�[��MR���6�P�^�trw���%�/h�ވL�I֡
i��0l`���u���
$�te1�ZL���ٶ����pB�%�6̴X�i��c����&B�TT��ebI!�|��Ms��O+�r�����.����������G�HE�Z�)�2�8��$���QNU��	�)>�H�I����~9a.���K�xԮ�ݧu�R_���ܿ/���^ĳo�8��Y�kU2{�&�a��R������3˭ޅ�J�x]�C�WtVEٔD�.ը=�TM�8ǈ٬2�x���j�� ���/鉴.�Dl�#m�ջa��8!@��D��?�l�,��h<6^6`�v��� �`e���´�96��y�.aŐNP��FAY�8*��"�]\���~c&]2bq&�x����a��V��e��0t��=Ԃm�e\�S�5yNӦAEA�y�vh�|��O����l�1!�e��,���h�OT�Y#��Oௌ������Ж:��`y��4s���f.�3>�Wov��a=��[Ơ+$I�)4��7��ڻL��;��7�6�5X��Wzw���s�KXid�F��m�Tͺ����D���y"

>&��
���#t�Fi>�@�<�E�\�0F�@Δ{�� ��x�N��e��������P0m~�nU@G�,Yj������c�t3�(Eb:��}4��M���+yUZ����nA����ı��9tA��H&��V���A,-`D��s�C���|�j�]v�)�*:YM���S�]eG?n0��&ҋWl�&��'��S�qૅ��ȭ�y!GN,Efe#���,���+gFk7"�{"��0]�i�e?�hh���Q��k���E��N���<��<����LC�L,y/���)i<�G�c틺{������^��ٽª���\m�w0��^#;�~���n����|�l!(u�|+�E����b+GbSU���xْ�-G�k��*�o��
(z<����P�����@���A2~r����ߊ�W1��\���������~ �4`/01����:����T�܄�@�)�K���B�J�Ձ��� ���$�苙j�3E^Z~�Mr�r�\���Kӆ���6�A:��x�t���IzN\�Yw\�>�g��ZG��@ҹr�!A��[�("������|G�2�xT�[����m,�q��#a��z�;�������B��)T~�U�L�l`�(��i�AHn"
,[!X+S��ddʗ_���E�H�a���Q2Ò��3c�� �D�g�J*^zY�Cqo�OfK�"�2��c�&�-��=d�Os�P1�����p��,t���4.e�-SL4�������x���m���>fOo�f'�l	��� J�x�X������X����j]w�V:�lnZB@W�� F1~G�g��n���E�o�����B�($fq���%;�tb�/�)�r��R�K$4�i�S�w�x��#)����X��z�,9���R��q���n�0d�oJ���jh���P�k�������j���4������';����:�X`��S
�M�N�tI�ą��ȸf<�_x�AًC`�-��$��r��ıL�K���ڃ?��*h�o�,p�#Y �t*�i����Dcc�&e�cп���O�p�%����R/�t����֖=�Jy�� �1�������f��	q��ͫ�7>	����HR��� ��m$s�eT��-��Q������
Φ@���{�5�p�ũ�F��4��Hz���"��`�g�s�5Ft*��7���~��OG�.����5�e��� ��-�9E}[�`ik��{�|'<!@��.��6ovLo�u�6:��d1��4f��r��$E^H%2&�|ҿVw�b� !d�tP'{�z@�4Q��咝�ݜ���%)����(�5+��~���X� �����XV|9�HP��
���Hޯ��x}���Ȫ��� *�cMcd,۶ߡ#
�M��<�5�M�3�0�m�}�yb�P�0B˘͏32[�֪&�3����ܱ8s�G� 8��~��-yc��y��nXi�y2�S���؅D�-&<��G{BQ�3�4�I�`��j�.w:�C ���H�1��G{6ħg����L�ʱr��kĬ��1���/�i �s��Г�B�����������У�ٍᘃ����-Lº�&�mqE��٠K^�!,B�5�a ~���-̛�n�a���U6�͚G^f���I��1��$���0y�0��	a�d�a�͎���>���hf��I� ��[Z��<TZ<<��P1�����GN��+!Ƅ�V�Љ�H�����=�1��m��s�QU��@u��mvH��#R�������r�[h!M>%m�����=���Vk%�>�������IJE����&CC�+BY�סW�����n����iA�+&�v�	�$N�Zª�d!꺥�ʘ��j�+K�'�x����Ei���J�63�Dk��T�����Ԩ����-�N׈eӝ�Zu�b��`������$X�9�wW�j9��o����A�<[b�ѕ�Y|\�q
�g�>�W����]ȥ��~���^�Ս�ő$2�]�ݧ��az͔Q\V���2N���Jy�ak{�W�F�����/Gsz�%�Mm�M��/U�nK����~P�l�r.�9?�ݧ�e�ǣ����
��bx밾65��p?�a���B�`^1R=���[�q<�i�k[^;�,ãG�e#��C�y8��շٕ��� �N>���l'k�D���AV@΅�w� ;���;Y���-c�A��F�Q����@w������c=��[I% "�A��y�܎�?�c�9:�N��y�|Q��	�['���n-���}yJ�9��ݤQr�I��G���#�#�`#�-�A-U��hi��%GU�~�1:ʠ�8 ��Id����O,��~˽�
	6�f�^�� ���gU4G�EI"��+KH�@mէ�b��p�m�C� ��Śt��I!����Y�Z�:Q�2����ح7���x���+�Qlt�� u�A��ͺ��@�8ʧfMz�R/1�7�DH�}7pwE]y ����J+��_a��3c�3�1v06�͗s�h��d<��f�60���?���,��th����Ƨ��?p�t����C�_�~Z�XX���`�I`x�u=6t�(+�����g�¨����]|�����ɖ#�/O��(�j���r!�����=��������j0g)�l��Mt�MH���z���ўE�@���C�e�1��Vi���ʸ�}�P�R}��KBz(�~æ��T1�,���,ucÏ0m�3PP�{����٢Ia������~��r��I��=0XP{��:��e�����6�B�}���IU���}6�砪V���#��8����χ\�*��ʃ�'lĕ�J��]��'��V���.��*��B4REs�/����SoW� �9���6���o� m��'��Ew��Gj���QI��]DJ��X��U�����PVQg(v��Yi%����	��Y͌F���Ȝ')u����bm��x+�=��o��J�N��>ad^���**X��/կƨ0rԔ�$y����1�		�yl5SP��G5���<V襖8ÿ�0jd��{�s�{�,M �nq���
}�9_�Uɼ8j���6 4�X{�4�p�?Xt��s�-�����BY% 4�6�beq-Hصw������I��g���w'����}���֏�`�z��'U�s��1�E��29>Z�Fc���S�z���G����+o3�򿃯
n��'[��-��M��^��ᩈU�����6��T�q?j���fD�(�彀��)T�wB���y&���_9���'DÐ��ku��֛�V����U6&jL�q� �yl�E#(�������<���;1�)quW�
,ȹ��]\Ó�����'?T���8EM�e��UmQv�h��ׂ������M����^�E[�bR	��x��۪;~�-�L�&�y���5���kaK����GQ���1�̕kW�X0N�`w�@Rۄ�(l��g]��$�h�2�nwc�d��?AGVY)���	�@Q���c���!}̴a]L斴�SL)7��bc;9���V,��r��� ]���+�=�	p0��g	�|�ξ�(j�{^���5,ƴ�!"�n4��J�F���ؖa�5(5�����F}�&�j>�7�}!y,4�̢ �͑�񤛗��t�f}�dF� A�{.�HO���vTO���:ub�1��tB��/9~����zbO����|��X�bؙ��7o�PBV�l�p�H�5k7��O���6T��y$���o�^��)y4�~�sO� �|�-����оbBu�f�bJ��c���vǅ7(���ӈYqK�aa�^<m{{t��?�L��%�d1�;C��C�y�{���v�?#��nl����p��~eT���S2Z�����
z"n�I��j9 �v����������]|�vɘ?Ê���rU�` u�0��z"�c����EG��s�R��ZB6��vd��[)Pnh�S���=�V�V2aU�J0s<1�4�gh������QA��l��6 n��
Q�f77T���n�x�>u��+\����+y�"^����bH�qRneZ�&R#��Fŧ�:T0���V��R��i�d�#�#w�c�)�%����=�Լ�,�m���T7�@_�^3���7��@�d��Ǆ+4���L��U<��xUU�9")�a�:�ی��kO��y"��H`�I%,�ӏu���9��s*<]�(�Y�IGu���z�Fmm�Ϩ~�~[�9= �e���xQyX$�E�7�\��ĊА��O���P��'�"�����^�Wwmb���F$%<�Ś��Y7%�)����E�k�{3����s��Z/��T:�����ĺ���Iu[YG#*���� u'����ؓg�"|e��=pF>OEu۹X{9�D"V�Q��5����Z/�`��ly!��EmP���o�Y#�(H��:I�.�k��TĬ���U~cC��={����;�(����Ί.��\�,��qg ����a¼���N�]�{F�<���a��a��6C�W,���HR���!���m�9��΅�D6�A�0C�K/��j�Wσ�dB2���s1]�8�N�	C�b���+�A�{���]�"����֎x袍�H�������P��T�r^!ք��2-5Z���Uj�LHO�#}�֌P�G�>&@5� ��-����<+�-#�@k�hH���_'�"��m�R��t�F����k��ԇm:C�r�;x�H`�1�y�}O��"MD���w�8Z�k��=,���%hv� ���6{nA��UVhd�bo�a7�܂���Q��'G3�י� N_O�aE)�+��ߘ�"���ZK�1CB�a�|7Ai�I�Z�~�-`�����!�E�RW����g����<a5ӳ7�������1��'m��^�v0�'��[�4@��������d<!#.cu*}��R�羠 �R{� ��%d��s옗 �L�zn"ꮔU�L�8����8O�Hںъ ��g�jӃ	�^��A$��U���>�c=x~9��P�Q�I/_�o� �����c���#Mɹ��G��e�)����%��J�Y�z�g���ci7�*Ϋ�1yB�%���q�T�!��-�/���a�Ī�n�D�wB�5 �J^,��.�~9��	� з����\0h�`]��[���רz��=���_���lyf+�)(^w��⾝���F+���"O+:���)� �cR"3!9���X��n@�<������G�}+�9}�����쀧^�D�y�x�z��E�.gsC<׋��.O�	�}k�Ԩd�$��>��em�JqF�6?�
h�G.�����ZG�s;���A4�w>��c̆�mf�����C�F �1g��l�S����đ����z�m�L�4�M���U��:��1	j^ �-�m<���Y8�Zm�م��I-_�?�=ϝL0�c�����JE
�����%f���#��0a3`����O���rM��O�Oh��h&�qS��N�����E����%�ǂ��~��B�pL1�oP�Q*H�8h��2�[|�r�Fy��Սi Y;()�E�r�H!&!��f0C��_��I\.����	�c��:�V`�4�7�;�HS�#97�z�I7��ϖ͈V/��]m@��
;��s���;D�!v�������/�����goH��4���
��[j�G��scB�DS��UI"A�?Gy�Q�I���+fLJ��LAxu`\C���x6�#T�����s��_l�l8�Om������I_a��Q��������N^r��D�7�}0�.s�^nT���l�Ԯ�yڙ��������J7Pr��l�^�S��D����?�H��y��Ef�K0 �NBU�Y��~7l���0�A�$��W*�r��r��D���OĿ��"���KYK�W!�h��r��$X�'.D>�l=K�1MTf��� ��{�<-��["�!��e���!أ��
��I,;3�q7���VG�1�������mH�c�=���N,��9l#�� u�o���4�ZW�3AE��Ӹ_�?���M��c�42q�df���F7� �'�#,mqxN�tifL.�����.�o���8����o���Iu���y8�O5����;L�	�cS�0egs�q�F`�1��%L�)x��;�5��#��'q�Q�U)���;L�8x-�:��3<�2��W�s�񭼐���^n���9�113���[E�3B��6ΞA��;(����h$�L�jg`�0$��8�תo�$tV��g��Rq��-�{������6�����N�c?aN��F�<���-���HU�W��|�W�E�,��o�60#��v¹��]mٝH�Ժ�wa�����P�s	�@2�T��"���ƙ�@���Q��\a9�
lY�f����v)��]Ec�}��K�!^[3fiw�I|s��&�3��*~ްj����a+�a�Z�/.�7�s�d7ʾ�s��^�G�*���H �����d/��r��Oe*y���\M�����}����.aV�C��&dp�b%���G��x��r���(�}E�wN@R��z��Ģڵ��7�t����}�0tO"��}�G�FG������\$���t��w��bg�
u#�����d����x���?�.ߴC�J~I��f���y��:�,�A�r��]\��r3�h��C���B.��	j�8� �O���'P�Z��Ҏ�'B����͈XA!��@ۇ�e38$�ē�E#e������K\�(�|F�k��qR�.$�H�Q�JxPjr;L#6�?[����5A0���c��P�cN�ƛ%�g���*��X����r��g5����������0+gy��WVL�듳�A��;o�r�%��_�^q�~x��)Y�$@���(�f���V��a|A���w껠��/dfm�d�R�]ހC��R]��5h
��IkU�S�I�'΀�#�
C�� 1����	K��N��(��Gr:q�/�sԙ���՜��Q�Z,�y�-�����@�uP+�Ts�B+�7����H^����v��OW~ϻ��;$�;��$@��u�
�l��g�?kGj�B�Ѱ�j�2�q���D�=ö���������x�]A�^��=�-���[T������a,���e�2Y��_�zaQ8�D+KX6��>����f7�q�)zA㾪7�6��z]�~4�����]MN7�h�M���M�O�xo1��Q���H]��q��P��ϧ��l�kn{�Ɓ�!�I���1&!3*�r���f%��-eO5���<�M{oo��ǰ�Wئ��:>�0I���F��0�x�xn�(ǎ��Rc�#��w0yh�)SI�k��:1���Q~�hJ"�WPǕQ��HR=�Kvc�v�9l���0���Ѣ2��-�;�"[�Y��I����%e��x�:\N�f�F+���&{a�Ԣ���Y=�r���P�8l��xhs��ΈL�/����ϲ��=�)��*'½�9|+f�%G&B�(�w@TP1��MM\���#�qg����l-0y��4$�.P�EwW��S���c�B���&>̊��޺�x���|=F9'R�6�b��3C�=:�>�F�;��tGa}KmYF��T��I}�O5�����B�F��_<��,�Q��IZb���������AX1f�dY@��JO7�U|W�����VCC���W���Г�fK�A4/�r+eש�نc���P�'$n��y��`Hx���_R�=��5�롭 ��Rk�+�Zh�@�_�z�MJ4�<}o��T�Xq�f��AA92��(-a��6f-c���,�zLH��d���G�N٨��j._�=k�#�j�W/��0��o�k�U�N��g+�m��;P��a������N�k��a���U��Q� 9�f���M��]5>�ݣ]W��=O��;:T�+1QO2u�&��<E	d�ȌpiY��� �bc[U�kO����]��I�!P߬M�+-SW�$���O2�a�z%:��Z�zסd�"��s�; �!@%�RT���⑿�Zq"`wf�x��3�iܫ�ܟ݊CZ�Q|A���*D�2��v�m��'��Iԝ��=́�*�qt<�<:x_$�%Jlr�(nj0�L�K^i6)�u^EK�q�A�󳭫ZIdg0k�|f~�� �#�u�Vl�����O���U��r�aA�!���X+�l
=R�i�*�]��>M%��C.�a�J�T�J��ڷ hp��`�<�;Q�B�暢����Z}�6n������)�JE�1	����*ж<�n~�ʬu�$���u�0�RXa'>6\^h����J�*G�PA���8�M�:ۈ�^�Kam� vz_��`gݮ����p�/��H��G'Z�i�4�����^Z�Ϧ��?k9쩮�!'�C��
H �eZHkK��!�>���@�8�>l����FN'��� ���s��p�^�.	��� �m6�P=�%�L'��$���w��E
��m�4&�����1��9�#��_������T��%p�A�MƮGb��E� �q�u޸~�����7�u�㯱X�H3��!����\|T�m��Q:L䯬�.QLBO��?f2�<tW�g;�$�IV�2\<���Y�M X��g({�Q��*$y�U4��/��_��<��hB�׭ܵ��"�%g�<f���s���Џ���G�*s�{�P��@S�H�r_�	{��&k��e�=T���شi�4��5���VHD�WQ�#�YG��<�;�e�e0�q��Cm�E������S����'ɉX٨|ߦ6�_5.YG�<s�3[��^�~l�b.��Cv+��1���V[�
n���{B�x�#�o�?�-Ih"�ڨ(�ƨ�6v��c����j�}Ǥ`�|,
@�=O�t,*aC�w9�����[��}�s���<3o_�o��H�X��l��B�'��?��ɯ������Rx>��bU�{�%�Q���|ňp�&�~��jև�c�Ӽ>�ųS��XR��8�i77���"���]��<4�6]����=��s�;��&Q��L��F�T��H�()q��0A(@[�oߛ��տh��ѧ��;�nR,�`7���i�2?�te�> ���5��9d��c͡hv��%}���i��-I�tV-a �F��%R5�<;KUy6H⾗���v)EN��5�QZ��AK�W�9��T�iV��������#�7k�_U���$f�l��(Ot�U}���T�'�rx����t�"P��'���<ک�C�5�2�T��+KM�R��-��
&	��8�V8V(���'�`��iqu�wn5nT��NF�g����*7�V��f���N���z�6c$\�������\e��"�A�B���}h����f�HO�������\UB���&˚*�Ĉ0A�q��q�*P�X* �
�扖w�p�p�R�"_�f��J[V�䜝�<�RρY%B�k'Y'TL�33�jbe)��!��+=������I!�k��K�����^m�½�rZ����G�*vCf�'��n��H&��G	_�
ߓr÷�c�)/4'�&��!��� ����O�!И�q��g��S�:�2���!����#��&�Ԁ�׾��y��vgr�t%�i�*��������?����G� _�������ci�ɼt3mٝs�2w{m����0��^�W$�nn{�X協���4	�ě�T\z�>~g)��m{��Kb@�݀7�!�_#b����K�S#%����	�F^@L��%��ljѐ�:ܐ}(��F ~�)��?u�N�-{Ŏ�?u�G��k��k���#1�D����rU�t�}pxx�:���'_z~()�}gO���nQ�0�9Ϧ73\F�6S��M&���x��!`;��Ώ�P�c��*�d�PKa�b-��0�&�Ėpe9Ftw�n�����p�@Ra��K��b�jhA���'@�]*��47B#Ѡu?�7��ڥoaPG���+�B��DUFl��̎rm����Nc���o�������Dh`�Tb����v�8'���s�N�{Y��B��.3��F�i�?D+!�/kA��c^I�`���pK��yDp��O�n��o�T{����Q���>qs�*0���_]ʣ��^K�����0ɮ+� &oz��;��F`(�j��|ҿ�dKi(x}zu�dr��)�_���(W���^��aK�����P�z��.Ch�I8u�P�G�7X��¡YL��o�/�^Kk� <W�=�A\Y�����Zҭ3E�J@�-i��3i�d!4n�1W��7mDN���-�
��/���5,H�O��,Y����N���P��d�.i�V�y���+�1�*^;�<!EV�)��X�d�&67q	#7�l��9���0^�����w��<J���g��o�,�)wm���.�@z���.S���`�RG�4�m�֏l�����ն�/hx��� 	��l���-�X��e�K�L�B��d����X�NJ��)�aɮ�i�v&���̺��vx����n;�&�����ԅ?(�q���>ѱ�/zT�C�H�]��`[�#sm-,�ʷs�
���k0���/~�el��_Q������U���l�j��5	�-7����_�㑶V#2���ep{?��#�M�G�Y�{8mu��U�5�b��9��~SY!L%�̖��:�S��K�zқ��o��nԅS]�;���E�8���8�!:k��|d\����������:7tB��d�b��<�;f`Pa�3�2'��Zavh0�>�X������T�3P4t(�w�E��An��+��:^P��E,�4�k�*K�
����u��6i���)��5��v�%�1M�o��Hش��zl�?��T��_$F=�Ւt�2��1>�w;��F&,�¾�ވ�q��1C�bcp��͍L@|��>�S�H,����A]���ڝ@�D�N�j��65x6�0S�m&ݡ�J8b��Vޙ��$]Ac��T³����!a �w ;�8���m��vVIs0G��8>&�&E��_�kQ�r��<�g9n4����ԫ<������- devn�&87˾i6	�M
�=�q�J�l��on-�񎌝$�(q�Z�*��(��Uy����[\�tl�1\fC>�o��Ǆ9J�E/��z!6(�a���\M'�"f�B l8�T�BIS����9����^�}]q�����")� i�vZ���RT�[��1���7�D =�e���ڔ!R�vyw���d`�Q�jG�"`)G�0���qipn�ZpbOE�'��I�x��mE�˱�1�HjK�4z�欵SZ�?���V��t�
��Е�Ŷ,��pQaJ����P1b��3bT�D)��6�d�	��v��q�S�眹m}���0��1γ9���w����`�@�ȚM��}�{Rv�R><��1����wE ��'W5��R��b�8(J:k�U<�`�B�ī��[�l�~�b 8 �oΓ��ٰP�B�#�J�X%�e/�&�P��9Y)�� \�B�>i���L)��H�-q�=�ފ��vA��p����zz���(Ie�B����!MY���m�:g[��T�sRD��p%��Ђ@���4���
���Cka؇�7Y��.�1C��2��ܭ����ӵ�.�O{�@�1l\簎N�^ȴ��*%r�U��81�QF���9��=��7��{O��%^��N���Qt6��"���8=���$*4GK��T}���.&��kZh�� �h�oL�����;�A��CuϹ2wV� ?q.������}k2*���p-n6�	���3X�=XLO��w��3̤?j5ɶ�!�c��Ji��~��~�ŕ�ޚ{m�_�G��/}����.���"O�H�lo�����X~_�j։�*~}r�n�����+���gk6�;@�=�^3�,�ls�?�n��/�D�e������1�آ��Z{�0�aX���"Rs"�>�ʪ$6��0�2kr�--��S,�����_��I�+`�E��^q;�?�VO�TUދ�fjgW�~
!v���䁯$��+k�w ��&�N��zX��b��x���޺b��e��B��C_��#㚸`O�W��-�:�>f����5Þf�;;�¾NM��n�?����c�'��d��::/uj�D���ɕ݇��w w���gC�T�6�us�9T%���a��[�5Ӗ�0���$����(�N��F8���_ˋ�I��?�bHZ�.ӏu+��Ka�Y�y���9G���d=V����ȮL���h�8K���^��X��ێ)�!���� �I�ƹz;���h�57;�W�z��_`��t�=��{���b,:�HOQl����`��*y��,�ﻨ9`w�sa*��sF4'���b��W��#����a�@W�e�5�@Er��o�,��ܞβ������q.J��%�
���F�����ט�!ԕ!�ש�\�$�o����R���<��N�W�Rzk�ތ�.�7f�J��Ch����G,��qf�=P�b��Y�EJ��S��:���t�2�)�F�'
t�;���^RnVP�*$�Tn�x�y�pU���¡���/��p#(��P�_�Ś ���SʗXS����Q�����63˧V��~T�{2�H�o;�ǘ���1��E�����"W���:�aR�\ͤ���`�����_�j�9f�[�E���K�"��?��M��U���@RDK��ѵJ=��[N���w9\] B��LҾI�ݓCJ�#��+ɢ!�x�8&���*We��=�:Z'6p�L�C�e�Ip��"�ˢ�+���>�	�b��N, X�9��tV�o�j��/�)�fR��} ��ʸ����zV%*i��K���C����t��bi��\�W�-�Jӷ{���.���Hpp��1K�=��h&>�d��f����]��2ʾ����f+Ѡ�y�ҊU�wt�i9��Ld2�R����h��,'�)(,Y�����wT��<Ij�XO���s��-�#���m�Y�����R3���Ff�p #���p�Z� %�lb0���������=u,�p���r��hAc� �ܖ,����������Kc�_��}��{f�ҫ������ds)k����X�D7=�5�/�k�C�&������~��lJDh��E.�^��<i�Mg��V�W Z�r�:�������>(0�h�K���C�E~W��h<O��kL�fs1���l�I������*����a���N���J���V�|`r%�sZ����~ŧ�v.����jE ՙN�ۆMM�mֽ6��-�#pFʝ�a_+n���?՗k�u�<�ayz��1ޒ8Ka�ֱǥUv&)�B�5�_ޑ=9i~"g]�R� {�>S�2����\��a�ĥ�J��]��n������e�~,'�_����[z��E�G|��w��ҳ�X����}��}�؁���Ik��)�����!���)��+#tz6�R����u�X7q�L��si�]� 7L(����B!�~�J�&` y��b�RKWG&�NXiDqA�=k���p�@;b�dң����Wk��ݬoa�M5�O��*�>�yx����A۸����Q��[���H	��(�y�F�h4Ө����8��.CQ;���Y]+,gF/2��*Ȱ����_{BjQ(4sWJt-u�ѹqU��\pv�������Õ[/�k^��(TT�D��+��͞�b��5��$s���:~X�}g����L=�8��k�F�����]�h�&�|=�=*��F��Po��nU���^����Wf��N����]�^N	d������̦5j�bM$S*ó��U�J/6Ec\?��Ld<�
d=o��fr��E7�a��I�9�"b}�l��.�`3�ì�7���Ʊ���[�^��pF����7s=yך�iB��/�}5�ȭ�8�K�0<�I�륍��n�-֦X��GR�~٢�K���Xh���'?�����;��O?���|�Q��6�4��ῠ��� }MR��&#i���c}ΥRs��n�g��2�x����Μ�ީ ��ԕ=�vGC�C�m�4�D�+�~ڱ6�p�\I+�5������VDUO�x�~����(�'����@"�&��9�C'Lƥ�mS#����FPr=�s�$����Z7��>�������Ѵ�[Y �bd��fVwY���R͜"�����4��$���Y$7!�f�r7�ke7ZN�2���O�$r#5�f�� ��h9�����Z2E���e�:I���vޡ�A�ސ7G��|�^���+t(��1Q���4pI����#�7�ŝ����8Y��c����e����J'�Zh��L��t��+�3�U�
��]%�j��ˣ� ����[_�A?F�ˮI:�yC�0?�8��yt��	#���1�F@��߾��xʾ��R/�̜ej6�	�5����I�w$��$I�17%�%��]+��
�xn&��ޙ���/yrh1���3v}�jN�T�E��0�@�����YF�[E�?��] �y�b���*{�b뉀D�"��Hm�usx�f���2T'�S?9��y~9ꅜFp�*dB�-�g��е#D_?���or���јG���LN��E�!Us���8F��m���v �	���FZ��C��w���e��� �ziUS}Q̧x�)�)�-ڇK�p	���E�����B *�m��]��Օ,)�C�/N�b��p���,�8�ED�z����=֥�?���$)]������|����;?���5x��E<�a>W:�Ԭ)-�[�Z��~�^xݹ�uN��-W(��T��aɬܱ�8��uQT��Qv��;Nk$����8T�9��Lo�Z����LU�U�ƣ\bSк������r�+ I��T搑���m�n�z�ه��%gmz@�QkS�)��-�$<=�����~�b$֭��2�a�y�H"���6
�u��@4��Vdk�ѵ)Й}��U@���Yv�Wd�O��G����]��2�n�XY�w��~p�0�����t����j�o%5N1��j*%�	��Zx����@邍��ׁ�Zdk�����yu�1�I�a��-��x�)A:��GpU�53�1��]	%<2`�S��4/�435���Z�3�+��hgm�����ш�(�l�
��i�>���[��:�a���H���`f,DЏ�T�/c�]zH����w��c`pW��Cs@�9Yp�[
�6|ui,^���j;/�|��BDX��>z�V�e�/Μ��F�����H�]S���o��0�T�~�Ϩ�xB�~�6���f��� Ȕ�P��6�Y��)IM�G-ęU���A�Q�-��H"N�I���t�y=-Xߞ���� ��)7� ��o�-��xd7�d^n�srZT��+�{���;]������{�;�r���:�����ͧ,sG��K�������pi��ڎ����e�m���������/�Iaa�9��Ģwr��^va3�d��w�:��>9��`�e �ε�Z�A�vkɓ�C݇��X1j?�2�#/����������P��N�p�<�j9Ė{�����{��!�g��եf���UX���'�6h3����p �&�k����^S :�=�e� .hj������� �*?	�@��;8��h�]}l�^���fI�=j�sM��+�"�a�4]nP<��o=h@�L����U�äG�FR����es�6obm���W�'Z���Z_+�"� ך�׎� aa%`�@��Y���2Z*��(ҭ�������"y���dd����x�P@(<�sء��ӄK�B�=�����uĶ3*|���܆E��迆[�<�Iچ �J�����{�|*�<f�\���)�+|uP�wJ�Yv��n�d��t��}q���B/e>��T#d��3X��}���r��k6���c�󾣒z����ŷ�}μ:��3�P�nd�pr�h�${q�Պ�<0)� ȌNE�5X�BL<%�x���c|>
4q-xe�%UIU�~wEH�$� �ސ:X�0Y�|�oX}N,��h�x��d�IR���*,Z���Y>���m�g�%A�"mɴ�[O�2���t�R���s��ͪQ���a��RV�0U}��R�#���~��[0�W�q�t���(�J�Ż�x�e��OL�`��[۽�T���wbK�ᑨ(,�E��
I��d^:����	�B�'�&yV�]1���iҵ��,�0U�v�� ����ӷ�}��Ը9,؊2��4�h%�&�BA�������	�\�Y遺�;C�����]1�H^޴x���V/��=��&ŀ��𩱷�}�C�5��V�9@:�Ps�R�56K��fiL��ektuK��  >[���U�:~GX�'�OYE�~tG�ys��R�}Gk�^�فt�, P ��:
�����m���M.:0�un�Y�5����[4F?�s����s�s���	]4�	��r�P
~ں2U5�� ��I3q��x3�g�n@���p�k�ո8A*N���_߼h�X���H���O����j8b�l�^1�2w_��"����`̝��,?��i�����w��<,�VJ�[�+�I�{R}��pM�j����c�tQX6��Kyi�<�\�jn�sT)ԅ�K,t�,!+ݑK�5�~���$��L���x���{�#�[�WM�Sr���?S�L�*S�1E�b/��j�E;��g�������/�Kv)�s.E4�.y�yE�,���� BZt9$�"E>sh�r�0������iȋ]ځ.�2�?�+�n�?C��|��&i�
	�,d�ι�sǿ�O�YВb&���y�����꩛6�5'Ў���Jw�o�^�.ٓ!1��:�W6�Ε��U1;&���8H����B�g�&��ܑR��AQF}�X\ɣ�G"���߷㹶�R||���Q�K!�k��ۍ�;��Rϩ;��]�zZJ�]�X	)ձg8��|^�~�qUӗ�(�HV����C�|F��_�P�P�t����7=�ö<a�����:�g��VCsC^�ȧ���V�t�H�_�_ך�yT]�p�]m��nDgi	�͎��=�Q��]y-/2��h����w���D��~! �쇔sj��\d [����b$���FM;"���Q��i�<f�\� B����Gu����6� �Pt����s��K�ʭ
z���i��&D.����MD����V������8���օz�\;�þ(�m�v_Q��o;_!L����F����7\x�.˼�C$"�[��V2�����L"��^�ܯ�/e�m��Z������gm�m��K���c��_Z�DI��h�*#�hx�Y.@�d���mq]%ʾ�.�LL�&��c�xd�Z��&�K��w�Y\�}a~�g��ıafL�H�s�T���s߹�.�ᑩ����{�Z�[��V�yVO��4���Z8��m��ح?���k
&J��>�:0����@��E��?��tM[%�oKI��3c=��B;ɏ�d4i�t߅�\��P$*�S	�vzNM���ֽ�iyħ=5��þ�L����፼��Ml0vJV���a��yPqE��QPz�!&s�E���X�¼��F���Ή���Т`I_L�6�(ε�^J�ۚi/�'7C	�o�><L�"��'���6EG��l���E�Ż����g͒h����ǁK���3R����)B@2���G�Ë{˽�kΗ�����]D�/��Wf�KU)J@�A�n�����xݑ!yMa��(KSL̼�k�%
�lR�Dk��Σj79�)��v�of��Z����G��dD��Ё���ʌ��~_�ȟQs?Z �����ҭ@�U�Ec����P) o��U�`Si���n��V�_���N�k����� �w��j�m��ޕ-,�&�<�� 0)h��gu]�5
���]�+�!�d��MX�;�ކ�h��U5u���^P�1',k��}}+�Q�4��C�Z<�����V(�(��h2�<ě*d���L���9b��n�R��Я�<5�-�8�P�#J-�>K�@p/�%Ib� ����7 Pe��c�R�:p�1�*e[�u�œ�Q0�2:o\��P������=�2��U��'�T�҂0(���29P���v�q�%��i�lim�Kg�Y���Xg@���ص&-��N� �S�k��@¬���-.�)�t�a�WP<����2�ꂜ#!�	-�O|��RAA>e�[�x������ɳ�ޝ�Q��g����r�d%��h-*�/܁��-XK�Dr�+��!Rd�$Ja�[��z�h_r%����%����e�-g�:F�ܰ��/ؘ���2b��a�q�FPIUŪ��q�*�Ꙛ/yP�Q�Q��)a���F�O,���Z��H�+3�'�#�c��y%�a�Ծ�kK*IP�5����������:_�l�<Ji@�dc�4�!Wl\� ��/�&����
@�e�ԢQ����u��Y��ь9!�*F��²~��A���"���.�\E<��;�ʇ�����JFB �qu�#��p�NJ����f�MN������=[ ��ڧ+�L��?g��C����۰���ib5_�p&p��e&���6��qʜ��@�w�>�&n��dPF@2���D)�oeo��Y�j4��y��⣑bQ����B�/�񳲸\K2��°f���N����A�"B��.�M!�����r�D��ܟ��j��/�!f��mܛM�I"d��Y�ٯNL��<b��^��W�g.�DQ���U:�m.$�7����:UYi6 �aE�kk��I�o�k4�G�p���t������=�H��%*pj̜rpn��HD��-����ˀH�C�z�y�	�Rw}��t�1��޳�Џ�-���Y#*2��g��RX�׾B��"S�(���C�v�R@\��Z��C_���Q�������Όǈb�%����37b<��6�رugS@�B�����9*����0�*X3�̮[�I��mXia�=~���;�|��ߢ���a��i���Q�d�gU�R�A9���������w������L���ǖT����ʠ�@�If�ط�*��oP����nX��>�I���!�9oŲ�RC��;6�{ℤij�P��m]T �(N6�<�9�Q]���R�[�c�e\L{DsPy�ĈN����nE*��1R]$�bM|�Σ��vF$����s����]"���[�|�a�j&<�
U�XG{g����W���{��rMn��\�0���K�]-�-T�v�D�/qK-i�2�IN�z`<����jKJx�ȓD���ch6>7�A��U#k��I��!h6�~���׬���$�J�U�|d��p��z�tY)6����9#�(�_)�:Ջ��>����E�Ϲ>N�x �EWZP��&U�� �;���f�}1�:M�.O��&��ȧ��=$6����M����I�6��uP�@�/�4>v�9���8��r����n��p���H�j@]�g=�3Zt������9�D��;��� ��U�麄��}n?Γ'�,̃c���
�M��1���	�z����*|��`�2���q5��?K�[҅�G8аǝ�O������b����hf�/A��bF@40��G剁��:�m���W�i�<H�2u�e�O�|<vY:�D�f<��p�Uz��ӋptgͲ�6u�������p����߸_[��3X?�u��᥮�71F'��'���!ղ�z������֯%���7��:��u�ۢrwK9�E������"w����G���A�И�M�Ei�m2��w!oOٟ �`j������ޘ~�T]�FZ�{W9	�Z�[UP�G'c��6t�y��~�*,�%t��4x9��f��G+�sx��r�˝{o9�)����Z&���^B0V8�$ �P5��c��p�|���:�h"�f�􁊳Jzp	̇'�1�׀nX�+]hv�Ф�K9[�)���)�_j Oy:��%���̯�eo-�8��{N�����*�%��j^R9�%  !�ۭ#5�:�k�z-zQ�4[�.����a7d��,��?� H�y��� �k�s	�Kw���a7�pw����.~z?���ٛA�ۃ4ͮ�D�!��X�+���5@ÛB�B�L��)���	pٯ��J9��m���I�r7�mX�!�x�B ���+�@�����/{�:�g��<�T����/���IK(v1	{~�V6��@p��@�j<f������=Z�2��z��\˚����En��j~X�j��L�oJ�WR3�nｙ�fuk�1z�P�'����@b�ơ��C���G�ҏ����Y�Ɲ>��|��Nl �k���w�{
�.�!�CvX�����'��]���ߠ?{���K���vQ�����(p6����1����{�?m��ts��Ύ��E������)�jn�� ��ò��'4�mE�.&��s��J ,xIw�o:fxƨ�YCv�������Y;}lw}4N��
S����W�K|�0�hD=k<ɔd-:�"���X�(���d��J�e/9�gѹ�H �����ӧ�V!���9�ڥ/˩����\��7��)b���Aܦ]ݏ����Y83(t�j���΂
�4&&q,|��,D���춒##��.~+�.W=�S�3�P�G���|�nB�:��5")!��[�t�'^����.*k��A���F�#ĝ ������p���0̐I��ϙ��S��X�k��"2��Yʳ����� آ�V��Ow�3U9p��?�(6wy
�v^b��^��t��o���o�`BRYG���I��_b+�<JM# ���'ɪ�.N2�ƺ��O���g�cq��j����R�W,_������	K�e:�+������?�d���n3p��u��X�~Nmz�	����G���ZT�裌$�m߰kE�� d�))�_��'�_J�jݝ�W��.���H�_@�m��eF0=W[K�~|]H���.G<��N?�"0���~6���4��!�w�M��+Z�i+ka�{4��\G�)��4x��!\¯�=�~񋥰.�]
�[W�Y56���'x�o�t���QaqN^>����[�GZ�?sE����A���'U:���_i����r�Ʃ�,�.
�
�5�����>�#f�E�ŋ�"���i�^������{���*��NeX���%��%A�n�
|%r=��6�
�(ii�F��s�r��[��WwF�X^)G�-��媰��c�(|F��~$T���i�g�S^ty��N%bt2��=
 �������
.)�|�wK`�v¯my���
���"��93H�ǩ���Ӗ�Omȡ0�*s�KSm����G3`��j
m*���nS�˰Z��L��!��MNM�%=ى~c֡}&|�Lo�\�[��*^���G�5�ɴ�p��U1��0ٴ5��F%qwf*��e�<��PA
�N�f��\�V�R��>�=���d��U�Λ`Q��L'�u�f��a�$L�,�teh�|���k�80�ҐR�94=���U�1�.�������_��Ŗ&�ŋ*Y����;�7�y_���m��`�1����9ރo	�d�^���@f]W�R:_%�I�)�W�C����Ƚ!U���2�u�^��Yf��"IVz��9�5�X�i Yq��r8��}t� 0.��9�����	,˪��
ݧ�!^79BU��
���� �a�Ơ�U�M�i3x�t2�?ó����ϵ�G�W/;�'S���2����s{?�|*�w;��J�
~���Q},�p���>�oQ�V�`���6*����5�D�x��ŭ_<��̢�b"�Ko�#k��N���*?7G��n��O���,B���R[�Y=��M�|�Β�[�ޯ�s�� �~r14,g��0���x���[��	yjW�,+��#֭P3�Z \��[�{����o*!έv��A�\>{��((���8|]�������h�Q��
�86gOZVze$WB"%Ѣ��ZO�����&�6̓1$P�,Yf!��՚8���"�� ��)
wV��E�	���2tk_@���5���u} �&��iTT��f9`$�2:bH�v�݄��V�nHC�x�P�*�5�>PX��
�Z���04t ��AR6�s��U�L�"��o�5U*�{�Ph������I�&k��{W.b�WLaw����ݦ�-�P��|�[��z���J��*�[F�<�M���GہS��t����N��.Rx�C���c�ecB�h�ڼ�G! C�l+�}e��ꨄTgW���g��V$\P�5�yɪ�|!��)��t	:��*�loٜ�4g�;���o�Kr�ˏ���FU[f��#"�D[��j�}�ߗ�,L�{�	_�;.rSV��O�'��Йw&�kGu��1��\�[��4W&�$:d,���(�:�^3N_����,�5M��VT��l'W���/���Ơ�uV 3�f�<4���y����"��7d:6������ٯ������(تS�!F�h,~� �\)6C۶	��7�>l���ҟ�(�p����Q{//�c��Q�!vC��0���\�(�G�v��ca1����L?1{��s�Ui��._ �o8K�$�'��P���[�E^`g�ĩ�z�'|A�Q h���H���W��I�d!���=����y�_�z�b�Կpp[p�Σ��CTJ#�}�,6�؅/H�����!h9��$�]�G��x�r<�p���K�qd6�g�ɩ�]���Ϻ-�}���Fy�\�����D�>o�C�/��";�#�2���3�:�:!wK��^��ӿ�R�"��
L?s�� Pв�����S�n:k���*1�uI�㭦��Q���8)%�� �L��i�K��e�>z)����H��A�>RZe�.���&�0f]��>��*Y7u�-H̏h���!�X�؅-�!d�??���=�I$iG�L^�M�~�~!@"��k�/ ��@��CX�Y�� |
o��6�;�Y�v�$om��V�q��I>R.j�Z�*M�_�Ac���fg��$«"�ˉp���Õ�z�_�X�UO&�q��A��N��Hf�gv�HP�kz�X����mbZٓ0Xf�����+[�����:��?�@w��T@�DU(���_֋�3�k8�j��'G���U�BQ9'�M%��W)��腂)��]7�z��r�I�m��03j��	�\c�u�&nd��8��S���w�S�&[��~�����&3hm!�o�ux�)��4��).�gH$�?�PW��M��k�9�nt��P�ͪD� zF6
-_��_��e:�Z6L6xݺ�.DL�_����'s���}x�+uJ`G��+=��������OR�9�ٍ�j2�ϱ�@���'b�J��YC���1�_DlgIʒ㑘 �R�w��N��Z���}[�2�)Z���E4�Mv��$n��o�h�p{��W-��4� i7Ç_�\ke�������h��uQʇ���K�v-Z��ƞ�4_JVLM�� ��Dc�@�bK)p���s���+�Q,�\�MaFa��m�� ��4�Ɛ�'��iP��C�B��M[�>wCp�)��#��!��xJȹo��V�}�e?�6�r�~�'ጺ����2�'�t��.�)QO���~kU�Hvr��Nҵ&���J������O𲚪e��	���?:��d-��Ն�~��[��K�3+��\�8C��D0x0�����e��d�U����=Ȋ�{�����`�<�ӑ�� �.�i��7>f��"B^zQ�F���r�([�L��Z37Dو&5�{]3�[5M�=l�VT��~A���:0���x����A�:F�2>�i����3Β�X��5�*��k&	�H�e?P���O_��T�ʺ���[�M�iX���"�e�5�yZ)�<�@�![�'p�����%tgLm��'��?����ʘC�gdey�U��q!=�I��脡?��*�f�����,&�^��Zպ���8d_QեN ꂦ����Α�zUp���CƑ�d��UGםU͡~��z20\�
D'&yԗ��
~d�i�vK�a��df�Cڐ�z��F�kK(���{����\������:�. $�n�W�	��D�]<��fT�������f�X�A�Z�ic�:�U�j��r�CH�>�@G���/��N\�f�D{сn��%I7�m�����D�D	gs�X��^�;�O��p0/y�̈uԦ?�.���r�r]	�pG�q��o��S��ه���vɹ�+6�fH����|ljQߜ��
�9�~���������]7��w��C��U�PQ�L�����*�}�����[9�ڑL\��H��3i�LL}��E�*,@>��z� 9��eQz{�;ڤ�Tޢ���޲�����x� | �F�ް�j-�".�?U��358Hizg�m$���Z���w�fp��E��`�+��� 	�zY&�<7�_�iJ��[�����(c�˜�k��8���>Kf%���b���+�lV��a� �=���K���4����<C��6�.��X�?�ٺ��u�y��]��V'��;�JeE��P)S�`X���3+���������5[}n��X��:�YO/%8T#+�X�BN_���HE'�;k.� �G8n��������
��C��\qp)����^��+�J���DO#֛�hS��jK?�K��w���@\��߂����g7��4���������z�^�d�a~i@obzK4�?�@yOU�������0�T�?=�R�A�$��F�2��ow�)?0��d�����`a�ֈ��G���F�e��aP�������t��J�O�א9��\��`{�	���I��w�(�a�p�d&��9j�t�	ex��pgt&(�*b:b�P��f���ۺͅ�-�E�-c��%���$���d�����������	{����Ct5�9q��(����r�� �.��{�<��/ϭT�7��sp��j�{k35#���~z��wD=�"��M=b�g#��/�\[`Zڀ= �[���p��mS�~��r�� t,����#����41��((Ud��5�@_�|�^2o^��P�@8M�ݑ��мjC\��v⎊bVG����k��G�)�Xi�p�������*�l��JӲ������ z�vW��RX0���˳4"�|���s�gJ�a��uЏP�Y�Pw� ˜?�e�t��x#"M�Ӌ����`"�1�Nw�}Y����n�bC������
o+t}5Y�Ô�@�X�oNc>���+�����^�$��t��2X�M����"U��$���;�&}w�JFw}|��]���
��R�x�c�}z��
�\����� �܆v����@�5��PXl���������v&AP��Y���U1���f���mj����"�R�\8`����
J�Y� ߰�J���k5[J�O۠��M������A��93s�󂔍KB(ɔExpv��K�[���}�jm0$5;�aRj#��E��
�?4=��o.Q��X,����]��[�&��=���L��(Sɨ��T�8�Mbr\�Ų����»��1��o��I	枃43Ь"��9�\wӒ�����vMp��G�����бS��#�5�D��?�9�BC�7-+rF����8)���e�[�Ƅ�2Aa��Ƭs -.��lY�'��;�NHR��.m`WJ��f-�֌���Z ����f���[�5�3]�Aa�J���řѢV��g0C�Dy�̕:��|�-~d��nWn��,�$U���j+��].�����sYG�Oz1}'p�{DM�BdP�� �K��s�0�9O"�i���jjAh���1����U3�b~�����K9��s�2~��խ��V�s��z���'I7�E@n�>���S�'|B ����ܝ��Oh26����ɤg�nC0o�Ag��	953�x>��ٛX��k���{+�V��8y4�
Y�S�.��oɢ�'8��M���e����2\����3�P����tF�o(W��tR��`!��rc�5w���bܝ�L���h���})El�Q�=	�~d����
1�&�w��7��R�[��������Ef���N��R��*ME%�!Ox���'�}��k�����M�C��P��Ԫ�{P"�g�-Z�G���%�&t��ʷ��#�6�g�=.��� �0�7X?0\ 94�J0+/�*\�FU��F��w'իYn�jA���޵ue���[фF,��4h�;��E1+��"	,}���$J��]��)ߨ	l�W��܇52r�JHHJs8�w@2e�H�ѺV�V�����s�r��-�MUF�#�;���p!-~ಶ�6�J�v8�<m���ߑ�5I9'��:Cm��I٭ʘU�����2&P�NP�����nc�hԆ�m����rĀd�D�!�a�PY�� p2^��>�{��-tx�����i��$��Nm'����đ����f���z��fc��H&����Q�ː��>��\x�$��2&������6�
�ջ*��5j��)�%f}D����g� l��Κ�(|���`]�`����Rt�Z�(�#�$*�8s2���.�_VxM���bg�<���A�~ȴ�~��:��F0�"�=�r�ބ�	5��i)�7B��h2�E��i@���P3X�P�w�+3>������B!�Sr=^l�W��Сtn:�
�uC�O�c$�R�t-l��G��ာ﨟D���J��IB����l�v�͎q /�oU�x�M��g)���П����K���,O��m�IZ�#L����ȫ��T.�`��x�A��B�N'�}e�V�RQ����)TKh�>�sn�Z�a�K�
: 
1�Z9��f�M�9�����T�h穳g ��,��%Zl��4�:Q4���l'�����d�Ժw5'�!�<Rj=q�*n�dCDq�[��q�B���B���q��HX�A��(8�ϼ?���v	&��5���vC9������y�' ��:1��B��'pٺ&�~�9�'�@���$Dk[��؀ވ)���։�H��!��}&@�M*�w�"��s��*���S�󊓽�9�|jl�DQ�?L oz��|��G�����_��)S5P6�rE4�۞�_��椥s��l�=9$�;��ǁ;!B�n�߬���
WK�h�݄J>lO�_�0�I�[�Ͳ�a�28��G��_�Y�.g��Q���QBL��P��1��0�!�XZ<�[�D�V��*y�=��DY8}MNm\bCD�^�H6����E�3#K	d����Wem�U�iv# �s3�2>��`���t.Z��Ɠ�d���M@Vk>i�Fa���b�{�-���_q����v���,�b������UxP��_��������x~����81���&���Ă$4��&�֧�b* ��6�35Haս�a6�쑈�Z�47�&�Mww�����Q��
��>�E1cϴT�)����lǛ��[�Y4T�LP����|RPM!L}ܨ���,�^�cP�!��1W���J��D)Q�/߶g����{G�� '5X9� A�W(�i��-�@[�wU$ÇyΟr/�O����rFD:֫j�������h�b�0�j���M�bgA,j���~dL%�5v�w�Njq����ލJX
Q%`�W�8���ZCm �����Q .3�b_��3!��������ݯ�F5�tj��ڒ�#X1�A���@�/���ߢ1߂5[���m��p>>��yOI5ЁC�z��?��a	}����ے������tI3�OA�N��S�.�W?���)�2��vu+Y.��kPU�����U�G�Sv��`��q�|C�EF7�so��/m]m����D<�N�n~&W��f�)W�л+��i�Ե�"6�
J�S�.r7���)2WF������ː��k'�m(�~�t�չ(R�jL��8��j ����-d����M�x^헛�������z�K������<jpn~S;׏���`����b��7N������`K�c�+ ]�qM�1Ӡ�;����n��@O�.<�`G�Ξ;����{�����ZI��:X��W�\��;�2����fԈ�H�NR�O!�-�b��fa��5��U�a'ܢ���j�.�� ��yvB��	0O�~
>�k-j��y	�P���D�Oܷ9�(1�zX3uƵp9��mE� �s�l�jT�1j`���4��Ȭ:�Vԝ[�����(=}�X�kZ��y���m"L�-иB1�b�lf�ε��1������-)A�/�Z�����8�m��y�P˭��"|�_���Q�f��/�H�	�UY�Fm8�E�
?-P6�����N�oV ��p
��z%�P,O����K��𠝖X ���D�C�����(P���9��n�h��O.�ћC!{M�O7څZ<��d�Af[�G�@�@߷&��{q�n�M�y���`��Bc�Tm	�=.�oǭ�46x��R�{*Nё��&�	���{Yb�WP���d}� ��$A(��	t�6s\��z;���'�h6��-2 �O��ޣXOy$)����11t��z<,�D��g� a��n\���5�X��0;��"'��5;�W�X�U+`�Uo��,�o��rf">�.��$l;ٹc�|�����*�8�H�Ɉw��N�*,�h6H����:��n�6҂����مop2�h-P�-�ʈ!ҏ�R w������0�0򽑪���Ԥ�Hӄ�_�U��Ӆ����(%V�&I	�/$9�U��8��`%S&�Px��ܯ�c�y����'="Ol���?�C��RJ (�@9|�\>#�����K'�E�=*���[s���'���+��#�ȥ�y��".�>�B�� ����:<4�tr ����u�#���s�E/�Jl����
Ь��)|=c�orq��%7�f"���6IH%"��_.B�+O�E��]��q?d�a��s�`�'��J@ŧ#Ps�P��Q�]J��R����*t�Je�`��n�M��,l<Q���`#E`*'i�7I����M�c���2p%;D�`T��s���A�f���X��1x�ggt� Ѧ�@A�-����?�n��"�h��R!���P�n��N<+	r�!m���uڸl�B��vC/��;f�|\T��rk},�+?�!�*}�*X�.����wm�Ǻ���f-�ys{[��7�����U�&�Q%ǿ\�R"��5������B�n"�J'R��S�E9Q�����r������;�BR�H�=������gKRg���#A�1ǳ�6z>䳉� N@������<��\���t]���T��c�y��6���Yդ�ǵ��^�����yշC�R	��ȑ>=�L,&3�ɂ8֊!|1�/��E��G$����l$b�dR���+Rs��������D{�2�/{����M�9o:@���0i�f4�[C{fG��}��?ޖ�0�0�x|�U�&���v�8�aL*wG�%,g�ǃ�0�e�Ҙ�pA�N���$�J�>9����js���Lx�uR�8wD���.��$�"z�3i���Z(`] .��ۭ-z��@3��nUom�ɩ]v��y�7�?�*�����	L��%b�{?��	 �����t[@�/F^3��D�S�'�?~���m�5w�=�@�
��=���ak�}��{Ai+^���[)�t�;�������j�<����$�Ux{�N��n,�q�����+�}(��!c��,In�EY�z�'��Q�衢"��Z��:�9�N7�g�H����z����(Y��Z�a���޶9��������LO.�G"���0�%"��d��:��b{n^�G������eH��5�����X%�1:<t1jvu*ҏd^��
�y=h�a���$��m���㉬QK3�ݶ�����~n�3Ke�����I9�J��6Ā!�������X��0�@����#�}LA����KΖ�x��9��Yn�v�4ӑ���?���$xE���b��Ї��p��u_b��7��b�Y_��z��k$��(^��"0/�7��ä0�<z������S)�ݕV��9O��O��[�Ab;����&��#*����nP��AĦ>�M}۠"����<�1Q��k�F�	ؙ��7���V��m]W��#\wW����t%������ܵ��-M���l-]����G���?i%�/�K̷J��ZH\�DZ���m
ಐbB)M:�L�q��e�}Z��<�0�"���ޭb���	��1�A
#�5��O�@O���-� �4R~/��H�hR�����||��&�a�u�Z�ƥI�8�P��nå��U�zZ�*C�-�i��"a~��j �θ�M�0�V ���*����O)�t��;[���0<.^�jYm.4̄7l�ǠR��%M�a�P/��
+�g���&S[ZE�3Y�Qr��Q�d `#�DB�_�Z����(��(��ov]סS{��إvC'�1��ƒ� QG��d�141dR�/���E���	o�1J=%]�i�����e�����N\Ad�fB�����p�Y5�r�<�F���6_��+,����2����<t�ym�i� �T���
A@m��лA'G�vW������;g�����A���r�H�x��5��pX�����K��Z����a��mR�mj��䱴�j7�n���ݨn/��m>B�^��D���P,9���ް:h���@a��,N��<���L@�4�N ��7/��_'�Q	�'�6
�ۣ����Q���b�ß�oӶ��X��q�԰�/B�%�V��H(�|dU$�@m�9(��RMg��,�)��"+��B�N�0�L�ԋ{��W��bB��;@��8�c�̔�\��
����"ˆ&u�Û�XQ	����i+"�� �k���;���0m��6&��I�0.�ޮˈԢ�M�%��`f�E9��F��4���$tT፵S1�!òg��Oܹ�Z�����)~8 $�c�`S�9=��!�HW�vj@�6 /�Y�+�?q�S[���J�h�O� 0[g�2�,��,i�C��Mf���w|�|��i�8"m�%������0ܢjF��ԑ�t]��(���a��,ǋ���	��+D�¹��A�
r��"�]�iN.�5΋;�z.O��83����6�/�p�I���*��Z�ؗ;�L P�в�?ّ�d�ɿN[�{� ]�:\qlD�3�������tFn�!):�g�7}M�Z����5��.���	�̀%Nn����� �s<�!�,�s���F�n$��z�-�e[5�8Z�ço�T��]F�z���1<���b��n��Z�g&�p�Ӥm�G���yw�e�a�~�W�K~K���!�ԛT+[�4�����yL64Ћ���_��e}+��[O��e�N�m�����!GIR��3.�JN�V�!���7�ľz��E'�	a�Q��{�����T�'��+�C��T����˥&�DG.�<���;=0v�{���.��;����o*�m��>-ͮ��(HY��:./%nz��Rĸ�TQ��-��я�ժ �\��A3�3�W˃D�Jɿ�`eĿ*��틘���"w�'�C�Oǡ8��X�~5X��$l�d@0�2�/��
$N"�A�������»�o����G�J����_#�Pq��S,��>�O���k���5?��Yu����I�zS`f�B��3Yt ��R��o��dﯼ���I�\��JHp� �����C]^ƿ$y�b�ޱľO^�V\;pv� �PեuoM�#@3�Bwq�uxT�K��k��]�eي��%�\��m5�:�4�؃"Kj	u�$m��,R���b�����m�1����s-D���Yb��۝'yT�_������*�107����
�>�i�^x��sg��o� �E���+�l��I��@ ��7Sn�f��F֗g�4�/(�e�g�ǐ��x_���?�Do����ΕKσ��	?�̫�w!����C���!�;T�F0�� M�G�`�����Xz�c�F�gZa�9Z�zM!�Ǜ��E�G���k1#����2QGu4�%�)�p��J��^����_�&+}�.._͇����;K3��f�~���N!b��Y	��1u̗c����}�ĝt�A]��@#���=�ݶ/�>;��|z��Z�nH�(��ǔ֎�ۃ�&�}��s�i�����a�]��2�!nѭ��	�7���}��x|�=t���w��*��t�p\0���X'h~� �����@S~Y�)� HOG4�|�e۰}.����C������b���K��#�Z��w�����m�x�8���2�	*K�`�n�Ǹ��G)}�{ӆ�z�h�w�DE\���5g,�X���f�_�%�����N�.j�T���||G-Rt) ��*y�����l@}��[��)Y���5�F4]_}�<$̵������:���X��j�!�˪m��Oƙn�>؞�����Q�y��w(����@=�c@�Z5L�>n9B��P����z-|�tșZA�]�d�%f�Lr+w�j����mq�}�뎲r����1�j���|�h�n�4��̏᜻���AN-迠�@8T^�IWŋ�|�m����%���d�f��Zw�w��4�a%ST,`(�E���ZE:�_��_�,�Qʘ&!n�Mk޹�����%`M�L�#��roNCx\�qVw=���K:D�p��	:�cfe���i�����C4]�k�u�h�E���2?�ڈ&���Jgqe75k�(?�GD�i����u��\g�w�P'.NJx�
)�px�����{[�j��K���6/_���?��Qyv�`+����A�^��~8�1�����׹o�h���}�e���`��t��^Q�������'�=X�#gG�B{���zv<�b�X).��t/G�>6��s[�wEw/��a����3�u�c�X��"�0��@��s����pU��2�⠛xl�W8��ɷ��,t=�#_Q�4k���L̅�.� ��Ŧ���A+��Wa8PR�t��Z!�d�����5�,}8�#�Jt{��z~�e��ΓD�:%�L�w��ab,����s��\f��4�bv�4F�@/���W�c��0�ڑ?+����Z�}�����l�g�%�ʑ����rT�]���ki�\@�aԺ��YF
���S�������l�0hK)�p.�/A�{�܉S�,m>3.d �B��!�xk��cFW+6��dB��v�|���@�k�ԠO���!2{�*���dU�[��`X-�\�:ׄ�h�A���\���$4����O����G���em�r,�X�JswJe�����RCt��,Be�X�I �:%f�3�P_�
��	E�߱x�i�7����g)�w�q���~���wD�U"-*�����Dv���yT�@{���~o�I�&��K"[o���6V���Y����ܼ�Xc�)�Y tͪ�y[�8:L�[.��ED�.O��m�3^[B}_/����xg��؊��t�5�BEG}ݧ�$ۮ�ё�����d�� ��J)��sֱH)0/6��C%�	ff"M2��[=����bXꛔ�cf��*)���Gy����s���������{����t�".�-�$������Ҿ�S�xd48}��NNց!��s�9|cDx���#^������Sl���ϲZ1���9�֍RO.���0E�O����}��<��I�ɇ	U|
�6���2�:���sT_��FP⽩��u�ILgb����!�M{Aa����	�ID�2�nl��z"�5�D..���$[���M�[��t PT��X��ďCE�V|�)(0Ny�	fId�X�%����x�sÑ�j��6�U����M�R��/^����4��0�b%�>��7|0Nu���_���NP��|����q>2y�8���#:�X,�L�ه8n�<���N��?�g��w�(��b6�5f�b*+������t9Ǧ�o�?pq_ `�����\���/$�O��8����s��`���׽�bh���v�"� ���j:�Tۄ��
����)�H�@�?���f�q҈A26�xBn�C��J��>7�IH���K��v��[?#)BS��
ᓑ�$6����y�p�d*U��Po�@FP�b$xI�c��:j��rv���� o�rM�u�m�V��� ���qXq *��8�0����+Z�З^�E��K�'�]ȳ<�/�h�dj��b-LF4qt<!R�J�z@�
�N#r
��H*�ǭq�E3�<�)�7f�i�(�e��9`�yn@s�zu�:5{k���MI݂d��� ����	���b #a��\A*�d��A�8��!�}H�#u��u��>�S*̠�(we�����CW^v�:�uT�!��R�t�d	�����#��y`��-��|RӴ0#O��G^V
�"���I�4~n������<��OM��y󻨓s�_��I �v"<�i�߯*4����Ʀ�B�)i�Ц,���%(����i�Β�B��4&`9�j!�U|�9�c�?O@Ԁ��WN�T�T攘9>WtN�~�FF!m��
#��,�����P�E�h:C	
o�p�y������R��X��o�s�\-�=��}��܈�ͪa��.{N3���ƥ^>:FӷX� J��~<%πm>w=�	��}��9�o�~�B@f�韔�vZ�L�Qy��|�Qa�WQ3�&�U�v.f�$�
��`�~'4�f�x^4��7t��wӉ������Bg�r�(%�0�q���q���<�ۣN�~�&Q�b��>nq]P�����S:K__0`�8��"qR�	��ά3��u�a��*����`V�_����!aH�(q����An�bR���<}CX��:�+��m)g?M��C�֦�����50�0+w9Y�Ǥ������ԚQ�kyБ'/��|T@���smI:J��gZ��j����S�c���;�N9��2-w%�F�n������1�(�$���̄6�3uNhK�T:g��9��������[x�E���`�m���j�{��/D�C��;[�Á�.������]��r��2�ݝ1�5��h��v���R5u������ó��l�Ŀ���mj�V:z�d72Du�
��wYج���MNjԦ�"��,��^���EK1�
&���S�T�)��ꜝ}�NOߣW������,t�zd�}��@��h��\k��~>��W��w5O�.Ĥ���O���P��C@Q�R��.� ���)���&�E�z|r[k�4>�F�:r��/���?/������?�>�&ޒ#�^����hTnB��E�e�����X�&7r&x���A��ߺ��Rq�C��'�t�\i�&.�Vz�~h��H�� ��LAY�a�⅟�Tu�������K����}���U�����i�M�T��(Q��:�8�s�HL/��é�5^��� ���5�/ϑ���6���o���	�;�%�9��6�@W��Mx�S�/c��(7C	��ۢl6Q-�������FgE��K#+���9��TM����ڹ�%�/��$$Hk&Ė�tq��/����ğ��Zj�����J������/σ������%�-=:��A�0�2&��TL-Pj�M/Q�lX���le��<�z§xE�g Mc'�~��ۨ4F&�|fi��pzڷj+��������+�h�(�-��.�ǔ�~3��G	Y�6�i$�ǅ�<VHs��I����Ht~�K`�8ó����h���SW���k�0�s&N7Q�X���\��Z���GpjM&VV��H�k5my�"c%��[
��[�f��	p>�h�bA�y�����X9<���8�Y9��I�<=�N��u����F���S�Io �Ըr��٢��������V�p�G�S���yhUJv��6���@�E�I{R5߁��Û<yP� XD��������Ƶ5�#��Ԛ~��؏u�Â\�8�A�K�xG�k�?�\�@bgPW����Vũ�RV�x`^%mbo��V6�ݢ��Y��yΧ�����~t�y̒�$Ѿ�^tB��akdb�]nd�������fx��;�vS�Z��1����E���Ƒ7�}T����=s"k�z��3�M=��J �1&����3�6B-ؤ�՝ ���5I7��k�����x*~t2 }�Æ��#Ӊ�2�ګ%�e��bÝ)�b@�8�n5�$�kT�������F�2�
sH�)2���
�������u�L����s�k���ݜ�f~�Y�=u�=�e�(�V^de� �=�;|�U��Ϊj�IRP
(Y�uu���$�8�w���= s��Ò�i��38�B�ؠk��|~ΡB��������I�2��rl����7�\�we�]σ���$�
'	Ta^Q���J���1�Ő(�Cl��!�+f��=PA 0�X6�ޘq�-8I�Mb��5��EĂ�Co�K�<Ц'�銎�����0�騄��� "���hrpc:n<2��!�_�g/޸�,N�3�d�	�؟H�kW�!0��@��'�y���Ų*��b2` �[|�� ��K�iE���/��pe'�`*7UN&����\l,��͓�Ž��0�y�#�0���z��<�"_{�#1cz�J��RJ�C|]7
�F.�m��v¡�v�&��6�e!����^wX�p3!�߆JT����^ћ"|��#��}�sp��86�iZ���n��b+~�:��O�%�1 �-�ֶ��H+���G�]r�5��C�K�_�p`���E��)L�9��lה$,�a#��Ȍ��˅��|#�G�x��/�` =���*�Z��2Z�������<F?���r�S��+�*ԁ��p �H���A�U��ފԥ��	
}B�g;����ٸ@{�-xI��ᅢvO�Xzk!�V7l5����,�}�u|�T}����}�[�+���m� ����U���vK�/�O��'�(�X��AL6+:��������n0ΘAN*Þ�\LW�P�=<�2~E��3�6�E��.�vDAH �l� U�@���L������#S����g&��Z�wz�"�#֔�o?d5n���0�l��#�\Ǭhm�8���==�IϣS��7�~��!����'�N��.@�L�⨢M�0^���8��8G�yV%�|�kTsO���B�;�6�����c%�T(�@�����3~�uB�<�Ǒ����"�L�>j-w�j�W�I��uR�6i�睑,hM˄[h�5�o�
���/��8n 6�h��)�Di���Z�ާN�ۋ>��@�S|1�S�BO��܈�
��$� �}2( i�2O�vd�,��I>���Q�AȲX��ٶj�ݭ�+؝F���i�<ٳg;���M+���vh�V�\�a~F�D3��v���M�HWؠ}O��ۂF!e E��!���Ax�����i_".���U���@D����!(#������$�Ұijs�4z�������S��	tPؕ�B6?�7!�6ڲ8
���`}s*�k���(�R����H
��@%��h����P1���zqVdB��s~������n�w;dVE�i_4��	��&�0�r��p��#8���\�sR��k?e��(��@Ǘ���<B"���m�'Io�C-����$�ԁ�c��������t�-�`%p7�>x���jsH��ç��}M��^�w��7qE���TMI�����%�7$r#�"�f,���Dgy��z��ޘV
���9$�E��^��fs$�p�	e���ྍ荂�����l}?V8$-BE@�	�H�|���As>xR�W��픧2Hf*	��h�&�팵�kJ?�������ș�;`�K����Ԗ�����iig�A3�z�BSh���nt�u|B^��<���e��I/O��-\[Fas���d²)QD+y	N�@�f��f�(�`n��8A.�� 0�6�����^�Ht�W���e(��+K��\(	�>�н4�B5%���ګ���?4�I\�'�@�+��H~�M<���E���#=!�>dk�4�y5�>���q;��C[���	����d��W�d��娘5�Ť*OG_��S7�@ɾ�c�	�x�ʩ=���6J_�;��-�딲���zp��E5qO�$���y�ƠS͛�QL+ �w���s8����UݑF�ot��ǖvYǢ�)�B2˪S�Q��Т7E����u�y�J[i�~�*�Iv̍��j0)��2�C�����?4���d\WTؖ�3$M���aF���:���
���9��qT7迉�b^�`G�DL�{b6rE��T���	d�c �0m��zvl���LhБ�6|�*:�����Vҥƛn����TJ�p�+�}�W3d�	�hTP�~2��D2��d�b��/�����(! F�).F�����G�����Aj�����	�2~`��>��~�!؊Z��$��1
� �z~4�;�k��=ۧx��8��>'��/���#�3��HG�m��G���ƍ,��,��ί'��8gTq����>�j��#�ɴ�M�����O�.uD�Ȭ!Qs��8�q���4��	TD��o�fC�J�&:Gi㌰(���q��$���I7q����8���_��|�c��]w*�1PS�:E1E��)�q}�?�@%���L�V�|���X�g�I�0���},}cTB+媨b|"f�[U�y0���k��a��C��cb�#���[��)���>z��H���i�Eso
cd��#�uK`Z���9��,���{�h��M��I��������[Ѧ����+e^�n�S�@[�)��&�޶�*�Nd6PN�"���'xGIɅk��f�Eާpv[�>�*w�f��G��_] H����$�x���v�q�U��d0Q�0�:�?�~�K&t��g2��&����,�^�Gu��D��LD9ť�PSp/[!���S�� �;vLr�(>4�
1��oiX��K+մQ �O�
0c�c��FIy�B�j_i�]�R<c٫��:��dV	�AY!�D,kD���E[_h72s��S��I�^E�< ?z.h��oz�lI��D�~!AЍ@*�*u��X���v/����G�r���|�+J��M���,�gT��'��H���v�$vF���r���Z�|=��p>�@n#�����;%�_�W����O��$�f?�e�'��`�
|��z+Ã��S�B|Y\��C�<M$�<7�@��K���*��A����Eƅ�^��l�4�Vq�ϒ�:Ŀ�8òB$$���e|���B�I�;к�и�t�@LP;B;Q'-%b�p���0�}2�I�,���j�Y��F�s��6==eO�'�oWw��56�w?�F�rq�p9SS�P�����v�<U�f�	����O�	1��u�<h1�.�2�_,�B=�x����\��)#�N�^�:�8���p(�`����3�P���a�Fp*�B^0U��a�ȭM%�L��vbрcS&�>A9M�U����Olŗ�d"ފµá��
�i>�����&�lA1�>�Ɛeq�!c��M���D�ԇ�;ί�� V���42&/�2�3�_t��@+�w67�ՏK��e�~j�`*��5s7v�ܨdcxbv��������d�H?F�j��s�w��miL�q��I��]�,I��h�[��`0� #`�I�,ɢW��������<���k�!4!)��)m&���K�MU<J0�=l
O����ww��Qib3�p�S�P��:Ut��-�xy�6�P���n�Ƌ�j�����.�qۊ�9�=�,��Cb"!�k�y��gҕ%)y)7�@�,ku���vV,&V�o+�H�c<���)�q2�i����x�77¤�+����l��g��ٲ+�J\������󙂷
�!�܇|�!�0M����t�1�
�{1�#>A�d��/�V�ŴĬ�]�-e���>^�c�Z�E˾�g��}�ϘJ�/hm�xR���U��l5��9��8���r�[G��O+��3 �"S�*�H_*��L�Ř��;�Eee{�.�G�6�V/�z�C��h̴r���85��G��������X��+Q�V��ʩٚ!^/@X��6���G٨=Y�X�����S����+������K9y��	�	��[2B�ߊTꫝ�m"�����`��w2�^�Q�6�_��23TV�"C��j^I
,GxWfM�?���IK	���iB���W� "�zëi��HP��ޓLw����U�~�ks�4t_�����c�U���[�Z"S��z���ˈ�؋�^`d�����h��W�̝V�H`R$D!O.,�b�<,Va兿����_~���L��i;]�+�B�Iǆn �����"c�]P\6���(�����I@��)ĸr����zZ�Hr V8o�
A�
h�a�vJW�����$c5W��JN����%L�͘�l��*�-rU��iMϦ�96�XE4GD�j���~1ɳ�`K����-u=Ś�%���M�N��	ɩ���J ���"�38�¶��j�H�&�U�|Co,k�����#vJ�&�@���f�3���}���,��ej)"�`s�|67;`f�"�"n��U�-T8�l�ǭDCU&wƘ���5�����S+s����g�����j�9�}!�L.����x��>�J'#�\��}�C
������:}����y��f蚽4m�ݎG��a����[(SeU�L�l;+�ȫ�e3��N���A�a9S�u��[�w`N�Aɮ\�]e��ƹ6~�	�9 b���4tK����0^u�<6��{��s�T�qAu�����}ϥ�.Ri%�+�:�Y~|�\*z,v3Өj���4�t�K~��t��v]�~2�Y��G��â\Z>�.��S����+�&��'�6�!���I#N����aԫ�;G�7���v�x��/N�	uE�qH`��^�;2�C�h���l��,����b7��jl���Zp'�Iߤ4�{�W9��ͤ?���P�tw�����:���
��4)��~�s���i�F�hY��������l�mfUu�<s1r�tdŨ���i���|씨6�Ӽ�9]������ecE2'�u\M�k8'�t�T$�uJ``R�s+�6�ʖR�{��<tH���"8��P��b����#Gh�R���P���J>�F��Bk4��L:�z!�����E�q�J����w���6Oc�G3��R�;������I��+��7���m��W�&�Z+�'�8=��F�(eۜ��<�m��༭�I��ﲬ�����rfs�:i��"]�����J��kL����!�ҟs�c�:τ�=D��_,&�{p���F��Ij=((�qlU\uɻ�_����{�a�*Y`6��VK�*"��F�Wapy��*5�ˏ��lw�R�檑�d$���l¢`&j 2n���Ǣ�S�E:�rœ
���yI��w������?��4�:Zu�_�_�l�h�w=���kV��� �Ab���ee��L��%��z�n��=جx�XR�e�n;�X���� ~Wz����[�a�>1	Cx��}RP$bYI�`�'dEcf���P��C������H
��5� �O��/�pi��9�ja�݆��@��}�>��;;��3;�k���ܡm�ɕ��#��{��!No&c�} ��o���#��E�9<V4�4L��9FF�k��-��b�l{����JO��K��x5-+m�mu�+����?J�Y}|+w�<�F8�ە`�;��	������뤃�0$�) _��z����E�Wyλ��A��|ʣ]�.�����yTv����8W�)J(d��5:d��z��q	�=#z�r8hh8/7S+�Z�lJot��~�}�>] q�Z,���&��� ����nn���ަ�P�J;p]4���?A�WE?i��a$�6�I���"3x��Pԧױ�,�H��3gn�SN�nקi�LR����N����g��'���.�=�7B�Uy;�P_$L��zqH��^��B���U�%�>&UM L�;:n�kh�A�	@�=�d�\�k(D�WU/��97~��P71;�3^78\��-������aT�\{�1WR�/�&Y��8���k�Ka�Yҷ F,�*Q)��,x�tȦ�ey)v�h65�dP�fȰo��X��>�3�%:��Æ�<2�R���ba�&�7��p����.���Q#����7�����f��n�ͩ 	�Y0 �[N�502��8@�}+��k�>����iP�p�u�Y�`�k�� ���Q�N5Q�D(&�hN�]ħ-lg���9�^�R��z6	C�QUP�K�,6l���_�D���DE�Z�B��~k�v1C?�լ��`���*��|��	C3)��F١gA xY|�-�[� g���}ׁ��z�d�/�8Ml7a�d���ٿ�Y[}�ME��X�$�u�����޲�~״�F�Shi����t�Ek'3)����F6m�ȝ��4�ʘ�x5��Ʒ)���D��#/ �: ���[k�ԕOkcNHo�>��"�2䌂�lH�C��n���4��/]>\�AH�i�ތͩ&��M,�pǵ�0����������[�~"^n��n�k#\{�J��P���9�<��iצ���,>��gm����h���/�G���=	-�>��{��Y�U'�G=�{ڑ�:A٠�q�8�J�\�n2��Ú�+S�o�7ka���~�krĭ�\%DI��f����=��* %w�ݪg�
}���>c*V�H�Y�,�P�@��H�ia��{D�&�NY�\�'7�V��G��rX���8�FVK�HP˞���K�h)�ZW�����|'�bn�-��/�2>:s��P��/ߑq榦t���2� ���.�E	�B]F[D݁�0��Z�L=��ܨ�A�o�U��r�@�?h�N��>G��$u���
��=c+Y�����M8����i�ŧ�P�-�����q ��y��^U��i���\;�����n`�9�@��GM��r��)x"�Η�����7��{:�>�����= )24<��d:�+��'/�74x�$P���x�i��7����Ă����u� k|Q�ouv�D�]��w"��b��n�x.�t�2JDA4K3�z^��W�ܱ;�Y�"gץ�
���?�����WZ��pm�04'�>�����K�ة �3q7t�ma#!��>M��L
�~��-Zn[�R��A�V΍����Z%�v�lP6]+P�]�9��i�ֶ�&<辂/
��T�}0�$�}���M*<����d�2mИ��"��5���h��k�p59pu�6�
��ݽ�a��P���{v��G��hZS���\����P$Pm���n������|��3�S��'r�׏��:���I5O�o�li8���w��%B�(K�y����R�8 ~�"|�� B��c��1��N/���7��726�l@�i��/$�s���CF�|9�4ѹ@��>�h��Z�RN�>�t�U�ޛ�߉d�(��ي�2\�=4D�+)m��v�ء _���D:IZ�'+0/"w&�yf����ӑ��SGi��V���9���������~?5k��O���#Tw7�Lmd��H�xfb�0b"���b��6����+2�?�˿fIR�=����Lֺ�׼k��d�Oeߦ+��ÜA���p{�'E|�n�ZfN��>�t�=U�p�/�y�i);��%�5��
�j�&k��b��ڜ˯"����_��4ɛ'����T��K�xfN�� �:�6	s�ZߜK2���Y=�׉�|�xG�/L^���[W����=��V�}��ާ�,�x�����I$TP�fGZR�%p��d�B�����z���FI�Y������Wm�V�\)�Ī�%CF�a� ��#�1�J�,N�"S��������t�4���^U��/�Ia 	�W/z���6/@l�t ����#b�}b�`��W�h��w�lzs��:M��>�P1�\4�+N9Xh�*"WP]��b`��34I�[�Q*�k��I�3;'���/�+�w�x�l�j�W�:�)mwN�~e	iJމ�k@������V��n����WT�$��ܝ��3s�'��nj���-��uB��0
�g���-�������p��tq�z4i�&\6��Uz ^���BQg�W�A�9�@�"9�Cc,��86,+�W�ڙ�Q��u�t�&�	�݀�+W��k7�Đ�K�v�}q�2�\:h�2'���
|Z"�OB(gv�[�K���� �!�<8v%t�<7��B;��a�,�׽[N��q�8}F|�2���m,��n�Kӱ!J���h"5����_��9�d��d���pH�{s���F�tϔ���T�9�N@�pJQ�bOfQ��`Ѱ{ϡ�>�Ɔʳ���0ף6+�X��/�b���҂����6�&��DK}	���79�$��c#�Ɂ5��b�����a���{� ]���#Յ?���-2+���8PgX�#(�RxlCov.��8��Uw�ø�ӆ��;��f_����r�N��my�n�[���&O�ԟV����:��#�L�T		4�_��>J7��W�j�Z5�˯�л@��B��Hڒ�	��y�A�X�JM6~���41.J���������c���ѯ6�c�J���<ْ�Ō�jb�����[��:�׈7�nA
&��B�g�ͩs�_������Nk-�+�S(K
���س������c�δ����=�)�e�f_�Bv�/V�Σ�y�����.�7n8g29{�bhy������vfK؎�P%�k�x���(L6��*��2�x��^;`��C��r��R�N�P�IH� /ß��B_e���p�ᙝ#uӸ�>�r�aO�]�����caw�����/�����z��t�:���9d�CƇ�j���0a��a�W[T����֡dj�܈�c⇩$D{��o�b>҈�Z)�F(�8I����$xe��__Ԇr��c�A�$Q�e��,�3o?Ғ�n�A����=G[H� ���}�PȽw�����C�=`��ɩM2 �({�O_�Gѓ�U3��!6�M���Y�
c@�e��d��+�,ހ�W��Ҕ�|Wh�b�(
�Sbpq��u])Ʉ��^F)s$��>��(Fc����
Uu
�i�j����%�P��0�
{q��*hhr�L���1�)sV���< |�h:���0����&Y�� ՘W������e��l��8�]�߸U�Ңј�����/��~ͭ��eN�{��'�ܙ��)�p���挃�Q�M;�X��T˺��F���Q�����b㒻��4Y�ý��.|+�@��4&�ԣ�Nd��S�+�X黶f�����Ʋ�8[\vӱ��9?��p񯅪�N�E�Ie�ݴ��wp�At��@��)-�ŵ��>mm	�Oa�������LL/�� �n-|�-�1^l��C�	R�ܫ����fi�}̅m��y�{Ts)p�ё]���3Cm�f�
�E�4\wԨNK�t�������Ƣ/����4�2/�.�&�l^�s��]��P}l��W���Wa# Mצ��K�ݫ�ar�^U����0��҇ԫ�5�7*�2Q����A2c��w@�_��=�ۣ�M����)k§h��L��3���yTW�Z�mA,_��*֙ȶf����ؔ�0�8H�zF�("
_2�5$��؋���я:� ���t.xs�V�e���:���hZe��&}e�Hg��=������?��w��Khͧ�����؝8����n�^{����	���q9an0%W��
~�m�W��Z��)���`QB�r�Ku�+7*���2��iю'8z�5*�e�L_>�H��׷��P�1$�s��;p�=����u�ɴ|�m ]5�nL��\��P���ˇ�uCaQ��g�����˖@����,�@֐�V��@fɸ��] #��#�bO�4u�������޸}�O��b���$,6b��v�gBߘy���_��j�. �*�-�Nq*ҩH�'�[hPޓ���e:��f�{Y^a�ݰ$sه����Ɂ�N�ϞL�#'�e�J�S����ح4<����s�9+B��'6a���U)�o��uTl�C(�D��D��Ϧ��7�p}���pȪ<{Gg{��í�5�~��k)�H�'�����δ���e�-��|]CWB�ŋ�ʵ���<��?�@w��9�	�@��oD�<�8���n�
�ID�Ԅ����hZ��N�f�T�A�Pw��-H�d�V����+>��D+Ç����Ē�_��M�ȣ$��r�.�)�o0���L'�{JK����S�;�J���4��0�c�&R�г�_/�n6TW�w���&���z"��֖#ZP\_.��
�b��dY7g΅�f�y4\��������Z�|q)��s͞��m�3�2o���*q�*��U��e����ď���R1>��8f{�����g��~.�� ���3�v��yab�5L(�TF㎒�,ſ>�J�lʮ�e�m�tw���#����d����ށ����wҤ�?o��uxx�puF�	�A����{+��jaR9�gS�o��ԝ����H�-���`�y�����l_)Xd��͉�.Gw��+�kK�6��M�d\��z�9e�L���P��h�2�� �ҒBC�%�J�]�9��҇��~���q:�~Z��5@����ay��\f���˞���S� /�G�YS�ҕ�0�ZY�P7�$D55� 2=�jʂC�\4�<��!:M��L�N<�X,����{�ǆ��T.���m�w�FT��*B�w���(��d��G+��AA�J�<	:�ۚa�SぺvRt�'U�-�*��nX	���x���[*ό��I:i_�aO�S��o��,�Xe�!���+�V2izD�c���dKw�j�?�S�_��*�&qS,��+G��o���,R�c�k�iq� �Q_�ܽ�*���q]w�T�t�
�6�M���E���Gcb}Ay}'�3�2v����D��r��;}h)�/ o�Z��|2k<{���]�e2h�u�{㍠�љ4P l r\�xM�v��( o|���Ws�X��=Y.���.^@��v[���>7 Ǿ�="$%�0�-|D��YkѺ����!/��'T�J��l�UV�ԿJ���+�A�MF��<\�q�M�p������tGbւ�\l1#� ��$*��@XG]�Z������V<\��0�@�ᡉY��Þ�kו� N�f+��#.	����
���|fPn���"�-[ֲ��H��ѱ�@�J+�K;�J�Mic�`�0T��a<�E��z�[�L.4�8�*P���5�w�1�G���K,���m��M`P��a������kWZg}�y���Tq�S?���ϫ5�]�!}�A�k����i�1��^�kD�d۪��o6O�w[�q�@�sZ6߬,�kP���%_�G�29�����V-D�Q��a����<�<����]g@I�:��a�1LL�m�`���q�G9Fcd�q8�K�}�ޮ,C�AA�1�@�h��ˀr���㡧�tZ���_��b�uf���器߉z(�jTS�D��,���Xq�u�]w0[4�gZ���:<̚F����fR�ob{��(�a]�x�l������g��A.=S\pG��x�EG�-������!Mu=������=ɵ�:�FS遒}�� ��W6�laE٥!�"ϸ�ِ�r�n�Y�t�>�q��Rt��I;o��4�Ė��8�"�	�o1>V%ywT��(\ʷ�^"'!�)�y�q�`\c�P�ң|�N���8�R/͹�5��r��4��*IM��J��ӯ)eG���4��b��ۇ��h&���޻�u���̨=t����v�q3r^޺���V�\�?Bb��W[4�����_y�;�u8��R"0�GQ�L��$�����y�az�wG��꓆�MZ���l����N�t��f��T�ʁ��R:�+M�Ve�U��ʱt���j:��o׏�i^�h�zc��|}�ի)�(݇�j��iQR�Ѕ�#���_y@���f>U��w=if���X:��㊔O��J�o�Tj)oSe��vYs���$
x,�D�w4���AB�@�@s� \�k�HO���k]+���XU͈M���	7c�;Kix��oW�[�Q��)�Q-x������bx@����Eb1.�C*>?}��w�j�������w����B�h(4��QB�9| I��b��>�'�t��*�u�8!�K>J���K=�V�l�t0pcx���g
u�Z���d~+�ﰺ�c��n�ey7�?/�a ���R)Gm؊�O�����{^zT̒��ilG��p�Qt�K��:� ��-=,bʮ�x [�����]a�����%b��*��}�<��*�a�.Z�E�ڈ?]R��(��k��@�=lՇj��Iy��F�6U�LUJisvû���NE���i��W��^�E����%�ޥ��!aXD�-��M�y�(�C$�B�Պ�H�Y~�!j���bX	u��G\=A�����/��&�o�O�v�������B��x�X�&݅Q�ZK���_J/�hRw-񝘐�z�vy	� u&�yi�64��(U�Eꍄ��ۓ1y��4�#@�j?�e�:��.\�����q`s�-�;�`J�%ý�9���1�B I����A����2έ���7�Q�$��3k`{�H��(�S(,f|&�<�B!La�l374q#���Sg}f����u)�.�LQV\��0&��]}`[��thQU��5$\7���'=�onq_�ɗ�TWF!�3������?}s`٦S���+��������+b�1[T�*<���v���I�n�7l��H���3�ŵ�������ٕ>QZ>�{q��ܰ�QI��c Q�E��8Ŭ%��1����9�	�8t�v�[oc��b�תБ	4I��и@�PͶ�ك"�ZQ�\�v-B���|����Q3�����_�7��qӯ�h�j.+�*�����F��*���@�=�NY�� ��4�_\�}�೑м�y��fw=�2bvT�/�����a��n��!X�+�����D����~a�􁛛�D��4���˹�[��
"�i{�	]m�Ju����^�֏�X�na��$|Wm�{#ֵբ��ᷓ�Z4z�7�[A��Uϗ�~�9��D���&m�%�C"���{_k����Ɏ<��ǢpS���S6m��-�[?%L�䠺y�:����>�ɦSW,{�����t��{n���9�~W�H���B�[�i����u;>�m�l&����1/�^���=�	�OO_1��K���e��B? 9n �U'i0��)�}#є�ԡ;7��*;�T"W�y�:�U���v#52�U�v���x�-ϧXJu��F��je����C��"�E�c��0Uk���ş����1��dÜ������5����V�lͫ���=2�m���*�����o�Ү����B��b e����ɗzc��iÑѱ���)7�?���h���q������6؋�߶�螨̒&L^[,�0o�|{���OU�\�Il�x0��=�M�y�n���e��:��'ֻo���>:*3�)zv�^`��Yh`���-\�)�#�oNH*���Z�W6s�ZA%P�F'���4�����>_�O�(9fw(�s�/�kN��I�Z�t�U�n�7͟��EXu|V��V<��e��Dec���^����g�8�� ���9Q��Ĩ	p������'���j�S)�to���u�yF�#^�Yy��hZU'ΑUz=3WJu��F�D��&%��D���+�`9ސ�4z,��U�Z�+��H�e���9I�er�N<}�R"�(_��^��<��1�'�-x��'�N�حX��c����rH� �$H�$T)O,{:�k6�\�݋�z���/ͧ"Y���5?I��S߫x��Ɉ>l��ݥPqP�l֑籯�SԬ�S��M��V2H�Z�`�p����t�R�Ö��N�z�40��b��5N�KS���{��`u�f�#���K�:X�`Uډ�XE��X���H��_�Ja	O�,Xg��4�<C��H�s$ؚ��'���6�$���1�.�*��:Eꥁ}�-`R�b�ˎ��K�^OJ��*�&;�)�7q������p�A�� *x�����>�`�n� ���+�CH�pת0�,/�����R)����9�7-�!�A���z��,+6��g]���[�g���~����׋���tlϳI8ʑ+��6u�3Ll`^��x���/��n�`��vi���Cx�`w��"�����u�D��RV�= b��X;�#�Jlw�X	�I��c��;<�
���"·���䛀���u�
=�1:V�	jvǳ1�gK�����es���r藘7�@�a��2[6�O4����D�����i<�ۜ�P��8}�|/Wi>;./c�T}��OQa��u��Ꮍ�s������������<�-DiA�5�^6�V̗����pT09@��C����sx=N�q��q*��x��`�Tw��e(�:f�Yh0�TyU��>��4�/�e�",RT��&�)2� ݳI���W�Ǽz�f�@G{u��mC�o�jܨ�c�dq�7��nPܓ9����!~#���<r~���*���cTy��{��p:ֻ�tT���6ж�C��jyB%pb6���H��$^�R���k	�|��lo�F�N|_%�pb���oQ�"��E�.*�`�K`�lb<}U����T�m��.]�TZB]��\�{�,�vg_۾:����9�~ր�\d��O�`���m�����18����xn��ƍը��{�H���<�]�D�)[��}��4x+���.8�w-%����IΘ1q�yN.��6�V If��m"kp|����'��囮{�}�n�Q��N@��\��[!�	�b=����b0�W8��a�R5�Kؠ�'��s����ll�eF;������� ic͙M�р�>�?"���p�˷�����3�[��ĳ+���If Y[2��7�6p�/`�K�׉����|�d��*n80G�Xf^N#-��@_���x���i�3,��Տ��X���u����b"2����־3.?�����MT�j*�u�����2�DP�6���q�UOnw����'hq'>�a����&�F�(��J��Bs*�(X��F���*����8A%<F(�p�0�K���Wt@��g��HԄs�#L�a�	2y0������v��m"���G����B�\+�J�+����8����#���'�ĿS�𓭛�Q��9$�
��R��v�t=V�m�C
�F���Ƙ��?�sP`qM���ċ���� �;1<6c� 0��'�ŷ�9�ߋ?��/��J�f�B7lYi�� +=��Ł^ɬ��-��M]�7w	�#ܬ��ԧ�pw}UTG&2��_y7��%��-|��)�e��P=�n$a���tЎJKzf1_�7��K<F�Y3`��)7l:S��R�(`#�}���w+��I�\�[a���Bz^=�?�*?�r��ri�ԋ�~�c��rB�2o��}����1���eTu	�e��XT��ա���Gl��:�͙���n��\��}k��>�;�c24���_o4�!��v�'�a�aREgI���Û�O��p�&Ö$@�P\$4<ꓨ�<Y�yM�	�����_�]�� �v�����wS��)���?���Vx<.Aˀ;��b  k��E�R"����;~��D�˳B0*zR� Β�K�L���)�&�Q��~:/�'��n����i`���4�(t����B�r%���	C^&2ג����$��55]pal|�R6���l�N����F���N���U>��mg����g���Da)���_#�􅧸����C

{	�*�Cn'Ya��i������1o����"�����5��c닡m�u!�S��?�i!�dƦ�թԳtaM"�>ĶV�t Z$~~`"��y:����:L�Ҏ���~
fi�g5+�k�?�~ْR8d
��hX�G�dS�OFI��K�)��r�Óy/�쉑2ͰZ4���)3C�PU�N%��4	�����RS
`�<¹�.*ˈ�H�;Ցi��$<A��P��s6�˟Jh����ͺ�a���;u���u�����p7_�Ը��?:������,��H�K�t�}������,�!� e���'�{©j
\A5���ú�x�l��6����=�W���j��=bؙ�P&��`�M�lmD��vW۝<�щ�8�Rx	j�G�������Y��Ҁ*�����#�Jj뻦�[u�3D4lZj�UY��`ˮ�����'2����zBB��F�J������@47�a6���z%(ɀ2���S&�pZn2x��X����"#��Բ�^5c��DË�f�1	,qnw�������S�á��ь*��Ɇɖ��<y2���"*�I������=��O��,�:����Ou�C#���dOo���2���%��I�@L6J�A���[�9�]�_ل�w��7��lȮZ�ղ��M	�Ǔj$�ϥc�|�i�&BM�k`�!K�N-stUA�)=0BQ�m=�+CH'�q� ܻ�|����Y�P%�?����=�J�� �
 ��$�&U��	�3�{���:��!+�t�I��%'��u���I��s��W#d=Yz ��<��䌂�Q;�7v�F���I�r���v��1w�CQȻ��9N=�uV
Ԯ�4��Y&�\��Д�Dx��{ n�y���q��e�8b�"�	;�YS���{-��׋N��VW|/J�����!�}�8��h��G�M&���c� �>�I����5o� �=��&���g��W�
[��~0Y�� �{��h@��ſ��|����2w����(1\D\���bBJBGr��o�'��̰>z0��ނ�}�J{�r3_��BI)7G���?)#��gPC־�m�0�z�ϟ��(�{��R�j�h~Ƃ�:k�f�H/9��DB}��f��}�=�Q*�,svCD�FQ U�:������#ZU��KK�Ӱ��%Wܣ���Aq�W�sq��x��dY��<���'s£��Y�y��c���3[���8�U>���{T@��e���z�/��x۳'F �i�c ���>�+x�>JY����p^h`����Q�&.�j��B�,U���c�����3M�D�q�L�
M��3ؐ��y�?�"�<��g�հ%)���3C���<伥��7�� ��r�@V����^��^��V��T����s��BH5"����"��� ��j���O,eqá�R�&P����݂�5o��2�Rpih�sf�L��@L���w�#���R�̃�*BNK�Ȼ���}�cA�0{7�و�J�jS�	(|;X�<rYO�Q��%AX�aO9³4GT�C� ���N���H���0��$g�ۈ@);���@���`��D�hyB�lQ�����S%����}>4�>睋�Ь;��Ϥ=�E��c�I`�yP�M��4�w�ZG��|/�l�����*��9�����[�fكO�S�-%-�O������5c�Ǟk]�]k� ��.E
�)�gד8p����\n
���:��ˇ
3�J4i���TnYy~P�1�U��q��B3���i���O����C�2Bb�z'@	m��u ,���B�YV�v��j��p�C�Żt}��r� L�6��1J,�9+kz�n��,�aR�>��C��hzR|7��^q����E��ӻ�"��A�j,����Ө9[�0L����F�LR�3[��K�`�Jp�8�/aAY�l�mB�?'= RH��x�,�a���'����<)�QA��\�t�/�^m�|7}�(�[�7'D�@�,Y
�����5s��4B�4�xmp�Ǽ��&��q��l����_�L�Z�(�u�Sryw�nX��t���og�!U�]�z����N�<�S�kgM� l�p{�Q����}���ӝ�\��B��`����0�0��l2�|��b+��2� 
W�ǲ͓�4�l0d�W��J�s&m���Q60��`NEEC{�b�$v�!�:�i��	�Q�j4.���|2hd~dw\
�iv�J˳T�㼐����s꟪-��Q�u��C�nH�T�.������מ&��Q&8Ż���9�O$��:�Hj��$kO��t(�5
������_���X�7���m*���n�S��̈́�((ti�Q��W�xJ�K���~����u+���r�?N	���1�qE�4����$�կ������� �F��`S�#f��J}
_(�?)�;!0��~,������\�PPk�M�p�SR,��Z8Y�
z��)/��8܏4|=?�q��>[Bi"\�Tk�cz��n�Ѓ���X~���g�w�c�yf�%қ���V~WDcG]�� ��)��; ,S,P<J7]ڿ�`=(v���� $���3��|>�q։�L�l��4�,��z�N5����B�����PL�W��g����*H��n/
��ʟ�n�R�&~?V�=�4{g���R0��K�8�?�tN8�߭��1��3<������E��ԋ�뽭�^��E�;��F�B�0�3�ű��&�а�E:����zA4�n��L�}�@`�5TDo�9;�z_��w>�l�7�$���4�����#�+bN��:?�V�NY�.ŀ�C�]�����5��?��o�I���Gk�MYd�'*[�4���j<"{Ϝ���6-�e
}Gc����=s�ٖb]��m(�s3���T@��kR-��4�g��hr�8P�� ?i:�?U�qx̂���r��$��f/��P�=�<2M��F��7��R?q!ϳ����\n�(=>�{�~���I�fwr��#+1�طx�{�ֿ/wp�k$J!�GܵA�z_ ��������o=�:N�`U<ކ��,o�-��vԫ'��'��9f�����E�*&m�hݸ���;��jϗ��~��O/��o�P����+@��1�M}�_z�ט��Lqp�;>�`��n�����G�
C�|杴���$��';��׾�Ò�gY���d1�8�8���ѤIK��WJCmPL� �AR��4��ф+A&��.�Ȇ`aDa\6��a�S�,SQ�r�2�i��M�i��S&=� $�}S���?;�#�M���,�
��UZxGy�G����K�i�+��Y�v��q�"��V7�d��Vy �����у���UZA)�5:m!+�%�	��E�[��l��Z t��ӴS��|���,*�>4\�$�����(���,���1�0ue9�0
-��B�vC�C��ZB⹐e��T�p����;��3!���E�onԲ��}O��*�i��6�Ax��dg�_���@Y�\�O��n�98�<��Q���[6d@��3��������dyq}�i,�F�=5��V��#�߫�`!� B�l�@R�d4B9Y���&i��f9)�w1����ӵ5��@'88�t��u "���0S������VI��pPIue��"�z��ulP����P�+x�]Jm��;���M<�р��'JP���;���5|ᐺ\����=8�<gh�F�������&�C���+�����Rxf��(���Z_���7Ǹ�������z�̮��
�u�(D����-�A	�n�!����U:^�)ˎ@��:��R8?&�M%Z���ӫ�S0��(^��PUP���ѓ{���Ⱘ�,0���6�y���� ��W�+n��4p-DP]yu�p���c��������(2\z����B� ���UC���J4&s��-����Ou��"�j��@��q��t0�����9�<ZZ�S;�܌-��3}r�]r����w��-�<c+k%ǽqc����}�ۡ<��0[��\��k��5�c+�dxR���;�B?q򊒹/i@k�B4�,��@�����N=aBxﳺ$n���V���N)�nrHi6q.f��lZ]��?����`$/�@S����^�l�y��7n�1��ʨ�"*"��ey�q~����x����ܪg��R��������5����7��9�]��<m>�n����#�ĵ�嶺�H�~5��j�4JN���,�,lG&[rv\g'��̬���-$����eԺ!��A�V�b�b(�/9.�rn�;٬%2�R����Rl{�'3ZC]�	��<�dP$������$7lG6���.����M�h�&�,�s.j�.4�����B�ΫY����fڄ�y�^�f����7i����D��2T���94�0���ORiëF�G��7'Ő����㉈}�DTb6��$ޟˀ݄�x�b����ɶp�<_a�*&}7���5K|[���%N�"�1<��譱v���gz�٧����{�FD֥�̖-�W��U��R>��jS�r�e��E��Xv_�>t��9�%��h
���cN�ڜ�}&�����6&�vG�9�`j��V��#������"u����Z���xp�!ڇ�_���~����د�-x�=�X\%�@����}�r�8^�"bRt�hX����s��a����>�s:�k�/��U&�0̢��Z3��|�Q�� ��I���[�R�f��g��#In7�@�<��ہs����V,�������"*�fG
�b���hne�G����{*��ס��|@"��T������4i���68���r4�K�ce�J��&�e}�=����s齌���8��P���� r��c��W7�O;
k����<�Hd�u����NAw G�qz@D�N�I��[�K�@�.�a�t�����X]�6��a��]���y~	���� ͧo+>��y�AƠ{�mZ�U��aq��P�2O��H�n+^h��O"���hԭg,T�Tl?�Z�]�U�A��S��dx�v�K��G��)�k�� ��d�a�Wi���g��g�δW�!; ��jt�I^��L� q�%/V��`�73�BW�Vݰ��Ē^�����p��?���|��Y���3��F�K�6$�IP5A9�Qr�E,���x��G����ǲ#��3�D������,�-`��/���#fD\pf�W��!�5��<�p���0}q���0���=�9�'�g;���|!��i4Sg-2���5�?�4� |S\W%�<�.&���$��w�i�x��miIP6=
�����i�:Q9K}��H����
�g�7GU����3�y����ڴ�ݩ�������ۓv�zBZ���E��%�z�SZH��hi����=v�iA_Ո��p�a<Gs0O�F�+�������`_�d5�}PQ��]�� �5O(��'�� ������A�M*�

.���y�N Em�9+�[!�J���z��x>�cT_��\+�6`!�o���qcٴ������*�RܔoZ�zD���}�M[u�$0�u��$ �A�i�"¢%5X��N�D���GQ�L�)8ۊ�]���6H?��0�&�M1,����v����s�X�L4Z1�M�|;'���E-3�q��z���c������u�ô3�4,�� (j�;����WV���%y���|�K�;ڌ2����ϑ����O���=����u�>�3ь�����G|_$(���e=|��tZ�3*�8ԙ����/�2�C���
]������;䠊�\�{5Iȕ'�]�2��Үj���/"bXe��A} =\��o���	�'�k�5���h���
Y`����Ԥ��:�c	c4e����:��g��
J�Yl/8o���3 b�^0�;���J��1R^�����ԙ|��I)�4�"m�K�+hp
���|�cF�$�3�-�S��J��#Vqq����iE D�[2��`��>/���*�2$ҷ����i愑U�Q��Ԯ9?�D�k/˟e/�_�CccCѸ�<����"�޺��z�ٵn�2c���w����:�a��|M̂��7D�PQ�?���m�bGP��"��=�{E	{�!Ho�O.V��W[g�K�B�I�L�^�db�{�}�^P2���D�S����x�J���"´����tG�5S�������oQ�·d�͎q��o�`O��o-�}�r��}6KHМ4ca9 2b��Q��`�Ȏ�q�	�p��8�agyf�q�p��)5.{�����>��������&�G)t�3uR���0M�G�ǎ谬ބ5�%
�S�3����2��Uy��B���C\���
�w�#4e��b�hH6������%�,$�M���u�����&|h�I�3�d�]��Q�3�Q��F���es�^s�?��&��N��w�B��O7� |��}���P�U��p4���6O�M���z{�4��Gx/e����$A��������'J��Az���Z��]y8��E��{�a}5����F�;G�#��C��܌���������faL�����7���@/A��b���x3������"�X
�K�p�B�$x)5	ǥN�3n��m� T�4������'	 ���XEh�p<F;�Ƒ�Tj��B��/��Z� '�� ����V�zG7�.�#�����ۘw�f�d�B2_宯��/c�8�m%TLV��i��%��D�j��l$�[ҧ ��j���@;�T�sgZM�6�s��̍��N$ ��*q��fe�X@8�#��%�ձO��$^eDGzX�.�.�����Vc9.H��h�L���%�%Zԉ�STO����	�Շ�@VL " �}X@�I�}+��Ɖ�6�������HAG���+�3.���Ϫ,޿�E;��(�t�Ϭ�)��՚�*dHkE��V�ثC�l�x���X8PC��9�[�Ǳ��X�Rrc�E)jl�1���)�"��`�vk]�P��#�4�����0��T	k��0� �Q&*K�K���7���m��L@�Jq�x=��(A�F�1��4�3�������&�z���"���/�}�wi��[�ۡ7��+�-��P)���Gd9o��#p���dhq�=^�H����Rb�:�,�t�2m��� ~d6��ҷc��T��\�= ���G�UNa���`-h�ˈƷՆr���bm]�ԁtW��1}>�B��t7�$(9a��w�ܒ�LO�&����@����<aX��?�-��&���l�*۵���:V�X�.�?���-k^��������}'�;RRH�N��y�L'��'C����^���B���X��/��4,��O��%Z�s�i��HF��]~/ښg҃��<	���d�8O�*�l�v��@���l��.�8m�Ѧ���?<".D�؃aKTśD&Λ|׺��2z���/+gJ�i��U�TZ@J&RF��Q�P��u�q�J߲N�ΰ�w�U�3/2��hZ#1܍�C��O<�ݓ^��i#>2Ӥzk;@S={z[�ٯ���E�-��K��X+��G2�
�m�T�a��������D�p�^" BT�8�s���9��ZX<��<����lg��3k��]���|R���\9��,����Jf��W�pJ����&�m}ӷp��I�~M��P~L�p`i������".6�'�/mj���d�E���5�X�T���1��jY�-�������?�|k�4�sx�����o�6Z��)$�X�v�4��$���J��ǈ�{��dܟ��	�JU����V8C/����^���=>譪�m>�e�3k���E��a�Ս�*���e�𿷹,���MY�d���
v ��&��w�c)t�!���嚵� �A�n�Wc;�*]5�G9�\,�h�_��827_��~]����"�H���#�3(}ىu?�n����Z���>�:\�x����}�]�1�������,�S?	m!,���{��W�4s�_ J��3�1Q�oL��d�F��.^S��K�4��;v��!�:���B���+����IV��V��|3���ʧn�d�0)�?�F���T;b��a�(¦���L��Śӱ�
����*>�`��Ě�?و��]��nR��^��a.�T����v6��T�1Sޯs�5�G�F�m�~7+?��kE�C���8��Ѹ��bS�`[݌-zz�[�,�n����h`�����CPA���s(߽>�{�=��ZY9zq3�ѻ+�%��<?�
�63d2lZ�(�_���� 7'Nؿ�'�oj+"�N� �|l6�i���!�X�-nMd��m;��ӵTF�#�ʤ,���ʸ�J��hC��z�����)ؘ���M՟�Z�O%� �W$((J��w���k"���M5GГvy��vD�7���@s:������!�[�݅�ߤ7�gTZ\�X�Vr���7��K�?d'x�Ny��>��Oa����瘍���c�>���Cm�-�{�W�H�I#����QFQ�=&���I܇�}�����4�l�k������w+�LX<N����Q�a���p�f.$���J�h�|�0�C2d�:q�t�D�2:+v��zg�a���Huԡ�s*������W�
sZ�P����V�:S!ǈ��p�Δ��W�l�WgՊ�f��QZ�8�B��W�����i�i��q�~*�����R[2�_���c���Ov`�1�0ڬE�E��lX��rt��uTQ|���nG���|����lO�`{;��|�C�>�,�@�N��Xg6�����p1
�G�s4c������bd����GlN�������r���垠] �|ۭz��������y;��kh�>l{�+䫇E�b���9z���7x�:0´�~�?�t��.ʹ缛�y4\���g�\�2���w��%k_��6����,��K�A^%'�(��i}Ǩ-ͺ'TDY����ғ�tـŤ7aLbmnk��͏�Pj^�h�?^m��t8���M"$�2<�@�G�RFD� ��r�D��΃�������z�I��B�Sh�:ּf�iN���vH2�c���Y�3?�"�*��M����
o��z�J���_� �Q
��0|c
&�����.�8�����8��
��kiǆ���䴐j�'\���� �+&Q�I��������4����ĭ|0į���& �aX��
�Ā`�g�9�u��hm��U�:�=��奡�g鰌��V�&�
C���{�v
��8Q��o�@���,E��ǿq
�ק��z&��p�e�ڑ����(�v�l�]��;�{�)���wk�M>��#GL~Zv����rc]�*3�yt�E=#�K�@Vs��(ۣ�� �'���<�b�u:P�it��aٺĂT��BAa�y�}I����/�L�D �������Y���ΰ���@��ĸۨ$ˇz�Sц�z��<�qV��I��Q�%��^(�V\,��ֵ^��*+��.rU��%���U(@��UT!�d,iѬ�P%�K::��F��������t|$t9��쥟��R����?ʌ��2��G�mS,�i���ay��w/�C�k*-�j5�h A�g�!�r��!p9��S��,��B�#B킂Hڽ�L7�<�*�5�B�\�Mר7N����fo+v)M��&�Lħas�*F���nE���%ګ7�'FN�h���F�.��_\W��f�>�ᒖ\Q��mi���G_��Ng��a��ַ͙=�-HBW�P����]���6G�
��(����7{�yK+�v|$�/�]�*W-#����@�8=גD�<�܏kս5��� y��oS���&��н�X|ZT�f�7�{mL]�[0��*�gW����8`�4����9��zS���{<?�;��#K l+����7'��CWԷ�e3�O�~��e4����M�ɜ�����o	�b|�uЄ�I�U���ɏ���#z����K�~B�-�_�i`a%�u0b���b�/�6��#|�Y�b�h1wT�N�R�d��u����2��l��0W�0j�����3 �����%�+�'K :�"��LܘG||,�U�%��NLMw�	N�srp���p��L����3�ٍ�(������q��s�w�)~���V���˱O'Ғä3Q7���t7׋���qr�w��1�r���������������5`���Ȥ��k��Q�NM+��+���ɬ��-_Z&�컘P��x��<a��(l�j�������l÷4=��lJȑw��g��k�	p�f,D�ϰ�%sΎ�����w�>��B�]ϼo�Eļ[�N�1�*��'u�9�M[<��6��~<�x]���F[8f��v��K�f��"�c��é�q����۟N�еLߜ1\&���G���g��ʚ�u�s�F�b ����@�����s˖�z���Ӱ�u	��� �����Q;4���=#�]f���
���OI����9�V �_�����ʏ�м-F����� ����v�x�� ?����4�l��=��6�1��4&��(q�l���(��v+lѫLU:&�����<R6i����H�'c��z��4c7�2�/�|�^���B��7x��_����j�:(�Ga���3���X�Uy^&��E����PQr+������{�=��Ü���orN���O�[�K_9��}~C�(�1�rw��hzk >g�*�n�'+��@�K�@e�*�'����Q�H]���V���HN�\��w��D�0xі)#��+po�96}�g0��m�]q���.�'X���1Q��p.�W���s��m/$E���3��`���c��O���5�6�M��LJ�����1���-�č,�]���8u�ꗔ������x0���c�͔�6�����v� w��&/\1�(&�Zy�`�KC}�?W��_�C��X�܁|�~��Pn��|��IU��4R�%�%�����$L��H�6>NO5*ĳ8ĤFa�(�T�q|�}�}��ccJQ��=h�����s/�]��R�i�������3xOX����#6c�=�V����TU)�/���@����+��$�fI�bZm����zl-۪��[4+6�K���X��N%���J��P���Ӻcy~��[��Ѧͬie=�=�"���$P��;l�5��s�~��V�8��?��+�z,��(&%z|EZڝ$��w8#���h�J��f|<�|����)�9�����Yxƴ\����#��x�������5P��A+�&9]F������@[;R��+C�A���	��S�`Rt:z�M�߿/��W8X��NVG�OGM��h��w�����T�n�Cl�YSq>�w�+;���?o�a�]�gzֆpۧ�����Z9���x�q���r�Y@��v��[�q��ϧY���] ��@���R�*
����I�Sn����F���N������#��J�=��z�&բe��6
��8 �I
��ۘ���0,�^ �f���t4#��?8Oll͑P&��^��䈞��DL��;���#�.��'�]q�$K�j�h�,ubM6n�*O�ɢ!~�A?ZL?b�_�D�d���M�������Y�)�h-9��v��I�C�{���t藺�뱁:O�Y,ꝡz�כ:�i$ԫ���a������_e�{e�l���m�3&�j�P�{T�E,`���5��3�G#R
�=Cͅ\���嵂�#�R`V2�)t�~�v�k��ޥ�x?�o��:�+BIS_�P'�Te����\z_`�V��^�Ђ'�L�O5��z-X�:>g�c
�R��tw�-��m��h�f��|d�+L1����T��fp��W<�w��^2tM<;V��5iW��		�6!(�R�_0HP++���*k`&��r5��c�J�
���L-e���KMݑK��;�5[��X����e�}L�SmX��%t�~Wf�6�w}���tUR_��L�*ҳ<��5�8s<��sޭ��a�Rj�����g��>Z~�N��:w�b�0�Ȕ��=Sf{Y?Y�2C��������_���IrG��H�:���>a��&~�)�ߌ ��"��	2Z��=!Z�XK�.o!��&�����Q�iZ�K��d��ڧ��P��z�t�����ז�k `U�4F��|D!_��˅�T�������u���t(zo�V+��J'�Q~��k���wm�Rg���إx���\�r�#��8LQ���1�(���9��˗Sӱ���<�x��\�?&��Gɵ՘,;�d8Vn����捅F��q������K0oM0���V�'1�f#5�R�C�(B��ƯҖ�o��)/T'5c�oO�o�`|.�ر	��S}n���*� Uy-J_5���uN�FV4B��S:��k�ϰW�݈�Ɂ�����H^��	!.-7���ju��I���S��Y�;w�0�t���Y.�v��d��b:zX&��c(0y@µL��4�B'.�"ΰ���;V���r$y�.��.�V
�,��'痫�c!�ոZN�Na��"� l~̖����ER�B�ވ�|�e�ϣG��(����3O=GXA+ڕ�O����WY���"�@��`��Mɮ>��l�
�9�0;l��������q)���H�3��:�SW�9� :D[$�����E�o�_v�	���9����o�����_	[����M��½%�`U} �ZrB��b��Fi��S���߲�I��'�o��~����ސI�so��N=�"ό��:	
u"Z빏� �i���f��R�섅3G��7EgS�:D�R㤸���H?ٰ�<��1Lץ�%Ζ�8��qᚊ�`�7*��yy��@.���?���X��!��!�ϳE�����!^�(>(P?ɅTOL��չ�ĸ�l��n�e���`��>���H�Yˌ���E|2�"�^L��[��	<��A�1�$Rg���Fz�)��='�a�S��#���O�)�y���ߝ6`?I��jb3-�{ä��pY��� z�y����1�K(.��v#��A�65�672�@۟2Vݡ���{��r	�X�m3���uyI��wʕV��z[T�q[��g@4L�^w�۽�s-/����-e�|���~�߾��g:�,N�s���W��m����ӏ�>C6?�w����k�\��0���Δt��r��LG�F�z�S��A���>f��Yc��`6L��|������?@Q|W��i�/��j��K)�W~���k7���L���eQ�.[�6wܞ������>k~&f���$4`u�pJ�ʄ�D]��2��G.���Q��Y;���=�"�J@�T���C�����7�2�gB&'c�%H�sxM�a?�wO�U��U5�X�uY��&�bߴ�ݗpXrƴas2��ku�N�rJ�i2:�x��n{�x(�-�d�f��66��*V���u���z�XI&~�t%��%:E9GY�c7"�|�f*FJ�x��ǯ�]5��Z5�.:�<qC����#�'l�����r���1f�E��]P�$��S@�O�$��6ǦW��� ����T�ҷˍ����³�x ֣�)�`!I�|�Y��]�ͨIz5���Q�<���AČ���t�{_Hz[SQ�M�~�̳܅dgg�fh�q��Ĩc	���D�ǡjN�&9�oJ���B�%V��L�+��GT�\��pWs$C+6�	Hb6�0T�����D�P�Vn'쑨P��Gv���3"K�<���] D�x�������gU	�.{�9_<d� �̳Ǥ�v=`a��uPl��:�W�D�*��3��a�q���"�Wfns��%�Jd���C�ǒ�W�_�%��~�@��l��̂��Qv?�K~0�͏��C�����l2R�&mT�wh����|I�Y�5��	b�4Ʌ��P�5��
V�1=w���aR��m�z7�&���6����ףe��y�/� 1��K��^��1y,_���1L8�����YYl�$�b�qiӕ�Y}l���Ǎ<�sO^a�M�~��32[���(c�0|�Ӏ�=ڞuǧ1!j8��4�X'uT�jN�M��գ�Hq�z�E�l����JM*\�v�p�:��j�>����6ƼK��i"#M��2���z,�4>��V;k��E���@�����_�x�t�Mn5ϱK� h�Ë�~�{T��D)rPH_�L�O£r)�iV\���e���i�X?gea�����b듑e �A�+xY�m$�;�M�\v\�@��F�g$������~�x�T`I�(/��:�w�d��o�[��R��U�n쫃	�%����7V��'n����
�~�U}�k�I</�hYZ97���'7
��n��R�_�v5���sĆ.�3����m��5����O⽳�b����F}i�eՂS�K�_�*��q�x��>A��~EȦ��u��熎0��Č&��L�ґ�go�ʕ�f��4�=A�@���[�+H��k��L<-�6���9��'n�mgB��׋ �ݱ�y�\x���9�I������O�M,�eg�(�;�WP|,�����@en�{���<��̋�x�X��Tl�g[�l��E��sX��S��Pv��^t\�A�n�m鎏*]J`�)�$����vI
%�Z��4�R���H��%����8NlJ7��c�iXԁ9�u����7�ԁqo�hU-]Z�7��bj�F葿�F���HߎFɩ��P���S��~;2SIw>��B�ʮ/��w,M�r��@��W�`�x��������CTjB��F/�Ee;
��y�QW��0�8p���`���RQC��D�?A؏���1]U��<�Y�,
Q\eȼ�|Wdv,��'ƛ�yP��H��8T�3|���pB�_�Ud�1���ӟB���ېs1�y��,�iWtʚO��tך1cP����h3��qgx�������Q����M�'s��&rȨ�K}b���<oA\���j86{	�ũǹ���s$e�]!_'���P�6���i�k��#Y'�L�W�I�y�¢'�٘y�U*�L���yT��h��Ĭ��T��8Y�BT����B�� g���u�ϝKʩ{������k�l��2^	�-��ڔo�U�>�̶��s�U�G��(���:^�I�2�
cb��)�y6��<]ٶ*��ރ\5N��a+�O��$��#��y�ݹ��6�| ��E?�Hۤʝ�]����PU'PԹ{��c��Շ�ћ�.w�ߗ���Q������zIZ�%��:�c��Ѷ=���Y�9Q%�?���v�nmw����\:�a�
��<�]��ki�r]��V�p�p������A�t�S�v3�f���KdAl�7f6&�93����$_�jE�:w5�w�9*
i�����
��&�i�5>g��P���7O��T����[�>��$��*? �ǆ�9�V��cl�H�e[d��`f������Rv���Q�)8���{������`�\�H�%X�)���1d���>w-�/zZ��P��'æ��r�cT�BH����#�CY|�� !�.��\��<��6��$W�V�z��,��B�U��P ���A������Ɖ��ͷ�c��.*�4��q���]wh*��Ek`����X� �e&}�G���)^>0�t}WB0JD�����/�_%x�)�+�%���d��T���?Yy`�7E�\�LA���A��,�������vↇ�G�����K��'�c���N0˟��]�N�%�<�$��X�Y���� KK�j��*��#|�a#����D�$�`��&p�ǎ�En7F:5�)��*�sT�}q���p�����T�TQ���6��X�/wfZ�b��p z���D�6�&:%��^�G'�D;W���-f�(0����y �[��vhL�����ŵ�� 8�2�78�� ���+�xx�o���u����;R������H��U$gLb}º�j㴽���y��P�=V'5����lS*+Ce!�5zۛ���������Գɫvt��$��0�_bNK�O��=ƥ���L���j'����bM4���
�(�9�\����o�CS���V�*�ղ��n���cڅN3_�-��ֲU Nd`��m��.�]��^"���1Zca��⛆!����J�A
�����M�o0(^.>��;_X-N$A�Q ?�*���M��Kɼ�:��������B�"�{�����2��a�����y��~�:-smJ4!��dD�x�Nܬ���ձ�zZ��b�)z�u�~������y2L������w+zp~�z6 %_�;H.u~Y���Ees۽2ž��0��������U?�,���!2&-���7�;g���Sg�$W�.�D"H1Cqp���4���v�$!�f�xs����P�%�	AY���}�b(�����U̿ �6���:,��_VE��TJ���o��E�J.a��M�UmC!}elP�,M����jb���e;�-:��5�WXK����� 'W�@�����t��ϲ��8�8�"����%_v'<@m�Tx�y:r�"����o����?������&�?�)�WM��
��}�)O#'90Z��x�`�	4n�H�f���0b3�z�r׉���x����'�mI���N8���S,���Y[�%�����T%Ӈ埸�`^�Z�ڨ;��P��B���j�3{��./���k��[l S�����`5�f�������˃Y�ǆ�K�b�H@�P}�z��ck�&�Gf"3� c��U9�Z��}+îI�%ҹ+<(@H'���)�Ƣ_������SDt�P�Ѕ"��t������8�$`�"Y#�o��i;���w�(�;8�oٚE2����TY[��[d:�2�&��Z�%������#cqx{B�D2�v�K*'��ҥ�ˊ�T[U�c[���z�,p�b|��ϡ7�	]���lr���1i�:$�F��������W0�h�'}q(���E�s�T�0,�Ӛ�5{N�3Z#�P��[jLDvB���s�h�`O_z���G'$G��B�%G�J��j��;��G���yv�vbd���k�[�2�HA���Q| r@�f=�W㏕��(�P+�����cI8K���G��9�z����������� �?�itH��"�#�!����@ӆ3���0�ܽ�����7�&tn8�{�K�GCv�n��13�ͯBU1��-{��-�L[eg^�d�<<����� ��D4�'$O��3z�Q^V�]|s}3y8�l�e���J�.�l'�f��Jg�U��e�Y6'`ّ�s�'8hAl6��,6��G���� �W�_����2J;��,\�\�搹�*�K�O��7�\�&rTY�x���	 �w[z݀��&!g��狞�\� է_b�I){���ʠ>�EL�<ܘRA���y�!�Y"C>-�����p.#�Ք��������J�����~z"�����3t�	R�<�O�������d9ە��F���TR�?�,s	�Ŀ:"�<���O���2�s=�2KY���Z���t��}�O��k<U%9�Q@��\O�1����CȈ�^i�]"g�`c���ֈ���<��|G�bZ��x!�!T��o��K�*�&����E+ɑ�ᙸW�ɞa�r�:�g��{�a\�E��,A����T���Ag���'��v�
���/�T$8=_��|F��jfZ���CThJ�9x�0�/���፳@�-5떲0�73����?��7�mr��70����,(β�ʿ+�)��$9>�� ��t	�=��U`�|o�3���Oذ��@{/��妸���p��O-[��3UD���h.��V��R�Qd�ݦ(��s&G�M8�)ד83�}�h��-�����"�e�ρJ=���HQ@6��w�$+�]���u�`�����>�x����șw�Ko��+��/�z�Avu�^�X�xOVFN+�nqC�k�N<B1[��zq�9nɴ%z��x_�cnjy7�k��Q[��뵔ٷ���IS�WR%9��kސ�d�i�&p�`���ay�z"#�^_�r`�`�Xq�v;�Nݬ�s#��.��2ן�����y!���[��"��/ AR)$��[=�|��.����q�@ *��=�|GPk�Ť�b|P�%z�=v��Z$0nD��f�}��7i__���gP7Im\���z�-k��wl��/%p��Ȟ4�$"�f���G�O��� a8���-��t��
�	�-,:r2��X��t1OΎ ��B�Q�S雏�T8�ڇ$�cK�#v۔b�g={)^=qn��=��8!����-K=.�>VU��k�U��
���Q).�Y��'��/%�潣�M � s`���M���yۅ�����V����"ǋ-U�և <>�y5����ȑ�J�A1�&���Bj=�\k���`���ƞ�A\;��E�8��9����_8�d��ʑ��Zc�2����J)eH���U$��i�B���rj���sE� ����XL�2���7*�:r}X��D�I^&̯d�BXM�j_c�z���ߎ:�E1��\�s� 4�G�6E��N�6Ǯ���l?3`^B�k��-�M�>b�����3��r(C�$}�mo�>��I8��1M�M�^�Qַ}|���k�H�H[a�|'~���Zn����M롑��C�-3�I��D��|i\m��q������!����ۍ���"1F#�䌗���+w�$Y6�P�Պ�S��4(%|����a+�Ě�z���^Ua�[	M����Q=R�簔P�ܦL�t;�^O�c���>�a힯MbU�g� �9֜?cj��K��#�9aP� ���3ە#�	� ��(TI�2>c�0�lND��:X��FF�y]� ĕ����� Dc_�Oi�ζV�/����(/R#:h�=>
�e��r�[�������@�{%%�&�p )g2��6�`����^��Y�E�p%̒�L1 �\wGZ�7α��� � ��k���-r��<�P�'nUA�W(�%J�kz���m�PR��<*�2��V'�ś��>8ĕC��}��"��t��#�����j�x��P��TU�ŎaW�_C���F�n?�i�J�>�劙�|��P(z��k�:���/q;���i��+� ѳ�'�H�	eT��Qs�M���l�9=����0d�
iU:{c�\F��ܐ��h�"O�Z�@������fe����D.Ԗx�i���ݐ�m�,�q;�IB1G��"y���%{��k��v���2�_��bkr��J��� �Y� ���e-�|����
Z׀H�šq�qp�X�B���a����=��HE��?t�)> ��Հ��]'H�Σ6�kP��#����?�q�z5�� pHP�,LA�:Z�o�`�ZM��&��:��#z��c���j7tU/dV<��
ψ�/�`�c�0�	 Y�Z�}���W� �šb�@>ơ�g"�)aq�����H=σ\��+�`?W�9-���D��h5#�W���a�*��gt�G\���U���E����$���������{,��<�GH�#V��n����H��&`�EѐQ^E�T����;��>���}�`��-�en�:��G��=�}g��c��D���M����:�~�y�j}��b���	E���[��t����p'\!aɡ'�ww����:l�!ʈ_����"%U<㷒�:�%r,{V�d�Ώ���l]cu��`���r�H�5f�T=ZM8P�3x�{ �z0�zk��?B�><@�L�p'������r�A>����3ލ��6�����Jt�j�hc���t��ͣ�X畆$t2�l����M
t�P
�8�0�S�A8�tH�2�#lT(�{�p؋A���zC/���$5g�+�w�ɜ^�W7 �Hb!������D�%��4�(����zb �
�G�&=o�̓=��ZV��6����MG=��߉5����_�O�6t9�1��r�y��6�X��*�DN��'Ow��h&M��j�,yC02-���SNǈ'_v�6KGYAS�;�=?���	*�1_us�-^~��Bg��U�L3�狨�8μZ�c����ܬ�q���v���+j�4�\�U
TD�YT�D%�Z��:D`u) ?��03�h�Ļ�<���6��Q���s!x���2�0t�f����_�f�@�a4����n�<�|M	*�n4ˎݓT�6Ǫ`���
m��)Ǳ�3��}W��o�]��#89���}{��ǸߗA����+j�I:�f��C�_]����Wﱪ���Ӡ ' e�1� M�'��<6[�ɯm��t8ڌ���!(�lK	�Z��+�$�5���M���pŭ)������]���G���L�S�L�����gʘc��F=�f��	~�D ��o�Ov���9�m�� ͸.\�aH�r��L�7��2ǂ<��4���#0-\tү���X�6ݍ�Ppx�R�AZ�v�_��j����˷#E�+�W>�όΰ_��G��YG��h�Zl5f� ����`����N�A9ܝ@����Y�v!�ļ�:K��'%))�q��+20
z�����^`bIߘ>v\�p`I�H,�¬�뉙�dR���=���3�^aI~ԲX[!NA�Q����p3�R��T+��:e��ҩdc�\�0���9GZ�Gl����@q�=�a��\r���y�0���vZ!c9���g58�a�F� o{o�%�ل��<�}aR�Z�ow�?��?���qU��?e�4��d���	�v,�����oxi���W��;)'Hc��}K���`Ee�3/��M����F�:�8�jC�j�~���#����ɢ�5d���tk3��E:N��]&#���H�<�}����=���L�Nq�;�9?PJ,VqF�v�Dkݢ�S��3u
5��ڪ)H�����-?K��0��T���}V��u5Y.a��3n\T0�n����{o��Ɖ�/�B͌�bBYU'qiĲ�/-����{����e��!6:Ux\�A�r����#T1�IN$��<*>���Ύ���5�vĚ����d�o�^K#�����?�#�d�I�3�� ��5��J���u��; �(�1d��~��^���T�F�-^g�􈋣�A��v��þSE1Y�*5D�d0;D��9��RHX?�����&X�bٲ�V[��6#W<tj���Ӫkp��W4���Į��l���o��u�y�[�<[mb��B퉛gw������!�ە��CQ�/���Q�3��@�ۤQ��G(' )�@�q�`��%TR�??���{����}�\�����l�� ������Q�3�^M���11�]�?����y�q���,���^���d�D��:���1�*9w�m��e%]��b֤��;&[���=��6e9�{Y�m9���9F�M�9�^�<�~l<��_=�lb'�DimK� �JX�Y5]�)�m�o�m�ay"M�xذ_�D��ͥ�$�K�jE6޸��8[.���0�$B��S�"����{��?l7�v}�鯣'��fT��	�XFnX:��g&:���&�"��fwyv!�u�=+��C���,�*^,�TY�n�˥(�[+hN��f�X�,���ikc�K��BЙ��*�@�����#�}�m��A̮��2��/���8)"f��8�p��@M�7T�#�V��{S�XeT�/}��"	ր �������"�$D}a=B�:I\�b?�C����c��;����c�Wq�<~�v�C�0�O���M���&ߠ 9�l G���泵M`PMkN� )N��7Tt��d�0fT�1xM \���6�
�`0��u�(I��������	�>�H��~���78�e#Ir��Ւ�B��K���G#�܋�:T/��e��͠ﲠJ�p]�:Fqx�@_��'��l�����uʋ�T���8E�i�KVJ���[�9�ݏ��͢
�j�V�Q��Ɋ��|��ڮ�ӡ�%��
�G:��F�����r��lt%�M��|#{*N��<�-[��=��{��&�a�i�b*�F���<֦�%c���A=mR�&/҇�P�;s�;��ֲE�߳$��� �	�2�s��V��ڇo҄��{�*�ʱ�vA�o��C��v4$u��XX���|�"2�ƟW/��V�M�#�)��.I��������:�Hd?�dv�
����ݥ�V$X���q\r_z��O�O�n0�v}w��2{�����.y�Jy�j�m�K��!�j$��޻�'W��2�ۙ{��J�S�B�4�����3��!TYc -�N��=�C��ql����#`��!nw3�� �&H �pޮX�3\-k����3h���-��@��>��u�㽸�٪_!�)�ׯ
�~4g��sNLC���[�3g��i6|t��u��up��b�Q�f1`��@�X3Pi�"����'᠓a�B��[,�:L�uipB�;UP�{P]�]M�J`�8��*�*,ٿj@<��X�G��ߓ��>�m�㌇��|��5����N��� ��l�S� ��^�d��;7�"m��0��L��f�H�;s�	�K8M�M����Ð�d���g�,�}m��T�D�g�.�v�-(���)a�=��\ɗH0���CQ���`��^.T��Bc}��/.��3� �z�#ձ*�l\�d���P2�k�0����Aq.)f�̚�r�x,�uJ~o��/Z'-�ݫL��ݭ�zs��W�O�	<,���}He��WO�6� gE��v�	��[d�M#�:80]��1���G�Q*gV�5�q8N��d0�*
�<�w�ZX]���Ǒ� tH�HB$Ry4�N+�
3:��GpF��-@o�l��@ �7���!Z���6���h`'�{y���/o���s���{Ō����;�<��Y|ʐ��Щ<����n���(8��*��G��A�N��fL0w-"��ͺ�e��i��SK�|�