��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O �ٝ�l�������V��fE��v�-�Q��Rj&	ڭE�����<��1`5��o"�l�&��3J���m\�tu*&W�N[��H��j	�����[6ҊZq]ս"�!z���z��r5����nk�/�v����~��8r��,��:ƛ���M-$��e�~4=#�g�L�C�� \3˂��M�~���Wξ���G��Iǎ�S��IhU�_J]��;'M�J�ӕk�g��b��v��ҵ푣�~���/O�ׅ���08n2�B�
|Rh�ώX�T`;<�/y��m�=q;a�߸h�{���ð�t���f��
*tLb?�S
n�Uj�
�J ~���lAoT?�!d$��1�-;�59�C@YO*��x6S�����0��*�?��'d�>�fCŝ�ug��ENm�HKj���i�@�����&�F�kZ�8���E���b,>�#z��Ƭu?�_ͥ-�BH�k>�K
 ���AS���+�����>�E�c��?$�*rJ>&+a�#PS\�-����r�٭|�!��S����7�9���[|)���
�;>(i�>����Z;C��>��T���:1x��L;Utu�S׫E���.�ޒ12�Ꮠ���Z��|�*Wټ �iVr�+��<wzl����d:�:w�"����:Z
�Μ���IU���~�w�HJ��P����#�>����2��Ms��_�'����~J<!�
?V�9�o���bM��0��� �E��S��k�[�s�L�O��WX��-3B��O�
+ʮj��"O��P~���Q�_����~�����ؽ��̍ϲ�=��e��I�n1Rn�YDy|�/�\��v]A�>����M���z�v�s+�a/G��TB�w4xnРCҪd�����iV�sB�郡�1Z��������0~��,K��|(�{�| B��\
)����b`�j>j�O�
��6����|z5&~萤�h�����Gq�/�!�`�'仁"0�q3�X L ��+ ��_�-I�<��ܯ����F.G��C<NdĨoÝ��F*�T����PE��<r�5��^��E�Jd?@	I���/HRd�X� 7��z�t���M����d�
Ƴ�%���[v2�5Zrc��a��b& �J@w�&�ٓ���ٷ'��·�mxQ���9�m+��Em�J���H���c�eYQF�ֆ��1�%�q�Mǡ�uJ��`jM�ש�|��=*�Ƒ~���-Vr���_�b�������]��!$<YrZ�KX�Xa�̾��"���;�ۋ ]�q�zR�nS�i���	h�R�X~��ϷrayE}^Y���L&�ݲk�#��$pa56�C]��\J6����f~}��|�h����J�<�t������@ô1Ջ�M��|�6�V���~Y�y�!�`l��UoB~�P�&w��#ߡ�Z�°�RC`G�nj�Lw��\��5yE"�Ť�"[�~��s�d_l��G�y��ۆ���u�b�Z����8��=а��5l������j~�Hzx�VB�Nضo#n�`�ff���iӱP!��J���Ӡ��~�f�r�@`p�F/���]q@7m6We�k*�᜺�o+�Ɓ/ar�v��Z6�#��_S�3�P�1H
��I3!��_Ne|�����
u� M�357�����!^#t����V
�#��t �^o)�Hr�#�?3�rzY��=���>v�ŭb����镂s�Xۢ��F��xOٲ��Cy��>S���Ɠ)U�P咸S��n��k�𓡀2�]�����rrP�JG�bp�gw���1���Hlx��1V��, ���9� {�����ĹI��q|���k.7�����^���ZD�4�-�@a+of� ^�����-[�a�l�K���T�?�T����
��,�qp6��E ���-X��$+�eo-�J�.��s	�uvb��Yi����Տ��&�:iŵ1�1����Fd��ŷ����B�.���:�7w�v�}:U�v6-��l����hFk~߮c�/U%����dͿ�w� *�Y'��:Y`!4���d0��R�CIg��QGe�}�h�e�-8�U���)��#�'��l�u��S� �Pt�"}��({
����^���W�Uo���w%N$�>�F>Ԉ/ɚ��'�&�|�1F�p˲@~�)���)�c%$���ꍳc�/�߭r[lڭ���f*�f(j�\�a,�z-P�V�a9�1�B����0�{���s.��+i��Z"c-\-�Z`$�U9!��a�0=okP1����x3I�_����Aoރ�L��UaE	t^274�א	�1,dz��gh-����,��Ao'�50e\�F$��\B����eb��<i��#�#^�e�af�]���6$h�>$G�;�r���l�V����.�u�7�Z�I_��mqe�3��7��ۯ�ᙼu��z#��ݦ����ȃ��\r�8Ѯ����0g�4�g�5I��L鐓����i#ZN�`��ř�O潙��FD�|���j��D��r����--�%��@�s�vŨ2�I���.`��W�ً��`/��+�����&6���/`�m2���YW�w�M��vb��~R�N����@�Ϫ����@}���iM�d��1�(�ǋ�jV�{��eY�t<.0K�Rg��M��1�T�?ڑ�7����B%��L�{SQ\�K��BB�S�}F���Bv�q���"/ϛ��Gҋo�W�9p`���[����J�F�<|S�.Kjs"���Q�PGR���r�]�*�j u�N�T����#�v�E\"�@���1p��q�*ޭ�o8�[��ËfT���5�$�v��&�J��C�tۭL��L�|+V��ZB��m�pڂ���x��
��x^=�����[�SD�> �HmZDz��Οr�c�Mͷ0�襲Ok�Mڠ�e�G�v�V���	|#�r�G�F�P5��Ƀm�b������J� ^g��
�,���|U�잡�x"5�+��3f���X�I��78g��U!���X����ķg cG���y��^�z� ���(�ڬ�'=IB��D-��_2N��z?]zX=����4�\Z%�u�� #��/�c'u
 �v�vD�F����k���&�C :G�����:��.�a�)�0���_����#�a���zXf�]j��-,����@��9)��v���͸�F�G0�Ͻ���_�հ����"�+L��, R�\T�����1 �C�h�A8X�����`:��@��"\�����g�p1v]�(���G�U�%f�.v)��O�c�P��x��R��)�uOu�g�����
Y*�^k��r1,v�Z�0�!���2{f(dR^����F�b;��S�N%���'�b2&���=|�f"H��BL����[#3|Y�ɐQ��Hǣ��s��@?�|k��uil��t)	R����om��1 ����=�GD�"��O�@��W� ��R�K��}(�M�J��A�&jT�6˽3�ȓ�w/�ͦcO �&�]��vrr����Є��C��ǆ�L��s�����(p���p���V;4����"�QI���WCe�^�,JΌ��h]n_e�o�q��o����d[
��r=v߶�=d�~ҩ��XVE��>,�Ja�7<32�;�y!�$;��M����J���rY��|n.��,ܪ��q{���;+��n��`4��x��4ĥ�
c�='�o�5 c�uN&L�������8��H���r�6I\��T6���l��W�"�E��z_`$��A��}�[=�X�f��薮��ҏ�&�8�	y2�p3u�a���y�BV������R���:/�Ȯ�\�tC]A�=���\�nAD�!����	�,��k��3��P�J�x�Om3�0����V�����Sk$d7���S�%tNv]�aA31�)����ԑn��I�>����#�E�E�lD�p|$�-�}�8 �6A<�4 �L-�q�\����_x��5��6!埪L�_��F��1����d��Sжx�q���0,���h*��>�`�1rp�.q�T��~��c�)��+��m�$~-�2�B����I:�n�0�0Ð�8�H���Ay�ǹ�)����Sq|��z̷@�:)�%��,�z[3�
O�#W��5B�#Z�өr��?�[���1�b�d�;+@�A���P��&��-�1�!�f�Yx��
�$��-�xYv�a*�wѨ�N��*�t�>�d�_��j�|��2�~/T�t=�����`MQr�ҕ��WkE��%�6���Ʃ��I��0�&���J����||,��O�a��*-#�±R^V�8�{�vݡ��A�beѪ �������W�הJ������U�r#�1�Gx�>|U,��h3ș�����h����?����P~���h��ҨR�Ta=�C=D�QJ��b�E;���AI�]��`I3�z_t�V��];�i�!���+z�ˏ:�ǌP��1hc�P �' <������i4G�sHs�3�#��:Ll��n]���0� 9<]Ԧ{{<E�S�|�(N�����:���Y�^��w��m�`��l�T�b/�{D�#	R]�Z�&Y"Hx��8o�
s�x3��q�z��C1G@O/5Rn�	t±W�G��]���押�-�b2���ɩ�`�fJ�|�ܩX;Rr�@�j?��ҼWY�4N#�
f\�F��:�=y���lv��/s�E?k��-��q "}�̅Ԗj�Sb<Q����NE"�߯��E��{	�;P���Q �� ���Ի�F�W�xÌ`=�qֿ�]��/S�!$]p5��*���"���8�J��VT�<O7Ob���s���/� E\�l��LK��9�)�$)4��U@���%�K�(���#�+��f���mg}�v9�����<=~d/�4ϱZ�����1�.�i���~e�q�̽8g(r�����!y�n��Z=�&�?uz����C.�}�"@�%�~o�J����(#�.܀�F�+�R��&�{�h��M� H%S��f'̽���I�p���L�\_��"`t���GG|3C9
 ��MB� �<5�C~��Am=�޳��3[=�ή.9Ɗ�8�YC��{�WH�2D���F�C�����"��G ����ma������}�L����ȯ��&ۧl��Xb�fz<S����k�Ud��Ү�{�K�f�����F�]�W8�~xF#O�'���TV�k��Bѻ�O0��w[���}D�͐f�7�ڻm��Sr�%5��v�k�A�%I�Q�JSC5��Ti�8=�W]���٪����C�K0�ѳ��KW�r������R_�L+�!K�0��.{x��-��Y�lpC��mE^w�x�N}��p1O���*;�:�O�x+X1x�3B͡Ճy���f��sQO��!.�%HU?e����N#r�V��c����X{!fz+6gz���ȰB���.�E���A�42/	�sk�����z�K�f^+��3q&��!W�'ѓ%n���p"�KDB_��j�7%tC���M��߻��"2����K=�L6a��6�0����Y�a�<�b����{�_ eڃe��L��fxU��_
#�3ދ5�G��?ީ�p��r� �q�!餭R��y�:nf���^�ym==:�YP��3�dk2iL0,�F��fݐ���(qe�؅o,P8�j����n�8��YF{�J3��\i;B��
V�S\�!\G,�P����%�ϩEBa�(����l������ПE�ǴC��c(;�57#�����}+9".eR�"ݬU5������_k�������<��;��[��J)��|t��B�og�}��o)N�{�w�1�S�.*�%s���b�#.�Mr���َ�mU�ZvXĝ+��Q/�@5pd��B)��*�٪s��.���0c��[k��pWa��XM���+�9��껝��*jo�@��j��1�nE߷�aF�n2� �L��i�f��� ߟ�c2ͧ�tvi{��?'k�/��?����r~�J"� ����u�����D:�`��j�+� Vk��P���m�^}�M^H:%�К���U8ED�`��¿��]�p��PȒ�74,�/r�;�3�>�:'�?�T\��3���ifQ�o8)d�������e\�Mm2��S%ّl A��*H����z�(/�y���k�S��?�um�(jRv`s�!Z�u����Z=��q��J};<�!�e+��1��hqg�\��T���^�&hE�s��W�ve�m|���hg!��@�F��I��q�W3�C�|�y�R��*;�ɹ�N��7�@�Xӵ�kN;��k	���7�7Ī|�"�?�k�Շ*��7�3��O;�p�D�!�=�5���DWr����pS^Չb��[[tV����-|��Wx	�0��➭Y�J�ZJŜ��ϹowE%��x��!������ACʊuLfS�r ��z{���?ԧUw1�@�4�7��>�M��<5��W]�y�L���D0�.f�t������r�bׅB�x��Z�n#�aXJQPny�s��)�t��j��^[	� %�$ 9j?��q�>9*�c$�ß}���X���2���u��z��ʺ�k!M,���(nPn9�	��ʣ@e#:�<N��z�j��}�b�%����χ͈rL�$��T+�{����b)���u�Rwa��0�	.L{"�@լ�m��8����ZrU���$�u��>��ճx�Cʄ�{!5�@a��߿p�Z�·�	8��Z��D��e$փ���7�P14�$��jܸ�)ۙ���}-#�E)��L1�����z,Q�	��0����~���h�����q��}:;Ȍ�:���7'�9����n�&󬓮��c:�N�����7�ֿ���$Ko�V#~�_�!^�O��@-(6x�:����j�0�� �C4�׳�r�]�@�d�<��mUǵ����b�W��`��:xdԮkn���(e%rN��6I�4�(�L�o4����C�PU��n;̘�t�bf>���Z�P"�w2ۼ�yX��  c0�͢���:�^�?��n�`N��[��ꬡ�X�E���A_I�l�5l}��,���cC���N��SL��?���<�����74^��B�9�\'#��E��)�VV=��2��-f
��s��"f ���*�n=XH$���������_�B�O,-q�