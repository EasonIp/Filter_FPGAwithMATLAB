��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$�ʫK�/�N�N�9**�����m<�&��uۣ���D�W�{ݑ`x�[Ǽ�:� to��b�M�eHޅ�u��ݳ���J$�w6L��O䳗�Gr0'�4�_l\����f�!IZ��q${������(OU�a<Tg�j������1K\6O��'o���z_e��6��q�ox�ʗrd�J3N�MQ��l�f���<�<v����-\cW��v.�?�sa�sV���q#��0J���t�.��Ѝ�&�奉2������7��oek���K\Ռ��`�����I�[���/
Kbe8;�n��`)���]�ʄ^���<�U�dL��J$�	��XN-	E�vh����suiP������*o8l�\����ϧ�
�X�N)�@�)�R(&b֍��>��E,��`���p����}ku:�#]W���j�xn�����|�K��!b½�Zn:�r�4�a\̈6l�!S,&��!Ac^�<Qf�[<?�~���e�3*s�K�b��	Sx2�Q[�!�Z�G�&��Z��0ޡ�[_8��Ţ���P�9���	I�E-���p�-�{�g�"|J�{2V0�Mf�FV���<�ã�L,�Wvm�d,z=�njS��)y�[]Z��x{��΋�N��yw.Vt;�V��޷��}�&�$�P��=���3�a��7�J�y��0�6�Z��p34G�(��2O�}J�-�R�'q���پn�p<��b���U |��'2yØ���$�/|>\hR	�M�Hn��99�C�p�n	�a���	L�g�@&*b��n$H�V��N�ݻє�MW�����,�li��RS�X�`����-ҧ]<�^v������U�|&�i������xy?쮟�+z]�3�)�����%t� ���xw�Vcyٿ�$����X1��&�Cc*鸃ܢ���` ���kY��B��zhh���	+ܩ���[Cu�IV���}3�6?+�c�X��p@���S�I Y�?+KP��?��Ve��^3FL;���_�X����j�	���k$�'�<����ԧM�V'�I�Քа��ݡ��h��^r"��3 �"Bd|��4mF-BT�<p.�ZP�a=Y%�B<?5ϱ�l�*o8�]���0Ja����#���>w��,kv!��6Fь�a4�	�;�G�'��h?:�Z���#�]a=`��R,�T�e�RY��������j�!�C2f�w��h�6�7�8ށ�D�T%!�����|���
�x�#�w��@wC$[��&����I����#^O{`d��k���g.�A<�_F:�H^b���u�V�a2|��C�Lbi���o��4ܢ�����y���摧k�=���B�C�&��q�}�@���I\T��m�Oo���o�Uw�����*���r�N~�p���W���=�˯��H�1�������^&l�e�Te��CpC�oLe�._V��p����(M=�ǆcc�G��2l>�e͎�;����5�'t�+Dp��ρ'�6���p��ޥ_O.�I/0���k��2Pw�n�	Q��̀�/ߠ�Xl2���*<�w��0�+��Uո��هv'�-��/�/�p3a�*N<aL\7�p�-���^#���s{�H��r���-1���HM5��-������Ot�e꩹앐¢�l���U9�z&���@,	��|D.��@�k�Dm;?pᵎL�tQ�q�6?���QEZ���>d��.������g�
��B��9.W�A�n��]ڔ�pU�T#Z�h:×�������Q�DT�ݛ��6'fV��<~��x�WI�;%(�e����S��#��jj��:��?-+g�sp�1�
�ݐ��Z���%a:�%��˓Y�u�%���-�yH* 5���[I����.8=���;:�,"�������u+�n،nێ�I΋�P7�1��w���A�A����muf���&�:2CԞ��٥800�~�2F���j<�DFM����L�,\5C+�?w�2k��.�	���ږ�>[i΅�nl�Y���.ϓ�Vf������m=�_�4�G�P'~k�TP0�f�я�Z�6L���_�s�C�L��ch�d��狰�FG��e髩��$�jlJr�v�]��M(JnM����U��I����u�uǬ��@�Ö�����r�@�kbh�Td�5p�b��PXR���a)-A��҆��P��*F������tf�_gE�����9����>�G!F=p2��O�p�z�f��C�����F[[��ޡX�?�N2��%����Z�Ɠ�ﮪl.RQ��f
l��m��I��`!2��G�N�aX\8����d��Og��G�]�/l��|�Y�8�Qԝ��
CK���ڮ��~]����	������X1̺�G�a|�m�`����
�ʜ�Fn��=��B!J� ��3�Ǉ-J��>?����1e�4�2�҈�7+��C��]��pa�v����Q��Dک� �>0���p���_b�Q's��j��שׁ��ΐ���˧E��W��#1Q�\nJT��RT�Q��l#>�Up�	P�@o��G��Hr~�f�ݘ5��#��`^�W5�؄�ta�@�Da�$ͨ�9m�w2>���T��3r2{DI^��'�x�a�e�9�HN:އ�H
�}Mh���uvmiC3�(���GP��	�U��&�;C���R�����y�sgw�N�V2G&����`{����W���q��ۋ6����6O�{9�`��#X� e��J�%���ij`l��#�S�(��x��D��r�I8e��~�S%�kzw�T���A�Y+7������Vf��Q����B9#�bx˵ӵ�3��fb����c����gI��U!B��A~A��̖�^�	�������/�-��-�M±'A������qi�?Mj�k���~�T���U����� #ȁ�X��fL�i�[�О����M�!�i�ף�BbG(-NM�rаSÆ>}
G.�ŕ: I�ѕ�C�0*vd5��n�ڊ�\�����*��?:����$�������4��
��!Q�z�-f
ߺ�k� ƻ먧Q�mM��G_�Ў�w��:��tfׄ?ǌ�^DK/C�Thd���Ib��Oot�����	F�qĘ�ഔ�n�$p��3yf��@@��d�^��u E9�=_�Q�G䬈��ɥ�oY�������i��Ef�j#�uD#��c<�>����C�+@�E����>��k�i,'XΫ�TZ�&���Z�HAťbx��|�yb˼S@��X0~fr;:�Cb%��H+F�.Z?Z������ �5�\��/9%�Ș�f��)g�R�����3�]��Q���lt��:.C��k:N��W��ݒ��-N�8܊�94�|�>��b
g��I~6�I��]!,�����GЫ@_o�x�$�+%�����+��"%�� �8��qw0�Mg(��RqWS{���I��|����t��OM*�?��:D�n�@K�|�%�Z�.r$�Bp��5=V#	�qv���6��%����֘Ղ��~��E�3-^��ꑼ
w�1B�h-�^�!:~�OYMp%8�&S!@�I�rH��I/����n���Q�s�4{�
��ˊ��S@����k�'Q�r��چ�ȿw�,=�����1!�L�v�me�����U/	ckr(;���
��{����"ߞ���t膗����۲l�5Օ�>�N����������^�_`\���~^d	��K��:h�В I7"����zr����6'�<Pp�s"���X$�$C٦^�="��uՀ�2�v0�d�h\�e�B���.Z)P����b y�×����2�����K�'ߐ�M2<`�wNj�o��7���J�GƜ͚�|iV���������u4.��vh4E?�Ɋ�[����-�����Z�nf}�W%�����W���|D��Y��dh�:�umo����U)?_��U�tu�^U�6h��2|q���HT����Jp�	]f�k����"S-�Z�mi6��M����L�^�%4����JӍ�z������i6�d����1\u貑_J�dy�X�ͿT�(��tl*��D�LO�M�Y(��[4�"��T�ٵ��B'��@��V�e>�v�wo�Jl;R�]u�-��a�������Y�����f̩�$�I�t	��u��9�lP��
"}4���r�9e��1�X��CL�1�Q�6��;f�כbl��* V����wCy�[ڸ���2�ۏ�*���>=�Ts�@�x�ָ�[��#�RGd�m���vH�t�������x7y�� ���iK��-��5Y��$XJ���*0��;~ګC�zR�E��7�;v]�[ܖ�6_�2��#��oz�o�w3����W]�����n����M�dh8����D�ø�K�U�xQϠ��B�B���JG�0����{�T	����m@�R4�~�1�^ʰ��A(u n�#- �8��F��#)���f��
X)�X9:����]�ȭ~F�|���vmNW�ҹ�9?ƈ�>왧��0]�y'�oN�,@phg����w'WQ6\������9����&�j?�G8�����!�Ĉ��/wj5X0����3Ҷ�РF������HJR mV��IݷY��ޘã��5?OS�K@B
��Π���&���ď��be�!�*a������V`aON�t�j�7�	�]��A����YP{���A�=�5F*���^,�?��H�.ʬQ��ORR,lӱ���J�[�������zh��9-Z��ͨ��S{Gz��J��y)ڠO<��щ�_<�٬낡3��z,�h��.�W�I�m'��*{%����g�
x�ý�^�G�C�.��ݟ�?9%���Ⱦ��3�z�q�/Gc%�uљ���
�ɚ>˥�(�P��� x�/�浯�:�$ c���
J�@I+�XdC��r�vͪ��>��q����k=�d�č�J��9��]hp��ɺ}�O� �?D=!�5������y�JP��ۡ�A�lԾy��.#I�F����B�-�~�|>r�?9l�rRҩ�R�w���8�?�Y���	�R����F�dސ?b:��R��O�dϛB�>�¸�-G.cޔ��ԞP���D&���4�2��~�_9�{}hN ��R��:��&y^�UL��`��Wg�Ƀx�>3�$��M/�o�P�*ұ��y����<��������� ���iL�����>����ck����N�U1�ހrv���NN��1��\j��S�ζ�C��V2��W:���+���N�;J�0��ɞ��ָQ����%gg�V6�  ���K"1������=�����cI&�
4�\i_�8�&א�XN��r!N�a����e�"۪��-5�|�=-#:y�
Q�:n��*v-Q�W(�ؠ��Y��T6�� ���� ��.� �[��1��|`Z� �83������)�7�˝r�q¾��b�u��C+_��7f?tQ���R��$��u�->س���~�#���?1���p�Ԏ�����6ĝs���<}zS�<���{��A �6H�2�BOf&�c����t���{�~]��ķ�xN�@x-5�"uAΦ��Čw? a��ul
�l��{>˂�Iv������/�@�SI@=�,v�Z��������A��!�ERw0{�h�۶���n����<|�{�(�A>r:i9;�Yb�,@�P��ah�6����D�LS�Va �)8r��a�qD*f�~]h+�b(� ǺN��[f��ڣ�G8ONJ=;���6�ӣo*�޳�l�p-�B��7r�)����Zx٧=K�8��襪�P����tQ�|�⋙#{H���e��������H�b���5�F�����@�V� ��S��0G�=��ɡ	��#�o
�5��bS>�_����K#PC>v�;������;;��+����,U
K����3����s�>�a��� ��	�����<W��F��߂�������{���h��:�����A�E�hm�{�^���X�1֩��e
�_�-�H<n����g���q{����X�֛xM����rF�z3F6'��0�=�^	�9�9�����T|%N�Q^������k�f�Y*׍ASm+d8��	�=sԟ��C��`�v�]B�[낕�Jf��6������$��4 t�}"�r��qS|�D��־e����"aM}k�n/�|�EF51��<WI��� Yk���*ԗ=��r⍜�(�/{2߯	Z�V���p����M��[���x��?S�Y֒E4CT�^��q����$��j�KI�׬!^�`Y{H�&ʌp*���Rv�>�o�t!R2EmB�� �AA)y�~���,�<h�9�G����9u�\�������[���`z���������4�[��0;4˓��ք֌�PL����I�%.�4����M}W���z������n[mB����]�hn����EȻ���8��Vu��T�$%��W��Z+���-��4���nuZ�
(�yƛ�pp�-��01=s��>�v��,六c���/R�q7P����oB�j������ Ql(7��x�:���S��qӐv���?��g��|/�I�Jw�R.�\ˣ͍l�D����
�8���A�q�E����)���e��:�i.�_8�_��w'^����l/.��ި��7��I����Gj�$��La���`z�s�tn�~_�R�"̹�����{Z
�TV<�G7/v�AƳQ��[hґ[�֤�}��{�O��u�8�3{w{�ϫ_���0� ��X��jt����C5�ڶ�p"����&N�B���v���H�4a��x���OnV�(��&��辝C�nv�y

D�F�U_��,iZ3�zۯ��2���n���:҆��	�,��=�Xw'����E6͹`�:�L����i����l�x#V��� e>Z�� �WUn;a�3	T%�B��E��@�V��T���0���:,�P �(��E�"��0��I�Ӕ�Hy{M�j4̳�X����2,h\r���6�!��[�i�0��g���,M|��-dxєl ����:vۓP�]c��h!L��z��*�v�a�k��U�5SD����]�����]������%R#
W���|�qs��Ȟ�\s����$���]Z���.��)��"�����Q�-��N�->��x��AJ/[�*�����ֶ���͈�!.�Q(T�����$��6��ή�Vܼy�͐k��D�N���U�u(�*]����M�F��,9ǷF�g|��	A`sd�Λ�ɔ�Oe."v�o�P���+om�$-W�[�Uī���X5��� !A��\{c(Xy�N��(	�L�-e�2ܙ�Z���%���m�[��"t��r���5�R_5�kP�m"	ŭ;��-%aN&���v�J��0��i��qlR�3
y!�If'T|�v��NG���N���UB�ZGnY�
��l������Ε�yl�1�.�z>3%"��k��H�	 Y�CF��i�!�p��� ���̅X'@��RbH��qL��"�Vz���[��HI�*<k�.)Ԣ��=)�k�o��h^�N��hr��j *�$�~�Y3Ջr��cG�/�������H�ǳiOO��s�5��O�#luY1qf4�F��b�/��@�r�A����SD���B�/�F����b���-����ЉM����Kx*1��x]?��:��;�|�*�RB�N^���JNi���֋���������l�{�M���:����Z��E �Zc��I��ݗ'���I7z�Рo������Rj��I������r��P>���ڡYOv�d�	�/���)P �����
v��W?V��3x_�۶�n������*�kI9�P���L%��1�ձ���,&�`�ZU�uvm�1��
��p����k^�w,h���x�b� �u�/LZ�|��8Q��1r���5�t�z��"�К�2��"*�V**	hA��3o�ZS����K�f�
v,wi�C�%@NQ�z�򠹚����f?|���;'��z��!4��D��u-0UĊ�^�ہ���'M�=
�`J��M�]����N���(��0ARu�J�v�Q%�����_�T�����l���`��<s�EA�P���V�?N��疚�xr���:G퇴�=�	m��TG���CD�ecS�՝��59��1c@�U� �H��ke��<+�pI�6����C>�R�aC��<�"YOЁ�M�Ю�"��ۏڭ�'TS<�!���KbcG�4��|�P[�Vk�re�5q*�$9-m��Kgj�0� ���c�~�p�1���MƉ��f�a��;�錬Y���	_w��wP�����~��"
�U�[V�/�t��{cf�P�2�q����4��+ƃ�R�l���W��X�0M�4��'��0 �Ӌ��fU&o�H�D��M��U&`�f���ݔ�4�o�U�ɸ#@A�l���Ϣ� ���۔�!!�mg�_�ÿL�[\LJ|f���V�\Y0}O�M��Z87 �?X�����L���SW�I�<�����p��r��j1�����&�}Է7v'o�N��|�%?��W6Y���s����f�iM�0�Gi{l�`:eb�]���#mL��+��
`_�;u?�J� #��kE�`�������0�GϽ���>J���#qp3D�kr���~e!�c��c��U�ot�;��,�5�.mE�7Ia6�P2��S�*�	�@��\!�i���z����ٹ��nA8��o��E%ء�Ct񣵋�]��k�W��ԥ�G�z��C�R|�;���kk��n+��