��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�J��"4�=�7(�T�JѺ�ő��,\��s���ӣ�F�؏9�qI~B?I��$��H˜Q�<)q��{⊞dh:1m 6C��LJ'�u�	!�^�G��wȲ��R=n
�����u��'��N&?<�M~:���,;y�J�������^�4�<��
r:d��b����x턧�]>�v���x̴���}$��v��v "��L��0"�@��	�i;�8ȴ,&mc<���Z��B_z`/c�4��۶����7�[�B��j�+��T��2�Ye��U��#�����-�=NP�K�������T�/]*��u��B�x�p��'!�^��WVJw:aB�eƉC^�8�Eo��s!h1��=GTZ�8���MM0�K�)Sղ/_�kY�Ć{�i,�uE����=}�2��]���6*�X6R
�n�|M�A�\L}ۂ�<��o]�k0y=��t}&v�Z l�%4姠v���@������r���SvyJ��U�Bסd��C�CxSO-1���aj�>�GQmW�-�}A)�/Ї9��I��xҰ��cH��Z�2��do�"����z��3�h�d:"�_`���\-?K�CI�37���::�޸b�Mz�L�L#�=�� ���0�'-�U��t��jN�'轴�( �"�)Hn� �6E�^����+L� Y�o�Kۉ�&��1D-6���!����z�>����>JP
�X�nl�c��ۤ?���w';gN�KU���o8���J���m�"�Q��!�u�+�s�����4osf|�*��C�L��b`�JS��*Xf���hޘ�	!�>:�#��pQ�$����{Zv�$ɫ��3v ����d
���/{L��!�)o��}|7�� I��l�����'���'��1���α�_���ګmS�4t9�7�����fr����j�j��,�Z�c�}otڨM�	ޕͪ�s"`�Ҷ��Y�.�6(�U�M�ȮOD�\$�U)�%ۧ�eqAf����5��V��a�����G�y���i�ͳ�uo<+��E���ym����(�k?%8�i��DR.1�$�.�Jы�훓X [|�k���G��r��U5h��� \	hy��`Ў��P��,�96�������(�D*�d�(}�D������U¢)��v�lJX�[�Rɞ�1g0�+^#"	�L��;��C�3X���l_���I�Y��M���o&g��D�
�8TE��(����w���d�JI���3��F��\kY.9��!Y�hЁ�c�������́�`�� �m}n4c �bD�5��`�]��L����9-�Gu��:��$�����5>�qy��&�~�'�a�T�>�L�����q�س�mlMAr���a�v��O��M����[���Zխ�b�H*o:ȿ���e��,J,XR�i�\;ҍ��H���V��f��27]�)�oT�)��O}+ 4���?���;�IF�Wk���]� �f��c��o�B���d��"��`o�����@�h��;C�䇁���?���pf`3�*�kO�*��ƿ�����z�G^����y��+����;:��4fHn�g�蕕pe�N�-W���fA�n�!�1ܚ�����O`(2ϳ���p0� �rX-R� ����#8-|	�ա�"u�o���Ӵ�i^�)��~)>�,+��5;j ~w$Ȁ ������@"W���x/٩9ʍ�1NJR:-��%�2�I p�8���vHzd7�R��ϞD�cC��f_)O����"��{��r�42��V�K���2�YP�~��o��ii��TW�r4�7��I���.v��oݷN`�}=���W�(�UT�� u�#(W*��m�/AAW�5�S��"x����lU�ܰ�h��?J^Hb=��GM�P�v���	����j\�	l:FqG��]� �WȺYErs�T}挟X�Pt\M�����!��D��d�*�v�B`���Q�%��6�9�]�N�a�>�h����,dãD{N�T=��\�+�q�$�D���:�u盫@и(�n'ډ���^�wӑ>�^�yc��׸�OU��=���J�i�a�;�V���n��Dk<P�����/����3������vԵތ�6��آ�:d���p�8ʚ�r����dr�w/��ہ#�Ü�#[�]�3h����[�og����zJ��[�8�����R����;v_)�K~֒�S靄�^NFw�)�p[�y@$�\�йL������x_%k�R��7��7Ѝ�g�?D��?���毈�_DL��5�Q�AW+n��^Q�5�Y�v��oR�P���PYu�'���n���^}�?hB�R��f����b��HѰ35B`	��� e�P�;�%����������,X]R�3�JRd���φ9y�}�����%`G��0���B4.��pe׼��?���طk�A~�79��6�e@IU���{.�i����ζ{��ّi`�֣��J��ϊK�s�"}�]��U�XI��ts���q�Zp��t�:�X�UI� P�`Ϟ��d��C&�Ѳ��^�̠����i�f�GD��)ƻ_��ei�$�L�66�צ!;,�SŵՓ(��0?%w!�x� �F ������'b�|[�$ZqXL<��z:�F���{K�p��;c�v�X�a�D��2z�'s<~�����#���Փ�%�٨�nA
���݆L�	4�9������$(mϤbg!X���Ѝ=o{H� ��2�W��0��F��l�o�
 ��۬�9���r��DS\�9l�F�i�7g�����b�u@��[ACBLD���ܜ�1�|-��C�>\n�M<ռ�^�|V*f�GIE����y��O%�"+�/]92C�f�_1��]����e��v^h7Zl$�m˭��'n�2��U�8�[�9����X�L>rȺ���Z��nT~;y�6L��ڇ	�Z3�]fh���g9�(P��W3iPHXL o�Z��.�Pl�5�����1��w<��u4� b#�UG�� ��5L���b���1K۵���uD��\��{�0B��6U^��e' �-��#���OX2q��CD�i#(ڒ�B�R�gwP���̌���t�2#��{@�lϮ��v���	)@�~.~-&aQ��\,�'�tc�c@3��A{�z+[�/=�^+,�RH�*����po��4;Ľ��A:�?shr���8S%��BM�Jz./�i@yX�
�.��	�R�'��\��R���-�"��.Q�Z􋅟x����\�v`����%G���R>5���C�yxi���Y앑-�£B�>KHz����X��Sj����32�t�KQ��Cc���+��'  ��F�×�׊�uƥ�Uې#.�Y��4~F�A�{+�h{UE�jitJ�����^�ɛ����f�xL��br`/.��'s8 �Q���>8P����1p��@YN\�k�Q~5�-���ި���}��0���NO۵�D8c�G:%ڷ�副ٱ��d�~e�o4*����g�2����}!�K�A�V�>t����M1�أQ��$�\`^�'b�S(�8\i�hM9N\�,ld�؄U"���-��KP�E+�M�Q_Pl�J���F�OT�>�pf����G}�\r?Ly��[�+ܗr 5uƽ�k�,T�h�hPW�&�aB�ٳ3K[A;?���d7�͢α�k�bx/�J��F�-_K|�7��֢���A 1�W��(�{P���"�<�l�Ծ�02�����C�	}�X�0�>2ox��)g�X�����\K(n�X<_lT�<�6rpkpTL@Ί�rͥ0L����������b�Q|�6�e��7=B<\.Տ���Yj��0>F�t�׷7��;��\~�i.)�����&�JҚz
��+���{�3г�!Yj��	��j&op(>�D��t�����&<�S���;��W����С����(�P(c���@�{[`�<���a�!,� ��B{j����fSq�-�W$�8��׺\��g>�l��:q���h\)�C���2!����3��u
Ћ�uQ[2A�}�$~zw����@��<pܫ��>��K 0e�D���s5疼-�z�B��}���ԥQ�r�@H> TbUʮX�.E�t��n�9ݿ�\�o����%8�RYo�B5�e.�5:X�E�9lG��m�+�hGA��C�p��,?�\jVS-GZPY�+�3��Z�U��7jv�1��:ֻC�?P���Fc5�����u������?��H�$��W�ʤ�� ����Z)k���G�4z��'��+�:+�(}�N��խٔ_�Ж-�����uy;��|V9����Н��!�fM[^>�C���_C��� �Ls�m� �+yX��ǖ�pt݇�$.��ӔɃ�������,zm ��:Q�CW>��t�0]�N�v��JI�_S�(6�y����:}elϋU��Ta���!�҅�J6c	�l�ֶ�/c娯bK}u��I6��z��������>)�v��j沤hI}�X}z�W�(g$�b��_\�:��l5$MS�_��4枢��w��L�N��3�� 5�R�/%�*����K3'���Grw�����{��܅-�ڍS�a^�Qe��-�nҝ��{��Ǯ�VCoL��=�	eV��4N��(Z�cz�G��KƏ6,v��P�3� �长��4�Yh��@Zol��&Jϒ��^Wz��B&R�WL�{{�͉�JҧBnn3PS x"Ab`q/D���]��`�͍�̡@e��� ���	��b�W�usF8P�O�j���k��=�h�$��$��/���$��؞6e�:O@ol�tTKzE���0�)g<�%��cƓ��\�^+���.�fb;QV�{`����H�l���u-�;ç@����#�j�T5b�x$��۟�Z(3�5��mK5m�m�+b���)��d?�M�������5ը�����?��v%���+0w�U_'����5m�����ȉ�1?�h�f��'ϗj��Yd�el"���:�!���JK}w�8�"�͵n�i$ȅ��E�����q��j��ǦM�G:loni�h�ޗpT�=�ar ��|�Q���Uߪ����t��_���s:��N�ґL^�gF@�u��o!�SA��v��WZ#z�>#�P������+5�{�&���n���4�熞Нn��zu%� ��%1�%gkb�n!�}�҉(7�����LcZ6I�*��D{��Ű���v}Jizkv�`Cձ_��u��=��Ֆ�x����v$�v<I׵8�ǚj?=����
[\3{�S��1��(Q�hZV�7x)�9�����pr����c�XA�Օ3o�bU�@5�!�:�M�k95��a�R�-�x����ac�W
?�T���A���Tf�������M��i�y ԣ��y���g�e�]�s]�=+:� Ə����O�oԤ�D*��Eߩ�n7�E4��yl�w�g@j+��'����GJ�%����Q
(P������U����{u���ŀ%ù%�8����P�J�}����zKg�G>Լ��i�ѧp`�]8���x�"����"K�[82B`��f�}9�i0����X)Q�'��
ӡ>�؂��[!x����5��ѣ�ymҟ;��3�$��#e��S��W�t#|ȋ��jpx�q���XzH7	���H�B�f<闅�����z���+U�`�s�V�dC�ŗiL����nn~�v�z�2O�\������r�N��hGjo~��!AXR
Y�6�wӒ��#�+����C߇	9<>�j9��.�]˷��,9���3���zI����@���W�1�����D�ĖL����$��Scf`!���`u���~��8����Q�P �ԡ/y���s3��4}��	S3����k�п����
y�d!�k ?ݚE-%n�}�����|n��{R��}�"��i%�o�/��F�:6Q����T'P������������rS��XV���K���άx�J05XيhY��3�P�_�i���TW-�n��/�ڧ_zo�O��z��rr�GrA4u����~k�{��,x���� c&��5�F�vEI�ν����<��XQ"��og��� ��BpG�@m7��+5�!JeZ�3��|���;�J�ٷ�1[����<Mm�o�m���gօ�A�yZrhw�t��O�b8;�.��uBZ?Aŉ��:�f���:]� I |1�U�[���Z_��&ɸ\������w�?_U߉֝:��J`c:����a��]~K� �N�]�f&�եk9,N�m����-Z4y/�Zf�4�p�?�9a�a������`���8Q�f@.&��zg��	Ohl�S�G���x��aBv�)�_u���mOf�el�y��T�@Ҹ������6#��,BD�<sP�{�ʋ�!8G�x��\�DH��jp����6Y�>� &_zɊ���vk��2���z��vm&��;��.I��#5���N�O�dI�;�9dn�mxk�Y��m��̵xQԋu�MZ�3��0�ĆK �%w����=<ӑ*��
��b�'��qk]s$�v�?�[4�1�g�� �Gߨ�QY���9DY��2d���8�tL5�㵛Mh�E��c�k�����j���,�p9��l6U��t+�ݠo.i��^.�H3�>"�~��6V��y	�H��;i��Q����iF5`���Ƴ*�`�X�cYd���c$��%���Q�,�հ���Rp��Q>ҙHD��k�9�Ŋ�l5��)+��_	z�W���id�X�b��@�������i�9'�/_�6N*Dʙ­k���f���a�� 
�Z3,b ���PI�'��;�ۤvᏈaU�(ϖ'�o�c����XN�^�����a�^b�&B�)i��fǘ�".����� PR��F&	[h2�Ԛݘ�~8��sa�Х�Q�
Ӥ�J5��v����@^�K#�^�Ag�Y`����$՞�'ؿ�PCڷ��W�m�:� 5DB�7��v8E�F9�Vc�����	с7�[͏����:����%)�frFY�L��A���5���lz{(�#�.�0�((��A��mBL�qC�#N�נ���::Y����<VO'B��m{��9��E@i>LL.�K|�iO��%
�z�� ��6b��h^h�,�zk�n����HU��<�g]�HK6e��Ի27۱������ �b!�TQ��>���<�ð�e��p�0<�k|���U����͍�֮r#�k47���d;��CT�M�M��Bv�1窓�]v��aO�ze޻�G�PqLo�Z׷d���H�a�ɘ�ة9��n�5�� u$������&�tN&x1��?��UE�Ba���]��
�$҄Qh�DB�Mٙ��An���H�LZ���Fu=���"�(��	�R)�*��N���	ķp����z�<�O�G3�/6�#4>[�LcQ&/�úp�p?�h�	��D�Q\&+�r��k6Mh^5�I������$]&W�v���p�m��V\�]]K5�����$��}�@J�S��UU�/�7-���2��Z�u���x��=�4	.zs<��
���^��e(bH
U�	���j�EX=@p5�<=�#�40��1�e1ۙ����8���f0 ��ȶb"�G W3ױ�A{�ޱ�	Ɏ�`�䍇�q������ؿ(�.��.�Ny���c��)J�ԃg+)U�3��@��VWCIh|bW���1%��[�|���%��z��n'ވ�gjZ��Z랦�n�_���[��>�z$�� JU��&-�ϋ��3�>��y��WC͟��,+�ۊ�'���nk`�̛���q`�WX�r�f���G��大�+m,QRuM��Y�l��Ň���F��PK
d�pϦ���y��؜���b$�����Sv��+|}]��e��r*��l����Ks�����E�]���y��u���E%���CD�c�AJr��U:�g �׎Yd���~�3D9�|�Ҷ^)%�_E��k#&�ă�X�wx=᾵�ɶ.����DZ�@)��T������;9z��zC�i��	95�$v�r����C��-��O٦�h�`���F/�PUkMY��PE:ǒ��)��m�H�琐@?��g^�����ɻ��OFp�+�$��<�gw�J�IL���9���*��@�'�N��c
�j��h�BK��,Q*�W/*���(���)Y�_��!
�Kb���H�~A�7:\\CS m�B�:U�ݓ�ъm��*@��@���v�C������g�����K
�Bϐ���Z�C?|�����%Q!���C،��,{I�3��R���� �����>�l�Vct�XA7��Ӣ���LĔ�p�V�w�R��Ȳ$u]�ԖTdx�K�����"�޸[}�J�D`\u戻�3;*�16L��҇�3@Sh���ob��7pp��1�<����$�owj6(���Y ����'����.p�>�sV�:&�5���ި����,^�v��Tr��G�X�n)f�~,$���/�~t� B̒o��h0w4,w���s�}������=�@'B��Bh�'8��W�X`�j$��چ3"9Ƕ'&nw$�V]�Ep��JH��b�F��E/iH2RPT)�N!Ep8����p�i�f�U�IЁ����.۲Qno���cS���x��C]BUܝ���9<q,%l�w��ɨ�J����(c�5< ,��x	:�cy*��
#Y���c�3P=�
�����������D_@�HEq
#Xܟ9��) ro��'Q����^�gY����~������z�e�T�g5�\m�Ş����C�_�����u�Z[�˕��u���<b�I_�/�/࡭�vc5�:Wob�^��h���l����f���Ϛ处T����y����&	�f�EA�����)�#+^Yf��l!�s!�9�/����[����'�q�:
Ǩ9�c!�%��r�r��*8�߬�e]Mp3-^h2dZ�?s�t BN�rTr(��z$� �5���9��t�v �"U���O{ o��/1k����wb��#O��\�7{��J����,z�����ߩS���M�<>�n�v$�
�R�"pJ��u>�?����p�D�`�qa��֌���Ր�a����4T� ҉rJ�Zì�p��Z���c�:�J���f��N��@�No�� !���\��F��p���:�t�R�Ba����4bF�p���7O���Uև��c'�J�VҼj��^�F��_���15XQ\nb=N�w<<mc�I��A��5$f=n�3���	j����~��-Q`���>��%)Oğ��I*z�\�*�Sm�U~Gܑ[hi�!��@��.�2Z"4I3P������-�WwS��3&�
����0[�1n%�v�UM�&wI��e�L"[�����=�X�z�%�s����:m�O�L���Y���f�,V����]?aQ�6���i
$�Ih8v��0����0�gmC���KA�Ft���k)f�~���ځK_é8�� ܆���2�߄�M���#��>͙oM�T��Ҏs��CHf�������-���#_�ؽ�HT����������:l�����]��c��]��z��ST1�3�#�)cj8��<��)���s`����ʟg����}�CV�����5�.	OM��֮�ˎ��[�6ў�ӫy���g|qn8�"h����:��X�ݵ��5��\ӈC}�-r+,�,�x@�cr���s��m�L%��F:�͚씰��-$�����^�y�Jޜ�<&P�#��4&ze;=�m>���ު���iŨ+k�y>9@F��}�,�%A,=7d���1��I������'~�Y�S�DsW���Xԇ����;Ō���@r�Y��1�c=���?	&դ)v��p߬6YDt���b�?��JF���u�1��,֑�< �H��S�����Az���W8��Ot��2����V4���bx�����	�e�f�h�(q��c�b
X����-�͜��q����
�y�/ \�µk�u��SZC��7�[�R�tVPS�it���ؓWF����_$V�[�<��.J}�#��g�Ӽ�gGJ \#݈����.ۋK����E�D=�:ۓ�,v" �I��A�Sՠ�����o@,҉���T�T�p��k:����m,!��k3�.��ik��`-M��Go�`�b�S%�2�����ŝ�/��D}�;�ņ"�0�$g�8��
M6�fV^��@R�0��E�I���%���A&�:TY�U�&�H0��G���s�@CTR���/y:�1c{���`����z�o��ߛ�r'�H��(���yg]�s���!�SbH�{����Gxf����^L�(��7������k��N*=b5�:S��������w��Sa���T������':���0ꆄ��n�+g�΀����"0	�����.�ګVGz4��p�ON�IǝX}�Pϯk|�a( Zlސ���u�`1���g�:�aG�:a���)�ojI�b��iJ�|�Q*Uwh?��"��p����ռ��{��W���[]wQ�s��}\�_a��"�WF�!.C����=nt�=◡<S�y!^ ) ���W&<��?_��сk�+ޟqȢf�8|7M#3o���ء`Z�%�w�(/j��R%�Ԁ5B�A��g�';���3�c$hN��v��>�W��� T)8�qjn��"����P�ZAa�_��g~̆��'ǜ�E�?�p,Ɉ�yI�1&i�DTWW%�e�X̤z1Rc� ��C<�\�H�6hl�����������z�X���dј�. ��Q�|�@%95�M�8,�@����L���;JOqV��?pG8f�?J��:L�!hQ���.0y��.� !����AS}%�l��M���
�-��R@[�+��Kb�[�#��pT#�j1惵 �W��h'r�:D�môM���i޳59��?��y�( �m6|��zG��qO�����ֱ�g���ME.�{��HVa G�7k�7Gg���&A�<�!���Y�f�1}h�W��q)�y`���N
-2��A�ș��ͣs�bT���Y|�&��c�������c^��˫��v��1рa�����]̳/�
M�9(�34�U5�M�Aw<�1zϠ9)_˕��9��E�����l]�qj��P�����	�`�"��l�p��f]𴑮OT��YY��Eol=�il�D� V���!i@��$ER����>� H�5����}�c���]sf���2I�/.@��n�v�/9eq��O>ͥ�9`�ۍ�cr �2v�q���ؚ^�����;�\E)�4X��	Y�m�
���y}YMe����Ԓ�>��xcYd�_̇ލ�ܨ����(��o��I�&-e�������2�[^�f&�+��(�jZ}2�h�p˼e��7$֯g;��^��MJg�vh�Bi����:WG����t��x��mH~m歴��#��3ͫĨ�1�0$6kP�* .�`R��ʤ����b��Rۀa��`l{�^A_1w}�j��ە�����P��i��ߋ���P�񟓢L�u$.��p+n����gA��� ����Q֤1K2����5*�n+��p���W�8����Ŵ��K4�g*{�����I����_��6�'�����O���˫��q��.�b���A@	�9�f0�\M�ݼe�*U�� ����%j�l��2Fcǒ��Zz�2���8��:��(����͇�"u�TکmW����aՒrE���Q#�T �mq��YG;���lIX�p֌�n:텋=^ۦBl��"M:s�8�(2�=��mbj�E��D��!�2s�9Ĥ�^?T�De"U��Ca�
� �y|�Y�"�#���pƫ�����w�.(T/�"������Q�Q|�	Z8V$��� ����?��w6����L)��F� ���$��)�@��iT�������PX�&Iξ�r\�c)ĕ��dVe�Xt-���h]�G�3H�~z{�_�,+n�qd���55��M��\�m �Q��}��h0���2s�z�G�˪#�_�������9>�HÊ�2�썆D^4PI��1%ypn'���Xӡ3t���s2o)ɜl ��Ԏ�i�3�A?���Ҥ?O����a<�LZ_�a��2�QAɟ���2�R�̓�0�J���/�X3�m5�	lSP���ROψ�@����`}��RO���>t�!��,��q����� eF㋋�7�-�)�1x,�pAr��;Q�ܘs���Y��Ֆ�h��a"�#���Q���G�����EI���Ya����֕x�,@I)��t�%	RNp�^^M0ޫSڋS�8MU�����P�B2t�@���"�W��e}1�1ę��b��9Zv��\׆Q�8�d�B�k)�~KOi)q��>�aäg(\��@9�+%���hdFhEo��t�\�#���zI�	`u�ۏۙ~�/�̸R��j�T��SV���:Ҭ�P�&�b#ً�>Y��l�_w�u�����?���h��q`�aR~k�s��q'���0X��Y�bd�H��q�of�@gq�) hJ��ܯO�o@K=>����Mr���%#�o��&�*}��г~�L���3,��j2�` �9�T�C���Ǜ��*qfy�Qv [ ����?h��l`YE�\1��%��%-1�4.yb.5 :A�L�S�=� o��͔fl�|��d1*��lLEଉ�5Ƒ+�"w&����gʽ�׋����#�	��;ОA�|���_�ю>���]Nt�Q�Yz�D����o��V�@�T�
;i�G��߫����kz"P�����o�H�8^"���6����7F2|�k�+�f��]��W+�*�I�Pw�&�zkO��KlF>2=O��!��2�˃ї���Ӊ�=����� �ڡ_5YW_��P�T��%��wj(�^SO��˸��l'⛄2�����>�P���N��[H�"�a�̈^0y��e���cm)���I�h�*{��"��.!������]�.�S��q%���1&
2����-�=S���AfN�=�x� +ĘV�5Q���g���Hb�sT��v���.ti��SR/f���(A���h��T�]fq�	�0���$��G� �f����VJZ�żj����@�7��r�~�#U%�&(s^�H��;�<��ա�e��Ni�������F� �|�;���Q���v�^U�)���c���­�����
D�skљ��&�/�)!��Z���gys�e�`�Q7��q����/.t�x`C��J���G!�\��L���I*Yɸ�t�jB�v	ԑa���"!^��ԱT�:��7UJ0���<�T`)��N��(��㊯�y���q���H�},�,�Wr��5��к�A�$�C���<�Nc?[s����G?Naʷ�@��(�ڛ�XQ0w4cZy�j�R��(����h�����_���.�{i������R�r�r�<�|���Shȕ����'�`g�B�#L>���)~��D��� q�5�_�nE 8z߻�UKʕ�0�Lۉl)T�L=h�����\���iQ�_\X�� �,g:# up��B)��0��8�Ր�P��[�%�T%FR2�͋ۡK<�jz�hE�S=J���
}2��8x|��O���	�eLR��]j�qH�l�m�A�#�����5�C
#.ܴ	B��>�u���u�_p�L��CX�"����8NO��w���ӷpߦ�.G�n �#���F�-��T�E׵0��Jș�䄼/�q�����g?g�j�XS�N�[P���m��yщ�q� "�}�!
����L��mM�
qq��1����N-�f���,'X��N���j<m.vK#=u>�y��`1%�c�E�z+�V�xo��ڴU�}�Mk���E)��X$%�A�7Å�	 �se�?<[�=l���cԧ@��p���۝��8��e�oeM锼�ذ	r��O�!-��eO�H9�����B��׋Z8�(�o�����9q���pl$@
��]��ѻI1�֨�1�r�&-��3�w��K��� ��y�Q)j��<�Bg�Y@Y�Z���lU�`W]�"�S�K��M���(��Ō='(�w����s�V�T�Ϗ� 8d}�n�e�w��	NoM��=Q(Hz ��Ȣ�@'y�*�=���#��\hf��	���EF`��6�-��yr�@�G�,��b�����@�}n�}�I�ư$A�)�~S7�P��Ur�fuU�<Z�g9�U���P��<�Hq��R9?=x����M�+͠f�/�#>5?#���q]�[���L��и Ǔ(c�-;(��mWS������J�f3�46pe\&�����1�R����a�g�[k�����lp^�E�+y��+m�1�J�a��/J�� ��B-��$�H[�o��%�K�\ͰI��AE~�,�/�L���m�Q ��^�={#��]�un�$�J{ Eu?�*�iu^����i���G����}��i���'RH�7G����%G	k����F�d�+�����F��V#ӏN���;�9�����0]ҵ}hD�DZdֺ�yͼ�f����2�x���Df�*~{���6�7)�}��J�tO���!w��ߘV2:0����_�=D��%�ٟEU�Ԥ��o~"�J_�.6x�8<K�,'r�?�9<)-�N�iu�¾o��8�:��nЈ���<��s�ڃ�ؘ��K��H�M���e9 ��A��N�����l�-g>Z~�阢I�S�[{���*�a�N�~��� � ��']N�s�CO���b5�o0D��4?�t\��|&���������w����ݡ]C��=yH2�J��H٭�6����/\�
��](mP��aB�D����ɓ�Lk_?#˧�y=*ɕ~�×>�]��?0`C��)���ćnJ[J��mxu`��R;��.���kґ|��ga��"W���d�%�}�9��fK����\nF�莃�[j%�2h�i
R��,j#�@5`��B�����=|���D��E\I
���ue*���tH��
\�@����p�S*�ȅQ�����tK0��g�(j�=�5FN���*b3q�o�9���a�u>�n'�o�M_W�(� �{��x�����mLG�'`�{�Sq!F��Jp��%�D��?�q�zF%CL��'8�W�� �)]ϵ���В̓R,�p"Ľ����W5��6�w�/?*�I,Hn66�#�tN�����x���hƑ���T7	��.A�."��|�������ÐG�[��8�$�jy�>��TK�ۉ�f��;�^�H��ް,����U2�X{�F��U���r_[s����} �J:�YV����O�u�G1F#G��>	(�u$���$�̧֢����U�� >�1\��~�;}ɬITۀ[�;����H���h�m�r	�,�n@ȋ���N	�ck��d��!�N�qp�~K{dM�PX�	I����lEyf#Hv]��#z<��_�7���p�u"6KYQ�_Զ}ۀp(���V��2b�b���I��20��I�֒��r����F�������𫿖�jTu�����K �M5)��uq���ꯞYH:ˈ�bnPѱ���#��jW8������*/XՑѮb?���z��"��9�붖��K
-��ȇS�pC���}&�ұF �5j�l��[�Z~"J��I�\��� ���aӁ_왖Xs��f���źt8���� �;�\8�:n�>�r/��.+��tDO$�v
CX`�jiJ|7��}�����5��@o;&%��,�;���ܬ'(�X��@���S�PՏ��b��o�Ӽ�FRƨ`�"��c��i-�n )=��w�i:�W�,P�����N_�1�
��:%��i58~��P��
���M��Y�8��s����+���Z.̹���/(�h�E��縧7G�T:ǰ4l����`�T~�:����J<��LM\�H���/��(���9�)d�ã\��i$ ����J�ҝj�r���ЈJJT�r%Ш���Ց`�� ks_�!N_��8� `#�;0��@�4FT���c�{�����k>�evJ��7����8����CcCU�֪������8��6�D��Ƶ�����L�_2�Y��
�	��c���ߠP܆7r����ng|�f����N�xL����O6�j4�S��2Hcz^��Z�^.�-�������C�W����h��<���57��qM�:*/��$�h��ϝ�i}��=cG�pA�r��"ΊJ�PU!�2�fZt��,�q���ZZ�^S<��x��ҡ�f,n��*�v�c�O�	T W8����룗�X<6{p�J[�"����Q��愾�N��&a�yŹ�&~qS$�G9��	��?vŝ������z��x�p���c�*x��=>�K��ɓ��1,�H��0`o:LМ���}��uE�=4u�uL$�A��
�8���?(bL���9�jM�D��]���XɃ�|ZI�
��d�gH���*�Ek�9�(�@i��,;Y���ȭ�B��!9�pD�����K�N�����|lj&�(Ӱ��/��L��dP�E���e��a"�C�d��rp˶ĤςV�M� <�F/n_U��,_�����Ò�5k���G�'����yW���(�Gm;���z�o��Y�J�7�*�y�<�>mz���lF����������K�*��T�@d�$��io m������YB�ȗ��B�+E��0�&q�Wx������	'q��5K4�C?o���O�sO���Q:DEl�`�l�L�W`���~A�퇭�m�N�D6��[*�Zq��N�Ve�����3���+�"�Ra�e��ca}}��$�}��|��$ɧLWkRA��:��E�G�SR��V�Xb+k@5r�����s�<Qj�2�$â$�h�2>	�� ������(�e��Q��҅]O>KK�
?�v����O"�D�H�~~V'��Ȃ�>E�A�,|�)n�SKry������~����4�X	���!c��,�/�x��c'�Lgeo��3>8S�*��~�0x���s�x̸�w4?��D=-m���/���\��7A.����ϋ/��B�z`���te��rd���6�*
-5����А�@�����]�J%$��hC��~�h������}��9ǉ.m/���Y@n8͟7匪08��տ��+�����a��Ef%�������E�W۷����u��u��{���r��M���p���#��mf��B�6�-�w7;�zU2����^L� S/}���=n�	�r��z���L,�1*+"A���ȆAUI���%���u˷)�E�Z�r�1�=p�_jC<����-��O(��p�?�&��!d8�M��7����P3B��=)�����ig�.�,�U@�,��>�V�J�\XT�Og�&U=�P�5�XR��
K��/K�y���aO��i#P��ܗZ�$P�'c|���f��Qj�#��6�z�+�l��Ȧ �����̜����6>�؅/=T��U��|�����H��_�N\����TD�'io󣖹l�/[e< �T�I8��g^gCxI�r�CI`�1[��F���]��n�,�m�g_����6�0��rnKK�$���C�S�en���~�i���cs+�i�Q��������6 �2-9r�<P��E�Ē�����|J�6������7Ѥ���ک8N����JM��
��ЌU(����FZE"]�-��Q�g_��!�u�29�V�U8[/�
��S��T�-���`��j�'P�&UPZ>������Sta�qю�!�xi�pO�4h�ٴ���a�G[h��y/W�ۓ	.yZ� g�o[n�l�Ak����4fl�Z�06=�Ɂ	DO�n�e��.���Qr5ў^�$�&�>�����ək��-��C$ၞn��|��F��!Wv<�8t�x[|�!i�kY3_��#��Y����2^&�v�hп��@a&���f������_���|="���;���D����bl!Oo#A�����,n�AKO�^�zz�q/�0]r��3���&�6�I�#V�?��օ�]�&ZV �%]���	z��^h��Y<�O��	#0*���yW:_�w���,@��b^z�ң2�E�S,mP�����:�uO�4C�,4��/���q�0�>����������[�(�cU�g �xy�D�u��}��D
�Nĩ8�J��j����2\���4������#b��C��:��̠XV[K"_�4��t��$��@�}1)��p	�Y�v8)(|_��^��� \d�[[�[�!�����l	\�K�pv�s���[`rK|~���ſ@Bi�73�ɶ] �"�0l���O�@���@���&�:���>뗖8P�h+���e;�%(�q�nA�H^�4�c�X~2E��_F3P	ۍ�b\�~�4!''��&�[�]���1 S�������c<���^�����c��!M��eAry�x�s��R>i��;/s�37��-�Li�%�:�gQ'2罋ԏ�B��6pk�'F��V����M��³!�������r�X�9����M�kC�4J�9�p�m�8�=��"�ER֔~�ws �b%�cdՑ�8���H"�'w�K��gXA��@m1��U6n�_�w�=�R��uI�	��`�e9��!�Aj;w�V�n���P�1*��S�0zwgTb�jX�I��y���׌N)Љ9SIՙ�y�W���9�Q	{��)g/�LQo�}8d�T��訡���t���$�w��\�@uW�#:����}_������0g>Fa�3�^�{�6e�h��놉5C[W����R韚��#5��cG��l</�ʦ��c����9����K.��󧋺���^{EorL?{ȺoEW,���X����<�(�d���A�l�$'��2:��ijZ��D]Afo��7����~I;����G��/�?x��Ƹ"�rO�Q��D�� m�V���)�P{S7(�'8��{C/�τ�V��ZW�x���H��j�7�T�a�<��h��}�)q������!���a�ȗ@N�j
���J���~_V7tx��o���rQ��%�N�8�N����L��!V��5�<[���x�X��׹�M��c�Wi�F��+o(���۔LM�f����xVs|��,�9�;���M��zͨɔ����ˁ�a#��;�����!��X"�1R2�COwZx�a��f��{�r�=|���z&�׎���j�"����H�E`�h�^�YJ�X6�y��i�Zg��ςGPN0���X}]��J��8��!��� �ޱ^�#֦:k$f�KXSQQe8�RM��gB?��(��%
�a]�;���u�4���@����YY�o�ڸ�ȣ��>�ൄ<�ֵP޺��,�p\0Z/C����'b�:�qF�,�1��v�� ��7��{Dg�֮-n�0!:��4-G�[-3sL9����)�l%j���y	�Y8C�LA������i���ܸ/&,�5��F��s;�,�f�8ן!7	�g��8�� ��00�)6����bꆀ�Q˱�U����T��^X����z��@߭h5m��IgS\�-��/2A#b{g��g��"E�N�n:�r7fU}�1ŲcA-��PS�l��-;w�Qy������d>?  ۔z��|Zo4t|��a3"��p&��{ĕA����I��t��	U|�o���:�Q�/'�d�����K��Olܰ@3G�ηKw%+�r��i��K|�f�O֌8��_#.x,ϯ�،�B�����ðTA��Ԑ���S%�k�t��f�0�3D!km6>ɶ��Y�fki�4	�����ez�Ǖ-Q�"s�����dVa-��>.����}+
�Δ�X��I�3 /s�3qC2�e�W/as'�s����e��m`��k�m��̗M�������E�ԡ�S4��O��`so{�;��Ow���B�x�pHL�.���v'��5������̂
���
a�C��֥<�Δ'FEZF��IL�A��w��î�A/�L�A�|,a�{N�H�Q� �̖^�v��(5����-'*l����fmD$�=�R,��s�{
�^^=m���t�3��%n�r_ݠF>�0���r�3�{f������x�4�
明�� C�fA��4�c��%]��'�O���;q{"��Մ)�>���+��X�����T$���n�(V^Uʃ��e1�c�%B#+��e�0��5����j�宍ho�!Z����Ol��c� "@�q�?��\i	����a`0�0^~�W�_
���+z�QW�dg^�wmU��Yk�ַ��l����	�@W��X�]ǵ��2���1�+44ޫ��r��U�[�jc��T�
��@�O��v�l�>���;�P�U�����S���p|Ϋ�A��x*U����2��?r|�<菁FE�v��^/W�]��{������q\�����z,<!�{4\e	XO�C��񄉬�z�U������/�H� ����1d�P�X�ʊ�]v�U,��V��%ذ�Jm�Z!g����󒏰���|�����g�Q}<�&�ٵ`F�_?�(�#�*Lő�a�$��1���TYr��)�;Gm���S��������g�޲�hnk|��+�d��-�&��ڠ�� {�|K6�]�W}u4�?���?��q��kZ�g����H*�9���I[��v��	Fp�$V#���J���ߝӼ���LM��W���5��ɻ�`�Cp2�V� ��\z��u3��OOŏ��<|�! �h��h~<��+��e;I����e+��!|�m�T.����&F����QBDk<�Ӫ��/w�kl��3O���VttM��n�QXL71lƦ��\ bc��r�_ejֿ����G/�7�kAChr��0W����������@5]Ld��32�t���S���#궦��t|K��0M���=��w�M��*ݦ
NV��C�斲�Ѥ J�`��8�`՞|ڔ��� ��E�A��-����,���)>�/�o�D���6��&H�;�|Z%��gJ/��7��|Kt[�¼y%X�~œ���i(�u�VOk qP�0<�*�u�ǡpb��-��1]@����T�U"Ij��?�rϺ��N�f8O�ƌ�0����f�
֌�B���G���,�6��]�o��_�s$��+Yp`�x�(H�y�
�W>4_E��-�Ձ�C�(;��A�x���������C%y�C�2��W;�.�ؿ���Q�:4�:k�tL�!�%�VQ���j�A�/푖S]R\��b�(9��6�)c�_l<�w5��9$�kPk�����/�y{.^˗p;�W�� qU�	qc�U`o�! U�JE]��ૼJ9���Y`�6y�*�}դ�~���D��;
�����̗,�9��T`�}��d���XJ!�ܿ�h��6�v�7��z��� �R%8����y3 >�zl�\��n�E��z��,����4��O2���If��>�t���ӓco�i��1�)B�[�a����WЮmK����	IQ��ڝ/�.�^��u��y��J�3`��p)*q���IkK�9�q.�-�!�����ba'deJ�ዊ4�X!��[Q��>�����N+���;��Xו��3�T�����cEp����8��;�L�f�A*9+�Q��`�w���a�fx)����V1��p�>Y�@����#���o*�(�v-��W*�]'��cV��?Jd:���?�^"��xaÎ��V�	Un三%[����4�*S�?x�7�������?f�m���jx��)G0ݴI�Z��]Fr)�C��Z�b��А�r�16����4y��t�Td#;a%'��yI]������a��s/�V*�ī ���rk���k3.���Hj�PF�I1���d@&�ba�� H�jI�Sc�F<�G��$p:��݉�X��`?�t�;Eù��9���-@"� �q%
������ctE��TKnMQ�XR]}�H^���8B��H�+�^E�x�"~S�Y?zNe���!f�(�\p����DpaI�C6}L�X��f)W�@�Ϯ'!� J�ͼ���~dqdn�+��J��_,Q�Ǉ6��`��@���\�����k��9�~Z��Q&�	�����`g�r���Z��*�|����b9纥�Q�*r\E\$K������b.ݙ�*�`F}������t��7Ge.M����{���/�����:v'�oB���mL�9#�s)�T���bfm�c�qW�LP��|��
C$a��G�$`Ў�BR��2������au �
Ӱ�Z)�[ck���9"f���G�d�Cg���f�@�<q���p���^�(ׂ-�Q��U�,C�3|�����>�����rt�2N/<�h��U�f�	�WMq��1?��]�u���Zi-��p�>,����}�����G��|j��ީIIz��tm}G@���[�pg�q���Lr�o�ž�=m��)�kC��xs���`ze�ޒ^{μ�|�X�I�f��Y�J.PZ�2�!���� �T�ç��g(�zW�x���q~���%,"�n�>�����&���s�*�E�w���<T�%���v�� }/M�����
��ztF����.+�����@���T<�Z'����ܾ�����{l���s���T����'���j%����,cN2�%Y�p��ن���0�؄���#�7!��rz�.W��"�ñm��	)'��_�^Ԩzڟ <%�󳞰|��7_���ֻ��Ox=��"E�Y�0(�����&o�OCCK�=L����zJ�`,��ԹX�h3������g�C S_�B}���;>�#d��{(�z�P�^?pz�"�J����m���yi��P(0��"�1��C%ǰ��u���Xt�P`]�u8�Ɓ��ǯ���`i�v�k'�Y`N~���5�yQ����T��Z��ܖ8?Z'����o���d�V�X��1�H�f��y�u���nB=Zc"�SY+��D�ZJۭ�j��i�E��E٪	��CJ�����q�u�����*U&��Kʐb���{R��������/yu��.���TA�`:O.d5���n��Z���O2�)gZ��(�C���������������/(6�p�2N�L�!tĀw��c�A��}ݱU���s� T�N��ã=a�g��M+(�HG�) �+�c.T֣ ��Y`0.&��)�[S�3�l��~Di���ĳ����\e��<�e��P��I|b�5 ��{�>�ڱ'l!���b�N��������c!��w�z�eiH���+��<J6�_7S'�$�
�E�Z|���ڌ���YE|��?M� �K�jv�����n�Kcd�Nς� ~9c5�q�F��{��7ϙ�_���t-~2��r��t��<���n~�ʄ����E@㊖�M�T�e����Mu��S�E7�ট��:�P�mc��n���E/v�p��ļ둉�CH� �כ3�˚~F�.�M�
�x�W��쎵���,��r3���X�NW\��N�E�Y�QV�Օ�j_�%���YU�B��n`οf
���i4\`�c�$>�E�6��&$*ς�!��8��=K�5a���IZ�Պe��ž��N�)������.\�l��y�$\R����l(��Q6�9�Ò��s�e�a�H�Jńa��.w鏲�7��ж�:���YRoLP�gw�57�v��y�����)�Jta0=��|Ge� JJ�b;O������F��-{`q!V\�Ul�n�E����G�Vo^��ba~�2R\�!�,ngx�[^-`����EŪ�^�w���;3������^|oDb��?4C����an�H�x7�j�<v�
iA�F{.��`��˻;+A�q�&��@-�;��2������}���7۳�u�Ed|��Kz��C+,WkM}
f�O����Db\K�u�v�U~g�a�3�$�I�/�T�Z�d����*��_�M7�n��<Zވ���mxInM�p%��K.;�Mr�Hj�HM�&���9@es��oZ���kPKWp�Ĉe6T��="�w+�N��x�w&=�����M榈�q��&�z+��U���)��w��W�_Q���C��߆�
=o���>�mzD���Ot�R�����7���*^�q$	S*���@�$�Rܟ쀯��Hꍡ��'�X��Գq
�;����}K&���O��&��-Iϡ����#"e�i&���q�T5����a�j���c����ָ��.�������q=/i��u4.��&�V�W_��ߑ�Mv�ɔ�N\�̃���A��D�x��!� RTF'G/"��܇[hi�	H�K&2�& d��d+Ev=�G��u'HZچL��zY���frTF3��I��%<k�T?k���f6s�����q�σK��`��T`ƫD/�U��#��]�ٹ�G�`�17�����#��F���s?�r6$���t1j~=�3u�F�8,R�b��O�[�S��YJ�tPO�Y�æ�4��⏌��'�����f�,��UM�?������"G�>j����k�/(���j��X�X�	P���,B�r�1�ʝY�"�Yp�;�z�GԯP8RSҸc��;�z�����ѩ���+�gH�62�:�	 8 @�Ɖ-�����'���S:'�"�y�Զ��޼���2Li��k��l��+�JA�^��h����QSut�R��x��㖬�8�87^7�@���h#&;���_(�WB&eQ�^g�a�:��=��(����J�8�Mx2�'��r�}|�1�G���7�KHc�s?�-[c�N7T"BL�H�[�����Q�-7���H��y-�J��u��l߇����f_~jg�D�C�<�$��I�C949���nq���ּ=�Y�6қ�x��/�+32.���8��%�f ;�;�ԶP
~�8�R�v_f`BT���LP�6�W=�W�]����j<G���X�]��p����++��7��"�A����g��^[�x�,��f�h~��X��?7�O���&��W��0Cbyv)ŀU�[�2��������v"9����4�tNxJ�*�oS�$|L�)"�(�����
'r������;xeũ"��:�'��:m��4b(�o����QT���٠���\�|��P5� ,r�:�$�y�o�9?K�������!uO�8���/���?a�3�� ��,�g~V/0��*����l|]��(k�`��=��K2#�v*L6��Z7�3�w҈}�3*�RDW����I�I���[8�f�(,�=!Ws;m�~]!?m$�66�[��.!����ߩ��qrK;BۉvwX1�I������Q�����.��Y��PnpL~A��C��*����bѵ���C��%����s;c�"�zY(��M��]�R�RV��\�,���X���|*k��`xZC#7�+�+0�>B���m"�������c(�5n:����0��-�Nm�����IP��|���0�r�,�2�X�r��K��.�t�xX���D�L{�6��/��f�$��a PoHeyWZ~�����*5�-��W�u�E���3��P�l�D�+���SLs,�ڽ���h������q	6�b{]��bp��4�,<�H;��d���#�\�v��ړa�a�(�����'��i���nL����y�t�� �̃M� �|F���z��x�V�a�+O�����@P�2߽���,8��	Ht' �(�*A��z�.btǃ��j#V:ub^���ʍ�)���s���W��/�B��d�Xy���B���$�Y�9���~�ɋ�?�.�s��Lv�u���4�����2hD�fîHl�`C��:'2���i�x|�����Y<�*�E;x��7Ő>G89���XT:,��Y'��};�|�i�3m��4���p/�%02&�x���($l�(�����!���0-7��E��S�Էf���$�|Fkrцp�m_s�r��85��(d*�[�ѐ�u^���n����#�+�҈��3j8�E��?�Z_!��T@+�{���L���U�Q�#rg����Ƞ@\����m۸�2_E B@Sa�"�����wyʂ����E�Y[�)w K���EUA��c2X���g��(��'Umw�O��D�b@��Xؒ�~�t��F�� ��0F�YȠf؝(�胙AT�8���8�����}�I���|�M�z��Csb�˂�ĝ<o��Ow�^5�p��Eqk߮���o��k�9e��x&m�xo0+��i������X�B�����'�����~1��;-��=���5{1�[;�+�+�F��YW&/B��Vn�3�����m?���Azz�>���V�f�}���j��]�P��	1[�ӣ/�1z��V�U�݈�,�1��21:�g�.7�|��BP��L���ǳ'��/�5r"��3���H^�$vY��$�j�|0�(k�������>$q/D[]��uA��p�H_��k��.D��h핅P���D��9� ͐Ug�X%���ܼ7��y'r8zRMB�օ7Zk�$��N�|��Hmi��Ԩ���T�}z�Z�+��d�a�U�ݻ�
OX�sL&�p֓�Y�$�a�����	r'���(�^�"���O�
G߈��XLXd��Alg��@t7��[CHW�FJnͧ� q�ǚ����t
F�<�0L��T�H~����a-�����Om^��?��q���R�f���Im���8�q�wY;qL����Br0ł�>{o�v?�ؓ�[f�W:��lMs�NSS���%����%�~3��:U���	sU8���H�Ͱp�"��{�ϩ�%LV��}2Ju9�|qO�>M�8����fm,8�8��߳Y3�Tӧ��u>���7|��]pλ�?�^�:�P,@&�,�Rz���G�o��Z�2q,sۀ���t�C�&�:�#J`�s}�&��R�-_�}vNڌ�k<���� J�!����?��	I�>��T��
����EOc��Δ�C�fU�ߌ��z�$��]��g ���ؙ�k�Zt�F���H�s��t����:�bAxqm&��`�b��u-�t�R���A��d����Q��@/�H�x�퍨��{n�'�}4��֬�93��5�j�A���n�E��nd�h��׵f~�ڋ�����tm��9����AQ��LD���N[��Z$@qk0nC�XV��x�h�8�l���w�'�~7��C���eӉ\&)��GR�s�������C<]��wW���ݻp�)�0М�B��r~m���8!�γ����P_!3"&����j'5U���%:�P��D���!���se�_��Ci\V���i����x%9�m�Cl|Mseʉw��Bgl��1{�� 7����3��S����D�ٺP������ 1DY_���EfG���;Oy���a��>v@h��<w�O��&�[��w�įό�c� �l�xqU����x߲O�=띷n�|jZm�HT�9T�Z��5�����ķb�m�Z�C(*��~y���r�89c�'̭vu���]Y��9moq�����I4w��_A�N�������-!yp��h�L,1��+hOt$�G��-��W������EK�a�ae4���3}DWbb_N6j���/;�\6/#xkj��j��Sd�'���Y^��ם�nnK
�y%_��R�9e�1��u��C�l2�҆͕�1�e-2Eu@Q�9��Rڞ�3vr�1R��\�ó-��Ւ��ق����;�t�z��r��\Q}ا�֚�C�l�(7��g�F�y|�^��'fg+�}*�U��<��ل�l��_o�y�4T�6%:G�VX���	���+zY�S����K��^��r����\,Ao�䕌�`1f�~�@�:q"��`Pq�D��ڙ��%o���;5��ۧ<����u��u�X��]��7*}�� �@�<�v�`��o���{Y��r����Sē���H�h/0��!�3�F��=���s
�b	�nԂ`'/��r8�i<"\/DTsm�����{)D�����lJ�Qn�`m[ܦ�0�@�� ���T�����m�@���7��2�Ě}P�����2������oB���$���?Wa��t�o���d�4��G ��#s��L��g�����C~��xx�ש�Sgo��4�u��E�4m<V�����v�HϏ:P�1��FKي!S�au�����򳣘����0Wֆ�w���rN!Z�R�(Eӷ 5D���I5c��ns=�kYqh%�j}��SiM�I'���h�(X�g�4���44�E��;��}�q�������c�|��R�u����z�9��fe�5y��=0V���0�ٺw�tjfU�1�=��1<�����% ��C���E3��S���Zj�G�ȵ;�W�.�?m��<�f�P@3g�k]j�Ts�Cw.9b�j��d-�~>�|,uy<��^ټ/��Z�w߯��з�:���;��q��L���%9�%�@aZ�h���d�n̅��g�"uzv2x�	��g��'P��N�'a��O���Yw��������(z���Ǜ޲WP�V�TeW(����-���u�*:�M�]��g�n۱�#�}�يS�
�b��d���s;��قWYQ�.��= �=ixR�X.Ih��dYΐ!�m`�Ȱ�]�rW&���@[��]�,�J�o�#d�Y�Y�B��2Ury�\�-$Va��2��U�l��'�>^�H�+@G�+�J6��rߡ��Z��0���@p�p���躁(���&bv��M~��xn0Ds����BG��2	 ��{�'���i�|m|!9X?x wR��k��C}���;k��E�X��ɫ�4z9L�$���/���1��$���f���|^��[B�OU�$�+��?Y�1���p`�Z(1�ʰ���G\f���x�Jd�"�&����L�]����o�����T�J���T��V��;��Q�k6}�=�ׯ~N�����ލ���V"�:!m���t� ���7W�\`p��C()و��6��.�����jY_M0atil�=�|1�����N��o���q6�A�Sm��@E��k�C����.��&=P|V��/�B�0/�vb1��R���L6J���E�Ff���>㮺�]e�EC��i?_?���{Z�_S�)+k��2�
��Ӡ楐����M��3g��֨�X�����4�
	r�-V�R�.��#��C�'��%�흯���������B���z���?t��,�e�6(�K��1*��q��p%��+;��J�MF��B}�+���kE�����ʐav��mY#��;ivzwQu�е݈���(�1�vTp!#�@h�j��<vz�L��k
͋���	��Ա�d���4�G��1�����s�5���#�M�l&ԩ�u��"�G�r�%�g��y��t�.�ּ#��p�r럳�@��G1�e�h��l��a*wq�`F,
i��{$��)M�0����-�����]�z�p͢C��y)�I� �y�-.;�{��l�d�<5��>X���1��BoKӶ�<7�����)DjAh��Ꮏs�6�7�Y��4]�r7�f�JLa�h�һ����X
��1|Y�=�Ziv^�<;-aL�~��)R "�lo�w��R��~�s-�p%�<_P.a�#��E�
�P�>h��?V�|��*iW�!���'�R>��J�F��Up)P��������;��O�O!B�0�'Q�WXڽ�s(P�� �����a��<y���qAe�o�s��D��xFBߌ]�.i�+�h���%�z]؄����҂�H���N��� ���4�A0�n����{#���i�s��S�uN��������z��!���)R����I7��WኔqM\��*5�Ȗ�C��5�EZ����Y����p�{J�y��� ]v'�:b3|Tڦ�<����f��r[��ځj�y��T:�f��a��NK֬ŕ��U�@��IR�2�������5���Q=ܼ���!�>����:���s��V�ۥ���:�`;���@$֐W4�˪�hm�5��ç���H��QX�(�����N��a�zC�e�pA�Zb-�Eұ�cj����Ou��FM!�}�^ n�w����D�T��I��a��H����U�1g��կ'݌^jܮ����q���\����V�y�)ӡ:�E�>�4��W�1�!;�o1������w'��U���j�e"s���d	gr�ͨ�}�� ��)l�?�ﭡ�If�?�h3�2�zj��[Q��y���A,(OҀ����h�$9�H��I�lN�RSB�|2�&��<�p9ɱؤ�NQY��K�* �����=���>�U��(�(E:ۊ E#Y���!OPB���P����S<������N+q(��5�@�	Ou��H����ԑPP�:���;��(�\�i�d��R.����#2
��]�uN��9[@n��;����iW4����+�	�M������VO#Q�k�5O����q�\d�Y˩ϭ�]^�%�+�9��Q�Mx�&����jXW��졧��(2�O�eԠ�q��W-3��]k5.�)���`w��4�k2vO�[�M�k�Fk�{��m��-���q�;�������z��6I?�=�=�A��v3��WF��yh�߉|��)tAOw�Ѓ��+^D�c���nֿ�c��Gv�'�=�P�tR�տҜ"�� ��/�kW��HP���ԛB%�؈x���)"_|��"�o��{s,��W��+�֧9a�Qxc��3�+��8gn��;�K;Ygk[�&gEvN��g.�I ��ΜN2�t�;� �	�$>^1�a� 2ʳ�ul&%��"��~�5���hX�oJ�{L�s��Vc7�󺠕�]+V�pי4� �ܞ?� �ӄ�^-pz1]�'���� g�ps�ASl@c�A:Β�d�{�c�5]�Ë���y�cD��[�K}��9��W��v�0�hW�f2sj:Os��#� S�g�VA��no��()K�bB�0T�]c��Ɲ��Ow.����&E�JW�����)�Y��Z�0���xr�n{����|I�hRtM�+���4g�7�!6�s4�WvW��YI�Z=�:N��4.�D4�ȅH�z�$�RnY�Zp9pBN�N���@��S������ո�wE��* E	xFH�Р�=�3���Fs�e ?_?���"�p����(�_�C�R�� 6��o��Q>��Zs_��e�#bGJ���Zw�O��;ƚqQ���@�!	%t�`�_����@����B!��ca�0���_��*�K�My�}�t-��h8�s~L�gH�;h����ܮ�I
�h7e}�5*'�����光��`�˺�lYh�bg�Z�å����Uz�i`�ur���X�v\]@���
KX�tQI(a�>=$G.���!ft|Vhl�e��W������'����F}qx<f2|dp
��J�s���y^��>�wW���Aq�`m�ϱӴ'�J�`ב9��2�&�G�5<� l�y�/����,6E@�|N�v�W	�K0����;��7n����dud00`�>,?����h%�m �DM�9`�+o~���&����	vx)����PjR�8>���%�t�t�r���筨��<��d�O�$]��C��6M����~�t+_�1oM`�	s�XN��C��{��F��r��B ��K��S5�A�;"���_��Ԩ^�y@�Q��Jΰ�>�e
�g�vw-RH��3&Ɇ��`�
Il���é_�9��"(�B!�ivЁf��s���dxҵ2�$���Ǒ�j5 �B��G�W���m�.�F�؇��������N��� ZVBa���;hv�b��f�F����+�O����^�ьn�>|B�]��lq��0y��?3�$���`�Ƚ������"M����`����5�"7a�T�����8�7����8��eP
�)�AP�s_��kSJ����M�]��k�l�Wq�E4���=A�� 8,n;�w���f�8�$�2��������M �[l�\��v�,��I�xbH!/+i;����OPx�?��+O+'�
�c�ݩ��B�.*`'aA9`���b
�bQG�����F2���TT���@U�T�! �s�2��W��أ���e��ŋ��%�ZT]���|�MG�P�'��Ӣf�x������e�8�/�l8��*|����/��|��f����,�6"w!���sZ�6��(Rj@V۵:�t���*Vj������g��z`�%~�a����
w h�w�0�>T�*:�dQٶ�Xu ;o�e.���h�P��i���8�m���N����3IL�{�g���2筿Y	T���e'I~�G4 �#��y�dy����9�:�#�͌���:C����J<���T�ߡ�g���=z��R+ٙ�׿�P���b���q��+�#��
�̵[�����[�.���ps�Bd�%�~��ܘ�e�"�sNβ��H,�i{�Y�F�]���^���g5�J�o[h���>�J�6¿r_��1�jtJW��|\�}'	B_�-����:��[�Yϕ��6�t�N:8�$��~�x��.F�d;�L�>��Ԙ�&�:��"���K��>r*�F�U/�p2���P��/�z�M^��J����Eq��8�y���Y�1[u�7����;Ik�	J[�-���w�1!������;=cS��/ܡf����ʶ�&h�j����Ɉӄ['�$���$��4$�O�@8y��w[�6�!�%��]�g�F3�l��ۦ�7�D��x�N��O�9	�z��e8�����2�Ȟn�'����Ǒ-۱b��3^�߄� ����E��A�,���O��lZ���sg��
���i�W�x �
�)�#$8V2ïjp��x&�
��o�L��w=I�v7�{��c�����{��-Q��2Qo^oIk�bU�3ߠe�P��ÅP�wR\ჶ�Xh/*���Z�N��h�#?��E��A�Պ�˲#��0,��t*�NY&a���].�k��k�B:�w*K2�esf}����	� ?7��|���7́w��ڎ����ouJ ��*���:#�,��]|��f��4u�ǚ%�_�����,��黪27�r�"�/E��/S$���ϭDm�,���(C;zQ�ӅkXu��ށ6Q�l�đ�KF���;�/���i����|v�r*���@��b���`��e�E2���<���:����H̶@ ۰���HS�qrM�Q��7��_�����N,�T��±��������m��I(�5�W��·��ޓ{��+�����1�P�1�:5e�h����~��	F3z�$1�z��E)礇1���x�"�]2����l�U
�s5�{k$�5�X���?��L�k��kG�O�0e~�Odzb�^['��)�\�h6{��� ��?�Um'3/jN��r�����t�m�K�K�57��A:��^S f�)���{Ƶ��5rx^�~6䠵�!v�}i)<��9ɱw��+�<���L������wS�c*�'ovO5� ���MM�"�po�O���	��rFQ�hAku8�ؕa-�ਊ���Sq0A�R�%Ox�7����OM��ȹ����y�L2�S���n\�����<`��@1����N�g�j�\�Oc�#�]�b���	L��X$�����0,eV'^w:�黭��'����n��@6i���F�����\r�㴒%�~*5'/L���HiF��E(H�s�3a���	�(^�C��"ٚ���ۯ6��C�|��<@���;�ңƻB1���?gz��D85e�x�f{�,��2y����(��G!J���G�)ȊC��G�~�9�����үs�9�Q.�������n�)<P
�X��݀v�m{�-�c^*uQ���VeA�%�\�ɛC:OW�	fB���@�����8+���/iAl�IR��#�����O�;����Cs��-zT��V7`B�/���C���2������]JX�,S0+o-��H��8$��"%0F�sed�.V�,�c�h?��IU:�&;�v�w,���\#��I��pUvV�0���t�"�_?��ō��r�	�ȏ�Ug9�@#���M��Z}J(��ac�;��b�!<#���
�+m��+�p�Մj'��ò>O����x��D ���X?3�t' 'F��V�OW5�ā7m?��u+��@���<Ja+�h��}��g$y�P��
_X<�o���1���H�a� �1� 5Q��)�u�CלR��v@u'�����A*���H[4��}!za����c��Yq�f����D���q^�'�D46�л�8