��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4dտf+����ؐ��7&Qa�z���m�ࠧ��3`����8s�=L��4�S���J�7�h��J�3�_�������p�t_3�ѹY��S�!����_-)�_�3s&zf�2<��h\V==q�/��Ke�AHk�s�zmE�C&�k��{�jc*ue�1�������PѤ��w^�&��{���w=du�@�S�?`�X���aN93I&���f���O"h���vu�DK1 ��7�Q| moS������L4&�~&i���v���/x�׶��N�U�_�����!e��d��]l�8�7"J���Q�����F��/tU,g'�X 6ϜJ֑y5�SP���G��������ǳ4K�q�#_�֚0]�,�ד�	��Z ��)ϒ��Q�إ�w�?�ڮ�+>fx��x��$A���� �TDc�m׆̯T�!���`�� ���c���0������	�6�+�0Bw:�h�&�ڒ4����]�����24Ɩ��t=M�0²#��� l'<�1dW�B~��U��2V��p�"���q�Uܢ؛�ۆ��tUK�n��Rf�iq1�=�v a8�H�G��M}e)e64%��-C�`7���H<&E��<7��aB�q3�w��z`����v��+���\U8Q�.��$Iȃz����9�y��f*W�&�YHy�@����x�fܽG[W_�B%Y�fɏ�0�#%��'���)����(ZN�ł5tPnQ��d{a<�� ��k�m��Dv�\.��۷�.8�{S)Ǘ.y�P��cc�l����5����d2�vw-з�-/C��d�u5�(z�D5V^	.F��b��8���l�T���E������R�d%0=���`�x���O⍫Í4LH�(!�Ar,�r�3�z�3����*�_���R���G�I���J��E1�l\s��`�����[°�r��P��K�/&>��k�����t(pA����,%��g�ni].�;k?���-T+7Rό&9
R�k�\%�-��V֝/��0���nz��&�v��50B`�����8-3��o��h����T'���&0����9 P��Rq҅���1�[VNe%Tk���~-�ۛ�`A`v:W�������
Ϛh�x�H�uﳘ���$m.ۖ�K�k1+wt��+3�_��!���i\��1U���>���翨�G��`TZ��i e�.4����o�c�ݮ�`##A�2k.4��S�֌�/A�ދa.},Ȕ���)���������^<f@C�ձa{͘����ͅ*��ψ�k��D�Pa>�Z����^�c*�&7��z�|v��B��9k�PO�AVu�uTг���ZY�E�򙈾��f^����>��Щ��SX�`AN-��!q��w��M#B���*�$h�eo:��iGT���F�\u��u��Tcu�0>�0��ED���Ћ7�K��Jԕ�f<�G�HA#jwK�^��� aI�=��sҒ�p�i ߌB���1g{�+�`�r4	����`y] Qk���=���2�;\�,C������-�փ�,j43�B�2%���l �&,�|F�Jxg>}���{���H��M����o�53����b;�*R �l��b,QU���
\��w~ ~\�cc����E��Z	�k&l�uk��~tyD��U⽐a���Yf�g鿩i�L����-��>l�f)�/N��!���Tӹ-��F��~c��Qz۸�	B���{,��~!��>8�ʶAR���N�A��T�kJfN��#%���K�e�l$����D�.�����8��<�>���F�w�J��CC�:߆r�H�X����� v�f8|yp�t�II�£i���ڿ���g%�:�XP������|�W����%c�����.�F<d:��Q��hd&�U$p� o,�i��,	оTX�, c쨾h.���Z3sa.�$�k!��?�ÔZ��J>��qvI�Z�.fi�E'���v�y���<�n��, #w.iˈ�Sn:�B㕘bQJu��Od�UG���Q;r��v�I��PFs��2�g���"�?l�e5�g��mb�,72��Yh�/7ȍ�WX"+5��pK��n���aN�^	�i�BG��E7�Z+�T�/uw��2�e?�ᑸ|�i�ɝ��<����k{J�����vA��k����ߴ�Zs*�6�͖���u�'v���ŖN��Y�F1�]' ��A��ߕ�a��+z��r����L4�֥��y�2�$=����%"�.��C&�Gf��^*O蠜,�A�`��*����[9���i<.�zy���yKY�&S���>�]��t	������Ҕ�St#������۹���L�x=�]Ԣ���}�A��b��m.H���N�P'0u�*���d<qع�f�"�T�-���2��P�Ef⟄�b���\�,�w~���}��(�F��4y�j)O�`D7�������yz%xx��qΊ�|yp�����u��,(]�p�O��O��f����Վ��\��bu"Έqr�7un6�'%c�I#���m������ݿ���XSb[�B�OV���"y
��-˜���VXȯr\o� ��ai'��(z�{!�"uL�9�,,�����vp=sRFo�Ճ [pp�����{Z�+��@�W�g�!2w���W�3 �j[�na��Az!�t/#_������?�i8q�[���_I�vI��J�L��}��[}U�	g��r"��B���{�I�9l���4&'�3�w��oa0|T�����r��a�3�.���q�I����~\k������һ�q<@�^���.]��k��Ē̼��lv��|�N2���Լ"2SG�2� R��m!�3I�H���Rj��	u�UU/ ��{�CZ0l{�YcΗޢ;�x@0G����+D�L�l�sڃ�Z��F�o&Cq#�?l��|��28M��7>K�����G�Q16[��M�J���͊]��G��ҊQ�	�%���ME��AO����Z�$L9d�6
i=CHH�ǀg�rJ��.�ށIa����,YR�פ�{��N�p���Ѥ`��	"��]�N5���
����$s-�K��"�XC�=
H��e.����e����B��`�_�/���6�l3m�yɝ��ȉGIlG���F�"Y����I��"h�yN��I��������[x�݀�[*��>pY������T_p�1nJ-*3M+�І�iOU%C�gwS{=�td��_*�o����{����~o���q���#���4c�E���K�:�����_qG�-z��Qa�9IďN�zp�0�`�L:���;����#���*�31&F���5RsЖv�J(Ig��G�Z���m|,F�e�tqÌ�Q� T��ox%<�o:G	Ţ��s��%���h.���R
�o7��AJ=/�{�Я��*�)����!1db�t����<�� �_1k�� ���Q�����K"��B�ѴC����4W��5&�9^��pF��H{bP9֭�O�1���X����q?ڦ6H��97�z$�^��_�{���&p��Y����:ݺv�;�@Mޚ���:㢿�83�.J(��'a|/Y���3�B�) @���`8�i��`=�}�����6	���i_���V�D-�dc���۲��"��8�]�<�����{�tl���`��u�1f�>(�Us��K�ܪ����Éy�v������2�g�����II�@�Cc��ح�2(�k��r�U�V�8n���p���i�^@4����fz��a�U��L�:�0�F�^t���%�<��Ƀ�juO���_���{�R�
�JY}5��������+<����&���ڇ��A#O4w���gPm�R!Z0�\훍ۤ-����͈�;�B�ُ�u��/P-!.6r�ȏ�`-sjJ�����d��Ks\ё,v���&� ��%��t�!�
�əO��9gg06�<�wR�9��J#�{���
鼡S���]<u��AvǬ��8��,��v@{N�y��T���V��\ NY��E
�Y�-�L>P���m�j�Oq��.9v�����1��2���#b�k��+�58?*�7��B�Y�*�:e=n�;�4��u0�3F��\�`.��0��xu�Z��r�����-��R�h�ʇ�v��X����w�lA�D6�&�^��2f��e�~�h�=�}L\�k�����.���ъ-�̄��I���w�D��}E�S�ݞ.������f�Z��;�;�pg 9��#"����d4�Ω$��y�!N�c�L
���_�F[.���4�� [8�-�Xu����߅#�}ӑ�uI$�SI��4͑��8�4�$\ܙm�;\I��;���&fS��z	����Vw�)��p��LH�9�ZJ5l?[.��u�(|����G�P�����"Y�F���%[�=A�)p�~_qX��Z�=l��V-�D14o�-���B����1�5�w'pa�%|���.�h�?�J�z� �2�(�˦9��g���q�3��?WEsVײַ,tW~۔B�%�

�o�X`E(�A�?��!|�p�:�֭Epv���
!�؃�>��xh�������0���N%$p����$�YM�DT��������]4M�A�M�-���ߟSe��I�ofQ5Z��u��0��7L75��R�