��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8SjfSު�U�.Փ�"o���Ol>�g�t��"��+_k-vz����;@�[k"W�3B�|���m�xbZ ����="�8 ކ��Wὣ�3��'��.7 /�ȆIc�Z���ja`�p�׭jO��F�����L�m�m(L��=��+��ڇ;��P`.#��١K�'|��
�Ut��e����Gu�J�#t�|aC��v���+�+�=/�ĕu7���x�_n+��{�s�����E/{�Z�	��-���m?Dc��p��@R�1�m���KBy:�sCC�?ԍ��cV	��(�(�ߺ��b{�Թ2�]���j�<�ಌ��%�q����(���!�%]����u��[�2��gFc��5�!6���qI�}����2�K�(�uS���0a���Y-`A�t8��t	%�؞f�H
SAqt�CD,N�YL\�t⹘k��0�[{,��-T�}`�ns�Rc�����L^��ڊ 2�=��uJ��^��O��>E&4�I����X/�L�6��l�#�Ж�T�'�od9捠���O%�Ԍl�)gb_ՌOw�j����J�xy �PϋR%��<��n�ߧ����*x�_@P#Rr��cx��9�~Gd\_���hO4x��; aچ��+wW��	�(�Im6�1f��l<�.ț8-�ȗC�}uI=�ȭ�ov�{"�3 �I�k����[Wy+_�.z�D�����0UŃj*��� Ay���SM_���l���o�0�a�Ô~[1�S�F�6ƙ��?���ř�1[I���8��vG��	xG̬�FiIĺ�[;A8��qV.}����Vn[��B����1��m�4�����[��H��S�:���"GI��PM�2�j�Ey�#L:	�;#���ԉ��&S��W=> 1 z'�h�	|k��S)R��w"G��A� ܸ�/j;KmA�R�AFy�<�%	��M�!x�?B@w�Q�ޣ��.e?��*�e��E~F��+�ePW_ΐ$X5����QYcT���;sk��AO���2IL���؟�q,����2RY0D����M��M�����
*�:лs�;k6�wl	ܸ(�O$���D���p@�� 2:���n\�W({%Pw��G�Ԇ�L�Z�#����ٽ�s:|��'�f����9L��^L>/�s��u�T��W���]��J�Ap��V�hC��f�0��<$y4X��rO&�@;�EH�˸�?NM|��ҘK#��9.B��YWi
���N�c�>�n����Ȓ�L���s�t���T��	1.`�!�һYA2z��/�VYi���jG)C
hn�j�2YF�B���x*!>b��x���) ���7����8��H��{/ƹ��V��O����|D�ۢ�U�?[��������������IH�'�o ����V�LR�A(�B��)N�^�Z}6Oǃ��F��1p$»�ھ+�������b�܃��]��'�����?I��|���gG�zḠ>Ņ3� %RV���J�1a���7��rt���4���@��S����@�����K�T���l���QH�,�#��2vG�{=�s�Z��S�z	����7�6�w:�|;�M��	-�ae����ߞ�L�p�����3��f��1v�X��RN�(�v5&H$	���~����/rf헭z���J !�	����t�Q���p;����L�q�����COG3ǜr&��$0/�J���Ru�X��ǂ�\^�F���!��ýΠ�5�<�1�>�<�D�W^��1�P<��B!&���Fu&bb�D������Ы��f�^�~���*�Y����Y�
'T������J�{&�� �0-�1��}�ЯCK�BG-��OZ�&����y+��Xܕ���r̵tM���o=����t�/Z�`ʫg��������i%k�����%s�#�:vY $�SV~`�@84���9���~v�t�u�|� ���r��~V���A�5o�]D{f�h��)ʣ2�RP�.�݆�n�^�A0�W�Xh�8 �O�*�}�W��h�P�@Z�rs�؍tW'�����5
<�Ԥcd{#�.F��W;�(n>�Ʒ�3Mb��V������e<_�l��H#u"`���$9�.���@��ZDM�W�i��D]���F��ֈu����G�$cHH������Ѵ Z���s��Rbe����3Ff��3Z�*�~3�錷1�s�3���a]��z�/�d��@�^~��C~��->PbK�n,�Qs��N-t��K9�x*�y��<k�vz(����=5�A#s�V�PlZO,����NB� �DtO�a ��G��Or�Eu�;�t��H��ZTi*�.�-�B��v�p�TݖqK��_ɿ@^�?I���)��R���P�u�E���^�)Ey��K7Ґ�Q#�R۪Z�
⬌����ꝅ�/�`:�
���	7�t�L�9�>&��k��)��Wz%��fu���=�D��k��o�����'��V
Z��'�򠨈��e����ަG�Л!���#�����@��$��Q���s(��� �DZ�x!�h�6 ���a��<G����-������a�09ǒ7K��_[�h��\^�U���J<M�>�No��!���MTj�M�?�vH�Rõ�f���=�(v]���s3r�,A銅����TZ�"*�������zچ:�Zn�,�]�h4�-���x�Uڛ�5a���Hf���;�s��R��x
Fo������_�XP���B�Rq7B6����lH�������� ���a�D(FZ�����H�i�93	l��%^9��E�qV�^Z. ߆_�J���pV`�����}�3�A�W�@��ߒ�(P(���#F7����T"�"-�p��c����غ-* ��Z�]����D���qd��7m�B��,8z ά��W=CG���U�#��l�-�"tB;J�%��B+���
��_���_��4v���^N^��.�a���i��4����CBɃ�e���V �����������J���V��bd���mt��玈�l 
���0�����y�7�>�M��(�
�Tr�slTz�h��R��d�nM�6�<:�ȒX��ٹ��$���2P�0|
"��'L�D@B$��C���g�F|�:#JTW��Q�,7�&Y�.|rf�ܙm�(�'$xK��}�c�q��hYBy���<�ƂyZ.
��l3X.�߯�L��:�`����t<!Y�I�@J�4��h�7���p�7��!X��� ·��D�Z/5Wo���r���^�(��=K��>�s/~�#� �5QP�f7��C Q;�勶?0?��)����b��<7oh+�0��*V���3�kZ��}����Q%M�k�:*��V&�Q'���̌�z
����mk1&s�r��>sl���p�𱈇��)��~����Q��$���9Y���T�8���9۸�{A�.$�"�zt�<co:P���p�;���p�Y��ISp�e885j^a�s*/I��[l�;9�h���d�c�n�D�ܵ	c|����d�(��[�G���&i3�Q��:%��7��o��bU�0�[��=��d&m�{
'�s�af�"���}�x~���D1 \�0<�Ϡ��4�y�"嗄����=��H%BJ��%#���aZfo���do�l��9?^�4c�]�Y��E��c{e��:�Y
Sö:�4��\�a������^��̰*��CTі�C��{P�.]	���B0�3�3C�fc�<�|B��}��p#?�ޛ�����Vć8�����l&���n���Sڶ�E��	����T�1���gN��g�N��dI�BN��w��^]ZD�:fi�=Y��� u#���~S�7V}j��9�f0����:�)yL�@2ƈ��F��{�N�dv��h8rC"��l/�)JcJ�dfVZk3Hr���~��<�wxxD���0<g��w<��I=M����:�;��)���:9)u֨�_�f)n��Q��_?�-�w����M9��b�|\o�*˻ps|��|n󼑂��jXi�S��B/��'����׿�'���M����q�]�rmF:Ë���j�z�	��c�7/<_Kstc=�b�z_+�X/��p�7=�7�<nuf,���K���
je�C�͌�|��o�+�6��1r���U�@�[��i��/4�d{su��I����x�:�~oc/��?%������k�H��,5���$��L|.�Y~��\ZT+ �b>�"T�q�3���]c�N^�,#��]���2I7s����D�}�p��������x�Cz4�q,�����E�\��ɼd}�_k�"q���������'����\NҚ*<���Z���x����R[��p*"�TN�)C*��N� �ϖOIL~j	絒���sHn�ȝ��W_:��G���1pE?];y'2�;n'�&���;�R d����tt*|��~�)b۲2��<�m���5u�:��%�؀?�&��IP�}����8����$F�u�	C)챁.A0�i`N�~���B�IpR��%�ɩd���^5.�u������HE�I$�$�WH��W0���L�����wޅ_/�l�ynW��8��إ��X\Wk*��������7^�CDX���f��Wbߢ�)��i�&�i����R��;^w�������"h��-Z��v�=��8����Rj���n[<M����53�Z
r����YǢ�z������)IK*��c�ZN�]�^�G4į��l��I抍�
��`p���_q�P�wF:���^�+cqjsμv�-��Avʛ�l�= ��$"x')< x���f(I�t7���^��k>��
�ߚ�39Y#y���*���`*T uf`"��am\!�w����N~�y:�C8�vS>a�B�����@������(�Oܑ���^&���o|�Y<DwM�)Z*Q!f����4I�F�8�v�D썆�=/\���?PND��i��A�'���8�_L=7h���}�v�z�����"��>��xW�>��"��( ��P�
�
�eq�՚�!�ˋ�f{fA6fS�N�_|:OJ��}�k+�Z�wv4@�H�����0|���[w��@%	���AƘ�kأA0�W�Vث=��J���M3m�y�Z bV��-S=q%蚝޸��v#Xt\����Y�� �"HЛ�QZ���*/Z[w�P����i��Y�d��r�2x���q�{�ZR���7&c��5�I�&n8�|��hN~�#"n������� ��(kե��$���l�?��s_}�)��cB"�ǎ��"�E!)���S�Q�7UZXe��Oy}��4�^ W�=�l���RB}($�m�Ǹ��U�Ǌ�|m--��RH��as�����h��3���&	{�!.:	5�X�Df_}�AG�Hh���q9a�P�	�^j��s ��s��z��a9�B�ftu`�|�Vff���ZP�w���H�^�_���uk�u��N]�m���1f�ұ�.�/�%��L��͚�V��{2[�+ɝ_�n�S��p��� y�YK58�~�T��D���ʝj��r���fq�h���1+l;�����pϢ�A� {�=,q�hi1���Aw?P0:�"��P�7�BT\���ဳ�Q�n�=�i�}�P���aVnq �`m���˓��	��|�H~� ��>�UE�6��
o��uH>�chdw�*�o=Jp��
;�o.Ng{��S[w9��������\����h%��=��m�n{�G�+1]��������7u��hG����nc�q�z�4q>��P_�����2ڠ���z����-
<�E�uvD>O�y��j@��C/�(:d
|���x:�V�Y�e�Y�ܵ�:��6����i&��L@y��h�ݒt7d@ W��֠m�	~���p��B�?ݝ"8��[ *�[m�U섣�vDHr��
��ƯS*}�ryR{�o�-͘�(���h�f4Ӊ��A�K5S�=!�n��'ib�*KX�
�P��<�5twR���C?rHQu϶��F��)p_C�X4^+��pr�,tx>u��򝳞*gXC�Q��ͻC���?�پ*�\S�}� �i�����O��8��5-�,�2![��~���t0.լ,b�@UU�쩋�z�X1B�Q��{��$��n����j�@�u�e���T�[��=F@z���c�W��X[d���o����VH��47�_p~#�$�x����'�´�T��?��k�{4
�o�r��
fPt&�c���I	㰟OYp����o�p��aLEUP�N�)J�l��!�G�9,��?�~H�pW�_;��{E��$���w��,���`�B}Lκఖ��Ǘ@�Ƣ�]#�p��|:� ���@�:;t��X^�(N���Jk����� ���<
P����;^��3�'�6Ǔ
����V�R�]&Aw_7���I�k��n�UM�����U	+ꥋ��$hOH���q?��CN���>nu��v^�XI�(����
��\d��~�p�F	�`��������$	C���/�U"i� �E�y?P©�M.H�;�Nf��m}Y��S_	wq�a+|e��J�"���v���&!{��iVo����[����S6ʻ/-��M�AK��ͦ�&:/|�Y3�u����JK՚��Qц�H+}EGY¥�x��M���m)^9��Ł��0߀�����������l�k0_^��4�}>�j�_d"��D	��\��"Q��M��*�ԦmD�+h�xy،�1�ex%9rGt>�0I]=��HM��'�(-��'%���v���n3 ��~ʘ]蝄�Qsoa��[�9�T�S������V�j_�v�M�1�1xoƸI�k�A�0I�$�Rp�s�r[#�WK8�܍�b��F��^�S�Ųz�7��p�Ժ����ʲ�'�כ�����w���C���,�4ϙɆv($���W(���</�U3�\���(�\����m�nMs��]ʁ8��=LjօUiy7S��3��(�ߓSq�dKםN+0b_���_+��AP5J_5���@&�oI�F�|�6o|j�;��xT̉����rI,;3����-J��bf�}^�Qm�Z�F�h�a�U�9����l����@��g�b�ѯ6<��5�ʸ�1V���p�?I���}�0$D�%�R�}�1�b���[��#n���E���,� �1S 	mOd��C�y
�.�O?׀ �҅�o|�һ�ji./R"�\/y�7X�����c-����Z�Pqڳ�*:P�L�U7s�h�y>?��5츕�I�*��@u�Y�=Hv#�1�%�7u��"�ؖў.���Ǳ�����=@�J{(�Յ#�A�#��q���["#�H�IW<�6Aת���MsmO�
���p�x���rf�hlD���_���x�8�nqBx��N[���/�,N��fL��G�}�ش<�u��$�#u/^E��{#a�?���X=�,[V~T ��&ۗ�Krf�审}���4)E���[��_��V��{e��Vˉ���;��W���8?��m�H@~���-x0�����݅s�r�,����{�}���k���2�:Ҿ�8���;�p8S/���W���9'&�,m���㑮%I�!������%B���f��_� av�#.-��4�q�y��V��D-���3wUq����FC/Ǚ��saj���]S�"6\�T%/�-DA���w�[�_~��ab�.lߩEc@m�Ϩ%���3��I������edPQ�sᢥ�z�p�q^�耻D�up���[���b����j!?��l��a��Z���1��aq�5������|�TP&:/%��*���9VC�p$��prlw�Q>42?Qʙ �j��y��e��f�,�+L5������Y�g#:A�(�4��՗B���D�z��N�����5��H2`�d*�9q7:�go�@17��IJ�������n���o��M H�q��U��4�o>�.��;�M�Re���I�I�G�!!O����
_�L�p\i�T��;�ۺ�/�S���,. 8�>c0ML%@̒Y�2$�w�,p=V�1[z��>e2�H�20=�%hf�&8��CZ9��Q�E�/��$e�Pzj"�n~=<�d1F#�Σ�)�8�� v�Zu����GK�R�W���-WSF|�]�mC�=�swZ�u�#���@��.��Rrw�Y�|Eh���=��4���^Q�����w�J7l��2/���A�ps����l��La�B��Ҟh(���R�<�S��%7�	�#�Z�5�0��1jW�{�'�@`n�%����d$�����3>�9�l��; |��qJ�O�<z<B�~��c�ζ�-��	��#������|�U��DI,K��&$׹�T���L��#���[7���0�a�I��[�7��Lϓ�_����h<���r��E�ϭC�m+��+`r� 2�҂��hIG*�>׀��pA��K8��sbU�!�7��Vܽ�#R2���}cMf%Ҭ<+� Ƿq��5��x���n�#�ns�L����Մl�=L�}��RQ��~J93I�7e��3}F�M��a�ѝ�1J�
��X���V�&��ԺP�u����	�t\.DewÅ1P(G�s:�c1�w��Թ����2%M�ծ�y�H���ȡ��޴���Ź��Wr;��ci�ȷ�����j<�+��יFX�C��g/�Kr�!�&�"��v	���R�
�V#�Ӹ�78���??���%c�b�������Tt��E�LL��2�U�꛸����m�D}2��W�̨j;��}����B3�N-&8�tt�/v���DR%�djvAN�Ԥ<�M1��3¬��PI��/Ң`��)|���!u9?i�Ҧ��3�V=��ml��.�W�bz�(��h�lőϋ�zX��(��Qī���T�	F�J���7D^�dm\$+���3>��Z#2�Fz9-����)֘v��T�pNP~9��z�uN�53�r!��%l�'����
@�E�꘥��2	]h~�0�%^� �L4�87�{�w&�C�j(Q�_ۗ����8q'�
���oɛu.o7���ă���Zw�"3�$bš���L�Ƙ��kgs���:/Z�=����C��#%��w���� �b��(!�6O·�!p���i%��e�ad��ڎ�?�		^gw�0M#����f��
4fk�P���,�P&]��Q���޳��c��i�.-��(Q�b�&mU�8�Z�ˉ��Ș
��1��X�Z�w]���q�:� p�y��n�K�d��g\���~�0�W���bL�(�`ZDf�)t��]� qĳ�R ���[�1ɚ�3��I�c��G���l@�|ƉA��ՙRC��En����	�z
dq����;6��^v@B~&��E �Y �󱁹���DtxБR�vػ@�~[�*��C;��ڛ^���%�I�rvJ��V�V@Z�=��k�:�l6U$��0癐%����\�^�~����� ^&��Ym�N�A<��J��v��G�-
���Q@�۳8�+<��N>rI�Q�K��2��Bl�(l�3�˿;[R�]p{0u~�/��Y��Fx7L����s�S�Q�iVP;sV�@�؀�h�+%�D�k���.�
B���s�����Q����D��V��f>��=Jg��1����tSUU[��Z�����w�h�OR��h���g�epXs;���_xC�C�"�e�F���$������^˚����3��n��:5r��T����7�<;fG��e�ʡI#̬鿶Z�{� �_2X4���5X��xG��p����p������J�XSj��;^����ReT�C� �� ������sfkha������������K�)R襤�n档�"�r9
��{�_bM��Ꝙ:�{a�*(d�/{�X�v��䫿ua�i9R85����Hh��90��y�L�@���٧&���B��;#y�4�ϙ���uLK/ϖ�FS�F��}_F��$>������+�Q�f�6�]'?̠ƭ#�F֨��)�Y�@�C{�;�����o*��p���<}���mi����R�=�1�W�E��~	L'gܭ~�V4+��ؙ�<C���C�])hJ7�r|Ҷ��Fc"���i��������=�AZ}%mgv��_�&	�� �����ٰ��P��ʵc��&�)8���{K i�:C��l/�� ���{t��XDn�b<�����jX�r~ݢ�Oƶ6���B�2��$~iބ��F��3l��j�p���L�J�F��ZzI,%�jT�OZ�)n�y�����������b{Fj���8��-p��ã��S�d�2�E��������%|`0��y�(3��L�b�Y8u�9��(��wק	&_&5�F4"��Z�?Ϩ,ӕƶ��*� �3/_��t4��9j�rq���,k`��Py� +ͬ�t�&��Bi
C1nra�I���se�,���;&-����C<�S'07�-�yr4�v����l�� ^�-EE_1����S�:&�H�?]$s�� �T@?L�4�k7� w� eUl�vT�.�N9Z�A�"��5I8b)�X6ă�������B\��.}�%���GTĞ��Y�2&z+FZ#��ь�3H��=�5�;�d E�~Z�=�$��~ob+�D2�ޚ+�A3r	�F|8[�@�q��G� �W��H�����]�'@��u$�%���}��,�Q����x�����W��Ŝm�Y��a!���
TO����!)��W���uQ��e�F?v��qvjʎ	*-�!�J��ܳJTأ\U�q�j�/a9D1�$���s��a�$�׼�������J��ܙ��Ec40TJ����N�0c#�)�h���p��)9q��業M5��*.#0��Q��"� i.lFHX���O�!S��$�\�)vH1Ai��G�/���<U��M7���r-�3�{��g�X�<'�*�(
��i��Zɋ�X?5�l�*CQ]���M:�L�z����,�C_���O�U'j[����R����}2� ���L�ao�O��g^xZ��`�T:�,��R�t���Y�B/��db=l���'��w��r�Y�2�n�S}a( �� ���[��U��9Zb�`w�/�M�������sB�~�ꇐV#��&���i�#�*/�8�'�����"62uB -u�n>���I���_!�E�c��lTg)�,�85�\��sS��&��!�.�u�{�ѧ�adص<����4��gB�L�(~Z�r�����x�$C%�v;�fT�Q��LGL^����/���j�G%�'�PNL/"��׌n�Ih�Š�y��W�@�I�xo=�Oj��`��3��6��6�A}r,�K�D��x;|3���+�j�leO���S%��h��E�J4O� �O�� ��Sp�́��G�͞z�Gٝ�uP�ϯ|��k����?
��8d<�l��Ew��
���=��0��!�ۑXV�9�?/��BXe�#��i`�,���\b>���!�5E"%V�*t�X:��m@�΁�����%¸�Mc��!A��g���,�]\v�������F�����##��F���/�D�k�&��L��I�4&�t���`_�w���`�'��B�Ay�~����M�2ܜRG&����U�|�?��;�@��t����T�稶>�R��oΌͯ���Yl�e�|&��ڔT�f3i�u�5b�(�6�o��o�4��k�A�M�o�F߱��Ӌ��c;�&�ѯv��<\�?�V��OG�PQ"�/��wA�G���F�:�����dc���
�8M��qr���C��#?i-'n��A7(����Pra�R�&���;̈́�ָ<4	�D����_sH@~�m��������[u����Z|b�8ͮ(6��`�>C#� U���<�3W(O��$��D�~})�|�\n@i׏��-w��JnzN9�y:��[��p>���kB�:�x�[������-&�c���F�9�A��t�h��	��<h�쩈��M��f�X=j������1a��T�?T���4ˢh�����}*�<�N�%"���a���h"Y�N���Oc�k)�󽕟P��~��|1d�5zZj�h�=+S@D=��/�(4�`�?���r�֝�h,>b������[3�gjT���a�X����>�����`�#TO�k�@�����W|�t�U���.[��T8����^���Q̦��>��P����HL��G'���0�7'� A��N���j��;S�V���+��3p� h��C����^~�iߺ�#�16�����Y�OVBs_�H 8���Sɷ��DzO%��a�KwJ�����!��x9W�ނr�c�͸�u��rp��g�����~ kT�%�2Ƙ?�J@tF�g"����u[���b]&9&["+�^P�yW�S�J�CKE�zR�t�nJY5����]��F&V�:WLg�?ܲ�P�TņV@����1d�գqQro�`��/P�=#����l��������F5�{��)D7��h '	��|}z"�k~���2N��
�X����Α\br�m�����U	a��K1N{sl-Vf���`��z'�H����Ek��=����Ѻ`�:���^��V`�^�G��K�o��ssɉ<D��Z��)��ʟ�]�(dU�'��OQ
Y��:ۗ�[�Ĺ0��}�K�6�	�����׆a�LgW`�;׫,�`+�$���וƖP����!���V�Qn?l�l�S<�v����!���.��#��L�~�L�[�R���T�mQ�Z�9o���ǷY��$�#9���l�C�Q�����A)�c�kH�@7�y�Z<3�5�a�݅%I!��B��<�;��6��k��_�̛�'^;���K�e�ת.p�����u��{��:f���,"C.���Κs���O��0+��'��0S��xߐ�EQF�"F*�	�}�2#�c��*.P	���n�% �t����9T[��|��W���d����mO�	e�B�o�����8�2�)��\�g��[����E��X���i>�x�D�SS���t�m�6p7N�{�^s1�M�n��������.�U�e�����m�2
�IK�r��<I�	��2J���t�_+7;���I�Kt�B_��<<H���כ]�XV,��	�t��"߽�E�]��I��s Wܢn�<�`~A9b���o�OϨY=41w|4%�
��۟�d������q��m#�I
ו<߷��*�8�ޭBA�Q��2��o�}�R�$o�{�	+�-H"J��(�DM�1-t�nu4��{�[�FO�<7mί�tHY6˪)%-KOa-(Y/_���G̬D��!8�V?k����	c�K�`�o�� &�U,G�l�<}����;1��|�ʧ�77�6@�[��v�C���%�x�������)�J�~��vo l�P@/F�pB�?�-��������Hv��dm��s/]#�i]��C갩�/9:�=.0�tu�G���G���W�k
%�h��,�2�>	s?�é-h�S��O��(�kոA#���ӗ�	����c�U�w�{#�D��1�A�WU�Ђ� �I�O��P��q�B��Y��I��AO��i�I�Eg�2�`i坵ن�//�y/s_�?�����ā�o�i����$���&��YosW�6�v6N�S<�� x�F5���&hA{�e��E'Di�V6��Ux^��}���i���@���*I~�F2_q�����M5(u%|���]�5�Q��T^*I�9�=�����v��hg9%}k���b%%��2P1�c�`Y���A� @S�B6D��+F�E<l�M��㢢���9�p����wӸ��Ҟd�����:�7�{d�>B�|2��[� ��d�Qk(�X�Pٮ��b�>���l�I���m�I��D���E��8C��@���27%��W������6Чw�D'sU��C�)�㇓"��:j��)F[�K$s}\��s�`_}�:�74�_�c�n�kX�BE�dF���l�evx1���3���:]�6Pk¬�ۉ����Ѕ�/
 H�7FaF�(�x�c��ګKOF3��8^F�#�7R}Ě���:7�!��v��K��紌.^j��~h���k��Mȱ΢����"�,B�m��1C���:�