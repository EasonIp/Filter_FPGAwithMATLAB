��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_�V?o6���p!��#��9~̢z�x	����M�8�DӅ>q 6��n��  �	���Oi����P�ª�ج�9���Q3��eS�&�ʟ۹����:�V�ۂZ/'m}�Dv�Cf��)B
�n�ݘ�I`���e,����i�����r���+=���%{��V�ݴ����{��L�����3,{���<�@�3��N�0X )b�t��~����=����y��(�l\�m\���?��B�*"Rߎ�R�ʃ��t�6
dw=y`j�2�e��J������^��ò��-ƀ˘��yqXy��1Ȓ��h*�׈��.�T	森�y% \PU�*AH��i����Q��w�YH�#�k:����db�s叢]����8�Q�
���d]�5�h�Vr�(��C�c���¸޽`f���Y���#�:D?��.Ĥ_��5c����D�Q�{\l�M3�r�������
n��b�������6AZ3���r���%���Ly����7?i4p@�tƛW "�o`α����n0��dv�qnh9!��П4��[� k:{��ERS4�ۇ1"5�E:ԄxDL��AFqDu ��b��e���6ϛn�?;$�=_�t�s�RL8��""#�Z=vv|�g�t�嗻CYY���m�n���
����|�E}������aS0"d��*�q��h��a�9��Xy��1uY-6��Af�����F_���Ԩ��|�Ч���_�y��\ g��H(����|�&�D��F���Vv��&Y�kP;T�7چ>�tH�w[���W|��5u�S�p��[
�>���B ��{�t� и~h�j,^@0��Ƙ���(6�ɉw�ި�Q�D�je������g�����M��i  ?���b��~컖�<���1�\a�/�jq����'ׂ�&K.��N%��=y^%�����?��$�U�?r~]����M�G!˨�T�9{˵Q�6�q2̨�.��/a���;X(��ѭ� �zu=W���u�pH�bn�/�i��{�v����Kn�Ʒ���% .h�U��y2�:	%{�'va@NinE6�F ��Ӥ��OjR�O�#����}�ϢQ�@�_��g0��q����.�K{�d���Q�P1p���3�u�7��K�_T���ȱ���򲞁�冠�`Y����gmͭ׫=���0є�Q���oe�T������H%A���<�8�\�IO���2�eJ��h�_|��j�SO�=��W��sor��[uϔ9��a#��,����!���E�\��Z	VNp:I ��U,T?�L�����=!��5�b �b�s�ƛ?$���d=y���,���������H���J���UfuaV�..sm8e��^Y�����1O��,Y2�YF��{��-�Q�]a��#�,g�I6��ݖ��f��衕;��oԼ"�
D§:#/k�	�@���y �!�����;���tkU\�(�p���!�mo6t/{���|�:t�Y��"�l>�m8Ϝ��#y5�Ϣ0>�F�c&��G� �֛DW���zE�P��t�)�U�������4v/<,pU�㦭���M�Ӛ`�A�Z��q�HJ����n��4�`u����7�ߚu��`o�U�0�;Չ�2j�By>"��@
}��B�҄�[Y��܋B��CK2�nd<4�� q����y(mf�J�Z6jOA���Bۯ�M�0�:@ZF�A�{A��(/��M;j*��i��/�س�/�$���mw@�^�J���
(40'�Ͱ �}�0�
Ld��o\�N�{B�B�Y��ՏK�'{떟l��/��hD>�_��R����0�5�"�����p$�>,Ꞔ��b8���X�$Y�t?�zɍ)"�a��$黑m�<"���:Bg��z���35�mN���S����|*��Ʀz;��z��o��~9=ɑ��'�ۧc]��.�������1����8N���v�cH��j�^�=.i��}�i v՗.�-Uh!ru3aK)s�L�yI�$T���B�w�P�>I�Ce&Z>	E�^��%;�Q��M���,|PP��j0"D��lּ}	�]�lݬ{��S ���[E~���_�X����@���nPb�Կ;p8*�g�~fKy|{
��d�d��M,o���Q�ͦ��X�t��H���EJ���}��	�g��}�|i*^=�-^��j�~S�y�HK�ǃ�`���Y5�e�����1)Ɔ�1r$6�Qd֨�!�,�x\ӿn�	�z�::5�� ��zf�`��y&���*3,倸��(ֹ�D�@,
̑3�9^��2X�8i>/���'��7öD�C�i�Cp�h���X"^�ɲB;��@\^�CK�j~���e��UB��saL�Hh��"��M��ǳ�7� f���W���&D�]���/8��PaX������v�o�
�*����^t(:�x#��$t�U�s�As`�j��'
�����0Qkj���n��R�=�o���x1Ud�%��<��U7�ڿ��c�y=�8d
l@~���;�l(�K�E#�ؒ�c�~O 6Ϊ��J�D��f�2Ģ l�fJ����%�V2�����Y�gU5M��^~�HA",LS]�A������.�8s��S���u��4��5���y&{quV��WCC�`�c;�������g`C�T3�^��5&g����z����q�
��l��ov��bj����QS��Z��3���j�!2��De���;���B�f�`�eD����c�bDX��B��R�[�]m#� �uR���&��w�bw�C�i���15��%i&~NYȂ�u8���9I�����T��,hŔC�D�.��g�2�X_�_atG#&��f}�n�����W%�;���>�D��a���h�Ԍ�2��=r�i���z.x���߀~-������P_���׻�ųs�<GR3��c�����\ �֜J<p�%{*������=�k���LP���Ό���>��Nw�ڎoĴ����(/�m��^��Znl�?���������V^L��s+�Iz����s�"���ϋT��Iv��]�Cq��4�¸���5ބB�ь�$Z�+���t��<�agȬ�g�ue9މ�$�m�W���NT}o�D�>]=0W��ɉ���K��{�|:�� �'1�sr��I�B��+����<��(!xQ�q���m�QY%��I�L4����I�(p���}�X@6�[�@��[n�Z�����"�ϋ�RŘ���9��P�ʗZ�8���-�7wg�Ss��ʹȖQ-y0wPs@B3|��x�,�K�CE��r�Q��-Nz5!��y��=d����M	����ۙ�H�}��fU���
�lt)���� n��A#�샎�s�O����lk�*vϲW��g���2%;��A<�ҧ�o�bhY'+|o;zT�xp�y,NV\B薒Sd��S�mp��=ۣe�Mh. ��+8ʘ�_�UR\G�Uyܗ���]>_����@�O���d;����L�:4u<�&u0��	�pR3�1��#ь���ɜ��Z�%�U��N��qޠ�X�[�w"j��&�s�ѬY')*���J��ǭ�`���h5ņ���s;�n���~,��Kp�[�����^���;�g��RS��|��~�eV\���i��G��N��{���޾�Y�!ϿiI4і�K���i_�"=��X'R%�]W��p�FJ�.Ϋ�:/�=�Y������z�Woz��,�o9����+N(�"QM�7��/����O�����PxF9���:��� к�����)��BA�*Ө�Ῡi� 7�a�
�2>�m�A���8�hkmzV:�U��H��OcВ�z����e�Sܬ�=�{��j������Ƃm�I��<C