��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��)sZtYzѦ�#����������^{���f����@,�B���ul@k�"T�z-��0��{�oQU�<cM i��CV��Ǣ���j*��>3���B��1����ݿGi�b�2g��8��H�2m��@�}
�G%�p���.�x�T$X�v
��;�b$C����f$����D�j����+���DM�#��k/��|�S��p�k�ҘMw�����t���3��	�ΆLww���LG�\��*B/qR�n�d�"O��
���<�[�ٮ<��?^�+�#�����\`2Y�Ϗ�cR�W�G���	@oU�z%�� �˗�#�fŪx��>��1=��&��mErc��ϿY>g#d����WQ��Q��h�.�8� {J��=}�17=E-�挴ە&0�3HFq���F�W]E:ń�{�B:�(��=Y��َ�o5qxE�~�4 %te���s�6cܮu_�b+�K�s�_H��м����-�]�Ô9s���f�Y�5@�(�:Fl���t�����"���s,*�D|�ޝ�'/J���v5�������n���4��>� W����� ��驣�֢�7]�DÚ�\�y-DӢr�X��5����}'�E3c�j��6�۫�����0D>��Tf�G3�>�~�0e� ��d'ɔl�GP�j0d�S�T@|�;�'���t�C����K�j������E��n1�$b9��z��!��o��1V��%��xh�Xy�����B"�u����hk-)���7�b�ψ�V�*�㿓M�}0K���.��"����6�4�yjᔌ �a�o��������6�1s���S��.��j9��;�;��|K��Z�n�>Av��)SD#�M�sYt��HE����J]�B���O?�X;;И�I�sx�8j���:tc� �S��p=:� ����sY��<�����W;�}} �A�a�R� ��T�LYYD�=[:��w�sXi-{���|dj�>ePe��q�.`��|�=�#M�4wD�P6���xU����]�����W��3�C����8�� ��4�������O��5�����Vn	�`�;�PgO¬Z�PJ�ˮ�&�X����D%F��P�`��:d��*�U�s/W�&A-)%��[n����t[�%��Y�M�[*¾����#���y�uf������V�}
��^�(l*�)ź�a�(ܦ�G�C �
v�2F�����?�n�e�&�j��R�?�-֯�a7��O�ɰ[��x#�Qi] ��`�_���~�ӯ>�F� S->"�HO���޴�>a��+8�(,�6�R��ԁ�ܞU�H3�
�8�im:C��f;6zqz��WS"�LLK��CR�8�p1p����>
��w.t�8U�-��;;�"/bUZ�t�~dj�8���������߸qT�y���^r>v@E��~$���Q�(�e �;����;a�<�i��f��f8���ܳ�L�gӴX���N��C�u�$�VF3�3oe�[6`*6�YY��4�W��*4V`�u�+#ڟ��%�Yd0D���gq�+�k��<��1�p�v��1o����v�4eO�]�!X#�L�b�ߣ�}��0+�+���� ����/��P�%�_{��O�S��Y�Z�}� ��f�x��A����ΊF���a��?B�����T'E'~�|J�
, v��}��՜q���i��C�x�Ç_���	-�����	�����Z���S 3 SZuV����J��VO>�f	�@�'�.Mu$�y	��0�#�'4%��>6�\Ci���P��J�p��� gUE��x57L8"���(;�nR�&"V?�6����궹!*3�&�c�f��m�{��=}�M4�&�(��e�pKb��r5eJJU:�.g���G(HG��*�����$}���I�=rz}��h���u)���&�RoT=�q�ٛ�i?&�}����P��x���09)7�݈�9�k6��avB�7sv;ϸ����� �[��R]���UQ�&��9Y{C&�6)���nM"څ�z��U :�>�ˤ��q_�H�䜚`�&ha ��)�����<c���A�k��"R�0���������.*���g\�=Cu=s�%�>Q��L���j�g��k�N�ɮE�n�E��a6ɚ��
6�U�rop �-r$�V�@�R��hj�f^�ŊO<m^"+j��s�\)J������͠N�s�qu�o#�U�cl�)o��i�)�I���NF�6MZp%?$/�����"[ov(,�������@����Y�X�E�U��_&R�xyJ"�U�rM�*���=>h�, ����#��\�I�j/~tݠ�5�]T@�����.���$�h�l��削Њ��_-��x5�1��cp
�2���<�\_��!��7|��o^���'��Ac�?�a'����s9m�RP�����F�z.����t��V%WX#>�7�N"����U�x���{���g����V�z���Hv59*-}�7L�De�x{C���I��ς��x��G�:��R~��
Q:iO������)4�I/볪�d�����M���?1�:#�W��Zj^/C���^^��E��k�w�9[*�Y�N���r��&7����8���0J����E��3�t��(U�v���� ��}tN4��1�J�?����c;Iv�'���S�D#~�M�1�8��#�3Y��xBJ�l�9����� Q �d�>�����F���f*���v�;�f�� ��&ى=���Z� �c3֍lEl?����cc� b	����v&˷�'nqIV�A�B6>���V뭫�W5t	_�5eﶒoљ�*�p��<,!	�繞9��2g1���"[�Ǎ�n8�M���WY��^� �e��T�tkͯ������^��n3c���u�kGI2M4���(]�qoY�'$8R���܃z�6:��ޗ�s��GL��'?<ğ]�I)�h����WU*�m��?h�6"f�.l�B1{UNA�}μ���+�d�@y�p���:���x�����>Jg��PO���҆И5�iC�t�G^���y˷�b4W��+\W⛽���dh���� �t�����)Ki�G�Λ�";w?kUڱ�E��(R@ܠrh��N�tF�)3��^����}S~l-��;�h����lOB�Y3S0� �du��Ϳ���O����lL=�I�O\�P�uKB7� F�V�1h$��X6�`7�s�Ϣd�3��#uI�vk��EMNy
l'����,2[{��/����ǟ�suYG��Rl�
jϐ�TȪ�Hu�R1z�Pq�P��Xɯ�'�v�41�gdg�l鸴�/�a��h��י(g|Z��4��p����$��7κ�U�OU6Z� F���v��mS�\| ��k��Q6�V{���;�\$6Y����֔��ظ)�hP	g�)����� !Zag�tc�(x���p��d:Ǘ�UL�$���i���+$�ֺ]���D��nytܒ�/7(�\X`=�v�s���94$���M�!���w��j¢�������ݪ�7��;��r�I'Z��a��t�8br���7��2��J�������S���Q�/i��Q�����I�)�8ؘ���.�ܙ�c�#�8jb�͌]SQ@Bӂ�- *E�Y�O^:�L��