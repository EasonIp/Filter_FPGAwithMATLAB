��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$�ʫK�/�N�N�����c���gb=$q%���+z�ۄcRΘq�z ��7��q�1�� �l�r�yӎ��鉮�7�p~� ��hT	��Խ'L/�!��<�]Ж�3-��W�ڑo�)��ߜ�@�W����C�<r�#�&��'<��\������=�k��ۻ4���b�\j<ݜ�_4��r�4+ ��:�f�=6�p��q���uL�7��?��V15p�Z�)�kMg{���g�u뭋(!��J��d1vx?ʉ��X�`���^׬���>-�E��8X�p#�Δ�-�y�q�e��W�W<��@n�ntSܪ
Z���=����4pb
�ځ�<:�Hnj��5*Y�v��߉+f#m�21x��Kל,4���g�� (?��#�z���(S#s���Z�W�vR/0x�.����0�ӻ�A&����k=�t#!�W���=��L�}.�����Z"T;hn
��	�_]W���xפ�	VH祆�\�P�� F�cV�G0b���Tk�Ÿ��5_�WY�=.f�����L+R���� �?Lp��k��fY䰪�������D���Dzu�
�f"�@��kO���F0>�z����`y4�6�bq��mD�V��P��+r��
A��\k
����D���ٴ��F�X�,�D���,��HT��YO�RWC�0�r����}gƏ��$p]�u��Р�����⮟A� �O o���`�V�'��(ɥ3vgHS
��(�n��Q輷EH�]�d>2􋪞���`�wҿ�t]Z�c�MKUB�+pD��"qY]k��/���2�<ݞ�m8iYN���ԟ0����N)0@��E�f�p��d��-fP�L��8R*�r+���G�v��:u���E��Cu�%���-��-~11�Ɋ�%�x��8�J�x�Iĕ��#Aߣ� ����뵢4Wܨ�"��B�������/��}X���q+�C9�阅�-����g�b����kAĽUL!#ud�xIF��?Bm�*�.�
�t����w����+1��|� 0�}����p�%�y�@�E'eb���Z��~'������{��������E(���l�������j�ߦ��{wS=�[-����AA��ߗ��G�����p՝ԝ����&b��Pe'`�1@�U��00g�U���z�������1�]�0�&�8�LI�u�¸D���q��k�Qo�0⸀���R:/��K<�
'��P���� ?��4~z[��QG��l8�jƲ���A�˨j�>D�v������`��J�6C�ۅ�A�P� ��Z�+��'.u��+�Ř�W��r^��S�b,?R�9ݯ@�����dt��t�ن�
X�&���"~A��#x_X�&IŸ�F��y��X���2��o�^T�
�W�grtJ�E0�_�뗱s5�<-�z͒kr�U���! �����mf�z�{A����U�E�gS{[v+�Tb��yZ�,��{�iJ��:�²a6A���`�_m�Mt�����dC���eu
	�g;���	E����UPX�{ (Y��\a���GȻߧҺ9�]�(a�`f�:��D	�wH�38IJ��.|���ُ7�~���ꥷ�o��c�˃��Bݾb���f�c77����`;�8k��������B ��dox�2H/�M����y@�	������g�.3�.��Ð�p.��n`͡恞c��'��f�A�%{ �����[�m��]I�hy̺jQ��(h$�܎������t���$��9Ґ%�p2��	k�T⾫B	��h�����v���I`΃�s
>+^	�δg4V�i�ڬ�6l1?7k0�%oڱ�n�$<�����(���k�A��B�t#�J�i�l΍����4�K8�rG�ɨ��"q�{*6AS��/�=P��wZ:o�G���ӚA���|G����l:�X��hK�o�z���4�9�yb����MJ�Ww���֊�L��Cr
��P^E�	#H�g'�|���Uʌ�ʃM�� 1H�i���LK	{��i��a�<�˟��NJ����ާuT�}q��0l�n� g���MMym_'J	���c#�7�{�1}RA+�|x��2�a�UX�೰e��/�]�?EoL� �:f�Ȩ22���w,n�.O���ͦ���(�>>�8�o�B�%fL���#�R�JŇےhg��M؇��.��fԖ�y���(/����8�"����S�/�˛*�$�q���S�Xҭ| ��d_�3�� SC�D������"�T�n�AWA�o�C% �
��3��9=�����ws�O$�g0��IqX0�6©�s�љ�P�T)ɶ�-/HҖ�����Pi���yѰo���E���'�G3�9A����?J( �߈߁uTt�yD*�Mt�����x�o�T��0��c��h���;��d�7��6��s~�%â�MƇ!�ǣ�9q���w����;s�_$^#����~���?�TTw��ԍ�.Xn���RA������Jg80�}�j*�D R6�8�=���#���D!0� /��u^oN �b��@C��!6�+Ȇ�!;\�w���������N��GTs���k^�b4�<�;�z>�7R��CH"9�O���i9��=�2�~ĽE������`{��G�!�v]q�t���3x�+/�p̜�r�	�9e�s%G^z=�@�sS[[��]"!-��̧��q≞���� Cq�,���_�)�Sg�em�f]�b�ܒ�
	�%?>����˰���W��S���$�u�TH[�˹�~֐C��R�}���fX��>l�|�"� =D$d�\�/&��#k2{��N��V��!�0ւ��ѯ�G�dy����~��%dT��;����[B�wp^���As<�lj|�~��'g@3�o
^���6�;�Кd����z<�V��9�$?!�K�m�˻�dժ��/_�o��#�	m�O9~�:Gr伙C��k�t gZp�U
۸�b�V|:+�`L!��&R�ŏ���U�Qb[���nR�xY0m �@�K7dU�#�f�<5������pMh���|h�K��!�`,���������<��Q!���9��Z�E���HJo�(S��i���`J����ΐ9�/��?R�l�pu�������t{��/1�ρ�6�+��\J��A����`?�t�0�h�Kw���$�f���7������Pw�-�9��tl_�ky+�څ�)+��`�	��*ndbm���˖��Bs���y��9�͍�� �?P�0��E�|\.E\D�$#�~�$35��ѥ��/9[�� 聹NF�6�"�b1K]���<Ӎ!lk}W��g��)����G�K|܃T�t�ee�e��8P$�H�vFFm�8��Dkt�����oL�����).��0�M�d@���j�P%+V&��� �ҥu���/4iNCT[������R�̺\�#+����c�x6��y�#���#Pp��GM��ۡQ�p��"�f\/�P��&�?P%���6J���&)��;��z����ĥk�u�¼�v��6q�*���X���B�l�ǒhп�l�|�F�@��k�y���kqˢO��g�m/��مY�
]EU�N�l飭uN� `h��f�`~�d[=w�c{�i`AE��z�*�`E���Ո��&������%5����eS��e�;R쑭�5�͒Y�?v�%r�z�I.
 ����[L��Ym�)�(��mV�T{$����$�I��P�����q�d۲�_=^�?w k�^#�2�2hP�餶ut�X�W�؅uf��#�@�mwSD����Z�FA�m���E=!8!�b��p�vL�Zĩ}�s�H�V_b�w̦ ��6�:�x�^�7e�{��/�i_J��{
Iز�ֻ'	ǡ�GJ���?P�G��;c�FO���xj�L��
0�	$�W�r�BSF�#J�n����T�"��ϖ���I�Cɖ��
�����������Sx!C�-h�X�]0��0ؖ$��O�� $��,#D�~S�
���
�N�l�hEr�o�,49�r+S)�
��:F�������.�� �%��L�.��һ����:�=J����)��{[��0���}����D�"#.��)�Sw /��_W-�gn��Mo7�����_Lu�_��<����]:��ⶄ��k�m���g����3gf7ZShz������������=I�K��^���Ӯ�*;5Uޏ���9��:��"�bK�{w�u�®�Gͧ_�p��:��Le�~�w��
�������'G�5��0�$晃`��i7�®�s��i-iy�c�C��'�20��l5�i�Of�M����(m鸹e�s��I���y�@�y��}O����?�Vi�p �����ƻM��n�tF�V['�l�(t7�#�X'�R#(�C���7�Q�0:�M�UCړ oIݔ�
�M�+�U8}�C����q9���h9;sO�_q���ξ����lS<��8�tBw�Zߏ�u%N�ӂ�zԙ_I� �i
�Q^��yPI�~W_i��|�1��BI�1v-F�u��	"ms�(�ieJg�u�k���}.N��{�np���<$�_|d�:L�E7C��b���e\&1t[<�{�L�;�!�a-\8t4�iG/�re#��