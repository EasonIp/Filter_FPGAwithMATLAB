��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$����������tϤ@�p�?8�c ����p��Jd���L!I^�<��B׹�Q �Q��
~�3�O�}��h�ju��Ut7`	��~s�ΉL<v�B��w�8�ӓS�tV%]Z,$Q#�T���NT��=,�l��R5��Ъ"��9��(9�M��g3"@��:���3fc��$��d's���L�ߑH�F�CRj�z���A�Q�"!���zE�R��Ͽ�D)mx�����9J�M��r�w�-X)h�Z�9V��)Mb+<�1�M�}}j�?�gtF�(�i��t��%�ID�J�U��ة_I�:$�&%���M��*��U+�޽S4QW�_�ҿF����%������i��]�E���O]^�h���?�B�j|��~����1ʜ��l����5��oJ��J,j�yY�rÅ�["�$�3�+�@�\~�ۯ�a�|���x�P�|gI����1���2��Ouv��{��R6^ߴe�����)]ou�2mn}��ݫ"
��rǆ��n�O�k�`�`0����������trx���̲��r˓+_�U�� ��X]�@�]�}M� � ׭6so��g���<[����-#�,�9$���d�d!X���1z���3T�MȄ�*�P'Y̍�X.L�7�Eޱr���N�č��"��?r8d$;,\��X��W $uZe����pPg<<c��1�����_[�'�����C�c/0f���(%v�:I�8x0��h�Vￖ����!9�z{�$#�)��HQGn�v���a�>����%�ACw��a�2'�Nc�փ�V�p�����q��0�o�-����U`��u[��/�u,3���&�'#m��.@$_���#MW��̈́��W�Ň3F�jߵ	C ~8<�K �c��T�F7zINR���/ҳ�g(YŖZ���MJ2���F"_�G�g1'�WU|_�`N%�S�54�\�X�ec1��G��)��N�~0~^:���������[E&o d��k�	(��I��ԙ5ҍ�S5�4R׉&��A-o�S�����:B���P�E=�ꅒʹ!$Z�ǽ�≵!���a{M�ƠL�1�R�z�g��(Oi��p��=���q�_�����Y�'4_�1F�b\���9[R)���~X7��G��lbJt-~�ݻ{Vzʅ!T2����p�WgB��R��ϔ+��v����1�`��m³�M�ˤ�kM�ʘ�Ac�n���4J�׭���*��I0ߝD)>}�"Ԫ���}���S7�(���l*f!�`��zE5����,A��+2���J���ig�e������tĸñ�ׅ��p���ۏK���9��-����� j�?��6)��t��^�Ӆ"s:4a�5�ȡ������#c%b%j[AG'�V��uWcJp�.,KK!
��*=���r�.C�]����%��͘DW3����;i�3��j��d%\�eP=>j0!��c@�
�"m��b��ٲ�I�Qޙ%Y�K.�)��U��y�kz���#SXg"y,�7���!6���A��թ�Ta���,!�C#AN�򍊍���]��p%�SJ���c���]�J�w��=�X�R4���gi4��������["��׍a��,^��U�(8f��aX��3������#�c� 	G����L�e�^
���H��1�v�,Z��} �E�=�����[���R�9u��Ju`�48W�����m`����G����io��؈$ե_� 6�8�caE�lI3��]�64���Tۢ)��������n`��� 	P�� �Cŏ	y�e�Ѩi��<�PV��Vk}7?��:�?����{-k&kA�:X0�=�_#@4����1��ĕ�S���A\�
���l�fz]���\E�ɠ�@��e�A���T�� ����i�* �ؐ����~;��8���(���
�����n]�_i���y��ӂ!�
���wI;��p�ת�]�gNԞ�Y����8?���]���.�*8�ߕI�:=F����M��J�`f���h8�D�z���Ft��+�.]ǽxR���;��f�^\���.��@P.�WdB;l_���-�͠J}x6�Ģ��E$��Y��φ�z��S&Lm�E��˜h3
���X�d�����r��%&��g`ן�T��!�ł����n�#���;�;�4�<]+E$�-��|¿��1"$ɑe�*q{cD�(i��Žo�~8f���m�P����~]V�?>n�1�ȳ@G��9�?�@�q �_��4>����;�@~�m�2� 
��u��u�C�2�n�3��>�9g@�&�):�9{i�	R��:T4�XK�>�*�&�����]뾏��O��Λ:��߽Q�@���ak�� :��6R�a��Յ�&g#]��o�,��LW�c­��c�RfA�w���J�!��>�U��ٍ�*Ku�fOJ���Y�v��y�x@��G��f��ϋ#R�n>X�������?:�7��֡�0�%}�?��ܙ�v+N�B
 7V�l�'_�';b���-R(h�4Ӻ��y,��&5��� �xˆ9?�?�$j�V��kc�k�R��ta(���ڏ����+ȁ@��@�uP�u���>-�+�,��`�V*��� m�����·``�>x�γ/$]�u�=��wO�OB6n-����ƅ:�d؀���ǥW���Vh�"l���d *����(�����*�$���W�R�Ď����Err!z�-q�������7|b.CZ�at�^�t<7
�B �3*]�7�B�n$/;�A�чW�@8�*��X;'m����æ�y0����;��ߓ��!l�Y(�<E��Џ%�����ӈ�~I]��_Ay�b��hp JA_�g�.<[d�1	��E]@wL}����@.,�5��T5z'�l�׏.r�����"�#�&G`��XN�
*��]��v>Z���Yߝx]��BTQ��b�}����qh1P�Q$�h��v�����e#��O���~!��kJ7Mh߼�,���M�����ҹ�����
�7�	\)�/{�����Q}����؎�"�r��Z��ߘ�S��{��ǮV��wT�uFzW5�u泾�p앍#�N��ҏ���J9�|T`�m�3ʕ