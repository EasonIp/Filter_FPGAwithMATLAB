��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�
���B�+,���O�t9�������-yJ��N���Z��?��c���kU��!�j�#�JD*�������R?�uƀѽnlH��߮ؼ�����3��G�� ������C��w�6��*ʺ��?�1��+��C����챇�LII�{>��g��<��9��bE#�؁v�"��� �:g��i ����I�%=2�s�%-�6t/ �5�Vl�ߤ��\$-\un�ֻW6WV�W��?G�	��!�'��33T��Xoa� �ْkhPgvS[ |%���^�uH��zu�tu"܈�Uh��	�%�l,\�������0��ŝ��m�)x�ג�?.J����o�q{���Ԍ��I
��XD�F�ʔ��@���}`�N�+��%�H��D�����j��~t/PCVyٹ�!e8@d��l�����ji�͒޻��*�3��sdD�ȨEw75�ߢ��4�� @5�ooą.�g+���_�	}+I�+��;�cKo]V�:�ꄹ���G2�O��x��2m~��͢ H�F�q��&}$��7�n�hy~����P@F��iBV�]�1�K��4n\� <6(�7�풿��"&:����Q��Z.�wcNDA^�	0�}��4���c����\
�ߦR���ӌ����=�3�T�4M��7�I5�E�@�-�70
���c���?-B%~D�īV��{v|jY���杨��=h��OLw�*g��D���{9fPl���3|`~HI��*�~�szS���\k)����m�R���Q�6�9ӑ�N:a{⡞I�s}(��B@~�i�/�w���^^���9�Q]� b�؎)�Pf�Xا٪o��_&#*Q�P|ؑr#/�pz]�{�O�O,��;��#����A��������Zo�Na5����6�-�n�p��G�b5�)��L��@�!)�"y�H79!���9L��'�@51�գ�%%G��w�pE��f*���.	��Y��s��h.����˒)_|%*���v�*���-��Gl+��m9-Ƨ��=�Tվl�+�2R�m�Y�i����}��+㉬�9�����A�=�*}ff=���."'�>JAMu�c�T�N6�������vN�!B�,�@ε3J��hv 
�_{k����C��lSF��K!K�7��ni(Z?:�P`�F�t@����E�.a�EvO7�/ɀ#P ;62t�hl)P+�"�4����Ӎ�z�_\��y�.*��s���;<�*g��տ�ä�7'A�z*Z�L&�ǗV�d�5z�3����[���/���z��3u�����4�z���w�z-���ǯjR� ��ª�������3f���?�ډ���%�bĆ�'��Z�����4��X��P���͍àm{e ��/-��O�2b/�b��r�A�x�
�B�J��N���9�������ه����J3|�U�h��P\h��o�˫����ޫPX�tN�>>���#8��P��K��.�b^�u1a�`�O_�/zly/�~oW���s
�Txd�N�Z��,!�
��Tl���k���z#��2ɮ0��ޘ��b�ZV�fՎ�Z��]V�k�����0�
�� ]i3��Qu��9�j }��&�J�`":X�,	��~�.E$��f�s�oÄ�N@.5��h<�o/�=�� !��Ƭf�-���?��C{��+Z`�*��������f���W1�ă�ă��]�
1i���ax)�ܚ�O�>��t�������"c\�[��#��g�9���q��to"ȭ�e�q�/V��6���A��Ő[_o��f�6=Z/��ٳFu�v:	�h�\~-GYQ-ړ)���)�D�
.y[a��#H��@D����+�7�)9�t&��X�3�9:� %�g��%EW�����j|N[����t@���yZ]	�����]p O�k�`b�w��5(�dܜT��p:��po5 �n���fӗ��Fb�W˪R6vuC�4Iѽ���7���T�R\eZ�v�����v��s⫪�CfD��fc�&��:ĿM\�״�i���#W�C����#灼y(����	��K���s�P�K0���x~-�=��Nb 0��z��֮��g�B.I�Ms���q���i���M4]%��&�k�hh�g��m���9q}+�k���-�5����L��~mJ�C��* �����^��đ�z��Sôn�2uӫi[�f�q�f�r�P�5@����?��\e>�qS��H>�`�����ױ��:��}5�Z�V���ئ�5R�[\�������t��6����8�ӝ�5������m���zY�?~H�6'��	�-C5�<#C��}��6)����آ���i�	�_�W�_�q�W=V;������ڎ�_��O���=�#fF�W�U_`���MBK]�*�:��Z�ɯ>�:b��8z���̤k8�H�h@?�veC�`S�u6�I���\���a�D���{��o]��Vf�N2�H�������)�D;�Vi�l�d��kl���#gxJga�
��vx�����VD�Q�q����RT�$o��g�7�������#�I|Wl�8�LJ�4��X�&2�Z����axw���B
VU�FX��>.Hfw�λ7�	A�*�G~�s _"ΈG� ���u�h�Z���?�GҮ��\(�j������Nd��s�| �7Y#�����t޼D�Rk�x�ʍ���<�>0��M�qk����ߵ��n'垾S���� Ӿ5+*��j��mT-"��+3Z��Z\�k*+�;�Uz�t��3�!4���ڟh���8�կ�P�cY�୪������2�~��/����8�tcU �g9U���(k�{�^��ʈ���[�?�&G�vMvMjFoz��������T���A��x|�R�0�V�Z`Tdr���_U�w�L�xm���[���T��:��h	��hVa�q��҆ (�ׇ_܌�N-?h��.ݑJB+�-Ԗ�3���x�ߙ�ʽ�<r�֬GZ��?P��(���Iҥ!����e�H�����F�A��cTl��ώI���"O(Գ�������u�'�5 �,q%,q�&ؒ�y�M1ꕜ:��K��M[PX�h�C��(d00yJV�$J������zTP�� �¨PW1���J� M�p��Q� �2�� �]��W�%R���y�97�^zD�J�Z��R��@:w�э�Q*>'W�o�	Ӫ�� �&D�x�x~�h� a�8]�B�� {0J2�w�	07�4���"��F�~N���:�aG����zӎ[ ,^�:B�DZl���d;����BX�T�x��_���A�RL��O�c3��C�H ^�Ұ�[������{�S��7wV+><;q��H�����?��+6�w��d|���J���C�l��;K��˟���G�Y��������k��0��z�5��!x�id��p`�J���Y��8G�ʛFq��IK�� �܇���5@t��w�+8^����8<�e��c�N�g��[�Θ9$�{f2��)~?Ѫ��x��%n��#��u��9�����Ii^���~�Q�����5X�Mo$bpaQ�J���v��l;DÉ���ZqИ��H��G��KC3����h�t��s"�;���|{�5�� ���Q�e� �+k��B�W��`:Nq�O���H�S��I��C�:���z����^%�E&�������e�-���C����s�f*��_�\;7q�����|�,���g>�=��z� ��ܘ;w����۸S�o�3���.�p�c�yF�ٞ��p�<�m��*��lU�\؛ܾo�����N������5��Sc5�C�)�yrb%KOp^�����Μ0T�������zd��m7�*�+H�w� �R)����`A��^�t!�,:6ȥ��B���#����1	@�:)ɀF~��p����׳���O�'�]��&^�H}�z�Ȣ<x#g("}�쁩&�)�WK�kK�A�m
��d��u"9FF9�r�,��9n!��]�29V��Ġ��� 4��ح����ҙ0� ��q	�Z2�;������})�W/n<��ƽ�Vobɰxw~n�5̌[���h���)I��q��~v5/��4�$�������Fr6�y-/��YI*����f_���'��ۿ5]R]}҈��&i; ��]z�Yհ��On��a')`;�?|�!��*��st���,�L[`R0G���6���7�����i�!��f+����_����WM��0�{��>��]�9z<5\�����Er>���Ǉ}�,8HCC3{N��4TdTj�Ry�6ϳ���j���u��ϧ=��-���Q\�c�4FY�f�͖�2
+�V�<X�����({���
�/շ�=������j�
ڟ��;�E��a��>Z�U�_���62+f��y^��<���ʕ��g��t���S��x�[R eo�=��������3B��S�*]��3�����������mǀ^�����Q�bպf�Ļ��h	&�K̈�3���J��y�5F��'k7�Žh�D�_ �a�Tږ{���U���T�~�֜�H�`�+���,:ĉg�rd|�c��a���|"r~s�'��$��G '�IC�Q��l6 D�u�K'�4wH�&�/,���Q�I�Y \�u0Lۍ�I����h�
��1Aך_�=.�B倣c Ȑ��ͮ�����j���@1� t5ޅČ���ÍH2����|��g+�槖���M;���� �xP�w

5���{
!g����a�`��T��	D��>��˦๲�g�����A9�꨽Z���1=y���i��E����j^��ء/�\���H���U���N�"�F/ѫ"(}n	F�h
cC�U�.��q��%�E�]���4�FR��G�ϋA:Y�����ԗ�@���!�K�G�t
>WRZ�J���M�Oq ��E��(��$}2av{��Eh���Tc-�?Q��u����0�?S�����2t�[xU��H%/��⠲���uюy�.��l�M�j�!�H�� ܎u`�'�!S��aY��݉���2h��smJ�rq��x6����i`�%�#*��3<Z�VK(߀�L��jJY4b��f�Y(z���z���a7m9����|�qμ�+�KȀl�m#�� 2�YDwa/g	HW�oPt^=�ө���2�u?���i��7��1J+�,,GY�`����|੒԰g.*4]ʔ�-�Q��#u�)�m��r���L�$��������k��ϯ|�coٺ���1��ç(�p�]�]�51�^�B�Rf����y�*˕3HF��G@'�!�z���ʍ�±�O���,�f�X�ş�&�b�H�X&ÍxR���i*֏M��l���y���̤�<��Jj��naTN���{�,Ʉ�a�~/�IG�z}���J�#{E���oH���'Yy��S�Ђ�J�˦˰�%�rT*ADmhK�:4�Uo�qܞ%J�V����G��@k��q�r�Eګ�wa��Cٞ?L���[Pn��4,�$0���ǰk$�(��gv��[�����dHJlb�fĆ����/Ɣ���w4�Z�m.��8n��#��֥F7�m7X<��p�{:��Ԍɼ����d��S�eǜ��Rx�#8��:��)*�u��濫M̈h�hhIܐL鐹�TN���?i�x�T%�'8�{�#ȁ4h�6#z�ksxp�/��tG��ѧ��2��ߑy��ږ��8pZL�ۧ�]ؔ!V�tf�L�⚆�<畭�.9z\Mz���+2lIeo�kM�&���Z{=�U���]�S���Y�ٌ5�'��ی3����ҩ�0��_"��� ɱh�r.��Jۄ-ܞ�����(ky��ȓP�&��6Pg��<ʇ��2�u�K�H�R_��&�E�V�l��9:B���h�s�|QWU��r�o�)����6��1�0����
�oFY)Gw$�KG�	���͕g�����>��ݣgo� }���8��!���YWc,/Z�]R����w�`��T�~WT	M}��短I帮ZxtX�;��?�mF�%%����g��t&j�G��M�;�4a��h�"㌍)T.��X�r��'\�N�vT��n��L����4��O���=��T��L-�.d^� �����M������[KP��uM���<7�g�	<]�A�N3)h���0
�hf�sF\�QE��yb�5�(�t��٧��Y�^p�?��r�g�z�N9S@�A��E��x_������V������ٱT�����!��R:���_^9A�/�{\lQ�a*j���m�_n6�8�5-�&�|�Wb?���&��B�W�V؋���E�-�+͂���[1Ño��B���ɾ��E8�T����ahŬ�g���ed�Րa�j�J��ws�욮��X��M�r��i������C-�C�ɩ��6u� s0�3�*Y0� ��K�:�8�����D�����&���A�Nr�>XR��j��I[QY��6��Ⴌ�琫�OՠP�
v��5ך��Ho���������m&��w������<�I=�C��2_��1��EB�u��шǲ���*� QZ�<ή��X��¥]];�4��yJ��[�J�"ʘԄp���/REp�)�Y��,#��\l0�4����B Y!lh�ߚ<`����-�^���3 �R'4�)hS�\w��e�h"� >��Ɗ��F�y�ց�E_��ň^Ӟ]�y��y%����Ցa)�Ujf)�����b�~�� 6��8�([
���P�~G6�h!Q
H�y����HL���삃 �( E�˼N~:�?�n��첣���ԒQS���Ǒ��	|=�;��Fr���7��U�³�!wS"��X2�+��5�O*B5�/&��)�9�nSt5���_3��u{���V�z7q.kq�'cC�'u�]����X��F#җ���}��/|��F�D�j���bzl��|�v�V���EP���i�P���]�PG%}�o?޵6RI���|���k2	���m���(������kۇ�&>��fqG�aB����9r,?d~�X����×�������k"�Wϵ��͠*|�ִ���3wr��[�e1����'"���Ya���5��U�F9>�)��i��%��Ao�?����ל���YL�l6���U����	Vw:3�����u��X�.xB'�����Kk"���(ˇ�R�S��'q�f�~@ĺ�k	��pLU6C��uT�IY�l	��
u?N�� )*��c	�Tb9�H1;زG�,�6�}k�)��ٌ�|ᵪp%���P�^�8!x��bDB�ߡ���?�h��zc�=uG�@�5O⢟h��Zz^j:g�����'q��mҝ=mX/YWq?c��L-4����NDð �	��-gL��k�
UG�e��r��O�u���c����G�z�5��%��n����ݞ�I�fx����m�9wI~:��_T�A��p�K��B��K YEŖ>9�5��ɮ�i�K��IM&D-��:�ލeӝ�ɟ���T�ZJ�wPi��遽X���Q�)�4��_t}�E���v���?�a\HyÜR��V�Ӊ��Nc�����f���=����9� �
@�,���|�YL,W������d�a��9��M��@-9��4�h%��R�ӵZ���\�a?T�PV��<,�!E(��y���$�}b$U�� `y��5H�	ĉ��n��O��ߪ�5,�2�1wư\|���qͭ2�-nn�.\�?_��!�v�N^�L�MAY#<�RXme�nf~���Qh��r��ϱg��Ñ_t��e�}�U�`������������B��'!�
;h�\����(��b�tK��[A��Ǡ��Q���l�K(�%\ä��M���A�R9[d��$�D\w�2FPa���Op�Ӡ��N`Ag �$�%x�=���}G�`\4�z!�CB�.�@�� I��0@R0�G�	P���Bc/����b�-�[C��g�g�}�O��=�Y_��H#,bn�f�fs��1;K���%�I)�~����(l!^u�Q��[��L��GI��v�0ʍ��ڞ�4��
�)hd�j����@��X�|V��d��A@�>+�Y�!Z.׳vt���2���\$
�F��5/JC6�ӱ��'��t��a��N���!�y�g#�ð'������<Iأ�׺k@�'��W焳�G$K��n�5�����R��L,������`�ƴ��ӿ���x3���n�_�m��v= �%�7��-�H���Ĳj�'z\��r�]�.�aj) ��_*�)�mT)�|/;�����y���U�p����,�dZ��b�?�(J��nW"b�"���Pm���������2!���⛷�-��>WE�v�˻??A�"x���!IvMG!��x`m�I�573�	%dR�_���p{40ҙ���11��hG�^�G�ͼ���n��b���
�bnX&p���8�8G�o	���ٽ��@�Iv/t��қ��Oж�o��M����q��Ux�Sm,��1.��<l�ɦ�W�g-�ɤ;F X7���bi!eb���G����̤P1����� ߩ�Ec�h^а���R��6���UɁ�����;*\�o�*^	���+��S�տu�N4�w�F��Q���z��p��cl^��=n�Z|E��ATݧus�&��1�L��hW]�AH�!~;��s�u���Tه�Ela3�U���h'2z/M8"䪴�1��������|���8p�Ԝ��\W��J�_�� N.�^���-
�[�
mzB��?��V���~j6���p*(�g�8���ҙ�H��JŽA��tb�k�q������:ե�?,�<:�/U��*��ůik��Aȴ�B��p���K�J]�i��*�`)��8��_5�~S�ϼW&��ɝ��8[$.���,��c��"r����p~���F���ː����� ����m��[��CAO����i̘��ےV��nNN�0�8��;RO���Nc���V�-!@�Q�w��Z�p�P@�³	w_<��5F�w����-�mFR�}u*;�(�P����� #W�_��b?�S�)���d�W��Q���y&�!`���9����Ρ�"b��7!]8���]ЄȞ�!R��Y�,�.|e0 
=�x���W80.݇.�mޱ�dd�����W��z`�� ��I�`Q��S[��ht{�0?ȥ2Ij
ɽyN�1<AǪ���e`��ú!_qZ�y��=�I�C��H,�1Ӌ˲!�.Ǒ^���*x�~9��C�a���~�B��@6 �}��فSp� A�����k<UP��ִ�(��
t:n�2$�v'�JmySɨD�6��x�u��I-�0x��s�7�cl�������u��Ez"��:�(#��6�܊�eH�$��\�),h��y$H��,ү���k��y�T �I7��"��v�f��6;ѓ{��0��g5���`�*��+4�S��4��R'X#��jK�v��M� ?߹�3�d��`&�e9VC�wE����F�oL=�*_�;Z����ڱ��汏O:r��1���OdW&2�ɵ���6��Mͷ0�{���g�����!�ᦙl��Y>^&K�#<G���իqz~�#<��ʄ�s���ו�a�8��|	��#6!�FXzyHd�`/�����''���5���&��?�����9Qu��{��Q��G=��)�)"�?W�WJ�~���߰����3%�\"�����u��;�=�{@�X2�����,{�#���v��7���ZC�:�h����xGy�Vl)'�*�#݋��z�����R� F��ԠXg*2�D��GkL���69�4�\.�~ꊾ6�r͓;�;q���9p2��1�PT��,��{+�_Ϡ_����Zũ�m_����z6P�T�eڼGH�a� o��z���U}��T�T&�t��1��/*>�X�s$ޭ+������v#��,����:�{�X4��`hfE\Go�(�س5�f��{�`t�θL5Bp�k����}MX�+���%��r�6vo�GR�4}�P�H�V=M!+��A�c��G{�k�f!���-D/󦇳�(:mI�LPt��\,s/�`���=(�Wp��&9o�	7�@�k&�%��c�ó�6B�o5{��P/H!$܃����*���S:&������ۿ�I��dH�M�֔	2c�M#���2�p��v��R��۝RTi��;&�W�Y�p:Ce����$�1���1W?��)����#kr$Մ<V�I	z�2�ěVBa�H�>*e.��yX�k]�	�����Zև}���	=�J�ؗ�En�U��o������*=�<r���9̼�g�HY
�i�֬]�g��G��x-U��^���HB\��B�e�(]����-����G�А���uRrY�9�u#}|�?;���;�pQB�M��U��81�Y�b��� ��O4��p������m���ɻ��J�D����w?N*���n�խ{!�F��$�t�����q?���\��@M���A�+��c�^MH4߲�~`�é�	�h	)p��Y�J	�~�2�X���Eh��rK�z�5���p�aŲ:bCq�H��w����u����\侴M��G�W��������p��Zm�w�廕����!\}:v�,7z�l������{��9?�"0��BhU��\��u�j���x�\�3y"~��<"�h�B������V݊�þ�diM�u �e����z2��~�� �{<|��G���*��ۊ�Hm�P62 �	��@9�!�l�ǔXVZ�#�v6��)���_��<����69(�->��g��������m�	te��5o�v�kx׃R�Y����m���ǧ��Ӡ53��#�`��Е�^�Ç��s8aE��=5;]ĉf#���a*��{)�����@�/휆��RB����Ӊ��>��YF�0��rm�%������'jF
w��!�}���O]Me�����_JWn�d��^���S!;��<�QM�4��-��@�2���mA$M��_��\N�,11��Gz��@Ax����*�s�WiU�X^��"� �I����2�<�G�l����$yՙ'���L��2e�S��/5�܎�`�x�20#�.j��9X�nۖ�m�sgrf�&sإbs��fZ��S����1j(^�_���� ��X��[U�����ʦ.�џ��q�iRU�L]m����u���ϒ�� �;M�Ve�C�����ʶ-�N�+,q90OKp%@�9E��JWp3�����=����o��÷4�Tjz/�,�mپ����y8��V��MԬ�� <〟�V|����DF��*k�(ܳ5�#��פ��i�-O֥G��Z�[S]����?�+0��|	=oC4$�T5�0����-_(��J?S�)lt�:.�����_@�2�1�`���W�~u�K
��x龯�!	Jttc��@���ӇIiL�g�L�v[_��
�`E���[;u�c���2��g侀aի`������#��b�Zd%d��:$O)�V���0�����Mc���J�$�h��xR���t���5�_ ^� ^s���u������rZ��`���;���]����硫����D��%�y>6�3b��:9��G��>%�NQ�����2�k	O��`�ƴ��y�4��x*��[��;�ln�˓*��W�2 )�o�u�N��O�`f2��LG�b��%��'��K:� ���M��V����zYF�\�I�wd�|?	ЎB(%�q���_��hEU�!�Ʉ�	���t��d�!�Ul��r��?�X9�4e$�.�9�����Q����M"�$ �[E���P4�V��"l�je�PΔ��_�6L ���vm�+�"�\d�1��_`nXP��cMJ�9+GG��O7z4�J?�2�ł����+j窃�E�?ᗍ̼Gˁ�G��$�;:͞���Բ4N�@�P��(`Ahʁ�ѐ�?Mt)�MЛq����VD��%R�҇�B*_vP�:��q�t����)M�A�1q��O5�5��xF�(�+\�uG @CE"x�!z]ܜ���T���v.�|DF^b�����⬸/�Ps*	O�J������xE��ی�u�k�{e�a蔞P�Sh?��$�wVN�x���L���f�;$U���.���=cz�̉;"]���[y��'U�[Q���AU>�ܔ��9-�J���"NC��Q��4#z�c���:���x�����&ޠ��I��,�~�4�D�3�	D����+~�tшTu��鿬�m����	��I �9�A��� B5��<�F�)� ���r��_{s�r�|X,�?³�,}H�ض�C�k���"[σ��!�s?�C>@c"f�}-�TVd�2��M�$BnO�fh���!�'̌Pƅ^EM�y�:hQ����$����L���[���>�:v�M�?Ҡ����1nGҦ�����Gy5`h�����z*�r�Y�		�l�>I���aj�0đ-.��e��3��]��yKtQl���94�	T�������qpN]w0?
h�n�75�5H�w%�,�i�@��%#�Ts��B�C����{e�$s��3j�ϳ��?�������C��g|SA�x푽xn�M�^��N��L)М@��~R��Hdڃ7��=��X�V�QG�zB�����K���Y�X?F�_�<��~'�"�U���D�j��'����b�Q�6�{�Rq�E���I`�PqZs�� [;�(RX�e;	���-4�V➊`&�� �>Lm�n�Ï������������Ng)�e(��������YrL����p�4��k3�U�:���`<G�/r��=�'��N/�w��T���@ ��&R��?����Y:��OQ�X���O��`�=��t�3�]��$JKTЃ�(x!���[WR�r�U���Si�к�,"�ﳹ��0�C�S�-�Dm+R����X�V2�QƁb�)	�=�0�[� �)Cȑ(�x����3���k�"Ӟ�g>|�hW��2�m5��Rm"�	�MY��L�)�ac0��`�a�b@��d�Z���~�����J�2>H�ؐj��d-�Jm�/.֮6��x��Zl}˨���Aێ �ס\)� �b��� Td�cW[�<��;�׃yĝ�"rV<�V����jҬA��E���<�|��Kf�sn��p��~��U��+b޶~Q�f���L���ܳH ܤ)`��So�-�D@+�F��W�9��ջ/I�g���L��l����қ���ب��Db'ONű����Dt�8 ���d���x���P'Z5�TzB�ɦ�Mqj�Z�Y�nA�4�E ��t�6�����n��Q����b\lȪ>�j�Lw#�U��F�~C���A�c�I�Հo +5�0j;���S���R�S�jD��S-f<�x��4�{n�򱪟*��~��{ߟ����;�Œ��G���ٟͨ����W lP����������~��;���_���}�w�T�zj?�@�����?�AՕ��O���Es�b�T=l. �pj��׍��BDe�������hǪ�wؠ�Lԯ-p"H�� 7�s�T\�Y�H��.�B�����3C�H�b�AE,�r��#[��7i����� �ߟ��R�r���Ͷu�H/���6�w�IL׸������<a����xq����ێ�܇��!�"ʞݒb���j<�R3�LRa����盨��S�'����"pK<�,��!��Vty�lg w��Wb�%�k>C�K#Ñ�Ӹ��$h���LCl�A�˗��ow!B}�V�Ɇ�&7���,�Z��Ğ����|Uc���g^G4��=�$���U�#YrE�ԟP.(R�2Zҵ�j�+7^�c��/2I�������^4b����a�ҩ����NGb���fq~_�= 落�dL��b�8�j+dP�8���3��&~�_18.Eᝅ�5�b��I��5��"�ʧ�K���>�a�5"y��3�r��5Z���>�#�G��{�{}�wS�G�m��:�ivY%�y ���nvy��c���D�����;�b}�
��q�L\��u�O�Y���Gk(�ѫ�ڴ����SA�;Y�4����Cϯ���[�*�I��\p�rX�!�[gr���_�Yl-�&�M"�0��aM�I�0���n���� 3D� +��~���o$�()�m[ˣ�t^<
�25b��a
�솤c���,I*朥hV�vJ��!%k'_�U�ij' i0ɱn �qX#L�QH�VSHoa�Y�Ns+8R2���3�ԛ(t�S�PR�A��l�ԡ	8��J�X��D �z��AN2�i�*����I��4a�,�)��.�+Ub�$_ۃI�ٮ�k4��#��	��J�2o�zs�r��
�E0���v6��s�w�N���#8���!��f�>US@�H�b9řRRXs��U��C�=���G�����ca)3��;����^�t�U�Ey/��V��������[��e �O��H#���\n�gj�=;&��Y��g���$9��C�_��>��}�S��׮���+~�~S�+�&�1"<�K�5}U�H���S\��-��2�_C��z���d�ݬ��&��V��4vz�%�s7�|���7�۴!�r��f���X�k�^��Q�M���}8��}�:vx�%
Ӱ�3��Υ�7+ BN��;Am��SN���C\�W��pD�g���s"	-l���Z��ष���^����z�W���D�������7X�/���Ѫ��ZS�1�x�����Ϳ� -tUNDqY�(�&7�^n���o���C���\��!~ie���ޅe�ji�@X�\Tr�/��Xf>�Y hOȚ_N��@��%���Eʗ�V8m��mC잿v<���s���@{/W���ҎE\0�w̿v�Q��"m�&�|H �C�=���hm�"�I���� ���y��s�Fb� ����Z}�Q0�S������6qpQ?�Oƽ���vC�b��Ci�Cyy�2E�g��ώEں��-�z H?��-�����DP�S��=u��6wǝB䃬�ҍ�/Ś�FH`���?ur���@dg�ҩ��]+��}��}1qp��R*�)}&��w�	͔ɰdQ]���Cp�J�*�-�y�d������܃D%��{ W8iL�=��m	�����E����G�w���N�cx�G~��M�4;�s��Ai#Y���1�En��$��y�"ߠr;���6����Ǽ�$
�r�D��}UP���2Q�#��Оx٣6D��ʵ.���m��hWD��L�҉܌2. �9��\L�k�k�?8eY��Lc	���%$N[�^*���0�Kq>�IQ�v�R���uW#̳g�ѓ�$|(I<�$o�j{�r<�K��Hd}�6�8��O�����v�?�Z�p������둄�T{GCB�M�� ��:���ד=��斤C�?/���G����]p��)��?��K�	�0��!��z�S�'����%���o�0�Ͱ��~ ��ZLy�v��>�_W��ͳe����/�
�c�i�!n�8�]IN"�fBjn��~$��q�=�>�E���ŵ>h8c�/B��`�TK�kFP��%�^��H�Cd��?�����3I��}��g3 �)}�����u�z��@Z���6�A��;����z����g#s�r���5�@/P͘V��(֣�D��`���c����u�%���*�.�m�����2���>U��Q� ��U�Fs���>3� 8�_�_l/�؍�j�.���%F�����<�=!�Z�/P*�a��a�F�윚�y��R3�?Gx6Mh��'�E���������04�|e����E�**ﲥ�B�j�&j�m��T:WW=����'��Z70
@j�ɀ���b��U�~N�o�)�.͒Y���J�Z��e��Y��]��f	�d��CM�eݪv�Kh�v�3��u�۸���}FS�њ
�׭��rC�cX�zBj�qvR)DOc o�;Z�H'��+���sa�����A��ύ5ZygR�x��1*%CU旂w¦�H|~j��Ja��Dߑ�-ے�o�ْ���z z����u�㠪 ��)��\)"�8���^Y��&!D�r�\ ѭ�Oa \zp���q�5L��_������ +z��Mw����ҳ,�d�"cN��OJe0'��؍���F��Eٚ@J��5��>*n�e�0���VW��gU�hҍ��מ���խ�⃃~|U�������V<y>�*K�-�@BK�#bWu<r���/���ђ-�&��ӢȄ�$W�Kװv~�*5߅�-�r����J>a�1���k�jc��e6��.�|+�Lk�ɲ��"��{��l�o�w�y:Oé@����}���rp�)A����=zU������Pfeb7��L�ͦ���;���GO�6[<!u��N���(/uY����L-��g�,�iP5'�r���J�c���a���N�n�'9[7l&)�F.T6��ѩ���okh�g(��u(�kBj(�&�	�x��>P��}A�2C�J��,�a�c�I٫�`B��)
l�TO[����g��Yo�DA��uq���8i6�`ms� &4��lӨ��5���*t�1�\8��ϺZ�m<䏃�2�2�1%7A�9��t|�i�E��~ڷ����xj��2��� ggE�s��� i}3l3�Ao#?��{��m	�p�3k��@Ƴ��0�^˳�G	CM�G��V��T��a�f�ib2��>�m�(��IJt�)����A�q�ק^��p"�b�a������3���q�2(�X��V���6�&��p��Ҭ�I?(�7��`����:��4��~�µk�κ���n�.:�� ���\r�I��9�NӬ�H�)�"{��0sې\��]�v�:e�!���x���cz��d���ta�#DQ���k������4�̈�p�6�@�Qx¤�:��?�?D�����h㮚��W��u��Ʀ�b�+���r�Ai�A3�9�lǀ�ʥMsd�L~��s�xJ�<�D���Ъ!ԥ�*��4�ZѠ�i,���uNs�c�}գ�M�ʔP�΀9�}@w�#����o���ϊd�w�*ql!��#d��4̾K7�gi�D��'��,?��;� �.�r�����G䁍���G�<���G�LBio���nvyz����#/w���r��D�UiM`-��[Z;����}��/f^u�\����E\CO�O
[�jkD����R���o�C>�B�z��l����۲ո�	��� =�~�)ȹat�Ep'��t�&�f�N%��~<�Q���DD(B�a�!�
�~m\���w绖��``唪�b	S���נ�P�G� 1 �-F��qα6
�v6v��.�ȕ'Yz���Sx��9��ng�M�C
i��01H �����g*G�=�*8����T�B��?s�v���T�a���U�8'6��Iyp��p��'��Mrb0s"���Z��ݹ��
4@���	��m@�Y70ֳ1ͯ��BR���ZVxc �-�8�̡�*��&r���d��֊5�Zj�*c�C?����_ݝ[��������6�����l�yk ��Z�����5��x�m{_���\i�a�t*������3���r�9�P�6(t�ɔ��;������5�	B�G=�D*lw-U/榐�&z=�Iz	�zX�u#w��2S �C��c��
8T);��/�ܒ�%����$�<�N�)�E$��,T�	/y[�p�&��d�xGk��KM�� �~	�.�վ+5e��;4��Ui'�O �Uvy��N|�2�Uv,M���E1*�kH[��Pe��p�5�à���	Y����/����_�#.بT��ld�"�#��Y)�����E��w1t$��,.s�#�]�#F���n6�������@�++���t��_�Y�L����硁ݶ}���~��iY[�[^�U����0����O�+~��=��"�.�j��g�֠R�����7F��+t��LG�O�aQa��āX:�!����!(�{r�
�z�&����x��	8��U��SA�#U���.-��)�;��xy�D��PIjB�����xo�����X���ir�ǆ/�$/�nД�/y��l'� g\�	�6-`[I˶�yO���ӎ~lW#`2��n�<��:�₯Xz�0��ڒ/��lܚ��Щ�ל<�[-�!�@i��X� ���\�����@NḐ�[�R�5:[spN� mva�/�RQ�2-(=7���X�%`؞$�m�Q��6��5������P�)�2C���*�K����v�IR{Ln�D��(|�L��7���E5!���\e	�r!��ԬQ]^ ��1)��6�n~|���$�}K��҄d�n�r6/�j��!Z���z�/V��im�eF���a���dOȫ0׀h6G��E��nL��Q��(_4��\#���/	 {��3�E{$��I���k����߀�
�J6R����J��o�k(�B �$r&��F�*��m[��x�7ށ��p�݅X��D��w������#���j��������������J�v�dh_3ze��#<�\�ձ�~�H=��	ǔ���S�r��ͭ%���L��h��a���[#ҥ�/�F�t8�&��
[����(��#�#]�+I/u��1�S���|�IPk�%�<y�'��r��Id#y���hA�t��i� ������*ɢX> _,K����ihM��$"#L5�n��o"ҥm6}�����+@��o�g-f)��ژ.�{2Ǣ�3���^��t���3��A���$	���#��bO�-	֟�:�A��e����]���x���=F�i��%S�,Iw�X����Ǒ/��zD��饊r�P8r�s�3��?}��?W���g�GB�R��*�(_W{pLl��쾡}�NԷ��3�=�|�;X�%��d�v<s0R�%L���NI�֔��-�����՛'�ƪnju�1rbg������m����5��(�U4*�Qֽs	��v�֌�[�%��+0,T1�n�Iw��jn��¬�RG-5��kDL��3���H��+-0�
��=�"	L#���Qt�Dθ�o���c��t\EYt����:����@��x	�7#nu��5���W�|���ڂ�v�lR1kd[��P@��[I�&���#ifC�-fr�I���6.k����a�#@g!0'�X8a��.� ��oy�&�r���Ov�����螤f .�ޝ{�۬�q�c�smn 9Kx#2��R�Ll��m��	̮WO���(I���k!]K��B�5���D6Cmp�(�X�ru<r������z8�]�@n��N����<��v�Ћ4�{��R/-ltbx��̡r�a��	�a���-���1N�ɷ�YZ�5>������z�r�wJYg_^�@<⠚��PE���ߢ�(g��~e^x��w�n���uiu��×xp��ED�Y�����R՝e�p\g���a5ˉ����ey��2��~�'��0�v�\OQU-��f�#%� �PY<nh�'q�ؘg1F�����N��3͏���n�Ȇ�^��E�s��G�{��a@���]3�_/���J��x\E	V�����x�?���}�<�{)��4�4�K�ZWp��V�˰�+�8�\��Aڕ�/������Sr�
�«�7�d�/a�Zܯ���t]1�{4Iɿ�ĳ�#�/�I�TfT߇��?f�R��Ha��R{*������7G[u��F�%TE�q�X�*e^�R�{�=���܏��,:��(4��H�'ͬ����Ofj�Rҽ�Z��Ql��)� v��*�y
E�tҴ��w��:�Z#�1����6 `Ⴄ�IS��L:<p�i������;�c��C���	`��"�%� o*&hj�d�i��,��xhx�5S�����N�-j�����{��9�����[�(����J.�Ѐ�B�B�)�.v��f��wfŝw}��Q�����Ӊ�3�_Fl��$�oV� ����|m�cg჻�Sn����1���k<A�N�g���`+y"B�xB��������x�*�a,��w�~��U�����H6U�	��9�X 2Ā7֗���[QǮu*���g���³��O�C���Ypb�m�n��?<je�x�1h��
�P<w,�N⋟��������ǋ>���,�׉�Ue�����7e{cMf"�{l/�]�1��*������[��X�^Tvӳ��8ua˭ZdQ� �`���FRL2�]*�r���2�pB��&�bw��/�cl��r��erC���g�"����z�qZ�2�au�bj�[ħ03})'��f]�L̋缄c���&$�W��m�,�����F��нC���C����saF�z��6�(�L*�f$izCb��؅*��:�i��d<UƷ%��f��ſ�Я$3�:��u33��m��%~�Kb=i���A�6�ےJX݌��\������J�o��V�+v��}iwK<�+oPXeԶ%oy�hd�ID*���b��z�e���vG �n�.U������m��81�O���}�.��m�,��)��}԰�ZEYI�(���-î�kw�#uK#�����pJ�#���8Ug�1����5h���Z�dhR������r�u7����H;ޣπ�Y��u�I�Ȍ!\�i6�6"�S����hҐ�q>��0V1�|�jZ��̧..ԒŞ����G�F3
�὾H�DE�|kBh��$��U�P�\���I�4h9|%c����[ȕFn4^�]��ϡO�`������<��,���n��\'��Q�)�(N��������8P�_<p%�d���m�Ŵ{y���.bX�b%^����5��dؒ��u�-�+]5k�fB8GOl�d�ɈJ6"�"���?2��.c��x?�0�ш=�@^�)�9
!��D	��/��MJ ���'�����-������Tr���#t���\ٵٰ�\��3{�xc	�nr�K�h�k�6'�����+����"yfs7!�l�;FJ�f�0t�/
��PY8�mA�ݞ/���h��I�wo��rr�X��A[�����*|�P�OC�ZS9k����$=9��j4J����M8�0p�w��r/�Z6Ƭ��8�5�n��\*��𩦹�N���*u~We]�PA�>ؽ�ܿ)�Y�Ӥ��<��C�H��"Nqy��U:�W��,�p�!J3^%���*��zi�T-4v���L?��
�z�s��)��d�ʟBȨڣ�Ɩ�"|�P�Q�V)1���ma�i	��O&�=*-�&}���?��bŤ���|�^gs��(��}9� ��H���tQ���A"�Q-�{5!���K${v�dUW����&�9�ȸ��Cߐ����od	,�z/Z]�D�����Yu��/�zQ&pr�!4��2��(-أ:73�{%��B3�Pͪ�\k�kC)Vu �fvxvl~�����*��y�`��^"S����\���C����)N��GED,j���{g{��thX;��C��-���m���)�$L�rI���(w� êZ���$ [�C�1�P�a�T)a�1K��
A����Hu�ä։�� ��U���$]<[7:oc���6C;�ߵ!:=�a���Q�� �lHż`h3�7��1`j��r��=��{f�z�\��f��"�rv��%�Ҙ�Q�f��(�*�m��N�!�hs�r!s���1�M�5!�/0n?ʎ)NDH6�ƥ!���K�U���LȾ4�2�<K�gG���5���,?�/.z�\��'cw/fR��}��ۃH^��-������+�C���3�jz+6��{���^|�M"��I���}�q��0�0�.�輡u;G��s��5�|�R��Hv��>���J^K-{�)=�������$�S�<@�'F>ŀ��S�w�;1&1�Ipe�n�����u�w�½H�h�:���N�\�-��u�?M�.���/��9=gW��Α;$a,�+����.܉�%W����ZT.{�r� ��v�l4E�;�+������\��RQ=�B��V���(ڱÄB���Ə���QP��4`��`��i<l�b^R�5��mc?r��D=eL���1dn����v�e�� ^��*����뽖�6S�T�
�.���xpɭ�]S|KG����p�s�N����v�#ޛſ��C|�_�鷺���/�V�09��^j]�^�w�#E���'������7P.�n�:5���k�ja��Xk�Y����p|fa+pͫk�0۲Ũ���V�+8��:UI�$��v0Ӏ
J����G���Tʹ�7˝:����~��w�g��
�8���TE� 0�31Ž�h�p�#{����,k�V,���Җ�
�*��*
膬1h��*����%�$ �w��s?�.6V�O�� ��ɷg�A�D��ԉ=�	�tv��4�;�+�E2{�qD�B��~�%�| 7�Tg�oY	G�ޝ:N����еn����(4C��3�Np�V@���?�T�@���O�j�4��4���6��ъ��=d�&1��w�[+Kv �J����W�E��-��yv0�eu�yi�R���$z�= ʔ6Y]
 �G.y��Y�Ci?C�[��o9�,i�
�3h�|����ۍd��8Z ���P�w�|��#b_�Ea�DAu�ǠY�Xo�џ�BI[$���2�AD��e����-a27WIљ���W����]�����n��՚x�2F������<Nj�m̶:K��l��Q���9���¡�; �4B�*�l�{���3짿��@
c��2.�k��&�z���=�t��vs�F�o�ƒ��+xz1�f�$�"i�������'-���Q��6�U�,b�a~��O[����X�_W��O{G��N{NSA�n��_���eBdb'֧�zxm�G����<�ߠiE��[x�]zˡ�9�kM��x��{ͭ�t�c��O'dj5���������# r�w}����S�#�*w�(x� r�j#*�T�@�O���a�Jc�qOF�L����S�����q:LI�B�a8[������_S���R��NgNؿ"f�
�>�*���8;��s�s����z$����R� o�WsO3��돟�Ld�zBsuJ�	{+���`�]	S���z�kjj=����<.���at��eS[�+�ڔF�W��"fI^�.�C*h������5=eX���.�]ޒ�a�a�����LM���r�f7������=G��	�7���wfy��21�����Yxׯ�\$U���]"z�vp�dgC��l�]N�
�}S%k�º�ӑ�8����%�obw�����u���H)˔���&�W�y��j q��W�t��.��H�F�����T�œ��X	B�&�D!��*.GD�0�(�fk��ي?m�<O���J�a=[��aǦ��N��t�~��L긅��V�"�\�f�h�v����V��U���_�������SM��Jv����!�������O�ˌg_y�i�4�M�Os+�6�Kp/B`,��T٘1S=8�Q��G����2�- =~����|�	-~an��F�<����0[��ÊP�6�9kJ�ok\�C��p���%���)�B���N�H�]�5������=�`\�$q�r�����1��rS)�T_Idl�w�@m{��:��+�g��&d�o=v��}|�B�^�[��	��1���5oϙa�E�TK��JF�h� Κ��t~�RuD�����S�{p1���J�w�g���p*{�����L!cTp��~S~���9Ъ�	8_�F�R�ClCh��#�����f�ۆ�y5���}��ĭ3x��9���wwUv#�j_(f�#�v3͐2�̤g���^�~ֺ�a��W֬���y�|����46� ��/��[(��B�\�D�Nhx��h��D,��Փ7�E�N%������~�X;U��h�%��R��;��L>fY²�������:��1c�Z�cB���D��O�P�JO�D�j�5/�i�F٤��.	���7:�ku�R?$#c_��K9rG#>`k"=G����o֢W-@�[��4����5��=�+��*4�}1 ཱུǩh-��(�y6�77�wTAc
�.�I��v�������@d#�=_u�����9f�3�c7u-=A�lnaPm���T�x��IA���8�7n���2昻�e�P���r��V�n
�.�,�K��SZ��G̛o(�rw�-A�ot�x��k �9x� \9��bO��٩I�w}DDE4����v�p"�<�KP[l�����VS�¿t�!!%SR۾q��h�Fʯ�(d$.���}��U�J-"ln��OJ5��)������4�-K��	�gz��x�[���k���.�A���N���%\�E��g?��ħ�n��3��ے�8�ӻ8C�Ws��NՂ�&4~(�M�Nh��˨��L���U\ʍ@\�}�fJ;l��\�jC,c�a݁6�֤�$��w��S*5Ν��͠�b���l �JW~���%��gz�XN��?6��\���]5tp�+#�g���ǜ�i�arr���x��ɯq~�Aku[�k�l	�?ܘ�&�!�[i���7$@���-�H��Y���x�֤��]��:j�7�r#V|,��6١�S��uXG�P�? 6o���]AEZ滁İ����0��p�k`+���G����������L�Ehk�V]c���v�I
���| t��+������͔*T���`�׷�WQ���*����(�>Aʼ~��]PnΪ^�N~N�v����|K|u��Q ���ۯ�Fx��z�Vl4W�y�a�Z���	�����.�FU�j6�z�q����n����X���}�(�v�Xxp<h���B��pZ%zo�
�V��a2�Gw7�)i��Ff$"�_���� �w;�_������3��рp�(blM�1Mcs�tc�����U��@i��-{���P@�����������9�a%8� b�E���񲜠{1n;�
C�T�O��[�z.I�D{8Y����&S�Z�ʖ�p7���:���.�w��?K��m���ji6K'���w�A����,4Ƨ"�����1��W�D�"#��m����g�|��@�)_D��i��s �a���#�@t�������W�J����M�M�:�����<qQwģͶ���8,�~���Kl5�I�q)�}s $�c=e)I�p]����B�
�4O�A��� ����׶�qRå��U���$��r͟��T��N�Y_��T�S��(v_���w²�h��J�[� ʂ͆���g	#�;�Fi�t%W����5r�n����e}�=�*�Ӥ+/1@�����F�9������M�Hgt�N֗8g��Mb��M̚V��v��`�0�=a����ڥ�F,��0�Q~��m7�R=�=�te�'v��["1���@��+S�Έz��[�����NXR��B�fѨ�3!�7,Ԃu��N��0;o����1G��XRe�	�3�mNx�_��sĜ
s)mBJ��I����ç� ���_�^��h��(��U�@\��_���{T���5PC�h����U���H�Q��	�h]Yxr�@�#W{��P,���QK8�p����1�.؉�������2h��\���1-��"٫7�a����|�P)�V%!6�#�{z�B�k|��I����V`�S�^>/��:N��]�7�{���9�=XLO�,�I�[ܻp�n�1�y�Q��eo�B⟍�e���[av9�$�"����a6����ɯo3��PWĴ*3���5�F�����G>Ґ,�~Fq�iĮ7�q�]q������vdo*����+*�& ���ܮ���R~t��g���|C�a����O�Wp�vQ"�[��I�I/T0�mOd�/��_z���\�I���E����H��ٮ�&�s�0��� <���x�zIG��6��0p�d9v��V��b����a�D�7�9ټ�-���좈z&��e�P�)3�F����k�P�KF�,�Q:E��$g��x$����D2������6f�j�ݨ�+\C:I+"9��>�i�Z0�zaش�I�"�!�V5�f	�6���Ħ���� �#��c��w��`9.�$��Һk�/���5=��G��/H����B;3>���_�֣�̺�
�9��0Au!��&�љ��w7z�G W��1_�"t�W��7gX9
�@�( �d��|��d��4>����t#��g�qA�&�n9����Q��]rBZ���Up�f�v@~��|���iLB��{q��l9N�[VFL`��B�@ic�E�X8r�֧����i�pr�в�6�od�d�9ep���壯���9δ6k��N?�q����aZmby0����n0�:�88�@���^�иW,���@��[Sl��x��ӈsuk��c�@�d��@�K*@J�.���6��'��ъ���>��?Ž�ダ��+B������UEd����1�JT�$,�8HQZ�5��4��3Xl�{:aͿϜ$���@G�A���6�B����*N�m�	��.��%[k�π�]K{� e$A �5�(�C��������Y.R�71�6̝�1�-[M�$���HRK59x��i��[oGy���_���a�<����r��e���(��o]�Q�+'�g����y*�uS.2�j��H�bs\q�B�[���\�T�u���pJ[��/7F�e����;�V�zdm�4ڋ
��^��G5
USe��"d�_z$��T���%�J�o�E/׹�����W�� t�М Ƀ<�U�x��(_���hj}2K@��|D�{��j\Ph��q%������Ï/�Tq?�<rnw�P���8%c���8�WC� ^)�����:$I!DB�%��uw�Z0X�`N�툤�����::�aD(�0���-lS�DEK ��F���ȤWx��ӃU]'P��L�4����.Vf��|$�x����:�Lf�_����r��/=/RL��gbW�{K'��kG6QŪ�dgB��=�'�`>����ޘ>�6Wv\=U�
,��^�45�}��)�VH� t�A�o�[�
�3�u+����h���ԃa�k?��j���43E҃