��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ��P�P�I;6��y.�R?* (�B Is.�� �AqQ�s��JV��H��4�b��+w9p���8ң�>��7BHr�3�t�A!���b|���;EܦW�=&�xiC���ցt
�y!�u.e��U��_�\�����1K+ܼ���������]���}JF�� ⒅g!�l�Q��gPXず�����/is3�=M��˛5w��o�C���Eh ���7�ٯ��[�>���i��(h�\J3Q�I��r�R�#�K���0�z�G�d�M@�SEFI��������D��/W���K�('��[^�.��Ir��z삹(g�^�����suȯU�E�οV��� ���
V��t�(�q�>�RA�sy���n��IJ�!���\:U�Gr}`a2�=��k������f��~Z6��L��c1>n	����X�i�lFl8i�" �W��_��f}��^Ғ��!D���EO��I.z��_Ԑ�J̯�U���Z��&e>?h�E_�&De���nTeY B1�gE���ɏS����H�����k�$m�Ryɔ����kvέJ*���u.s��\�{�&�Z�D���[S��:����*�^CC�YwO4ʠ�9_�Jz��ѳ��Q��i�����'���$���?�3��Si�_���/'���B6#���~����5�/?!N��w��%ƝU���,�Q8����}�i6X8�	HӤ��?�8[���u�:Bj�&��Db C�etJ�#�X�E-�K� `U�(�*I�ɼ�������#;Yh˓M96`��k"�.�z�r��O�OӈoW5m��m:
m-�7{�:N��������S�O/�0{"���1��&ڷ�d��_N�aE}dCT���No�S�7��u�����DV�G&���	��A�?�y��tFa�6��#m�p<1d'R�0ݏ�C�)�P{h�V�t�-�s�5�ۦ�(T^So�8L���<1�Rg5QO��[f^���r8c7Y��Ҩ��X��} *	�6lS������"!�>�J��ߙ� ms8�N�^"P�Þ��eR���D�J?;Z|4�x���b�L1��0*1�As�"����4S�/��u���8�Z��%������f��D�?N
�(��f��%��u��8�:�����d��~�%[Z��/9���*7�C� 5��Z���ƕ� ��y�)~�\o����I�|e�J��٧Gtම�T�be��8v��JtJ�ܒ�	���<W�Z�K��b���5�jŎ$^��&$O����[��x��ag&�X`{Q�������NW�A��  s�z�#�&�V�o?��u��6$Ƅ��d!���*��c��������]���-�E|�P���3&�٘�U�sA8C�1�f�w��mKTN��ƛ����1k #��S`�(�ֳ/woY��3���Z�eq�D�����V��$�I���n��=NMK?�����f�|O�c�J���\8҂={�0���hS��o��Z`X�q��K�J�&��3y5kd1�|GP��KG�V>�/8j/X-������=/��z�����_~\i���pq쫔?�SH�w`l���\D���-�OcWH�����\�8qq(��o1��!;������x�S��9�nJ��{�?�97Z���F���f���2n��=v�Bpәb',��� ;r/�����kO$VnK��(_ŘJ��)dZm��;��>6Y�B�ia`ξ0ӕ�+T��ں+���oU�/n��%*��5{���˲��?K2A�C�#q'�(�L��t�scR�8�m�`,��]%^� �Jp%���J�xӞ���R��1��i���3sZ��a�i]T(3��"�,$�F C�u�i��kh���!�NuXD8A)�zAQme�x�?E�8���@W��Bo6E/s���_��e[8;N=���!��z��NQ�n�F:���k��-0T����U�E�sg��h�.ث�*������Z�:�5��YΫڜ\�}��F�м>�N�Վ��M��fQ{)�e"|��(&�[s�n�fx.���n��έ	CU;��O�2U4#����u���h�K����ɂkh�!@�5�ZlL��$"�ȋP8�蚕*
�;�[�V�І<G��V$b=�J��v�es��< KhrzU1��m�h�rV8�tGL���W�I�����qx�S��w�5[��#5��82t0\XA�P$��T~�K]������[N;LھL�qīcCo��X�P��K�`�U#�y{��n����1N���_M��v��S��J��V5t��+�kS��ň)��tB��������"��6<�K��G
�Pt
�����>q�5�MXɒ���$z�m\��k�������r�s�?	�S#�����"��j7>r�/�����9t�߯f���hp�Kj����D"��`��S
IM�^F8H�8������������K �0 `�}h4�>�M�d�WD�l��ތ�q'�'\Ռ#�i#��Z4�$2S5���A�m$(� �R'�83�1;�l Xa��#��q�dn�	�Ε�o�f��݉|t{d�%W�ʦ�gP>e���A�U����H���/ڭ>�/Uvi���
��7p�f��J8�@*�rl��M���4�G}UVR8�ԁF�;b%���(���j��Q<�r�#�l�����rC�{ �9&�#��FV,��Po�G�`U�^�X�Iw��CE�̳H����wg���������D�mU#��Q�E�Q���e}�E�w���eL�SI8���!2���rB����C�p=����:<W�0�<�%5����c�����oJ��4��"�ػWK�5�ŷ���=2������|��ā�"�
�1�R=�@�'�i3c�ܹ�����̮H�6�Ҡo	�=�"��w�i:��!���-]�-��wm�?�4����2b�;q����I����Ϗ�M�hb���CZ>��%��@��B`���\T"��;���L<H$X�Wh��y��`h%a-O�{B�np��D~SyN.T�YO�D�'����l��.�J�o
�׍�����g<=0@wE���,���
ݛ,:��/%\R-s�5W�N�{!��K�R�-	u�H��V�$��c��2r�u�;�a�+�V˓�B��)�l���m:57����\�R��:�H�g�t�
�����g0#vē�.�5���}�ւ��m c�<V߈x�Nf'�MH��*�)���:OY�l���_0����1q�?@7ʩ�2ez�K��9�tglNB
5����I:틴�D��Az"^z�a����ť��9�����RNʭ{�� *@�o�����Iz��~!�q�m�[\�������4�)�9��̷GG�����W�e���y�үoj�����N|�#��kz�	E���R,LX��A��,F3E�;*�4[ʒ�	:�T�յbi	`6Za����լ@��C���]�����|5��צ�qyW
�t&���h�'�G�|0��F���ۍ�B�f�F8�6��I��I�M�v|"��؈O�W�Y9����-c��$1�����B`L���df���� �)��*"���M��Y���]�Lm_�R����p(x�i����KX������؟����4��p�>�a@k�SQ!��3��9(*+�N|�wUz���7N�[W/Rpm���k;�����xV&Tљg�Ȍ���&6�ái	��7����ڇf;J:��c��=�Tjݸ6{<�dvi��K��}���&r����a�n.�`R���s�b����qY/2L���hd��3uT��`��l)q�[&�JB��N���]�$�'Y��9�ʯ�d�ΎN��U���P~;h<�W�����L&�5C�]��3,h;��~l�2�}�=��S�c!�;.���$M�*����_��䧽�,s�}��?C32���"U/�vs81�:d,�ϑa��bZ���^ʕa�c��(@�3���2�h4Y�d��oaFB☻�IVl��m;Va���!�JjCx�U�<(�"*<�X�ख़ҿ392m0RPw�@h���?@��g� ��w藿"�ێ���if�&�δwM��ʢ�_�F�#
9�lo��]�Mցr*��
�\��gJa:CD�/ʃ<��g�g@+>?��'�3�֊�Ӳ�Hf/8�"��M�$#̻{C�}(ý��yS�o�Ԭ�_JQ>?�
�`F]��1����d^��<6G�G��1�=�=���.UJ��m`���@�\����?��H?�r�N�ĂB��ۂ�Ѵ��uX�|����U�zVr���	���_��jr��:�%����Ip5�-*���()�Wa$��E-%�����n�Ɵ[���<��\�|R� �|���H��'�e�p,7���)�������YVqF��p3���k`�R"��RQ5}�DsO0�[S�f�*|���*������/��Au��gE��^�3_�Hߺ?k�z��E�e �~j�Ƹ�ZJ,�3��:f�&/1O���}���~�Źc����gO�U,~�Y�Oj_'���!�N��.�Fd��'��񂲺�T_>n���Te	L���d��W�ͥm����d�q�M��& OѫB��
 ���t��w�_PN����%�ec�@�k�{S42~�<���ZC�u���o5�r-�o2̽��vԣ������G˵(�� �!k�թ=���vx�Q��E]��MV�M�e2��gDN�]��ad��{�U:���\�XQetK*��Fx�/�$1·����7�{��'���R"웟�i�ϰTSɒ��R�c�_N<����'fʨO:���>6S9�шD'n�����r-�z��s�y
�u�znVO5�tm4�6�����()A7�%Ľ��shW��X�G ܺ���ڮD���M��5A����F;���@�n�ٸR��m3��m>ǾmM>���f"���=�gW�Hm4�̣i�ud�(�4e�1m�_�29u�y�9f̫�=o�-���{���"��2mW5�ݒ���m����g��ҩy��!{(a]d3�mr�e3�/GsD�TBx٭��L�s$�Q�-��ͣVh^��"�yA2�� 1�q4�z�RK����Gm�[���.���ג���\UҸa�X_Ig�7��E�����=�� ����~�I�"	�������|ш���U̚��l�@�UY��c �q�v$Ǔ��Y1q
�&}1�r�Cd#��<ʜVn�0�p�X5��p�g% �K�AD�q1��7�@d�Cf��f���o
�u�7Ɯh���3��:oŸ�m�ER��"��������&8jJY�n��';6�ɸ�aL�W}*�iTd���R�ُq$K�/d�Y��Q=�z9� �P��wIf��d��x��@Vhi6�����4_�:�4��Q�Ys��RdLc������W��R�S}rg�Ne�ĳ��[)`C���<��d ��c�=T�bV��o|�\Q���+����w��u�YSO��S�Q|Wu�}�<|O��Ǡe������4/����2J�69��%zeQ�(�R���J.<ǈ�%7����˔s����t����	������6aJ�SÑ�$C�%�/��B����y�Eځ�����&����`>�`���6��p�軏�4P[��|��9ɰRN����?�	�e>"���B����S��)�%��G�Tspܳ�:��'�Nc���X�t��R���+>�ն�iu��-�Ι~}�_�hW<�1�	�6� ���i��{��`�c#��X�+{gƔ��N3��Y��Ɨ��,Z��w<nL�tI �(�6XNOk�b����/�jyO��x(z��$k<:�����i|$W��2׼��R�(]jӐlU������f�>�m�U��@b��.|��h0_Fsy��K��j��6#I!��A^S������a��N7�f�0�X�K��B�C�HmX���5D�}�E�U�Wq�p\e�C��{þ���e!Έl��u��L�����h�7P6 -�}T`a��yJm^�9u�3���XiܚE5>�B{*rR��k	|���h|g)0���ޞ	Inr[�jD~>O�}es�l E���M�U��P�6�\�Va@�5���l�� �ϧiѡ=�6nC�$!����V�@�> �hg�QƶඛȔg�0+3�e�Q��ꑿG�,v�U6���o�8���TW�������V�y��}H���~�xxe�((4B���$�%Z
�mm��1�#�;|6�(�#��Jޫ>��쑯���ӳj+P=���
HgE_�y�Y���Yo|�#���6���%���:&�i��K��^r6)�o.*���S�gBM?��G."��oV�M�CGJk`R�{/��O_D�锋��L�h���d��1%�1@a�s@=��h"�6_>;���2�@����G�L�����Z[�������l����B��h�_-��kyԀl�Q�D"�+a���o�"����F�z��Ӏ��gS?%%Cu���J]�(;���0�-]�0u₁�R�v;��aA2�f�~�٩;�%̏a>��GY"W�y\\�;0fQ)JQ��S]�gߕ\�Qr�
l/�W��0��M�YQ�������P���#���5z��	�z��Ã�O��B�������Ss���\m���Zԏg%���!d��/t %¢
���i��ZFo�vB���k�-�mꅽ�����N�q�{�&CC=�v��p=c�4E�o;^8�2��`���#�r���(��v/���6z�{� �j�:�(��x�uS6��&���#xE(Se��V|�;��*��l[؂|��4�k�V�u9��%����`^z4��^U�)|#��C?"���Aě錺��+v'*�f����[-�`��+_]Ü������?0j��5��$���WI|��x�O��!��k����	�4س��`!�c�{�G�s�g��ӽ��(��u�Y�s�97B��1�j���!T�'���0[ ���2O7�x_R������ t�/Fƣ��x1��;��6�:��5�uR��B$�I��hd�&C)��""���Ǝ�ZyV�����I��\b��B��������ﵬJ����HAn�[�[� �C��n�?YU~�^�ʱ|��79LwF�jdna�w������T?�e��O$�:gX�1�19o��,��9:@����)���Ͱ�!Bp�ԪX��\����=��B}��������;J#x0W,a�X�u߮��M1���c�o�8<��~�ĩ���,t�-����Պ���<�&eB�f�)�k��g�#�K�D
[A޶X��K�
K�Ҏ8�ӝ���8|���d� �;!m:pۏ���-�q�M;iY=�gU�]�<�i;��E����$c�<����"NL�<����/�R;�����b��YL�r��h� �9'P�(���}<�&����P;k;��q~6Fvwhb��)������?�e?�$O���L�����HU�LF�<��@�0�%O�f���\s������Z\�kE�10Yc�Zn���:��l@7`6Jf��������
Ly4L���K}3�����ux��1��w�^�"KKD�����Z%J�/�=�����,o��D���EF�iK3�?�T�ش�@�ִ5��r�*� FY�A��� 
���.��-ݓE�����[�L[Q��i����nZ�jN�
}k�����ϑɝ����#���"�I�2m/�1\�����?��{�����K>c��K���͌ţ��]ҽ�C���T���pV�L��5@d���eE�E@{ 3�A��vw$����
�aF�=z ���K���I���Qw�����	�,����uC\�v�H�|@mQ��=0�*��\�aN�ě�fY8�}�k��cs��ET5���z_ �W�8���w�ez���E����Q�R���8�%��1�%WG٘jF������v�nT��6�%X�5.����g>M�D�ȅ�޵9 ���Rq��?�ļڳ���#q�@X�R���x� gT]q�8��1>�vH��g����a�J�Vk��֮&�4߀�z��EkZV���ǅ\Ne����#�tla���3^��z�����+�|+���Z���ͽj�=i�Wp��LW�A
���% ���VI��Z����"^g����p܃LL1��Zw%;�l�γ��_@����T�mtq��f8��%��Ra��Y�sa�5Ŗ(#9v�ε2G�P���UH��M�;7�򽺨�u�	����΋2�k��^�������۵�I�����:{$�le97�Ct`M@Znv8�0R���
m�]��� �N��0��a?*~�'x<n˟�H�ɵ�K~��c��m�;�ǒ{dHf��p�Uwj���m����z�e��eF Ȁ5l�	|��R��GJ��>�����e����g;~�w��jn���������cw�4�˺*{$�=�8M��K���H��|��5��]{Edx�\��?ܓ�Λo�{��W*@��F╞Y$D_-�
Qܳ�M�JǞȕ'ب���}`戳��:��*v>`J9D=r���X��
�6����"2�b���1<�6�dP�a�5���vq�Z8tEWj�	ڡ�B;\"�5�V��n��3O~�Ͽ'Yb��N�M�#�ȜA@�g2�Q8ƺ8	���q2�l~`T�NMG�w �Aڜ����J�D����?��
�{US�f>�'����	﹆{ �l	<��.��0&Fثc8 Q�'��i}"M��O���D�A�z�Ӳ�ii��M���z�m�+� ����[~�ݛ�� ;�s>���"�x9�Bu�7�'@�G�bDdoxi�
��K�Ĉ��P=jΖwUeM���H��"����M-�����7��W�Y�0����E1:�32�
z�G�v�T�=[���� ��z8�*�@Ѥ<4hå���YKC�MK��E1��P# PDޜ��T�=���?�FUFí����[ݶJY���J�D�+����8�yJ>J�<�J��;�EH����v��7����� 
r����s������e�²�JnV��[����5��v2F�w�1�P�0�#�b}�Y���>�z��L���X����R���=��L�	%އ��x���zb(�� D�k:f�eЖz�L����Y1��Pw��^w}����mG
�����g��v�l��ïtk�gs3��i�	�D]���+k[2s'��є��������;�*m�@����To�] ���+(��)6]����{!�d��d�%�l{t`<�������L*��n�&�޶��,��/n�VO*���{�#��x�� 5x�pw�X�hu����j�<�������~j��0�{��L�r���%oQ�>$�y��ȝ�W����x1�R턟 ��=�������*�R���,�j�^��d@�~X�\���!z� ��Y�f�g�߿}���]{�{��s���I%e,�@j�d�Oqd ��tr��[�(4O���rY��/^�E��������5×똢�a���Z.`~B�� �J���+��P�Y[�����u}ksz� "I�g,��7��0��#vC����"f���cJ�Q���'���o�=�t������L��Yч}0r�$?�l�^62
A]O�D����D&��-�@�ܘ;�a߹ߖ�q��s@5���x�F��(vNAʼ�ݸ��3�PIұmC��?�Z(�T	s�=�)i��i��Yf��mBX�~�5�g�@I<�,�cW�������{�>�F飌��6��hFU ~P�Z��Gc���s�ݍ���s$
�?�����ك/�XG�,�����Ԓub�`�s��s�]br$���gH�J��Ҽ�zK�P�v&��L���y��];����\����-$yڴ&�-FR��̌�qS,1\{��>�p���y�L=h(GD�d��	�lg�
��{��Ij�5�����sBT6�|�h[m��a+ ɴ���=��l )�G]�^��h�����)�ٯ �#n��7�[R�a!�CrX3����S묇-c �̩�ғ�D�+=]�-p�B(�3�(�6�s��{���ə��g���j���s����=
Y�������Qun�`�.y���,W5s)�����	�j��iW���q|A�д�����l����-9��%�CUd��@��hq~�KZ���W�uŤb�4���t=B�V���;m!rڼ��N��u�􆻏�M�+V\] S��-,��/��sN�-:%��?~���$�S�O����dV�ͬ��8@���d��k�p��8Nc��nHB}�,��+N��#m�|%�-qݬh��F�e�,��	ꛣ�i�C(���"��V3�y�"J�}�K����ܯ4O=P�H^Y�P}������#��kϛ�w#�h��D�?���3?r��C���[H��h� ���M���ي��� G?��0�CJ`I��$�<�O��nהm��a�z�U�{ۓںL���+of5�2,�����l����iciJ�Ϝ�����H����Y<��?0�F�fD��y�H��
3�%G�|�"0@gr�	�t���k����h�!�e��S�M���_�%�N�Գb$����m�p�5,7΢��ScE9�?�ܩ��d�ǝ'��P���g���*!Lm��6���k�dVq����6�X� ($�3)8e�#�	�b.0�cY6�[��춥p��;fzTH����	-�*�6r ;�	�1L��AY�n^���8�82�X_T�$�lT�l�����Ekf���_0*\f"�I��c{b�9:I�+p���.צg��0 ������ ��
q-M ��T47i�AovBmDt�A�8`
~�Sf����*�	�Av�W�;�����-;Ua6Z\���a_�YHT�l��rDs���|��	��B�N 4�Gf������sO����B/�^�6�a5ʹw��N���^�#���ew?gc\��\��od�|-@�QC�XI)�{�-�x��dXt��Q@Pi�p��M�&z'F~P현�1:�0�*�▭����$ig�(��m^��,�n��$f4j��S��MBn��ah�>[�rk�8�ȬK��A�ش��\&�u.n�u���;q�8��Q��L