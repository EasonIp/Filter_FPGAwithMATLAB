��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$��x?M1u��9$fu��6R���(-���5����� ^ �8��lKш���T=K�s�[g�ͼ��<�5�?T��,�?�QB�J�r�i2yӑQ�{µe��w�UX�����/�4�N�/�:�NIc�_aBzo:�"�DTح�����S :�kg�NN��xt>��aR +�Y�����֗��}��D��<�l�4}6�o����1X>�u/uڌ��01� �G�}/�h�ɏYg0�4�&�<%7�b��xp�.J&X0����t#Ja����@�8�.�F����)��)�s�E+ӧ��Q�̬XeQ6h"���6�dY4�8_GY1�2eQ�C�7y��j�W6��
io�����o |��F�V� ���c�w*�Ғ)��x6��#n� �b�������U�t��x���5u,ًY)����'M���T��`��?|�c�|�RM�%t�j: &��h�v�8v8Ƴ�'�ef����r��L�>�#���]�}��A�'ni�_����Wⶺ���ٴ7I[�#s+�rZ[��&<���J�Ba������A �2h���%h���w[�6j�����ŧ�#�

�� _}��7���!(M�X�)?V}`+.��cP~<]��[�?�Ѣ�i�+Tx�U��ܱ���[I��`��b��
��x�yU������I9����P�_4E�[T&��)�����۝�Ǭh����ҵ����`@k��x��X͝m�����ځDO�Y�v�����f<��`��g����X�K~�t�7���(M�#{�d�֠J����ԡP�ݕ��^�(��œ�zP�-�7B.[���;c�aq����*����7m�m_�U� �yP�R�I���%S�z�Ȳ����%�t�i�6��5���W��ﷷ���5�����<��N�H��Hm��#�ѭ��(��7� ��4���u+�Ei��@=����A;�4?e@���m�'`Qq�(�}K�,�B��)��	� r#�����	��m�aj/A%#�Ac�f������l��P�[���GR#��^�;�0X���hY���$A�6`|��B�{�{��@��ʲ�B���q����*�( /ڰ\�ATZ'�#��r�_�T�6��G�i{��]�j`;NqR/>[b5G=���Iي����	6b��WuX�w$I.�Q?�_�e��b�ƃ8W�`����b� "�%��"����b��K̟>��Y���x��h]AB=]+�h�#D���S��X�b�ڞ��K��R��g���S��^E�:y� ���X8}h`��}����.sYL~�����;������%��iH��#9���+07�.ź!HM���7E>S��Gy{R�@���̡�D���o�K�q��:�����DẄ�	^�%7V 6x�$�C/D+N��>!=�������;j����`�؛
�h�s����4v��&��o,au&
��F!���7Ý���=�G���i<Ȉ
��\����T���e����6���,44���	R��*_����>�'��"2b�u	�E�L��"ͳ�&��N��W�A��]v�1�$�O���u�Ӄ���[M�CG�=���<�D��ղl��Hq���b��]7���͂Q�7��/\qha�3��	-?}X�,��"U;�:�������F��{{7}���.EmRe#�����Ɲr�U���  ����r��l��؍~��Ϟ��O�R�S����0��t����K��(�G�Ҡ;�s�[����"24b�jl@D��+�<�U���>3U��V��ZM���R���#͇�P��2�#������l_9A���5M����e�ǿ5b��V^���N�G��V����ww~��
%�8H��T����0�q�*^.�R���� �����0��f�����S��?���*|y�j����!�D�`�M�ĶkC�E؁�9�&�gG!!:4~y� ��2�}�[-�n	�C"��I���v���Ȓ�!����yOVJ
�4a!P3��JS���&c%�{������5͘�:�ť�7���~�w]x�U�S�O��G�o�:CQ�}���6n����F��1����s&������`�͵�|�"ת�YYt-���m����gs	?�@�4g���@N�w�7�*�s8��}?z�>#ƾX�����#�VI)Lؙ@d��@�A��دE�~Kf{I�ZW���m�xD�4+�V�?x��/�"�T��P$<u��u�^ǝ��H`;_������Lypm��Z[;��{�uR�$�Ēb[r4쵷P%�ZP)�$�w�S��!_�J�I4=��	/����w�J{��v�k�3��'T	��b�����	�"��!�:ғ ������Cf��ͻ�c3���0)��_f>�x���I $p?#{�3�6)�q 6N������xb��㹗8Ab���4-*�7]��u9�8\��{@���p�H������E>�*}2\�2��.j���+�zh�z:�b�h�:ֳ��`������%1�|�����u�)�ɽC�̈=b[�Ks�B����Ԓ���d[�f�<#/O�,9ЕI2?��3g��B�����E��*#�<=��۰^�^B�o�����٢-*Z�� L�'bz��/h.��k��փ���߻���܆T�`��~Jj���1}��=���oS5D`0%����V4%,n���ǹ������;[���� 6#��Z�D�K����X�r��)��.v,��2c@c�ii�bR2�1�Y�Пkp�����גڽ�BI`�=}؜qJ�	A�fiϕ����0��7�*����ꅕ��-D�<X@׀#�ۄs�I�{ԟ<�r���J8�6��F�20���I*��B�
�t��K�B��;}}�F�]:��~-�e������ݙ:D7���Cu�Jx��39��=�;�qJ<!���C�w~�|C�R
�(`@��J]ż;}�1�]���g؋�A����QQ(�����o'e��/�q�P�')9�^��ި
2-דW����m�'��h&C][~�;H^�Җ5"7&��}���w#<���Y��\��Anf��4�mpx���Y��pR#�\����^������]�7x#������,�4�Ю�_yܼ􄼳w���p���(�Y5��ז;��G�"�q-�m�J_�6a�N�d�-�.zP[�;��?�C�L�����j��H��~vw�P|Acܺ*�#�?l͹�ګY�W��|b��)�J�|�מ�W���A)3i8�z7�v�>ԏ��3�L��׌f/�7n��S�F��������S!���3�2%��E����1�k)`�`_�&h�I��$+�Mv��w�������w�L���j����g[��F�B�z`�ʢ�ح���o?�꣒J����e���RG|IK@B�����Z=�Ñ��hݔQ���
P�VU�p�����%;�<a����"���u����A��e�8���Y�e�43�3�S@���:��p��U�/>)�~�v�7��M�pQD[TfP��!�S�,xW� NJ��uDTo��0�F�}��ȉ��N�!Y�Bl@ȹ		��"����K2J����H���I�k)�7^%�tL2\c��ќiT�7��6�Ȼ��W���ϑ��s[>��)SY0H��@t�`��_�ӑ�ԫdz���W����&��~�Ye00wg�*�#7��6T�bM͟��W��9e�o7:�w5܋t�n���v��%V+(= ݁�!0Y����.�r�_��^fs�@zR�#��fMc��>!7���^)��rgrN��ӏ��B۷�0㻪1�-��yY#������;^�K�����ʕ��Ä�9l]�[4�<"8O�}�{n��k�:9���L[�R��V����+KY�	��/YE
�<�z�A6����u�=/-O��֯�ſƷ����'�-�'=�����9ccl��ܬH`Z�^i��o����v���6���b%6�2'90�y�	dUv���	��l�l��
���t��R^@�G�B��u1��`��l�����\�kՀ�h�t4���Z�2��&C )�l��\e%}z�Ѫb1�"��.��2*d�1;,0!�K�:���9'�؆8_�cuỤ��Ϻ�g�F�9=V��q�R^3&=��Z�n��ٯO1�q����]��`��/4p���ٓX�~���C����]�@�h1�n,q����u��P���?H�oJt�eWb	�Vue_z^f�IvQ�t)7Pꝿ���L�6��G��t����cE�HrQ�69���+�r#��=߫�*�8m�<��@�G{pI�<\�dY}�їVѸ�nx@�o�|���oMJ#���(�!*��*��ܭ\��j�ɡ�Y�3�����v`O���m�o���?�(��밟��le���r*�'~xqV�
�Բ@*oK~����j�a$sr}�{�a	��L�l��w��s�8iu�+�4����6 t����[#������G�@P���4� Y�w�n@�E���R�����)B�����u�K�Ń�oy+9�,f�$��Jс���N�����=K�Z8'3}\�
���/�$c:vgr��7^G���ؽ�%��Q�
ЖeK��u92��^�F+?��R���xuU�_�!�A�s}c�o�:�y��CF`�*"5OD%�ECd�<0D���Iaޑ֌�!�O� ��*6U	��ea�ߛ̿��;~�RC��q���^�}�n%����feJJ4�<Kxh�a��s#3͌�} Ҝ�zFdj�eT�'("�MJ�����c;��L�c�de:k5'ab�\!�M�q��i����]E�7���ˋzj�|�Ι>�N*-�H���a��ȈO����`'4R��~K܇�ZUҕ�^9�h�9WC�tE?���a��|�?�#��F%��7�M3�"�%D�̜����\�Jj]�V
�_��(����@��!/�4��'�6��$��Ȣ$��x��_L����s�	��y��Kh?�w^�K��)'�~�.�C�8������0�8d	t�N���w#�'zw����x�~��2G�;��}֚wY�7AzW�Q�����B�JbL�U��v頽V�L���%�؆��(�S��E�&��O��T%��P��TĔ����$�2x�T�y�Rnc���v��^�d~��0�*��, ��D�L��I����p²^���������8b�r�%�V�D�ꓠq�
X8q�>�(��7ed�C3�z��_j��0H_����:�Z���W��z��{yj���܃'���D��g.����޲�l#{����k��@I����!���r��(�ɼ�I۲���������%�F,�!;f�IJ���c 󺵞+��H��D��g���-;X���kC#�8d��Z�	�5�m�#�
���]^���^�_¥����� ���4e9%�Z��ԝPB�����O:�V\F^F	܈�L" *Á�/k*�
�Z���!+fm��`��`h>�}&c���x�43*K2�������Y�Q��q�>*�%�>��%�kԧ1L�7�g2���Ĵi�[
>5��S�o�>��[��,K��	��.��(�����S���X��A���Lw�o��sp�ϛ�,����s�;��o��߿��Kc��  �3$?}�8���"�5��;�*��&����9��r���W���tִ�@3�P"�����jh�
$Ҩ|��"k�zt��L�XY6�˴{	V{�(}�����e)�]�����\܀99�hw��8��yx�,L�ܲ�c0�e���L,�?��_tla�`ii�G;(��}�-I
�;����G�b��ݲ0��!3�)�V��U��@��a+�a�v�>k'��ei��8�������AqZ�J5��38��ҋ50�>LT@����F�{!��t�k��_��n�'�� x+�W�P2W;w3c
�G��9f�2xu�_ ���ԼO�ITzR�Y �6�Q 6������h���K����'�(Ua��\ΏE�HGj��_���,t�π�����Vx�]k<�N�.�lN)8�j5�ѻ0��c>�vi���T�8�ʌeY����x	R��$;�����*�\�+�CJ  �ttS����c�"��#�:yQ$I�L�h�#)ըL��:�΀�'/��L6�5�J�r[�:?2�Pxt_���P[��8\��P���#%�fH�ġ��M���	�W����/���7�\�B�*c���O����q�<<!�El^s!_t�{�ɫ���|��.;�$۸�Ѹ���ь��Tr �[�ƚ�mC1���Oˡc�����)^�#jr�|2����~T"I C"d�R��ڪ����0�ca��Y��ZU�����N	�Q����v!@d��a�٭�!���|����^9�{ol�>��1J+�%f]��B��&�1��H_wƱ�IP�R�!��?�\qt�b��#{�!�L\D�����}�b��q��8:q��.�נ�Ny��*�,�Ҕ�����H��O��-�#��|8#���q�xs�zQJ����6'�,e�$wf�6�ӍN����sD����V 6��'ĠT�O��<����[�_^N�ϫQ` �2�d�F]�:좋%��a<��V+��V�p�aH�f�\��P���΍�����7HR��j�Z���(�!$>bA�g���z����u�!#��L�e����}�����7
�5�މs{5~9V����������gԕ�ղF�;1& ����18��[�~`��h�:�Hg鍾���8l������<����i���rh2��!�K &#;�sҒ��x$[ �U�b��:ԬGz*�V�4r�j�@�ڕ�@�♔�	��A�p�D���՛`s�s�����س����4u��2�J�^��o���+���u�-��h��7� �ep����:�u��ӆpJ��Q�@p.ٝU�o�Wxag���b�}��
O_� �ܠ�
i�1{�����nw(�7���EV)nv0�R��`V�>i��ӑ&�ѫ:�x׮��~д��_A3�&�Z�#|7����=p��ȿ�_��A�8�x-1f��$\XL0�	=��d��V#��+�U"K^5 ���v}��hR_�歹������=d6�����;��R�@Μ���U�'�����������@���wk�?��B��g&��~a�Mr�*��1z����#�)�����F_�E�ƙ ���~�$K�E�Z�E��^m�F'؛S_�
,��$/�䈸9����ˣ����z2� �^����3J�>N����B������������_Z��;΄�����`6��C���OA��c�-w@֠'2q��h՗�z�'\~�U��+q��E��������r��V�9m�(��$�����jD�"ji���1���[}�Ư.	�p����%����Qa�-'�lQ�1�7�<?m���	�%}
:o>VS`�K�
^��k�4
��ze ݕ$�8�n��G����J��e�Wb��Z�Q����j�j���UJ��*>F��G�t������rh��N⼾>|O����e�͆�� ���{-_��ok��}���~���Idc�EzJ��o��S��AiL����⏨1��I3�Z�cs�a��A$�����e=����u�����,P���Tݫ�+'1	�ͭ�Fky��t��E3k�c�Q~wvNpH�w������'�"����F�)-,��r�{�C<"l�EA�h��-6����E��6�%y<���v^����x��|���\N{R�~��p:ǜ�gl4&@jp��^VAN3�	١N3^���#W��naC<���
e3�t�p�J5=�X}����%�v������ΏWo��^y�^|9%�����=9����4�ړ9<ǭ/�z��y���_u2ww�܁}'0�0��X�
�)S��7Hh�6�p���Њj��E�X��LDcΣ��)c���ٴK�BDt�ѷ|6����Y��We7�6��]�9���6�/�0:׻ӛ'�O ^��:u���*^p��y�hR��t��x�4�ؽ��q�'j�Ɗ�B�EA�Q��o�w�ey��VY���aQI��/��̅,fw��mt�g�pB�_���_���J�kA���َ�ᘫ.�7-;��B�X��|uHh�����.�_:�U3nY4��H����7���Je���7yU��k�lq:9��0䮦��_Ò{����)Z �`F��6O_G�	GL<j@��J�c2�☈O�`��\@x�E�8��]��{P
g��gB&�̠�|����M�T,7�r~=N����~!�I�e�J��1eao�!�}���[�;l�"L�/�l�g)�"̫�Q�Eŕ�y��m�&�x��� n��~1��O���\�꼧_V��Z�\�
rs������!��]L�1� ��c-3�Z�� �v��#Z]��/E���_���']��K�I�;�\�6'c��~�FO�ZsG�1E� ���\�7Ď\xZz�� ���3�|���1����B��轙��r��XE+I�ug�
��N�}%*�Q���u��U�g��N:���w���I����2Bi$���)�^�>�K=�D�-"O��|J �Z zɤ�2��� ޏ�f>1MJ��I.L,0�� �SJ�D�`����� ��x��V�#O���y�u�t�8[��ZѣD�4����'J�>8�W��fK��9��# ,��:)���q}:�&n!ͭL>�$�5ZYB�_��&y��s?��ڟ�pj	qǀ� ّ4}��J���:#
�G��X*,�:| �[!�S�fN�Ǧv���?|�4����S���������B/f�װ�Ã[�7��y\�=��٬�u�9����� �#�/<��"�28Rol�@4wQ^�t]D{�겙�߲(4�+M����S0:eAB߇���e�~�V�����&�R�R"зp�6c4m.�3oV� B�u㙢'�A��x[�%fr?��{E>�����;�bmа��˓-�A�Ӫ"_O�ߙo�M�n�r�B�W/�"v�j�Ǖ�Ew���<m��a�Wf|d���7�m|�?�q��&����L|I�ڬy��"��:��*U����f�}��!À�'}��<���MN���v�b�ڎ�O�r&�(������"?�/��Ar�O�p2�=ud%S\N�����hc��o|L
$�$c�%*K�d2�$*���9�do ���NnҞ�ӆ8������r�ן�Ր�P�I�r��������0_!��(���jKD~���~�J#G��-vL�J�j_��;S7�#��ldyM^᏿�?�I�e�%����5g����TZ,�P�8K�ȏ��	�/��+�b�	i�ֻT/��	��/�fi�ρ`�t��B�l��Fdg̛KtOau>��x�V�P��UhMP3�|{����P�}�����P�F 	�u�Ͳs�vS�T�[ܰh"m0�'kE�x���������g��k��=*��+��ML�7]�C� �ZXz�6��c�brC@���wq�N�#�Lj�����I0��Ӣ*��a�� 4qػ��FY�!�TӒ��o��1@�@�m(�{�D6��x����� ��yM��X�ᩅ|��l�hw
x~$M�Dc���)�:$��Ȅ��A�Cul �d��E�26_�m�h2�L̵ud��;dW|C�6O䪭� 19P8z8tG���ua�C�} ��5��떖��N$��r�c|K`zV�3�Y�� 1��ӂ;��bװ�0� �A�����⋂�7��x1�@֠���:�0�AؗXv�U�ǍiyD ��W/��Z���⢜��%�[��Z�^�/	p�ӣKJ|[z��8	0�d	3:YVwj��F�At<��"b��-��h>F��xk��><^`�X8��8n�ظ�A�"����$��*�zx w0Od�ײ�پ,�D�.���7�� ��*A|�M��7\�0ـ3UM�j~�穓��aR
�j Ve3U�uqG�[��H-�P�VGY�R�P�����ۮ�*[�z�ݕmc@=<y�v��C�!�~2��LNЬ���nV��<��&B�c:��%LQJ��"�1���i,N�]�H3l�K2x��_��U~�Yܵ�EaP��?���7,JUU�{9�M!첬S���B���{|ޟ.�6�����0�CF(@�?���{y/23���v��@§�m��� ����7;���7K!,��A�E���]�̿w��`x_�P͝�9��;�ӼeƟ�~:��^ѕ�6��1M��s���<���h*�ů�C�0p��!l��Ȅ�i�^�����B
u�^����>8&��~`:��Zs��	2�Fd^]���_��w��o)��H���ۗ�;�֖�%����O/�>��/�9u�Cm�-�ݲ�96���hWC��{���##������s�P/͊�Y�Fj�U(k��a�S��IrJԄL2���Fl�~I��^8��ƀW`����.S���r�R�
�'c_fan�O��lW���5yn-Ƙ�(����9�tMP/ڻ'���Ӛ�\~ǯ�{m��Y�$�� ��fO�����X%Gh��y�$��D�pyF%�����@�.	�M�J����Q@��LXS��F�8���&�����v�m�Y4ܱ�����4�8����#��&p��{t;���:$6�u�@���f���y��p~A6	�#YY����QѽRsBZg@�
�<�5�}����s�t�����0�Uқ�R�{����z�M<<�Q+�\�l��R�:�B~tt"��/��k_��,N�|ӝ�1n��є���Q�����ʻ��I��÷`���pi����j�OB�B��#A���qB��4�7~�N"6��izquFQ�UAa�x�˃NdO�?��!�{$c�@��^��|�]�>�0d�P��3����1��C}�0�<���{=�7�}=?����������?>`C|�J��� ��{��reI��Z,A�`�&��`E��,�YQ�(���Þ����h�9h����,ZS����>Sh��#