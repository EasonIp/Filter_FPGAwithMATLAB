��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�J��"4�=�7(�T�JѺ�ő��,\��s���ӣ�F�؏7ޑ���L���r����C~��N�[ѫ����xE�/�&n@O�R� �e�ߟ`_(���Ll����q4^�,m�K���ґ0G�f4<�!�#=cZ���3��QIzR����2[���7�SP�Qpz��xT��5`�UG
��Fr�V��.� �5sF�����,�UF�a��|c����O�����p�Uۊ-m�q��'�\��QWEJ����c��x���J���n���p\n��H=�!S��t$�,C��-��TNH̹�,ytWӞ�}�B�=�,��e��=�[=�˸'g�tW��9�Ş��@��M'�q�v:<̱N���8t�i˕��x����i=N\vy?X!�&Ȗ�l�ts�v,xĚ�{H�&H/wȘ?3���"�Ucq�4m��'MCQ�l��������b�~惪AM?���ע?ɋ�k�`�����r�Ԗr7t\8�G����L�H�����L���.���6��Gw/���L/u|NN����;p����5�%ϵٸ�l~�Mޟ���	P&�Cm�Dı2�HP7����g���kÖ��w��#4����]���a��W_���[�޳�(4���BWo��٪E3P�`-j�lN��j!y��=�{E��v/�痶�I�O������*X��*2x�"�	3�{Ɓ��4�P�6}��J�<%�"�� [q��Nћ2P���yj�i��Ԑ�J���Ϗ^C��;�߅Ý�:':��su ^L�E��.%������I�ʛ!ǻ��h�3+��9O0;^�����O{ƿ�|��j��^������aLk��)>���Z�)�"�q�&k������SI������\� $��:��{�3��ҐT�]ቅa����$��'�����|�3-����5� +�&X�\K�C�$z�7Z=<�RT���QQ�_#�ֱ{B�56�Hv'4$O$��baI�{l�7C{Ϝ`�3W�!�cnF�<V#6�7�ЎE�'�L�.;^�t��삂懡ܾvL�J�KH��j\�-���H��8�[��7<�~X�/�.����Άm�{����]�hd��
�4���8�?���Xɥ%�ELU��.��}��E��yŉ:�)�=�Q��w�`�J쐯I�V�:�@y������w� ��gD�,��Vg�l��6;���l�X>Kq<���U�"�����@�`������'��gnc���"�b������uW�{��h���C��ap���.�R��ߘ�1aU}�k�,5�L���l�Q=!�u��:]�fHň]����Gў� �ö�,�&X��6�\��9@c�{��j�Y�t�j������q�j�4��e�Q�)!�R�4���HS����m5Uλ?sa?V�Da[��$k�:GLYkN��!��<�w�F5k�í�g@�	�<���^�bp���We嶸XV����k]��_8b�b�	�B\V�$��4��JR��A��x����'n��P2,��KBV�uԿ�n}�����{qu��Д\��МV���'0?^�z�c2:XHf��)�{�����x�&�y���1�P37"���;�V�%Ea�xA�?rcM��&vs���W_����Gr�xM�:�Y�ұv� �{k��~�#83KI��g�p�>8dB����G�so=��]Gĵ!������>�������S�83�Ͼ���l��	�`�_2��J���A�Ĺ����3�3��z�Α%���P��2m�M�,r����m"�'��r��,*������nF����Q"_ψRKIf�����N߄F�~��-�0@ĝ��:�P��D�wuH�����dW�5t�m��V��eW � ,C=�)�D7#��	Y�hC��� w4g<���Mt��cW8�'�p�җN�V�L,�Y'�1�⽅qyǹ{�`t�{Ѥ!:˅-�2��Kn{H����ڵ�ї�V��I���k�z�d�:��9��o;�|�󸸇����dV�HS��P�m��z�����,7�`Iz����������b�V�[r]�C�jZ�N��&߷��J�P�KD�q�8ɷ�|Hc��
�r�4up%�cNr�ٿ��?H���`�0%�����g��]9(�I�-v��N�Q���}/�_�I~q��@[1zKQ�#BU�B��}#;�S�Ju�� �F�w���,����3�J�Q���(�Z�>�ɜ���y6X�{����rN;�����)6�x���A"�Y6�ِL�����f[%迨E{�ݤ���d�h��L�4,�9�g�;'r�Z*���0Uq��m;�����,I�����+����8��p��7���j�G8���d��5�����x�]f;��Ҍ2HZ�w� ��T����a��QB�ǻ�ǻ��^Ug���7T��+���wMl�KDbe�;���Ӈ|�T�"��W��y�ݏz��H(���2 ��{��s�����t �zeȳB���t9W<U��N�+���W���w�t��c�c�c��i\�R<Tu���
�"ʣ�m#8Y���˔�6��/®Ő\)��2�Q���$�)[L~PIQZ��|�� �t���<JGH	;��ó���u-���8&�,��k��(���d� 3�q 4�n��sF4����$i�����^��Ӟ��Ͽ��׍M�gv���dGPGѹ��Z{���=��Ɍ?���[�yh�ܯ�$Ԙ�E�����*��<Իs���oޏt��D.]�T0��ژU�bUL��i�+0b�bo�*�@���3�B6�&��h��#�o4wJ����,$2V.��m�fc��  ��]�5�d�����I�mr�)Gj���}!R�	�ѭ��M�$�׺���O��)��(���d4�K#T"�F��'#��K}M�$��h=(5F���Տ�!`��I�8��o�����\�J��n'���
3rԾ�-$�}\ޥ�@�+Zכ�H�N�c���;a)[
2����'�!�9�O��W�	f�i��{;t�JM�脦}-"�kɏ�R�����j� 8uʽ��O�*�Pw4��͓�L���sP�!�'
wH�e���7xq�)\�ۢ7q�^�<��hg]��\�/R\�E˞	��21)��C����|tiʾO�5s�|���@�[�����a|_�e��Vdq�	�hh�+��i^΃���/.���]����}ߋz;5�<.:�da��b>��,<��������p�ʹ���nuo@}�Fd-7��=�/����@/��f�%�!(�)��@w![�O��^�d�vs8@
�f?~O�WB7	����y�ގ�׭l2�
��O(��,k=��b?���(Z"����Í�[LN��t�y-�6�4{�a,��pOu�O�lOEhK�t�wi�Ѷ�E0Hl�1�V�w�x��O�4� ��cf����9�ф��C��[Ȑ���f�Dj���;}^�ɻ6m�_>޴�W���<!Y���(�`�i�����yR#�Z��H�~�q���J0-��Eۛ�r����k����:�)��z�����5� &ŝM���c#n�G��d����r�;Qhf��s�/Ű��IX{��z���~�����'2R��/Y�=�Y]����k�������?Ƞ��:�ipL�l�"
-��Cv�l�=��
���y Y��!O�}��FH�\7d�����0���|���y���Q�~��f�1˧\��� �Lj�F��L�y��-:��V�q��%�(P�Q�����Թ�'7������>*�,_������I`c	;�2���������N�5I�c�h�(�J�ڣ;�=��ߙ��b�'��=��Z�3��^�����-��l����	���F-Y��S��J}��)6�B<����$)��b�E����V�oU>���&�!��V}���=g��3�fP0pO�L�Sf���M2�b�#x#����b��B��ݽ�'��XF�p흛��`#d�#2�'|�9`���nꛜ
����d}��O����(�_3մ8��u�?�Nr���,��4>�:�ʘ�T���ٵ�yf�w�۬�f1-,��T*:��F����_`��n)UU�d2�#�#8/�+��!����;�ڙKfAw؏�.x����4 ��@e��<ɿ��l�N���e���jF__�T�T�D�g�L��Q�ho��qq�����W�
P<����_G�̓��JZ�\M=��Y��
}/<���o,�ګ݂P��,
o�h�iYyK�5_����ohp�mՅ�6Z� *3�MW�U@t�O1���>�o��,�r��F_�=ʙ�}7#�u�y�#����߶]���Y=��݄%��g���]
C`���]̨]wj��5�C��Y�A�\��ح�X�Z� -�;,�R�����lQFP;)���l�?���8yN���� L����9?�Z����~߂0bV�e��8����U�IûT]up��J�-N�:i
���=�Η�����d3�ɸ�� ����w'VG&�A���>�}����u��9����xMI�<ę]�����,������R���$�x�5���v7�ۚ������	�ڑXo��%eV��ˠ8��s4��鐚Y2���/���Kм�]���R�%�������<gli���zz��섯FK��@���z2x�O��Qn#�x�b��Yp�j\��9��R�
p��n��vU��}�aB�u����L�X�4�&>���n�[���䤀.���*�M�����V��a���	�����t+��ͅ�k ���Ԟ��E�F6���ߓ__"|9�����1D�Z�'�F�MM��%����g�U����w��r�����8v�=*��B!a�%�jy�Z�H�)�z��s�"㌴�4�n�6E� �~���4�x�mr:�fWq�����6S�t�F��pt���bI�~����<��$�	��a�����}�đO�!��!���n��^���J��J�\�02r�	��nh���c��G���)��)���&V��������w�=�L��y���H�N�Ӣ�m?j5$�=��_�z��I%��-ӣ�y�w�3Z�p�]�0��A��$��!���DS*,W��H���*��vZuu�R%�� h�`t���J��Nu�2��
��+�DJE�4��tf�^���9!�����E�	�ν�����R;)����25�mv�eޔ�~8U�ƭ���P�nM\�G��	��?��@>|a��F#�e��E�5�p�M��]�G�Z��r���]���1�h�֏N���XGx_�U�A��+��	uӥd�)���5��&�DW���3��b�Qg�a�
�n,�w(e�U_O�� ΁:�L�C
b����J�ٞ��{�Ժ0���s�������=*��Z��3� �Y���p~����q��J��u��ϿYzΈ�x�"#�*�ҡC���*�.ь�?���`�&���ܟz3m��#�y��"aZqkV������N��mq;E޴�>��O7LÍ�;��E9v�A��%��l	��.�E����#�27�v��w@ž��bzk��Tu�O�?�XG�`�@�{_Z?,�=��ؚ7G�ͭ�Q��֕�������� 	�T��c7���8^�RcsI+�k�r�(|~�K������dm�l&A�+��������K��SoX��]^�(+�����,i��/�%;X ��p��:�,_����B�G0M�5�`^�R;5;�P�l���������`Qʚ��FV�4KvT�VQ���n3B��}Ú���FQ�v�QM$H��a����2}��U���aT�bg���un{���70�w���<��oK�Y�������� 7f�N�F�p��H[�o)�vI���1�.����B��y�Q�_�`�2
�Y������ڝ�#�z?fΥ\�db��D!-�N2I�ȁۙ�[m*KJ%y�q��Z&��lD���c\Y�JnV����$�v.`1�g!�ޣF�}�~�J�֣�
�ꐎ�����
8č��W����͋vg����|oBi�a�[dš��o�Q�������+`H��w,lO}\T����z�������i�Ԯ�Xh��5\���ϑ�!��p��R��x\�&6�J�t/�Z�	-��^v�2��y�,��[[y���
�C@e9���@����ӧ���t�鮩�'�K��2QJ��>�P�s���f�&�����pj���^7K�Ũ�갻�ά�9E�%G����(N`�-�<ᅿOo�46ƕY�I����Xu���Q��}�r�Ҕ�T�r�$ܩ+��R�pq�ٜ�ҼV~w���֙�ۻ����ߪn1�Hy<�Ճ�<��Gd��(������ˋ�ȯ��'���k�:[�2$�!rk��� ����r���r�E��S�BP ��Z; h����,%p��pι%�z!��[[�R��w4]�6|q�̽�(�g{��k�l�E��P����j�ݎܣ�㒸�6x��Iƴ�W��Z�@�15����R�ڷk|"~4�0�(�٬0Ro�X*�^����۟9�!.X>^Yz�j�P�w��V�����=j��ݞ���-rdr�Ҹ�GN�2���W��p�~��nr���v���Ԗp����Y8�Ia���g�Tt`gr5���%�[�Р�$]���ݍB蚤�����0����c3�qw�T=���rO�`��N����	�@w%1��F�{3;�ڳTl����`j�����ٜsT=w�4�� �>M4�'�IG�+p�?3�C0���F��c�Uc��z�y��9�����}A3�7B��p�⇸�u(��!*,� �V\M�Ȇ�K�9%�&����]�S@�����]��J'�,aE����T���Q��X�h��	sM��%��q(�+G�>QH[�y�o AUcsL�|j~@�O���\Y�M�h�XE}N�/�/4�<�^N�8�ɺ�S��@]%.V�,��`�`S$[?�{�=_���.�j2�`%�@u��P�h�0�4 �����o�;%��뿘�������]��3�xl�R�ĿH'*�^ҫ�m.&|�1�!��c�	��\�OD+����+��P��D�?�V���� t�")j�'�Lr���H��X��v�I����N��a���k��y��Vs1�V����;��f���x��ı~�f�̳u�MW�����#��E�xG���&Ϝ�B��2K��K*lI�)mh�Z��V��� hAj&��