��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������"0F��}�h'��8��<���9���-�j����,W�_/�H: 2���x���CH�^�g߹+�F��0�tw:�j��{�)�0��H.�'�[��'0���ck�D����L�Lq�&��IzV�G;]V0~ݭQ�����)�47�gP�ILO�"���tAf�?V��-8�/b������$�9~�
�l])V�"q��&=��b]��[��rL<�\��+��1:����Q_��!>5
9�͖RT���/��Ől��W�f,���th��sC|�o�lԾ���3I�*�)���l�넢�}�����'�x�nM�Y
8SE0����K�!��I�C3m�G]�3�����v���:���fT�~��g)�������5-�& k�9A`Y�	���ċgB�yF3�mӞ7�n|�s���s�#�E�k�䋂�1��q�ѭ/�d;��АZ5ib��Ku��e��(�D�u��'Y2��!��j����s���{���F:����t�������fL
#]�ݮ�UTD�5�;� �]* ��׬�m�Bb�q�������pW7���L�_#Z�R�'�d�}� �x��^`[Y�j[��-<���[����F;	sֶ��i|~��/Kd��0z��1DǢ�7�D���I4E��F`,�|�3��
\aaN��F�2��z���a�'2����tF�N6X��/��K�I�����HAQ5���0�]D��>1���zc�k�{,��b�@F��f��}�9K	����W:�g��CԄ�9ٛ?Zb�7�u�ɛc:;.�U���	p@�&�Y��q�1`杘OfI 1��ٯ��fZ���Rc��x����I:5�)$V5>ǝ�i�6��Ϝ��(� F�i��@\��EO�����P���X0�J=�
��t)Ga�����^ޯ���5��n�i���1:��/��1Q�p��񘇐�5J��|�p��;w���j�xO
� ��k��Ӵ�EI{����(�3w^WAC�����W>�Ux�#�6�U�cB�H�,�-�Oj�v�k��k�kY�J� S�1��T��}5�1k��\��ܲ����\��8�`t�	��&D�O�N�6A9�9)�dB缯�B�3��ڬ�5��n.����О�;��i�%�
cC�H��V��ǇQ�S�����m|"�"~5Nج�6W�m�i4F����y`���ɧ�?>�����p��S��}�J��;`��`��rT�Ь�M�(����?i'�'b�nS͵��?N����f�-Q�!�D�zq(G�#�փ�(����A�xi�xݨ�ޙ���?��Q�$꣠��ީH�K}v�"�Ҍn�~]���Z!�Ї�:�m^EB��mE���.�爝�t��0 /u���� +�����~��Z���80h%5�hj�۵��1jZlR'�`2��:;)d�$�Dy�Ii$ۀ֠<��N��mn�[ �J���%ˢ���n�~�(��1�n)�n�PVPi�n�IOʉ����(�u)V��)%�Ъ=BcG�z��^����B�S�(�<.�)Lf��>K-�ѲO��R�H��������r��JS�]jp��s���E2J9B �<u�4D�u˲�� m&��/�Y�~����ם�Z?4�Y��}�|��j���t��(d_����e;9}PdH��~<��yR�"g�����֑�v��vܙ���Gڹe\V���5�`GT�^���b��RS?k@Wvfؘa�Y~�w?|{�thl�{���v� ��좝�ʢ�h�!ߙmsC�|����CN~���Q�6)Q��
D8|Z�^��*���^_@D�Z����K�oT`C� �][n�+�o@�Hh0p
�B���KS���Q���Ʋ����$[�!�?��&�
@�	���m7�h�̜ћrsG[�^h�R\Fo`S� �:�Q��I��B�P�J�[�gk�/����.�(��o��X�ς��x�jK֮6Q�Y��q~��Wz#�@V�?L4T>���%����i���jte����++�;���I���Y���b�l4[!�f�f�me��z�0�c����w.4[���Fs%�!��;���Jz�E폥m���V��_Ư�՟[�)VIkL%��=��2Ģ��� �`h�g�{���mM1�a����_�~dC~��)�9:��F�%*���x�qw�"=ck��x��:r�d�	d�&q_ޙْ<`�@�e��ԍ�P��}�Ǻ,)���Ҥ��1&囦
&_m�~L�O���B�-�j1���㥹���ɉ���~Rx�)�,f�R�#�!S�`JK~�i̲)[�����X)d5g��x��$L��Э�]�4���OmX�Pcff��d�$r�����~�Ĕ\��5v,J��TLz�ز�u�TO,�{C�� ���I<�)����Г����y��_Ti1©��	�ć�-�J_ҿ�nz�>�Rx��ãΆ�y��i�8q2#����	��o��[�_��&��Í\�J�;/���)p�O�~e؇m��,|�!�����/�@Dg�:ZP:?YV�' ��D}l(k|BD}����|��������C�3 �;��&��C짨���������ǹA[�����:0��Ó׹��A��(L(l���m����$:d!���_�D
�5�|zH��Pس%RR-�mrX#p�aA�Q�ׄ�u�i��4:qR��c�qT��D�5%R�v��h��#�Lߜ����}.6��1a���{&�c9�) �lXO�#��k@UL�A[����4Hʕ��D4�j��K��K��G�z�4�TU-���º:�*����"@/���PFXϩ2�9�B�N9�:gp({�^��fq؞�����C��F�B�_;A?�f^L!�7��pK���4y�*�:�]s��gE0%�4\�o�VZ �EK��/��]7ek�/X��T�-a��mh��^�wv���*�����j��N~	Y�����A��3?�v�J+W,И���g��t��r�p�P}3���j=�?�UJ��+�λ��tkx���l<�9��\6�)�C7�(o�V��M��Z�lR���ys���=o�x@�
��+����̌ҙ}��;�Ij��ɆE�V@;�7�(+��O�GX�E@\���Q����!K�w��}�?���g @��t�G9dIW�@9�>̌^E�A�Bݒc�e��W���]Mt�<�Vq{ϱ![
��<C�mq1�J�U��L<�i���ƚ�2:�E��˯sl��o������Q���CR݈oC
J�k�=����QZB�����D`�#��s����_�|,U�/ _�en��|��䬉f�X�/�H͟�⟼���5;�=��v7t���z��~T|hw]�tJ�YK�_�cn	cS��
��!\9l}�N�Z6WX�\4��汝b2Bǂ�J���P�θefm�x������@Btv�A��G6�%w�V|�j��}����[�T�=�F��OD�.�
�p��g��p��jZ���9�U5C0T�N���{�4�K�U#Z���K�ۺ,��ww���ava�����1(����r����:w`�$ٹU`�?/�}��i��:��Pἂ`�ai��cH1k<��'��v�����!}��4�S�Dn��%K�h�1A�yð���L�BAZ�^����rX��$��Ē/5
8N��,ɔ��t��8��5K,��T5lx+�����uSS��nrsy4��"7�Tx��^��s�+�כ�콠���.��*>c�[��Y( / �:���8�\n�KZ8l��,m�[�ĴO�L2J�>;���=J�e*.����+�,�4�d���.B���b������9S.�E���RJ�.Eu4x��>B���Z���H�wyߌ���i���^بV�fu:�6s�Ms�	j�W������c�H�B[V]{���Ű�p����1��v�5�Wy���ܾͳ���p��X����3ǔ��	tֲ$5�TÇ�pTD�?��Z2��5;4o!�a+�ȞT�!񣭱�#{�`h��Wo�Ttq������:�D�X��U�4��A�<��B�P�Q�Q)w�3]�a��	{�0yC���o��G�h���!���V�Wϛ��G�R�)����\��V���bB{�_�1P!��E*o��v��(�m�H8�r�����THƃ��Q��f�~HbEQ�����#�9u��ǫ����^	���^��%�R�W�sT! ��$�q.4����˹�vMd�� \�sxzD!��!��k��Z�S��5�$f����q�/x��̷w��el6eoƃA� ��)�h�X
rُK�GH� 8Ŗ�XM� ��HR9L�HK���-���l��W�+6��ŧ��	ڋ6��G��Y�W(e�f��W��I��p�[��1��l�&˰(�`{�Y����Y�Ba�p�)ϓn=�@���e��

r�{�+Af���l�BꞸ�$Y��n����ƭJ7 ��A���N|V@O�~|בI���hG ����u��m��5��;��d"p§�JaOn�M�Yo��z�kzx�!�9�C9 #���ݧ������ȧ��O�?^Xt����/�^�x��/5��f,kY�K4�"���u�pgP8Ϥ���S�	��^�m�m��)�8myO���|��T�'�OoL��M{7�C`���|������5r<�0�>!��kfH!��
/�f�.>��4��p4x0$�:���$�+��r����Z���k���a,Ln�H?�ν�Fn�扂 ��m���2��U��P'5t�6Һ��ϱq�JY|�/�޿�݌��:&����3*�`ݞ|Ǻ�0��aa�gn��V� !�]�Y/�����7/ �Jݭ���P*nt]Z;I>��w����Ь q��$�1����r'�6~�X#�&�$;4����s�r�L�K��>�-jEU���S�'��Z��K _e��-�K/���#�h�H�w�BiK���K����4�0�c�_��܀��yC}���h{`�תVp���T�����l�v��H���'��H�;&�������o��;����ug�yh��
-�*4R��Ҙ���Кk�Y�{�~������p�!�t�M��?E��4'o���-U�������wfo���!AjNh�bxu��֬5p�jD_?pp��� 
{����p;�O�<,D���� �n��2zS<(���5�u *����ΐ��N�W�	ښ�` �f5�3|Z���G���Q���m�>��]�s�W٤F����:
�)�˧������>1Zi�%�{��|D{`���ʥ�P�h[A"��\�[�!I���I�~'�l��H�)˞w�=嵰�w	��.��3������L�D�W��(�T�(P�Yqg�=:�+�����5�*�{!i���0,�x�H�iz�-��stom���ޥE#a����s�.{<�S��1���a�@���s�i�1� ��w<(�0���:��`�`�⊠)rur�� �Z= �)�&�q��q&�*ó�&a� k�Ѭ"�Aj��)Kç5�-UĬb��絏=�6�����v6r��{qx��Ub-{RB,�^e���_?�����51N �Ā=�����˖�.��љz!EF(�a=1�UT�t=h^��m���J6s(ˡN�����>S6�49Q��j��X#���v��� U�{n���rF	<�)�'�y� eV>%)T4j��W��e?Hȉ��� ����4J`�Y�Z�8��sh���R~�v�{�����V�����z�����w"������Ҏ�^�l��V�*@�@�a%:�Mc�Rw�!�Ѐ�a�����,3�lu��F�V^j��[X&w27���}�ˢ�Xx�lپ�Tpu7����i:z�B�K��`�%+o����y�˩G�{F��0��n�	�K@��>�lb$*`�u��B�|�e%/�R�S���/Nշ������uѷ�}IY^�^��y�0���l�x@W�k4�(j�����d���IN�"E�������uk��CR��E'���z���L������޿�����Fe�\� �F��S��m,���"�G[c�i�W��|��jN|�~H�q`��=�8_��l����^}d'�C��?��R��Y<\<I��C��Rx2q�c�)%9���CS(�@�Ɠmo�W�;失�&��YD��}�Iw�e�6R+����k8�M۽B�_�T>�#{8Q3�dfCԯ1U�4��҈����Rp��خ�/o`�=�g� +�6j��"��,݃%��i�4Y�Џͻ)�o��� �J\Mh%�+r��^�O���N�آ��m]5��V�ЯQ�*�+Ž�U+E�5�[����]~�v8d?����^�����}(�g�S�9BJ�V~������ ���˸�(�R�5��!L�_Lmؑ�>��0����P�z� n4!�;:�q���?���'������q!��(��ԕ���mft\�,�ߑ/���_rp,�>����E۵��d��f۞��G��HK�� i�t�!tEZҪj9�����b���1�N3�*9���b� Z*�����p^WS�芆�|�}#C߆j1�X�׬�L���q}��GvǞ�EIiBO�6����N)��I�f�ʅ���p�b#�)�w�ל��'}g)�mZ�M�w,�`��X��/2�?]��fo����1悍ZK�bH���y������w�<������O�N��)�f�������cԺ�GY�2�,@���K���DB�|؇u��g�FC[�Cz��cQ�mW�[���8H��X	K��"B�H����T!��������.�y9K�m ǏeF{�O�zWdt����k�7��&6�O�n�W�|6m�P����mRNY��Yr�,����\�8�Yh悵��"X����>���5@=����3�6��s�o/�&$J�~E%��0J�yp5<�?�K�F!��|<������ո�ժ/@:x80�s�����MR>���+F3��!�AAm�!��8̈́!���1���@~EsiGgϸ�>�b�p;"����a%�x�Q�q�@�+�|��(���������.y�	�F%²�($�݅�8�V'a��.Q�����{�_D�]�i�����֋˞����v��������i!�E̦8-|H�^�:�Nh�������8�L���H�������)Բ�`l</ܶӹN��6�h���ЂO
�Z&�s�ʖa��6ɔ5��#k͞��@�`+�k�_���� �J�}��i�w�<E�C\pi�G�X5N��E�����%6�V�J��d�戓���PC &�\�L��g��. �M�s�H��L�|�����K9��ݬ�2	������z���|f�2v�����/�b�,�A@-���+�'}z��̈�7t7���Z0џ�ksbHN���/U'k����5_�<u���GAэ��K�^�޽�0q�eWe�q$�'�7P�w !�ر���SLhf���I�V�Mj�9�=%u�����q.�bXJ�S�N��m�v�ꘋ�\	�8��aU2�̡K��?��4�1���J�73n���DE6�u2XQM�(��9���c��_�:{q/��H����Y.j��I��Ϧ�����t�sH�>%_�	�x�w&>��o����Ceik�Ʉ�iD��8[�z� �Β���]��lY�J�Dy�w�N}�r��@���"T�����8�'�b*���|����wet4Ӳ��O?��y����ō�]=z9��c�ka�2�y�e]Y��~Cs�ԇP͞�x�fj8?a�$Gc1����:���V��jõ&?3>>�>�(�z�Rk�]�F��E�����j�3A�KV[�yL'!n��h�&��F��rp�~�����E�G��)qI��$�5+'T*��*p,��r����� !���hBV�	ƎɃ@#����t2��.!��[aG��� ʅ9X=4���ȸ����u���@����n�%�'�j��5��^�)y��Hmǩ(�W#Z7�9�0���dn���ـ�sv�b}�ɺ��GC.P�ӑ�o��Ki�������@�Z���1
9�I�Cg�D� }D��g���]�����T_:���)!��0!��e� ��K�xQZ��A��d\g%xV�ȹ�Q2k�zh*���"�6b [}���� `(�7����|2m֡�j!u�Q�S�x�Ԍm�O"z}���mD�����=-��S�Vr��O=��gUyygJ�{����V:DE�j�#�����J
݆f���w�J@��p��;p�B;at7�8�G���-�.�� &�;��(H�Z%&�L���W׀@�͗��>�<�W�,���f��?��bEz�P�V<^e��:�箭?phqutg!C�ȓ�h��M��ϦF��ئ1���pة�P�R��X5ζ*Dj��Wz)��l�(����(q%�B��,�G�,N��ʢ\@z/+_mV��{`��)�<C(l]@]6h\�e7�>"�a9��5�ƥ!�W ���;r����'��Q�:\��|��Bg�0�C�{"�c՝*��8�����x*���WO�QB}��Ίu�������9�pH�Bv�X�F���a���0���.��-f�۝wM�
!c���:��֮	����eR?;�n	�F�^�[S3/�*�R�`�˃GLl����U},,G�ScG���gޜ���&V�sZ9�&�棪�[\�]�x<GE0�W�RZ`Zv0��sCJ�h"O�Qի5.n�2��P	���R�������� ��v槟 �"y||I~�ڝ�y����������O�c�wp�	s��X�j���D%�wY����|����"Jd�횉>��u�!aydѴ���aǝ݇J��7Z�VbȆ'KcN�e��IT� }��?¿�U5`"es#���?ko �L'��r�q��5p:�E�W�+����\��OVOG%�C7���ܷS.OP�/~[�"|ݭ	��������P�.v&���X;�-��
1�E�m��Fb�Az��{��G:(:�H+Z.��(�{�6Se �¯gi�$n�~ �r�5}D��/�-�}� HB3{!� ��"��?�\t�n�ѥx��,%���ă���%i��Hj8s�M�2d���D ��%
"��Of�nswT�����M�S�tk�G������a����R�u�"��U�9�c��)7?H�����x�	 a$��pZhG<@|�M�L����tʎ�Y��3F�m����{�zĨ���-PgZ<��ҷ�>XE�)�D�f�7������em���5�S�e���U�GI�2�S�ܥ}�eK�Ώ�EP`�ٹ"`�e���0�����c���Pޙb�0���3ޔ�;�s�E��ha�gVN<�
c)���ů��3�r*�w���Q��x�{����]�{qss�5ױ�ڈX��?ظ41�����Y�B ���X��I�@*5 T��h t���uD��߀�5" ٓ��x(Y1`�g�r!p���N�pa��g/As�H��
}��3T�$
W�ȕ���k�]��8=j��H;�1�W$�Zo����ne��F0G$�7���`�E��Qϗ��4<c�q�Ei���Nw���a�$�TLR����#3�Rh��Z���a�%%~�v��u�j���J4йs��k�)i7�����h#0���6��5��b�Z2�tro]��Bpl��d_��à˗�Z:�B݄(�{���)$ۿ\�h@��#s�b�nC6�vIT|��P{s��ny��j�Y�@�[E�'�G퐀)�kJݽ�1�Zu蕣��q�О;v�]Q������0���7�u�~�ڌ~�۔X�z��8�Aǳz�.�M�ZP�V3"�Vl1YɅ�g�Tɍ[��S���qJ��G���A��{�I�sUu��? |�@�~g&� b[--���.�#�~�QSR�ta��>�x���T~(D�U)/a��]�	@���柭e4x����)�Ƽr"��Q����Բ�I�9�l%��C������2;B���g/�:0��w��A����ȲG�Jvi��a��-���rb�7�|�D6���FV��3�/��(�$勽�/G]�X����)�ka��}�� ��d/ycB�RK��đ�0��ޙ���uw�γ�	��b�س�^#�>[�*���y_R�P�5j|���\��hy;h�'"��|����,;�_E2��Mh�tmh���
�q�;����-V�����$����4~�&#Ė�W�k���6eM�Wa��
���6����ނ�.�4�d*a��=�Sb�;�C�pdXi�B������8E������j���!ȼ���)�O5�8�l\����|���=#����ha�杔z*,���x�)�@r��K��OR�T {�9�:Pd3�B�l�1��7����+�9�*F<H��Y�I�[H�}_ �|�hw+^1NY�j����bd�X�#5!䘈SV]���7+=}G3��`�my�V���^Z���,&s�7֑C��_�(���L_��e�|�<7X7�g�c.��ߢ89��c��DԢ}���Fl��D��wJa;�k�������aˏ7|� ��u��yY�H$�Qc�N���5����x8$�����b��F�myY.iPA@f!�u��ſ�H��Y|����I�eU�Pj�c��D�q$��tU�� Ȫ���*Ct�yl1\��Bqg	�;"�Vkl�L4�L;f�-��-g���ĚV�	�33}�*�R�)��ϋ8���/ <�v�)v����Vd�[��d0);��Q�9���R{��eFs
���/rl7�*��[(��Ӕ@U�/Y����&�~+#T.�ž���-)���{��i�9X������S%����=`d׺j��gx��z�/������v�1�9PKsV��(��L��Ļ�j�CP�� ������ݖ�5V&��Wء��9Nw9ǚĄwrhŎ�BT�����D>�{�#8<p�� �`�k<���a��[u�)����N�Kd����e��E����~ӓͿݍ�UĢ^ed���� K��t��ɠ����h��~��T�R�� ����T�F�7іư�2k&����~����j`�j�]E���@��p4(�YT��T��?ͧ�"WQ���|T�pc�"��xRC��}��9��Gx��vӛy�$l�����K�:��c�@�7�3r��W���1l�J�G8��X{/�Rr|B("�<�l7��/��$�>��u�p��XP	#F����h����3nǭ��:�~?��>hV�L��*��B���m���H��V{ƔI&��}H�E�f������["�ҥ��i���^FcQ���!�R��C^�BKk���;
�q����)�<�M���з�n<��I��I�(�&�v�f#���t��˖ʁ�1k����Hɗ��/�U����G��f����$8w~ޒ�eóA2Ͳ�4B啔� z�ک�L1\`��*��˗>=��C�dYCf3.]ʔ����BSDס9a�X�|F��n�" �`枌]T�*���|�