��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�x�W��$�oC�Lw�S
�,h�eԀ)�CQ�_���o�E�'+��l�����qz%�[LըMū��ş��Yz�g�#Vz���E���_�����/��'�w|g>ѐ�=dC6����	NwJ!�
�PΙq����F�<hŚx��#��aT��R��`v����*>wEb�3�4��	ηto��b���RQX_�?+��M���C�ӛ��/�7X�FՃ���W�"�Wa�'_ ���0��a�ߛ߈"�|J�0�g�w���r�~����"0-̦_DoU �0�,���-f��!3�!
\/��M�;�P�[ni�s� R F|�h�[��UtNi�qDۏ����F�N��Q+�9����f&D�����Ш�q�v�.x�a󖷮�]g$�3��|�jWu�m�lB8nB)
�
:�$�y]��Uhֿa�dfp ��:��b��Y�ٻo���i1߾x�B�i��F�"�<0A7l$&������y�Vk����1 F���C�l(*�]}Ԓ�*H��*PPm�>�Z;8~[���Z��{H���^��-���؅��ʫ9di�����K�vk�E�:�3^t3Q1F"�K����>@�H#����]է��檹J���7
W���Z��c��<?��_�[d{�ч��Ϩ�lB�����A�捳�pf4{T\K�:j��.~�����l)��r�^��y�u���s�:$Hh>���	��'xN9��yEySSKҐ*���L+C�4�]j���*�ŒqK�KYeU ��	���X�Y�C�v����]!'XK��q4"�cE>��q9�����2įP����?(�"�{�����,l�{�?l�7�`�@k3L'�����2u[�*R�����V�YN� g��}&U��KG5��[![�@��bH�<	�� "����ޡ)8��0>u�$�U ��F�Zd6��E<b� &S�|�� ��c���i�ڑ�A�h�'��vS��y��+,a�OG7M�ܪ��̮2��x��y:]�/���>5t(m绶Q��
NqC�M����a3�@IHb�).[T�|���L�ʻ@��rk�6��˨�S.xU��x�	��uo��Bf^�-�;��J;���@^��I� L_N���̀v,�Дm����+X��h�߶� Nm��`�6�+�9��`_�	�3��ҢV0�[69�>�(o�Ȅ	��_�o�˽���քSO�a�u��1�]�rcy�;{<���"Sp?BH�/�٬�>K|��$W؆�ۙ��1��(���r�w���Ƿ�+����S>�K�%!�������[E��d����O�|;#�T��z�>!S�;.����0���f��y�H�Ĕ�3��ąM���FWZ�V\Cw�e_R�����5���S[	=�B@��x�ː�9x7��y�!�� +/�FS4�ΚLQ�9�=@|���ݐ�V�I!�-��R�dԶ�gr��%���Xq�?"�%��	&ğg��nNw��~¸h�ޛ��p�\V�NJD���j-P����|�cP/�C��)=R�a����H�ׇ&	�ub���
�_�*<w��Rϳ��Ã�u��h�`���"���m�o�bL��53_�tL(�^>�qL���9 =E�B5c+��T*���I	����A�އ{�2ɉ����+
�1��,�;��̤�t��Y�z�%o�Ʀ�8��h��1��EO������o�Znb!�����^�o}� �ŧ���J�H�Iߠ^�SE�]ރ��'Xε����A�`���y��ʍ_�%���(peʃOZz��Q��^i���Ͱ	\�.ݣxFO��3J���V���4��/LS}+0��]G�9JH�IB����px������B(���Ox��x��R�$�=�Dmp�ђ]1���7јj����)9]�$��U�^h.m��8e���v�p�Gi��0�;9�tx,���U�(0a�C�yʀ��d�m��qj	q��������P�oȎ��9���;zJ�.3!'�#�ҽ���^� �J��Х���ס�r^���a4��N0�[�XbG��O+�@�z���a=ɾ�ߛ82
	=��*a���)L]�T�8]x�eIu��r�b��{�eV�!�c�//�lJ'���A�;%���ȖR5zq�mF�I�)p�<m�0i�,	?�0��D���G���Μ���e���K�'}�{B����vX�7
<f;�
���n,O,k�ብ�A�/nS�iK�u���/����&����uNJ����59��������X��`�Z���`g�~�@԰�!��^�p	ːd�C����u}C��X����@/N*�:t�P+���T���q��I��k��܅A���
� p?wk���妙b��_ㇾsq����@O�x��Οi-���.��߆Ld�~��m0�[>��aqt6>Ʀ�^R�ղH	��H\*�,ZiG�謽��,�%@QT�?�s|��'�2��"��9������=�����Z�ܵ��B�b~>\V�aNY��܂#4F�Ckx���RmF�=��h�@ce�k"��C���:}tT���o�xx�z�	:��:��Ԝ�J�-/^��Uc��b]�� Uuk�?G��v���5ȝ�28�U}�NFc��;�7��2� �`_Hj�3�-�L��9z}#
6���(�����5!XA49�_&a�Ki��؜V�gS_ߋ��Q{���^��8��hO�V�ԗm��jQ�-��o��#��(�ί	I�<4t�Q�ʑ�Tw	�P&�#+f>��Oz�������As$��z��qk�Q� O�b�A4�~��:IoH�"���mݔ�9$�)�O&MZ�q�&�ט�?�Bn��c9��|� ǅ�/~�ľ�1ۙ �+B�Yӥ�\)�3x�'��	���?����h�|"�T�k��L��Ȉ��j�'h��!��(��X�<v0l$L�W7�:�T$&x�����Aq>e�OG�Q��`�=�
��Qqؑcu�.�i?���!��QN��'=6x���ͿJkE
��J�{�s9h?���L7���x��jS����f��c�Q�J�������4b�*^��@��;�t�^ǃ��
�uƟm^Z�pp�6=p�w�H��<����|`�z���o_��������m���oW�${V����?|�9�Puc���@��?��Ծ�V2����8&qJ�JU�ՃtCCL��4C���̀�ﲰ�vmoK����ܸ�yF�bC�퟈�?EM�]$5�2�.���
�2���p�z��ݑ1�"���'I[,���%g>{|=l_��Uc>�V�}pa��t z���tw!N��܎w$�T9$Y�׌Q����'�`Œ�*`����8�
�!M�w6ß�k#����/��9)b���9���3<�CĎ}�Zt�aۨ�ۅ�7cY�k�6)��3N�G�7����5w��_�v���|����6�|#�7kw�!�S�"�Q��'�(݆W�i��x����I���t��7x�hs;e��2 ��3)*g󠩰}���@�/���<�#����I�K;��3�yh�%z�S�Ϟ�y��
�DdM-e��@,^�<��5��,��2���7��M� T>��-�o��.������A9'f�>���~I��xfyVI<�'�$q�W}ش�y<֎��� C	��$ݙ�y�׸}x������+�Dvf?#�ė�ˁ�t�oa�U��C9�g�7j�c���
!e����*�ZI�7���9R��å��:�7nVo����C�K,t������J6��t��m/��l�!��\0*]o���]��:��映i���D4p�+f�zvQ��v��B�@����G T|�p`���<��)�|�ϡ�L x����Y�H���6���*N�����G�ěF]�^����r, �t��L�NҤ���R����`�>*V�n�#@�|4�=�j�����;-���҂Q5�_0�Q/��A��������C�o L�2`�lD�����}��n��� ^;m�+O$���zS[�^oĹUwj(��/��
�R�n�	�*n�r}p����c��bߜ���d=���`���vǓ�TU!�)�~	m*䠮�,O92��ڗ׉��h8�����v�8�b_ǜ<�d,��ŵ�$"����OG�˴縀���[��WI�~Z/s��o��]���[!������dk��Ĝ��,��e�@�o���Ln�"6rԣ�� ���H|���h��$���/!��ʞ1���?�3�G`=���w��T)�8����NGl����UV*H�l��!�x�����"���Y���X�#5u��� 
g!`[v�r)�?�F���Ϣ�k.�e1﹙_=��J*$�'��[������dJe)�]�0Db��>�����W�`��9#���dfwnt��O�=E�_l�����U����NP�
��Z�rʺm�� 5ʰhB�%:pܖ��\���3F������u<��D5�p��n�x{�M�h[��`���k�V_>;M�.�k�����c��{���}!�>����/\*DT�[��j̍i��!dи~���ڹ���~��ԭ9�J�n���YԾ� ����͗���D���?5
k�ؖ��"�`"�Ü���K"��,�Nv\�)=3 c�e���]b=5q@J�;�C��!�/�<�u[p���{�|x�d�����&zO͜��g�,�;.��2^����{�s,��(����7*��#U���[�xlUbO��J.�R G�zl���i&��Y]q*r2�uֱ(�NhZm���ϿS6���|U�C��0=�b"n��7uk�Ѕ�Yf��o﫢=�JS���?�Zi��61��4�`]-�'��'�^E�fV�c��_F���͑ǭA'n�3�<�p0W{��֠P�ʛ,�L�����Z��S�
��-���Q�p�p�s�זp��9�h��AJ��-� g��w�¶�#�S������i��2(}o���O��i�0zʜ:���W'��ޫ�������Oy��|