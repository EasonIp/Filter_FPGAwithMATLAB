��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����)n �n�NP/x,�Fu��D,�C�)��j�vR�������|�]K�U;���A@A�qY@@բ���e�̍�gF<E�0�z� n��Yaex�1��p�+ [�B��;$ţ!
�_�c�>�Ή4�k-�e�M�}Y.tצ"[^`㻬Kg(5�f��#��D-s�q:�0eP�%����+���ݐ��j\�8��n�p������xo��|�v ��o���o�4,٫'.Kq��$�q��\�6R
4�q0����R�R� :P~�آ@�����Sx,[��0�$���E7ٷP�g����w��Ϗ?\x��%�2Ç�n�Z������eʔ�/�w(¦.o��z�2y�m��#��S�F:�..!U1��#U"�SF��A~S#��?;�
�~&�Ҝ*��N*D��bg�K�JsL�ql���dD���p�1�79F�ryσ��zp�+���W(`$� ���Mk�S�<6����%ү!LxGp�̓\�J7M��d��$ �)�.$JxK��\)�ZU�<!�R������#_�r-q�HJrEѢ�*�C:�&�D~�/���F�������^����S�C[;�Z�5����RŤ�Q�a��ߺ�b����+t��h�]�*Ԑ�;��C#��]�r����2���?]�g��Ϛh�D�;�<��l��W��4hJ>NeH.ř�!?=x,����p��dAdp��}�X�=���y �w�S����0C3U����&;5E�� �����>�ݢo��Vr�����m�4��q�=��Ҧ+$�HIgKp�PB�F}6��GXz���x��b��)~#�_�U#�=4����q�ȣ�&P@ ^\����(L��V�:�������e��`�R�Q*���=W1&�ݳ��C��b�k�,F3��2	]�]^�-��ʯ;fg��GG�7f�.��~i��������Fچ����I$�Y�@�Ӈs�d7h�)~.���0���t�h�:�����8m�Z�"��Oޏ_8��n�B"kk�|�TƢWv�S3y?��ߨ㳦D���2e|
���Z��"ĭt҄�X�����Z�W�Z^~wx]b�[�+i-ja�T/�"(���Ѕ�K<e㹌��N9���Q���G���e<�ˉbbN�ۀp@��1�s�b�����ۈg������g��eu����7=��m�S�]Ճ���P��M�;���zO�/���K5��N��#���xWls4"ZA1���#��[���._�S�ʁ�E�]���ʅ�ڬ+Br��Z���K�k�q����\��4J�B/ޡ,:T�[�E�7'�}]`B�*Qq��S��<�d��\S��(,�yMQ���tH��0J���$k��(Z�r�nS 8�/!���5��������Nu����S��+��%F�,7�y@(%�9h�R��k8ĸ,�\Ĕ��>�_�J'%�{}a��#���Sl���!(�yG�G&J����1���M����~��P�Z]�3���*R����1��M�~���@�$���,2x���$�g-7�&�Z��Li��a��x������X��R��"O*�Ō�Z._���;�8�yT�G~�kL���GZ�+&v�6�V��~�"�4,�g�&��On�������_1^84�68��:����tՆ�����z*��N�ިx�C%�H>Q7
`��Y�5%���}�D�������N9b&�.1�&�gƬ
�'Z_�L
��t�`��	PHW>]�,�qW.�;�2i�N�NT"���_�P��Vn=P�Z�s�/�V��n������Ɗ=m��>�Ke(�TA�>�"c�L��g�����ظy��B��p���7������S��$���h���Z<Y�T��9ܑ�U�Z����K�#+^&������놗�T��	� }�}Mͱ 7��O�������P� ��k�����u��o/�URi j��u3`�
Z��` ܵR��3���l'V/�
�f8Ǟ�g1E�9l��+c�r!����D���`+���4SA�!m/]MS�|z�|�2e@�{�vө�_�~f�E���k�A�,�5����ˁ��4y"D
��\�l��%��[�Ye}��F�LC]�ʻ`��Нm����c5j�#I�,f�xͰp�u�<�?M �������ٮ�F�Z|�9s�������E?�3M������JÁyz
��;_�ͳ�����L|	����+�_a�K�2�e�����tI�F7\�Vf�'E	�����JR����Er��}asH_Q,=�l<�f8 6��E!�Q�B���8���e����/�h���&�d�U9�b�r2Ĕ�.h�U�X|<E%ɝY��4p_}�Sv�O��b���<��cǓ�E�w������{;��ۨw�p3��fi� ��I����ЇX��K��}��y�<t!�i��t�^��:Xz��i�p��7E�{ �*�٬�6i��A�����lwuZ���:��qCw��w�Cc�����a,k�d�	�O����Ǜ+�O&������� Y�uU�q+�j���l+�MqE����0H���7C��U%����B(�\�$�f|�_�'cKï ����OK�����;�/t���|��( /cB��39��s`՞[A�R>/�9]��^g#�zb��Ļ<V�Siɷqm��.>q�u�ԒX�K_�"�#�.��0 ����p@
]z�"g�������#2�n�F�xgh�@����X��2[c2�pU������ov�Ou�;�����yl��2Y �;�
	����C�N�|p3yW?7�`6Ef�Z�++L'O���T�Y,��%䶿e�{0aM����$.So&�8�z-�����ƥl�����x(~n9e�e[����=�Q�Ћ�S"g,"�����3�.����E�ǫ�ǣ!@�d<%v���y��mBV��2$��f�L"��d_���yx^̡�4����%>�M���B�Hba� uB�J��g?]����5:Jݰ=�+��>Z����;��mD6�?��?'�Ү>3��<�p�p�m�h���C��$�No��\9��?&���R����3�>y<?���q�;d���% ~R�u	�s��I{�A�r�tF���W�_=�d�Nzt;�*le�?*�RG�:~���ʉL��'L�k�|b~.����p>d�<�*����+e�߸8 ���ڒaw��]1pAm��/�V����8���q�
�(��k�*�d�`�f�X�S�֟�p��aج�4W���vlJ����P��%Vk���+�W#�ʕ�.�O�kP�7��?�O��}��(���9f+=����'�B��Ox��^�����y�39�;��xR���-�����EX�L\#eM �)5`��!� 1�1�<\q/@�HRJp#�@S����i^R�f���$KJ�{�q��V���~G�QjL��l���h:`�1��#�����դ%s��瀟�~��W��&V�@@���t��0��z0�!��"ˁ��T��������)��[�:���xX"&�>�y�'[$\_��\�JV	�%�h�	���f��}i��O����i�Bg|������,�+i�G<�:+��*����N��f�"ݏs8D������p�)x]8i��xaݣ��7�1@�f�Pkfh�����ߤ���/%���;�#�ḟ|�N��#΄���2v�"K�?n����E�~q��@K�{m��P�Ճ��ф��w<$�f�6߱]i.�ƽ�����h��`���64(�	�#�!�Ϫ�Z9;Ҽ$��q��m��d���{��e��e�kbAjb��̱E�y�vF��3�H�Sc��h�ݨ<�������3@�L��+-�w��&�pN(k���i�o�/���׳_����ϝ����U�|I�o���iۗ}��A��2��m�I�H	�IK��+��aj��Ҍ�A�s��b�@Iʧ/�ަ�;!�*ӛFI~�<�CY�W��|���}	���� �Ň������N"�!�	U�1���|L�s��fN���9r�q����oI��~�׺(��̄�T(2_��&8X 4��i��v>��-Dagb�m��7�����Yj�^\iEޟ�V��b.>�}�N�R�������:�m�l?�Ja'[k�Ƀ���[B��ܱ!�&ږ�2�������cE�����s�j1n�y��e\6��UN�?� ��2�zxFHP���g�������
b�z�'d� D�x��o�3U.ZUl��o���L.+JY�R�������|T����