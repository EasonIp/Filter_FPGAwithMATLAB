��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�7ټm�lQ�חY����C9�n9%�A�iN�k7�r���D���v�O�P�V*�d�����Ρ����Lޖb�lP|�����,yvJ�O�;Ҙ�e��< _(�����637��k�g��t�+'�����m�@��5֔�^Z�mwG3��p��s�Ư�W)4���J 4;]�]:Aq�A�Oր��$���D��q�=�dm-$n%m��;��n�'K�+VȰ�~B9i��X�Z�����sCaM�,w��ն=!���br)3>t��Κ�zoR��U%���a5t<���߭Cベ��2�:����)�\Hߵ�Qϼlp�8loO,�3�fE�B��h�$5A��Ս>�������^�ӟ�����qkS�n`U��5{tz	#�呤�2d)�!>�����P���(p�NP;s�E�T����8L���w��!7l}a��a��̇V
!5�I��y�8�4<��A��U.s�����@ac�`������mdLK����xw0��/����N�j^�ˣEkLٱՂ��"<��^��M���]O/+���3�uᷕD>$%���+����)�*���R�� L`�@_�z�h�O_�TS��T���V�哾�)}B_�+�*M���~����Їi��P�uL�! Z�8&׮4���F5���gt]0�p�x���Կ�f��4�q&76T3�:aQ�F�XB[g"u%�����V��=�w�-W��o/�Nr����B" ��o#�y*�!��|!��{�U.�����A���^�A�� >G�is(h�ި`d�&	/��ej?LMчG� 6U�3ɉ�8��p#�oiT��C5(Y���͸�$�H�b;�Ҍ5~9���=����u���:��J��P������Q�D��&o1k�%�"*��/�߈#��G�)m� W�p�u�9u�83��*K�j�M�tuA��0-�sf_&_�#.�lK���6�S6�����h��*��[d~)`�\���4�F�T��K r��S��I�hh(N�1�R��0uuB�Ej%�LyC&�%��e���)m�+m��]b���ok��g��lO���I��S�b��Jڦ;��ߍlO����=��u3!����;P�f&��� Do�MF�qV����i�	r>��`�2�Cޱ�9�9�8U�R�W�	�P��彾�׾���]kQ`\�u*��%�v �P�c�do��N�@������Ktx٭���\=�M��7)�E��\���+.,:��a���F�;����v��Px(�dc
�-SƸ}�C�(���b����Ɍ�:���m�QuIjΔACx[q��`an����������5Q����X�J���.b>���kǘ�؜��x��9j�0ݼ)�u�}���6�0�]ެJ��Jg�o�w��QK���%��\L,}����;��\&@/�����~5N�a�Y��XlwNKjFfC�$�f�[Q�N��s�ZV�1D�\����4!�r뺉7�/��'N"���g��󿣆}y�Md곽��?�A�1�hC
k����L�P�ڱV�����wT2	�Y��pq��f���ȇ��U@�	�U���~�M�E�L#�W�.+ݒ�����xW<+ى� ^�5��Kޫ��g�*�'��:mN��35��Ihi����-N��RH�U�/��p;��U��Up�(�w��mJϸ�&�F�{bu��k
s�)>e=��f+v�����xʐW'v� ���-��s�O�����<����0.����	�p�'��P��B�U���nx�<}� ��Nv��K�L}q֕[s+M�"�̫2N���>1	_�����r�N���v){�f;C_�s�+����-gBt��J��x!'bhf|=�����-N��Z+/��k���>�_�/=v7!ׂ����g[�v�ֈ�#x3\�L�8�˥Ym��'���d�q��B�DO�GJ���}h_���� �y��=�E�>�X�Ҁz�K���F�$�GG���1c)����@;kA^�o����T�g�3� � ݍ��{,�ZW`J��1yg7l^�Y����N�)���͵�Z�p�AkD0���@�"e9 ��>�����z�c �r��bV��D�k���&d�\`�D��@�����0�N��	���'E��m$|�E�e�����ap��J��Hg����W3C�ޕ���羮��6$ˡ�Ӭ���n^���W�����6�G�u�.��%l�'���c4 �*��H;](v4�Dj�[��F�P#�n�j	��(�<�����4����p�;t!P(�TEL�9�'��S�@�6)�Z9q�rp�l�{G�#�,��:��	�����u��( q(��o��9�ygգ�qB=8Z2"��
|��']j� L�Ճ^1�G�)�R�C�V�qA1$5�3�:U�A\�/�H�:1~H�?��&�I�S+7�y*���A��:pQ��B|�^����n�UZ"L(���K_����f5�3�j�jx�: Ed>�ʲ�[A#���������$5�n:a0�����=�������W�E�:�%*�SY9b=�(�{`�d����-���'ǔ*���Œ�1#�mI}��v��P9�ͫu���o9*��	���	&TS���:b��%�]���;ŷ�D��YW*C�1�ʡ�iQ=X����7��QV<����˳YOw]__�D�����576��&��}��e�O�K�ٸ�	���;��4����N�� Y�3�:bf��Ҵ��R\4X��T����K�sbv�35�1*b�mk�NgvX�Lp#?�7�l0��F�{�}�9D8����9��YgSy]f��fZ����b��w5I��L#Gg