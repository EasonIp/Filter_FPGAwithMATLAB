��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
����Tӂ���^�2����+t2v�g�VU�r�H$�\%8/�!8�1���1,c���'���c l	�� ʁ����h���z%����\�?�;�=�6����w͸>/Q'\p�~����|��k﯃�`d�C\br��a��D�z)*�&fV��X�v��H�F���i$�MJDK6�#r�n��'�>ro��K��[x�?���IÚw!	�K�D=2<�x,�kx��s,ŷ�v�QplC����R_)�|�m$�L	�cߡPX���:�zI���H 
"k�6C���O�^8r��	�RؠN-��~��-���5>�*�hbD�c�D�Ma"���BRҪX�F���P�wy�"��=�댣�����
��KY��Nn��o�o��\�������-��'�'�?9v�i|b-��g��R��i��x>����	���Z��,��G�э�i�ʫw�mDT1E#(/#<S���c#E�E$}A;F%�K<��`�Ɖ�o��<����9 Q�ӗ�vg���$��zk����顛�Jt���>���.����U�!B��'o�{�18�>���ƽ�:Ӛ��������!��(�!��`X�2�3?�s��;!��f�	�ɉ�jԷ������o>2�c�z��v��
·�{��S�_XSw�h��e��o�o��߂�K�Hi���mb���ܣ��M8$ő�V��B����[_v��@u�ԔV���.J!���H5fG(F4��d��ثeS
.���T�����V3��[{�7a
�[[�wy��e��^^`�2��� ���j�9�Ǥ��O�,W�x`���f]�o��2��dPk��ESq�O����Y�mM�Z�r�<oȯO�$`q�z<��VN�, ��C�|�����jt�ė&�0H��6n��������_S��������8,h�%3��l/�f��P=�q�_����X����`�4�(��D�4�}/��POXR�����Ɣ�p!�Ù�́RD�J5W	�D��'YW�L�˪��z�C�(.�X�5Wa�f�+�T^��A�P�.����� �O��M_�=����C��C����Y'�p�� :�;b�k���bo���x1ƽ�7/ /��֢���HӜDÉpw�	K�e�& J��ӷ�Of���.�� hk$|��W
+�L��$Ff,�MxH7�ԇ�3ٺtrӺ|����\r*+�\@�g��������W[�ʳ$Y.Q�[����h�)�ҥ��(?9�?縒�M��l�\ҺO� C|�|�oC%��3__c�e��X6�2��)�DW1��U�<�q
����U��
O|��p��f�c\�����������w����c��6����'�5G�޵�������/k\_�FzȜ�N/:FTc������a���Ӊa+b���3�Qs,C��Þg�O,)$���h Dpin�XEpT�%�ָ�$Ϭ�QaFZ i���,&�<b�e�v���C�t�^>{��%ar-o� A��T	��Hx�Yv��s�0�ʺ2մ{*(T��z��#Z5�E� ��c�6T}�N��h������)�桂�t`��/kl���>X"� ��e�k3�6D���$/�����idR�#�OIZŁX�JmN-��q�ۄ�a�SL[طh�r�� �2��*��@vͰ�I����`����ɫRN��#'_����4N@jŏ����v%J�=Ed6Hə��z�����K�lP.����r�y�ߺ7f�7��D�H��yB7=�Fx5X�
��E��P����F�;�\���S1��w$�v+4����T���s
M�9�ƌr��������/�aCd�N�r'��e�1��E��vy�lN�粃Ķl���Ƅ5)������FU:s��Nњl�g2m��8M�uյ�8�Z3x�oɳ�(�?���`��T]���`D����U>���$�'ě~���ɞ�ݳd�_�kJ_mM	�oV]1G�5�����F�sK�Ҟ^����	}�cͲ$F�����NG=�TJϣO�����g�&H?�c)rdODO)��C'e)>r����	cQ��$���B�����8 DXYOI弜^A�����܈��Wմ{j2s}�sv�Sh��j��]�L}�q ��갇�m{��t�=C�XFNӛF8/���B����CTXjg���a{��~t�]F�<G��3���d7���T�i���Gc��`�;;�
;������UP�.u���[=�ϸo��57)I.�r�z���	��>$��S�~q�QtY�U�'��i]^��Č ^Z�����%H��V��<�����D�A4��utTK���U.gg7�vh+{Hf4���f	�=Ä�$��~':�D�.���7�bg��e�_���;iD����N�	Y	;1K��G�B��)D�]�}v~��Ė'A�l�M��A�c8����7�h����E�tfn!X�_>�"CK���6�nJO�_|�=���,�M~���c��ύ�t:1�Q���oRN߲=�� ����j��!"�=s�-�B�.�������'
�~jw��0�Ⱥ�26:e��S���& ��l��(໙Zz��|R��Vw�����e���\"�)G�Ζ�	qp��
3�ĒkD�2�Ȥ������\o���t�M�04��S&�)P�P)�n��U��Z�o��~�׌J��I��'�� orc���P�#�OI�_Q�Iw�v�O҄�,5ψ-��ԼR~sY�������t��a\��o7� �q�냌�D�B��y]�^�0܉#+���L%��A�Ce��~?�ĕ��Hn�N�I��h�����|(m�^�O�v4�"[�e��.�,��>�!t	��!f���9��X�O�����u����,K��[�����x�y�������}���.������{����j�JUմqmx��ɵLB!�۷v�8M�����Z	��MF��m�~y����)8�obE�������/��ty�O�On��[��U_�Bp�S��f�����h!��n*;�����t4�s���˼bo��d4�*g7��pG̛�a��܊�A��#Ѱb8$��YBR4��3�S~C5,0]�OK	��v��j��%k�������yy�� |���?Mv����M.��}�Νh���9��V�.-X����X{	��߈����d��_��I�H�ن(��
2�L�s<��`��l��0r�&��ש��t`��}�P�P��M�h�e��D��1B�g�Q�
�����&�m�r�a%d���E�*p��*��՚��B����=RÓT�K8{L#k~Q�̫�t%1��,�(��_�2�|o6�/����ڟ�#��� gιr��C�o�g���#!(�K����?��$Ud�ZGՇ��:�݄���
x88����C+�����4\�|� T�����@����M�Ȱ7`}|֗��� H�����ϫͩ��#W �ZO�J2$=�~1�7��,�_���
��l\�~w,�U�;?��Z�9�����mu�z���~gڲt�Kȧr�������^5|�a��c��>7ZṦEp�\w�=&� �ڽ�e�1��T��Yi�S�&N~17AB�՛��/�8��o�����v���C�*`�r�3��E��{o� <R��,�sT��m��F�l�q�.�  ��wn�U`��n>�㝕K�8��E��Up&
Eio??P����R�9t�%#+�b�sT�>�������H�� OpٓOF
 �;��&�R��9�n����<��W`戋ܫd?x�.�RN�,iو�6�����	�B�#�e���F�����)�ر��<�l���3/M��3D���5����o57��%��L2/ 1;h4��a[w~Q˽�.{u�0WM�2n��7��8��<�)�"���D��
Ä��k������2H��I}��=Z�g�����wk�,�_]�)!�ڹ��/�pl =�q������\btZ{�<����T�ȼ[�zߙw��wq�g��λd�^����^�2�f����D7��n�i�m&/_`�Me9-�i۬�� Cw!	��3��9��Dʶ��������H_�\���
�w���G�������ҜQDDӏ.V�3R�)�{�])��r�:ɭ_������]��u~�����J��N "�?��+q�	5~�丏a�ET�xms >,�T$��7H��F��l���VD��e���H�����x�>k`�Yƶe�W(�g<�$�q�뵇�<	�a1�	��B呀�E�H]1:��WZ~�ٷ�
�����}��<�eȳ���gܱ|#�Ќ:��'���2���0�WǸ�l�e�}���WP� ��UkQ��w��e�	�\�U��R)P��Tv�Y-#�9�-Wk>���ٵNU�@
�ҳ�� �X]#��1$]�����;M�1�P�lĊv�����=c i$º�'�XGދ9 ����Ml�%{f�7`������}�rW�A<��olD�BD@�=�� ~=vIm9�.H��s��Z�D�����)"pٴ�rzj��K�][�b!��m2�('G�+h��D�������Ø���̥�a�B�c�����M�O3l��x/��۔IR���p:���<Hx�
�e}�E�.��a�YF����SߨhY@pV̉����3�!��Uj�����Gݰ��!��DW=���S�'N��+�2�k�-#�ͧ�[}��X�o�F�p� ��T��b&'�r.�~0�'���7���.	W�J!RؘD�>&�� ڛ����C�p��L8��)��6S��VL#��е��[����iHn� ��x�tb�v�*�������Y�˳���"��_^{�Fs�1�y�>ƋKTXb�S��%����]��E)�VT����ſ�OT��C�Y w��}[����=�5O��i�!�%;��5k7�sh����+�?&�Xm�'�J��W��FT:ˎi��睃�U�r�̨����WXS(�^X�Y_�3Np21|���KALۡf�e�P$����SS*n���iS�_�c�h\�k�X�ǧ�c|��}hsU@������&�*d����A$z2�7�d��j��`8�C>w�N[��\�t)3�}D(�"�!�Q�%OQ<6u��,�n1��8_o�5J{<�J.�U�V	���u��^����9���Ep�����ό߽��1�WI��	��NN���4�kx�l�L���q4'�Ҭƙ?Z궳pM�?$�{�:ҫJ^���l��`|��^.q$�el��K90��[i��vM����t(Q#��a�_�T�(�x�j�0��<���6U����1��jG��L~O?Q��BFz��V��;�Z������S\!��C��
��6*�@,�GқB���,n확s�+��{p��67�|�����"���m�\6҆5��U��a��������`� ^:�ҭ��Ld=s�N7�*;[5�a��)	��[�e�z���_Z@�m�1h�H�ڥ�Z%����u;��0�T��r��~SDK��_�	,Og	{�_,�xs�S�� �M;A{��ŉ.m�8}����~1���]ƾ��Y/AP�Qu���P@���
KfmU/s�G�A��4|$�_��t��R{'�Aa��ɬ�/��[m"�����o�l�^J�bŸ��rQVҰBH�+0���|�������o�\��X1�]����V�2�J�INm�=��!�8�	)�4xȰ��3G>9���2e�R�L��Im�o��qF�s����Jf��"���G�U�i�;繍����P�g��k�А�嵊s�'�����Yf����,q��4@��������f@����e��{B;�p�*T�GM�V���J&�iqDfYw�5���&{�e����Q+�fl��NE�c?�z���3�RL��8�Dx��OT�m�}b����^k5�Sǲ�+�i?���t�?97�N���R{�����ܱ��D9C��f�����ۤ���uፆa<���A��n$ܒ_�&�ũi�0��!,<���	|'L{��߬$ �yŽh��~��O����.P#�vb�U5�GfH39�k׈7�+nj=���*Jn�4ш�!��+��e���m")�i��DiO6��E��IC�'W���˚b�@�Q����ۄ����2c`�
�逷�i6wV��
't�~�p-F���.��$�Y�_����s�az����a���l��)���ᐷ������UT|e�r�Ѣ^����JMu�#AMތ���{hrn�n*���K7N���/[��c8{~�K\F9/�c>4�K���6	S�)�1L�G�!O�ZDV��\$��2�7�{|#�-z���	�<؂]'D�o�x8��_��m�"&�#�rb-���d�$J��!7���*��x��ߟ({E��P9�Pr'b��i1�ڥ�)����Dw��R�v8�%��R��`��*h!W���_���3�:�����!��;������[��w`=�k1��WD�\a�Ј
�&�u��?�(�5f����e��IKSOC�=&�UN5����]�<�aUZ����Wv�cm-�{I��]uWl���u��������Ⱦ�C��?N�*9������4��s&��ǖ��s�<B$Wͥ��۲� 6C�S�lqy5�H䱶�ᴿw�Eo�siӒ�@��,MyP��;j���K0�	1�≄���$S��Z��D��۠;�����0р�Y �q0�1��(��i����U��C�׽֐���S���e�{���#Rv�"u��z?w%l�^��`���i���։w99L$�^\���W�8m6p�}��F
��/�SZr.Q
,ԛ@��2�%׌~xL'����~
Ϩш�V��;����/�0���ӊ��ݙ�l�!Ѿ���f�vڒPH�
K,��)�H#�0�4_ xa��7��M��E.���w95vh��]�-4�S�Pa�4Q��i�=O��Ҏ�v�9Idƚ.P�ns���7	=W)
�8��_��4'x�Jjm�<|�־œ���#r+\Z2�D�5��Թ�#��iǎ��=�]#���:�/D)]���ٲ�p㞘X=���C���.U��&m<��M�љAPf����>�2��29��@PA�f��9#�B��1�<0Μ����P�F� ,��"�KE�M��.������ĳP�܏�L������>� ���[�S��;2���V��t�X�7Ս�)B%y�h����3X�
8� 5����'�`�>�i��8D>q8��q8S��*!ʦ�7�7���_������lQ�E.�E�y�M)�8�Q�M6��wG�iT�WiB��)5�sp���m�z�i�����	�6J��v��kW�
C���������o���؎,o��q����n�������1'��s�z�i:r�s���d=�'qk]�%�*�pa�ڗvT�� �> ����h'�S�Z�n1�E8�(�\	�er5e�Dڦ��CsF�\���4�D8��89)�_�|��J�j�'޶*C�jk�TD��EF�,R;�UYi�/Of5� &b��G�G�3~<ד;�[Dܓ�oݛ8A.|&^w�V�Ml�}�������{��W��\_f]����3�7�T��0�������8B6n� �(��"u ڍ���z� ,4	��������6��n���������U	�?��ֹJ��vFd�VX/�I�
�uDƹ;���b�tG���4w��q�ZΞu�ҏ��DW.ħ��e�҃d�%��!͔*� 6:,�?��+.��܊�̔��=�>�Eq�2�f[c&�ڹDR����P�G����0�Y��7M���|{#��<8kf�b�*�?E�Um�GxXyRL+�[}Ձ�{��[!D0gZ4"cb�9v�Q�{r�
�׋Z�����_�0Bp��͛��uq��5�-�C�D�轮�X�P�Bm��0��q+@��r'|А�����Jm0)y���|P��L]3��do�Fh6���j����@Oc�V/�w�9���I{u.��izV��0O�0'��TO���9� �-�7^+�b^�&x�C������\�.�ۦtS�ֆ�����^�ғC^�=䠱Y@�w�F�vg$���ٚ��ۥ��.�d��4T&���m��Qg��+���F$�"Ē��Z�;�Gi�G|˹ݟҞP��+�]�h�U~����'��[:���4�H5y�^M7���� �u�/]=���E�4�5�۫`�B��6VGEx*��u�'3������I4����`x
NkHմ\��X!�(\�)SFңZ$�n	�r�[��%k����.�;bs,���Q&!�ft��`��9����E��A�I�k�a�M�MQA��w1��"��q�K��Y���]G*�ڟ�3��%�q��Ĉ�p��"]!�(�HQ���[Q���`��N_����g�b_���	kS�f H���߃��3�!�I63z~@��<��AMݠF��.�bk�F���1�ѷ�B1��w&����I!dn����0b�K�A�T,��1v��Z&g��Ҟe�Z������E/��p,�H��Q+p�R#��z3('����cT�o]`t���*�\��.]��͒��A�P�.�����ݨP)��g�h�Wv� C]�V@`|ؑ���a养G$�v��)���^��s����-�����z�𫯓��3[/�� �*�RBj�¹mo��������$�T��aXO	�`��k���ւ�W�Щ�G��q3�km�{�:'��|}!��}%˚�o���y�������|B1F�Yis�Y��	���rq�ۦjh�=�o�l����Dy�B���?į+�Z��������	�H-8VG��SG=-jv������Tq���Id��]�����NSRC7K�/�a��>�˜'�HR��_A�����m��Ĩۯ�l��ز��,O����e�3�F�/�����n[�����`�+^�&� :y7�-FL^L�o�@/S��)�	!k��*8Z��2��}a\��te�{�nt�[�7Μ7���dK�%0�\``jWyR=xݝ%��3�9����Uf.����F-R��Z�"��@"/4���`h��߸޼u��(���i��E������5?�,��-3�(�q��׼Zy�J+�Z�Y;�?�C�K=�TNQ�}�)���>�$�me� �(��1q�1��˼����	ǈ(q)��D�����h0������[���;����܉vl���w�[ϒ��m��q��m��DY`:��&���į@���9�v�P��9�6m&�n}�j��������K?������?�.[7�(��ΏΛ=ެ>ex�FŬ��p�ޞ#י��yj�.Z�]��[EY� ��~��;�˜�J�Eyq��] n�G�"�M�%�)l*�Q+*?�86�t ��1y)Nc��R��1_z���Œ~��Ç�ǩa?�vn���`r{��p��k�,����g�n
�z1�4���eVk#��Q�`�u|#9��F��8C��3o���"?ղ'���i�Q����O��L|��0܏ �H���ߌ�Z/S�i�$�B�;�3������ɶ�M����������z/�'0(nx8�S�/��t	��*x��];�R�D��<U1f���$�n%�A|M�Λ�Sɞ!"��||�i��ӏD,�0akCk�v��߼�ʴD>��n'�hO���<Ɇo�ټ��!:l��ɰd�[��3��-|�GW����\���ø'��;A���!��];`2��T:'p�i�] kX;�.C��X����<���f�n���m����<X" �[g3s��j*�>�Cn�G&������-���<=PP�?|}�?d9��{�������;�ͺ{o�A.�-�p�Do�G��v"�<��a�s�������X�)"�R7�'_Ib;(�V�_�C��k!���A .�L��^�g[	2VP]I�{⺍>�KZh~������M��{nx��מ9�:
R�E�Q�|G������+���M�T�)���7(�B�W3Đi$E5R�/���5ސȄn�=��3�B���@��@-�7��u�`D���1���GI�-���բ��1!��5IkU��lۣ��ML^�� `�s�tJ��7D���j��V�<�8�ٷW�(�(=b�LG"5˝co�W;�Zs�<�����:�CZ�Ih���y��fw�FU��h��u�54 �hcSAL��8��b��t��V����8�P*��K�@t|��5�D�"a!wT=��e��*S��tw
"ev��l�p��r��:�� �E��ý/R琉6���"#�pLS"Rn�v�'닓�	.�r���Y��N	I)� ���;i/��O�v��N�#��֪܃�q@�7��`5ͥ{�y��<��x}#��h��*��o�`��:tMn4�H�he��諭BOߏw�
��&�ˢn���bk���k�v�y i��?=3/Q(Լߛ��Z�ihi��������;�j"�ۺ)B�fD#�ƋQN��l���}� r������4�@ ���x�>�j�T�(]t��R�����L�����;s1#3!�<n"�xU_�lPL���o.�����S����d��[
Â�vO $)F���&������C�HV�:~���GSLREdsr��xo�����*/��(`��ӣ�6%%0��R�)��s��+�y���
쎧fB&._
�J@(�z�n����?��@g����3V�$�7�$�VU��[&�����@\��k�T��1x��ǢԘؤ� 9����6b��6���m���;_�Y�m�?5� ���{?_��9h���<�uS�tN��,�+_j_�`��>��-���5���{і���q�semk�/CzZ:���{��fIb�G�W�i�m8|���9�������(��tGb���c��e"���Я�0y7��	��l��m6k��n���9�)8o��豖Mj�����u��K����Pa:DwW������tf�04aw}��ѿ��oP,>(~�y>kn	�z����X�NƩ���I�72	��M/��`�y"2�����3&��ޮ�+ˇE2ow=,X�1��� 	�/+�l�
* o���5t?�s��k����d�����2�� �پO�HUeK)�Y�d\�&O������yd?�|a�>9I��Z(��	��^�*�:	RK��Ѝ�|��� R2C\�şf	���y�r��+���Ĉ�{�Ћ�U��{���Z�~U�K���P <R@��&*�<�^��t���jp�����ʞ�qU��j+�`�=u�a�ˉz[W���]�R��7td1:���Y��2,F+r���"�8]�]����>��A�Рb�
��0��%�:2x* ��֋ _�GC�����e���`��؄y��Ԍ��T�<\����eԲ�����I67�m=��<�b7�hp��r􂺀���9!�"m>4��o(_��V5�Q<$Y�+��pIM�X4<,LFHK���n�F�H�����6�:�@k�]k#O���/���B��Rۥfi�lR�u?�u~~Lg���g��od�;��4YW��|Z�D��e��,B�����
�L�x~L+��%�4�6��'�fs���x��
C�fY*'�qED��+�> �e��3��˲K
-�+f���)���B���-qS�#����Ei%P���z�s�]O,#�i�T^X@���'M�c��b��ޖdL�E�%Z�ޠN�i�i���='Z6`_�/�j�������.dk�|���o�E�ډܫ�Z� �`H������k�D�,�XY<����A�nl椃e����q$����k�̓E�(��b�ڐ��qH�Մy/��k-9#l�����j�`D�fI�Q_sҕx8�e=��4:��do�}��������/��j�ı.
�|�r�l?ib��ô�z�#�&�W-���X�F����_(����wܕ-��}�ŮH�* �z���]�r��UŇ>G��� l��|iۯ?��5�_)~���|��ٛ6k�=sʖ��j�{I�6�(6Y�T<0š�����2�j�w��	T�M7�c!lf��ڋrsX��6�X��Ϲ������g�+�<���'uS�U��pT�*���e��aB{���,x�!3@�$�93��~�!X��%-��&2n�o�&�u���$�F��De@�uN��%I�N24{�;�Ҩ�C:�W�[�|{t�ڝ�̱��O�l(_2(�1�ur�����?BF�ԅ�7޲�4C��p�|�>A<0AK�>X^�u��n�lQvg��`mt��#4��}�t�͋������E�
8�\	������Ϗ������*�P���.p��� ���^�����z����B��Zfw����d��zc�,$��}�s���\l7���U�w��1S؁o�_e�� %Ǥ&��2�~�E�GB��	n�C��u�<��B@�	?&��9v� ���9l����z��M�Vp��piIo��:#��P�XO���>�p�s���
�f��osI:�$�!ᾠE��_���������=���&l�2N�f�X����5�W�Y��7��|Y40�4V��&r\4J��a%�>K���r�-DG�n53uU�-�z���V�ܪѱf�c���A�z��uH�=N2�a*,#W-�//��skG{/�7=(ѽ���X����DĜt���s[z�Tw.Hh��fWqX�R񧼠8�F�b�L�&���_Q�f@W���8�ui?�q��Z޴�x����Wx0z��0��_�P#��H��Z������'�,&4�n���H8�ۡ�������^ގ�x����8�A���c$���ؗ$�5�h�E���{�M�V��`��|	�5J<��خ���^7n��8����<�z����C�2�� "�\}{�v�5����a{�ۀL���h�#P�§��(/�'�)�A�+�wl�M�Wm�
�\,kr��������ZD�����`ŉ����v�D�w�JГ���ʶkG����*c�����+:���Uf.m;���]@�4��˝ʉv�ډ��x��"w���ߺ��S���5�H�Lף���35G��E�E�y>Qkx��Po��O�~x�� ۺ'�B^�����TT#��iE2�1R� �w KNF�<�J��o��Z��p�U���j�]�iFZ|ԃ+��{s�FV�5fr�n�-����`:���d	�%eQ�.]XN�$�Sp�"Z�,W�� C�b�b���z$8/"0{�Ff�P[1�"�YC����1��	]��=�8U/�Uޖ.��^�v�mm �wl�p��H�i��"�z��d&�jr��ӫ���� �������mw���a�	�L9���>������@2��i�$��C4O���-tk�N:��ԅ�`�`�F��;�7�򈥌UJ��c���ǒS�������ρ� �?$��$Q)�|@�Jf�� Cw�..�������o6�`����:De��Q�w*0���m?��x��g3�X���; Z}�$w�i�Y�W�=�����]�f���j�Y��L6�����Sc��k��d���
�`B�H���V�;��|Ʈ��h#�Nם��]��!$��g���T�c"��9� D�ꧺ����XW�Bj����8�x(�0"/�}226�B�B+���a�Ql<y�2��k��J3�.낇��_�au�r^ros�Zí�9�=��&1<d�I+ �v��ہ�6���fM�7^��J�� ]陀�z�	�C�?�W�mK��0�^!e�‥����8�H�E�$(�;��+`{�g�e6�cN?�3�e���-�s�@��v2������i��j??̔���)/A/σ��W�Wq���7�h��`l�q}���#��*�wA3.��-бd��W�+"�<fm�G6i�����\Rʠ����o�����a�`!7�ikG�#��� x�4��Pn��ǚ�#�5G�.���3<I�$e�|�o����7(A��ؑW�Dr-a�<��K�����}`cQ�˺lA�4r��R���(�r%1Y��"Nc��LИ)�,GM5k�5���ǿ|�lLQ�	#^�����^ �J&��^���D�2����)c�_����{���I;�~=ځG�j��ܫ�Z�A��2�wS����4�����u���;��D�#��w7�	J6V�?c$��X��c��^6	4��R�',��sW�a:�-��f�����e��Qm�����t${3�Xsj�撕ZZR�S<�$����x���Ua�􏼝e�1����XA�,��"gd><�p�vP^�'%?5!w����1�JQ�B5���!�l�����y����;��5M�`��N<�p+���4�B��/Ć3W�h�A=�v��<k��BX��6#�,�|�����RV@�}�`�/t�[]�3d�(Ru�%�lN�n���<���5�^
AI��l��	��;wْ |1���nn��Ȣ���NG߆x�f�?���U�	���L�1oE`L�'L���RZ�	
��2�Z_�K)<'���?�$�����&�%��%]���V�8��h�YKv.x���)���� @��A��J`��xu׀��qwyFç^�c�iY���7M�^�!���+�*�g�<��j/��RG�NM�V$MMl-'
]�\Q�5�%{9D��,B\u�b⦭�%HC�S�Ow��5;d��q�1E��c��D��ϯN�p�Ь�'��8�L:r��1�&Q�	�RE��	Y#�d77�fb�8���[j�.y�=tB_of�s|ב0L�~��o��\o��*��p%䦟<}t��~{�F"�Ż� k-�ҳ�ҟ]ן�n8����q�7K��ad���/�����=�\y��̀!6��$,�H�ea���HC�ȩ�=�MH��(�-�U�!��"�=���R�O�'��������������ι��Ls@�&R�Q�N�Z�V9X~܎�s����b5թ<�����T{Ż��"�]�J�M�����p�,���0G�������2�,t������S��Z-�P�y5����*�^~W��]����Q��(Ϝ䮤1?ʳ�+�N�$��ݡ�؄ȡ�Ix7�3Թ��G(PS���׫]P��HO�K�i����¼[���>��^,��b��0\��ow�νU��}{�jhvޔ['fq�@/�-Oj��q��+��ﻆ����"`�ѕ)���뛗�a����5P3��.\����_(En�,�<e_A�tpN�����oi����A:��d��<�{�+�5;��?JBdn�z��'�`��1��+�!�%�2��E�qL������9�wO�OvV�s^5-euE�<ĀG8������K�'��N����
��_��>�Ìne19�l��;;�}�����L����^]����62S ���H�*'d�}��Y�
R|�PU#���i�Z�k�T��%��.�}����ƌ�v��w5�@Sޣ"ғ!}k���q\��`/��yQt"�9����F�Px�(��jc�VWUy[�����I�+���;X{;�ܬ+�o|h7��,&v�K��A��66�]PT`���k��o��Dh�b:�^D6,�lC�5\cޒ��zA�������z��즉TC�Y�-��E�D���U��a� sa�ә�b�X �)��]�����y��x�����>F���c/frd�5#���^6B��@e�6��q�k�M�V�	�rA4Q@n�,>�)�_��<T{�⭁OYhQI�'���L��W ���7�t}_Muv�v6= I\�����/_� ^ɇ�Q����e��9}�אޔ+��_	0�Tc�SI,7I�:����L<�z��i�,���z�O\%��h�<!)�aQcbBZ��^��!�� �Dn�h�n�n�:i7K����W����>�O�ݥ��f��fD"�͝�m�b�y+7�ƌ�>\���^n�2%$��ۼ��a������c�sߢ�����t�t��8 �Z �O�����q���IsJ�*g�l	��`y����u��l�ʅ�dȂy���Sfx����^�8��[���������C�l��z��)�6�]/c��ָ��l����S��^�4��d�^2�����\�x���p�IOÄ����U=A�Sվ���&ə�7�y��k�m���N<�J�e~�U�� �J�N��F�il��I"�?��!�dgPѳ���N�(��	^�~�^�2S��횎�`%�D��.F1W���;��Cߴ/躋I7�a�Q��z�/ݧ_�-r�C+>��W��G���$���p�i�
���S�p��\f�ܣOUc�U���Kh��!謩�~$��~
Hd�@s0k�I`
��?��W������N<p&�k����]�N2G�����G�N���� ѸH�W��5� 6�8hMMi�̠gls�Y]�^īa-:?+�O=@ܛ����[۩l;.�s����beUԙI��Ҳ �b9V���D��lޥ��"%k�e2n���9�^�m('=y��\���^Ꮋ!yyYР�|��ø�֊�5I-���:+��䧸.z�x=�=�ы#���m-�����+����)�+����BG�R�~�φ#:4�3o�O��/��W�s�Z��ɔe� �C�Li�{4�;��A�m�b�����ar�^]�{�
:Y/I�����~�M)*?&��'=v�T��bG����%�K�D+G�����̅Je�YR��!MȜY���x���`M@��64>�5(�л�R:�������_~q���8��:��B����U�Y��ws��w���\�G����˷�O���G�#�@�8A�40x�ř/(��"����%�}$��4�}e�%\�}d.y�yML
��$$�*�v0px��������)E`)�z�"Ff��!�C��&jy���K�sAޑ�S\� ��b|{��R
���%�M�����87�� *�o�T��O��R�+񸛯w����p8���ؠR"�P/��_���+ſ<�@�b��S=w`��NL߁�{��Hk���"k����!����˼&���xVw��3��$>��8Ċ �N&(��ޟ���Pt����g�Oݗ��5V ��0d�#��he
M��?�y��'���[۝�B���w�ɫ�xgi�Ua ��n�vO��D��E��Elڝ8�R�o���T�v��`���u��#�=��U��j3\Ic����X�}>ưI��?S6>mw��y��>��[��H�4�@�/��O(>|-��Fn��#)t��Ӹ.}r�,e���c�����+d����#Ԅ�J��Uv"�l�{-؈=�%��F3��*+�����g+�:�/n8n����	��N�:,�B��*5��gP���u�fbV��t�q�,����or�.`%��?Ga���.%\Do��a<�,~�֋ZX�7��T��cP�H�ܳ�VX�����ſ������-k��Y���C�J��?W�{���˖�˽�IDNgK����䋖L�h�ۑ>�^��h��D��Vp^AD�ax�s����sٻ���Aǂ1cB�.z�p��#du͕��*0��GEI�r|^��bB
 �X[��l���c�'�0��0-ՠ����Y*ļg����ל�gY���P|�>����!�����)YZ��Nz��/*�M�&��1sQ�X�,��%��e�nQ�_��
���%��@�\�u��f�B���.q�br,�dS�G���-��a��+��ah`)QQ��ǾT��=F��r�	�פ�W6���G�'#��'�A���.@�����G�Z�j�E�c���:�=r��:J������lEI8C~����j�'* �������/���c|;�W�Il�|GW�w�F�G0�Xq�Z���
�l��l��3;0�F�e�+�?�������!D{�-6 9�E!�ez�r����r	O|׈�q[�Oᄫ�"���p1#��Ia�iàG��s7�[���=!Xr�b��qz�s�����oD
'�8L���#��o�7ޑ+�r�a���V��"�S�6�_���cjx��*B;
��r"ml�!I�i=��젨'm�0��#�WI��Yێ�=9r�3�Yz�ʰ�!t�>؏�\�X�/=r����@#U�p�F�P� 0�:�ޑ�%�m*o"����#��G��e=N[]ሴ���'J������ ȏKf䖎R:���	�:k�g����W��4�(�]�Z�e{[��6"���~3r&�Ǆ�����ԟ�������Kv���^ȯo��UFv�E��4[b[�g<�P1����TI��Jl+�>ł���#X>��1��Z��˱�2����� �RC?j�Ik�]����Q�/%<��,�d�g�Dprjh�M_�@��%����n��@��-dK�f�3I�����E��O�n��=֠���G�K�|��������<��l��ˬ^k�Ў%ԃ��/��>��Z=�����~����K(9w]�8�6ѱ����M�RS�Mj�>W�ʪd2w7	���X�Fj���(#�g�4�7_��y��X�n��m�G\F1']N�LWܽ����c����Y)DL 7�0s=I��\k7�]I�0�Hl�����Z�˂�B0ɟ
tY��Ų�^����W�8	X���{�j�)���b��`S+�Y��8����N�Wj�����I��%>���>������\��;�|�T�f��Z�1�������6�~XG�Ƿ�|Wk��X^��4|2���ه6��	�����ӡj`Q����0�������Hۄ�rS��?�
�5ye�/��i!�k�Dͻ��^��ܙy���"N������u��	|*���LHC�yi��d��t��q�l�[�Ou�rK�n�c�\SW���y_>I�Z�2Z[6$�?��%ގ0єR� a���Ѳ���m�ngɑ�*�-���ҧ�!��T�S� ��g�s��+��kCRV�wn=/��d�qf����n�����8�����4��H�����!g
M�b���۵���0h��"@�{an�D�TC��<�����_�f]ɸ��y�ss��f��	���6W��o�|N�f���#\Bk�M����{>�и��u)F�@m����������߆��@Pq�4�~/z�	���6���;.'���#�y�&��m��<�ia${�;���76X������DQ����\+�$�m�A������^��K ���H�Y�epﯚ<?HYv/�&ݸ&?ے��dfUK�/�7ب�����ECn!]y�
Z���P�ȑ�u�^'U��e���N3UT��*�*��;nܑ)�?����TB�Q.ɗ�b��ںAX�ٷ��g9	�����*ݜ����xi���mBd��Z���������D�g��eG��>�2�)V��?4q����WB�G����ܜ�_��	��镨�ٱ_d(h�6
|,�0a�3&;�֒%/��PP z��lM���\=2�r	%~�z��ʳILaM�b �L���u=]S���<�H��TPE�W𑻡z!\���̖��X/[Ѓ��	Aڱ��%F���"�n�f����
$���+n�I�@ �D%ٻo�?6&t��R/Xl�8��ҁ�]�Z���'K}��P���+D���3Ƕ�tL�W>�����E�K��}�}�8f������5�_ YUI�L�wW���n�ffzJJ�t��j�O��6�oR�H��b�cF�S�<��E�S ���wx%������A�����?]�Z��0}��̰ J���ە٨�0�K�t��mK<���,A��Jr���]�� ,�-��˼��k�������=�1&-�xC�_#��B<0;;���7�
Q:��>��_�k8pt���ՔdK��q�~�HOVw�;㍜���X���[������n��Xz��)����P@۝#L���V-�8b+�p}j(bNH�x�]�������ߩL4(����-U�w�"C�L������ؒg�$ĎV�΍y�u>�8+X��b���Q1� ��|�A�)6���d~��D�mm