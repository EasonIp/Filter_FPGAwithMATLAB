��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+@e9wR�܄]�-N���w�Tf	��%�9��#�Ac#�3��@���q��#��e3(s4e���^oV� ��bF$)���LĻ�R���a��V��:�V�)������7�K� |��'�y�ѹ�i�^�����U3����ћ��A��}\gw�tq�:�]����I1�I�=�F��1��g���#�1�$R�gx"V�@v&��d.wC/��A �Q!Ǆ��F�W����]>�q�R#>!~{��6E�d�B���z�3�ƚ�'�+r-�"zS���[��7��;@B����4<=ӟ�����<��Q�<(���;�I>�n@����նC�����R>�r�u�Z/,��	#�w�TAS�%xM='{�3�c.����Q>�|F܁���VaD9������Vf/�f�`�����4�c��;c��Ƌ.|��5�!�s�dMDk�� H�ߘ�t�-6�V��+���-@F�(�]��5'�k�^���0��F��9\�a������g��ӤNdy����Ңp�x�?��qZL�\����3�&���>��I�߿Mҷȣ��S�
9?_;������t����/f�`���ӥr�{���Rv�2Wi��lz�j����t�N�e��\^R�f��AuJ�]���e�һ%���Q�6��֢�u�J	,K8���L�.埇�hfh5pN��^i�~R��+؎V��z2:��>�yTY�O8��:/�h�j���L��o�B
(���"�:�T��f�X����;��*�H�(����H"͸�r(`����`��o�W�W� ���+C�A��'m������W�&d��:u{Sݥ�a�j�ř�|& ��`�Һ��roDn�|R����
�d�X[��������Q�"��)vM��#Yc�o0p��;2��|��t��#QN	 N����V�j����=_.[ړd3$b��۔�|;��&]	�߅��rU��V��L�`�?�'�s��9�(Kʋ��I$Z��q�`Q�1.gZu� �gV��h����m��I$YC?L����wD��	e�poi�_�B�-*�Q�[�u�toz�!�F�9�[bk����/>h�T���������s��+D�ՠ�
��s˵����t�rIE��v),݀n5���ffQ��GӞU����ݵ�����;���$�RI��]�-S�[�rk<���:��g~B��hѴO�DR�>O6�< U�"�i͂�ڂ�C�{����F7�$��V�G��0Lt;.��-o7��ٸ��/sp�XntB�~�b��(��y �5���X?�a"6��[Bs-��W��͘6�a[���&�J5���1��4��dm�0�r��a֍�T�Y<m ����K���B�.�e~|`W%�w�K�h]���j.�>�9�S�~���e��*-/�#���9�{�'!�l�PS��f��)�J�V3��;��h~9�jfa2E��&�~�V��s�{�n�c}�m-S35��h^�Aes���"ߑ�Q����j��d_C���8@��V�	BJ2�����~�޽���3 �-��}�܍d;NGo͢K8�2`[��� /�z�W�w]���V#wlR��jBg+�L�>�B�X��Ar��P�֋��T�Q��6G�����3$(-��?xi�W)wVBe�)��C��l�!�=�J����� ��9��>u���f�;'�qiĕ.:��G�N��j���=��9�%J	��a��(�U���BI��j䀜�1�w��\�}1)��V���'.�Yy�x��vs�X��ml� ��TEhVG.���\p15��?�f���=
t����b(&��( 0g控�~�����o^%H�-�o~<����R���Fe@bMW�2�5~-�©���[U@UmR;�-��Y���[�����A�/Xrc.�f��a�?��-���j|�`?܃�I��7&əD�#7*��<��^k���I�ߖ�V>��f��`�g�L�@=�ٷ�JYS����+%7oxt���D]��L�U�"{$f|�}�k�&�R^ԓL�tr�O�, l!ƈ�D���h����t�W?��bM�B�}�jec�}׋�r[�_+�<�A�Ү-�"��U�q�%;()��՝����H���	-�2߫S�fr)