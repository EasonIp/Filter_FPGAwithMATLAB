��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0]��?l
�4�!�ߦ����"�p8"	~��kB�J)��NbM�L��\jO��#y��r�3wA�y�}�S�{�����X�.m�lM(��R�g������B�*�NV�X-?����$��$�3�s�`;��y�@�u�ߗA�R�|�Ԝ�+�)]f��������҅i[^�"[��t��00��6�ĔR�*[�]�V�t���9�c%kz�Q��*N�| ea�z ��@������mU���h�$}���~�k��'C ��� Z���>J����ׯ,�'��3@akCc�U�U��?��a	6S��K󊀧uh���Z��&���9�+�)�b�В���ɀ�t�]z[��z�/`� !g�!*��P�����I�<V�� /o"�����@�g柅˳���.���5����9�i��)�!Ҏ���f8�vh�3�Z��ZC�:3Ϲ@�+��&�Ư���	��������Ϋ< �����"�����!b�'G����Z�!�R�l��Ã���3�����y���H�>����/{���?R%|��n6���gJ�2!b/ΧW�}�/FM��%����� ǜBk{�.�-�ّWz�*J`����'29�05�J�NYŪԚ��N�F2���������q��y�-Y�	����D�0���7��%��,�-.�O,P�y�w	�	�JT6'�Z�Ҟ���4��\��י����Ə��g��y��E��q�"�ӊ��N���H��`����=l�r�Ed�tP\��� �c�G�����/�('�'˷5����+��3]ʸ�:xõ|D,"���V�d�@��^Nm�D�dK�+l����E�ȟ��_��O�՟	����ȢM�6��������U�²��;偐&r�+����q���_j/�/3Ew�?'�Y���7ϓ,4���W�X�`]���eop�B����nIN�_K�����+�-�J��^��8��c�.)��+eR\_�-�/��?���}��@�|�VBp�zq�4���tsT������wPφ�(�,/��3�3~����]4�_x}����M��t,�Wv,�,�t����#���ιXz�^U��#|n���q��LlW�'_�@aQ�Ѽ��Սu�7�q��"�u$��NɌB�ֲ��bWE�i8�q�q�mG�It\�!�Q�~'���!0��G����i�A��h�¯=�;��x�F��H��s�����z�l,�������0����� H^�`8�a�Zl�߰��"v`�UB�u�1�5rk��d��Yu�F�� �R(��x�L�iy���w��<�DO9a�����GT9B��	�e�B)���ҍ����K���YjY<�Ј����R��yf�����F�����w`�a�&��qdMJ �%��/��H�4�Sқ�����e�2�>�YN4��r9�'U��ý�{03Ξm���d6�ͪ[�Pőz;".�l�j�ȹ���=R3O¢�2�cO��Zç�����
=�^CV���]m\����w��8���:��7Y�}hA0����!;4��P��d:Щ���Y�u9_c�|�w�l��N���Ը�� �����������o�V���8������3y'�s����P���<�Є�(#��B+�y��Ư�d[ܱ2���)]�+�,^ڀ�@3�]m���Q84/�����=�����%���4�d6d��z��h�B���V��I�$

29?��]�AK���T8���j��5͋�w_Gjڍ��3���B��)p熛�P٦� [
$�sŸS��؎B���UI�<	M��ٙ�H�qY,잸�TQ�h7�Rx`�b1���i�����
��a�4,�q����K{B0.���g�2p�.�\k)�^�(���]��8s��m�P���d���=Mr%�����w���h`�@�UqeJ<�hC�}��>�:�n�;��="q�|�����$~(�,������Ұ$j��she�F�u�D!�W��Y�}��0c�*� ��C�ؗߍ�?��MRb�����g��e�/;�#ܒ'
����R�eO�y����:�,���u�Ӛ��R<YZ�������?��U3�ɿ�ƹ�ښ�	e��`������0�	�wM4Jc2���2bM��)��c�!�Ӹ���_",�����tA+��E��@�+��[�&����K�\���՝�7TR4���.����6��={�g ~)$�D�:�w?�s[�X>�T���/H&���)�"4����0G��<Rc"��(�Z�Q��*�ԕ�&t���D���o�IP�	՝�I���{����K�<�%����H��)�h�^h#t�l��Su�"3C�v��_�7��i�J�i+.4Vz�Nvq�7��{s����W1M8�V�*G��g� �C���9-A��e?f=�$?�ۢ��%��sv��Rw