��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�J��"4�=�7(�T�JѺ�ő��,\��s���ӣ�F�؏!:��xb��[�S�8�$�8�0�A�l�1؆�h�{dY���4J������(�ʳ0�3U�/���{s,�E�OTR/!��L\�7v��b��UQ�"P:f�v?}��ޟ��j�m�Q��q[�մt8T8�霌aL���G`�@&���C�K⹅.Q�񴦙�r���2�p���i}S��%m��[�6�\��C㢝����O��eU�<̒W��Y8hܩ��8������eu �ۛ篶D�'	m�59�X�<���}�����;��Z��@�@�$o�A��4���o����`���[���(Z>]�
�,�D�[<X�5�3�3@��q*�A�9tI�i��_�@����������ԞB!9�ї��8q#�q~'�2����J�?��ͅ�G�B�
A&�^G����]8��o&>�Z+��(�y	��d��VN�+�0��6�oWؼ�a��h�5Ƕ�h{�ڿX�Ĩ���o���%&p�!��H:w\,��U������NW7@�At+��ڦ�4x��q$_��w��0�bh�(�_hL􎚭���d{��O�	���	2Q��7F������@?���� �xݤ�3`�4��Fa�V��vI�����d��>K_xd��c�ƽ�����Xa�K���+��*-K3���qU�𫞤�kq�R����uc�L��Mkb�/m��Xn6��#��2�/vc[��Cƚvŗ�(�㵂jE�X�����V�z�����xȈ���#������U#�2c,����uc>��NR�����I���"����%N�*H�A�|+�95�BD����,���қk/����/T m��Y5^�oŹ!��^�V̡?�J� ��}B 7�������Z��r���T��P��v� '{l%Uq�4�whY���,6�4�	)'A�5m�YJƀU�@Ak	��x�����KR�/+!�5k�ހ�K�f�j�&2�{�y���Lk!�"Ib���a �6�)P�K�K���֥����� �R���Tw�1rZ�����t�y}-�PUF��p��N"�����k

�/�4�@�Zy��l���R�{ ���g~�pI}q�Mc�;œ�c��9�S���I�-S@I��{��@}D O\��:'ɻTC����i�!��NG	ê9H���:��|�l['PH��ٓ8>��&��O8V�&��_Q֗�1��N�W6�_ڔrf��XB��r�8ψg9�a����ˠ9h����G�}�n'L�X�Q�����T_�DB,���7Z�����5!�h6X:G���0�/�,c���+a���K{��Y�&9=,c�@2wנ�㋜�̺"�}��89�Ԛ.q
��=,�w/�G�ZC�M�*��׮_��~�I0�cLC|�>���,���[�(X�Y��4��LG�
@�2��Œ��d�����â?ևɵd����`�%C�������j��'���nոvO��0֞^��z()ҙk��S�~��+l�o���P칲��� ��J���t]�|�U�e"��>5��I����har^�7=G,�1��G�	i����%32`�䄭�QCcQ%03H/O�
*	"�6��1'?�k�P �7N�*�VV�q.U@r�C�p��#�t5P���[ŏZ���y467W��̇�z>v��$��3���L@[n�I��q�I&�!�m/��	���9�t13-�Q�3��t�����Pm]p_��I�D�����^�y�&F�� �}O��:=���aj��AF{����'k�n�F�A��8xQ��,���6�������t����a�$�L���ZHw&�f{��~&lt�t�Ņ�H:u)b��#S��GD�U l�K�HiämY�WEen��D��<T����1⣡�n��y�âd�IP��g�A�֡I�F��ʘ����D�ѡ����٫F�/��)���6Is,��\��_&�l���=�]� 3����(���kQ-ܒ��w�������:?��ޑ��� �9��d��"���@�Ff�ʸ��O�X�Z�{<R_\c��-����|^_���bf��!L0���a��|��5~��응�M� .T� C�Yu����Bq���Pk��ivAy1����52*
R8Q���^	�s1%P8Em�ě��Zi�%N�\�Ծ*�w�?|����H
R翗�	o{��:�F3�:�|�c3��ҍi�pg�#��,x=��Q���c't�@��%>/bn�vnj����p��I`�~���̆$gS)D;q�I?Jk���+5Z�O-��s��aXܷB�Zcfq����)[��?p_%��~β���z�N�,�� 3?�S��+��fY���������}1z��L�Uj�|�N�҇�'Ҡ�nӴ?��1�#�W=����T����������F�X%��hĔ`P�ޖs8��jt��y���lF�(��sv�����y�L�L+j2���E%G[Y��p6-g��Zʚi��9"yY<��a����k[h�Nd������xi��o�� �������!N�h���8=#�;��;8D��Us^�wApBp#�	��'d��OQ�oO��iO�V,���Љ�9�1��t�\������X�agn'�}�tZ]�^"G� |��}��{��6~�#r8A{E��0Q#��Y�^���s���3]�ԓ��9��5��ٷ���.�a��zA�+�ãP�~su�]WLW��;���*fu���P�֮��<�ّ%AЧh�ccl����G�<���9Hc� ���fw��Ex�m�.׻��+��j�cV�x��*ׁa����a�x�R>�u aR����>T�v-V���'	4|�
�wm�
�W�BO�O*f
cښ�*�Y�a�Y�-�즀�^Ob�X�dwi�� g9�ʅY�s�����"���yV%#��Oz�^������JTd�q'��fDL�l���gI)�����u��e��~�;�x9>Ui-H��MDN�Vē�D�<ה�����{Rd���P�/bhY�5��d/[H���Tn���{;*��ć��8[T|��g�n^S(�]�@�.�G��a~�}��&�6�)� sq]��=�}O�����7�y8�B1V�o��N��%2	����n�U�АNJR=M)�h�#�5N6	��-�� VA8B�9�u�D>�W
�(K�y��Q��S}6
j�r��:EgW�c����Њ��^'�؆�O_��V���Q�g0�_A����Z0�M�1Jq�P�V���s�A@g��!�r�Qov�G�7�����׮�*P���i��_��T��"/�a1M�7�,v��w��uX��7�!����x �<�n�vk!D��8�� Q���H�R��le��'hފy_��{"[�nH	��p�^�(2�AN�$_�Si-w��	�)��){D��2�Z7)]l0���q�����p��(��p�Ҝ���)?�h�t���[,���u�J�H1NRژ�Cr,�3��wb�f�C��LϽ��(b'����
ld���Eh	�y� "��/���O���E4������8D������e��KT�ߨ�j�t4Z��`�Еq�H-���L���RW쀭!Pn"{6VmԞ�&���>:��_DA^R؅�,wR�<��^������*�����	�W��gs����	��_v�S��W�~�X�n�<F�r���AiN�&���إ�
�c�*xהGP`p,�)
�?��+�+�K7�[ X���Z�q`q�י�<%��kpB5ͫ��8��g,)F�r�Y��������<�HI
�4_9D��i���a�M�����[{�ȃL���IwP�`*F١�a��)S%&`D`�?��K���Ldί]�j��� g㪐1���P�۴ָ^�	9O�vR��ŝ�T�Խ.�k9���$~|[�����|7V&z-�N˥N����v��s��{� ׫��X��B��n�:�C
"`����������X	cT��8���R�7�Pբ\�*�ˢ�ݣ��l�U�4T�^Y&��v��-�*eĝ�7Cy*���>O�[z��Pʹĳ��@Ǣh7����&��ͻ�c���n�ױ��)�O�z�G��?%�7��0E`L�6����m��AvwS�un~(0�5��������h��u��M�B��`���+��b���c_w�|E1��u�7�~:�J@l~�{��_��cK�}6�YC	@u����;8�`��+��A�4�MR?R��&}Ü�'u	P��|jF���)X�qfq3��\�k�&�sq/1�U���������K��X�^��	f��u�A����<�,1.��yJ:b��~Й*���P�eb��2�WC�#��-N������)Mn!���^�PY������n�pmx��TO������o.��lU�M}�p��0_�u���P�g�~�W<��)7�`�4�L࿇�G�N�����Rn�z�P�l��}��@}͔H���Z�0
�#.d�3��~�KnP��yS����L�^��<�kL��7��#�\X֕��+�:g�$]��K��5O��R$�cA���r�;vl0��ߖ��y�5&�Ɯ<"Y �%��$R�1��"_BȖ��s�$���?��7a�։�p4B�u@�;zߙ':x�!1�	e<�HU��G��@M8��XphN�r��jHЫ�AAw���W�i�-nNA�gu!�
*��T��+6bP�:r 1�:+�_̀�
!��^�$���<cn��l*xX.�����f��d1�Ċ���-k7�r��)+Ee�i�N���1��X��;_��� �K ����Gq�(��ڐ�xO�<��{���wiQ�/��=�T'�m`y���� 8A�0�L�:�[(�&X�؏Vm�1h|���*,�>�<���E� ��w�h�R������<��Q�z�͌ �ݧ��[[r�b�*����T �0�;�	��Ub����Ty\4��m3��RZ�s 
��q���]�V۳��O���#�˿M nZ&.�U�;�7��3�'��v����u���V��{@�_�����Z�%��6�%���b�}ԉ!DȀ՛"���
����b�JQPD�l9ѐ-RN3 �������f���L��'��󞥚E&�I2E-:oGb�6|�b��i���i�b�-�ݏsQ���yˊ��9<Hn4��]��z����FiM�y�~İN>=�Z~����*�-�:Diw,eR9-U��ztE$�� ���\$�O,�hhϠ5����μ<Ta�˽�φ�xOL��򉿳�8�W����9z8��ݼ�w6u�ZǱ
d�nQ Ӑ�j�:���{����HN=��� ���6F�5(G��dդ���4IC�V�P��(�&�A���fA���9:0�.��k��p����KU���=��!���n>�F�#�p&����.|����dqm�n��%����i�0�+z�8}>�a�?�^�s���eԫ�(�Ց��RD^���G]U����q���:�gx��-PY@�s�/]��]H�������w΢Ev�a�-9zʓ�������R%+k�Ƙ��`���B�נ%g�6�/�����%&$�@��᫒Kn����nu��Ҵ��~�"I_�`�aZ�3~�~�%���B�rdk��m�~�-$�]�u\c��J��T"����C�U�zI ���΋Ez��4�3�ψ����Sf����_�}M�״)�2Kv��5�`�l`����j<��0��r�
�~y�ckj�S����-����+l�� �%���%3��1-�sS(D��ά@�k��?��KWO�;:7(��i3��:	4<X�n�An����ݵC�g./?�i�cɧ����#����K��Z�cb�i�#��*��;b���J��w�,:�*THN�Y_u/�����e�@��z�5hib�A��0
&�S��z�!}1��mr�jN����Ft����[z�����f�V�L�0t����g�`�	�)jl��6`BWd�t��Fk 7F;�k����~�Buɐ��t�EB0%���1o�S���f��4
;�������*J��~0�������rG�9ۓ��rrg�nb���J���1��"��!���֝�����.��oa,�xn_:BU���8VF��p�{�/���U�]l�̖N_��鲴BR
��1kqa�?�8l�e�Ί��?zD��g�/��n��Y<��S +eJ�N���8n8\��خZr�]��E��ڍ��~���%|c��fL�C��!��]�?2k�L���sC3ؽ�w�M������U�
b���PqȊO�H����Z���}�����.F~���Pk��'��?���G3a,oJ��qM*
i�h��u.M�@��y�z�1���ӄb=�J�/�F�Z��g]��ʸ�/	J}D�2S�����u���Fb�E&��x��O���z��*��{l��Hۄyt[7�D�29�]�f��;��KLc����4�J�v>����
5�#`�ي�&�6T��:� �Y�q��4����\	�8\��@�#�ǒ#G��1L�zՅ�}(,�ގ�?�& ��>��W]U������G��CB]ʵ�����q���]�	��,��$/��x��(k��^�B����FQA5��?�d^o��(�/�^�D%{'�Y,S�T���=�������={4I7�p�=8�z�zvy�\��@nF��~I#����*��P7��HD�'��D7���:���/`�)�d��Pm�I<�A%�2 pX#����]����o/�`���������:��m�⭞��U�A�na��U&mB�Zӏ����p�/E�]���;��oZ�t�lO	:�Ԣ͔F�3����2��"�-��M�߇���r�%I=mp��',H���������;=<�2rb��ǈU�=��2��[Ŋ��gV�C�X.��}�: ��v�N�H�(�{����PS��+��b�L-iMc:q?kρ��rukN6�QE�&�-~��b*�� ypO�AR%�9_�`���YOaedU�ɋ�����o�vnS+�eLh>���΀uX��(F]�%h7�P/�R^67"KL�������pV���h������+0�~w����|^"��^ ��z�S~���so�*�4I�g�T7u�	�7�W'�y� �z�ša+��Ɖ�ذ�CD��V���!��؊:�ޟ ���恓���ш}��09��bn��Sn�1j9��%d��5tpp0 ���ln�Nl����;��H��}�y�.ď�r�73te�/Y�d�u��Y�4%�&QxF��U�3x�ҝ�����+�K8���Wk_J	��b �zG$�u_f��� O��<�8D�ѓ����㴟�sH?��緘��[����M�l��e�3]�<d�Q9��z�(D2^6烠i���DB�&�k@�u�����'P��H&u�$�`�t?���՘*��ׁHt�j7B���`®X��
K���٫ z֠cT>0�"�cfo�w��↾�Wь�\{i��Hc�p}���������p��m��\������_X:��\���&�	M��D�<��I.��2��<��6w���K���H8��U��~�i��EN�9hr���ݪ�P�j5z�(�%/`�f���s�U��x���e����X���00 ���9:b�O�)�7���{Q���|4��3B���Ylא!T�Ӷ�������>�0��G"t�DosUd�`�_oS��7�B�������c=N���{Tz��a@G�Y����ޭ��{	ʖ�I~�Zh��14+�XI�b��s��+"����<0�13`��Z�CO݋��g�7P�岃V'-dP<WZx�tb�8�:��OO+�2�5E��S7	�|9}"J�Yﳌ�-���79��s�L�l��Ec9��h<����.��i���6m�_p �^�p4�}Cma� c����g
�-�K�}F�e�j���G��Kǐ��]i�8�#���e�\��|I`�fu�B�#�Y�܏�]����N��3|V����Ԥ��GP����"�4-�'qZB7���Rz1����h��d��]���������O?�O�1?Q���Ѫ��(�3��i��AU�qJSy)�����<����b�WV��;x�R���ּ�**�u����i�\#��fhǗ|࿙�l�i�d�z��?fy��{(��@0a7w��]Q��V�}Z�2o��Ԥ����۱�b"~/	ӼUC�m���u�K¡/6�G���e/�$����q��|���RZ}��I��A��ϮB�k��`iZU�7S#���f|"bm$���ց��AH���,�KxƩ6��S��vŝ��ͺ��K����Bu�I��	�2}��4��;�9��r]���Y�s|gP�<��?DQ���s�u{���'�~�)���L&��wK>����r��/�wV�û$j�S���a6�� �Cx[�i��zu;n�1P����h(�4lQ �K�D�Y�r�M>i�M�+ͽ�2�4=W�7}q��\���2�F��Ges! �f�<����4��o
[��94��`��y� �B�ϞҫPJ�ȼ;/��]%)?�Μ�ƪ�W~j��2em�N
�$��fƹ$6�є#D�E�x\/V��2^�Jd7hq |mC
��IB�P!��W�}�9M��� Fh�.�����h4h�&�0�8v�6I�ޫ)��x�vA�s���0R��� ]= �j�<�!�«"Z�'��m5eBͽ�PE��*+��B;�yn�t��+�LAY���X��G�cܾ�[HHp�n�'�\��{��ތBb�㰋��-�5�x�\�#�9�E�hگ�?Ap�ȇ	�LO���Z��N?��
Z��z?w�wcW��+�/v�	
Q}̦_���0�a��^�P���T.	[C6s&oB�4����dPE�*�{+jT�ܝf�-��6�j�]0Fe�9��6�e��y� y+="�$
yj�՚i�SN�4��IО�,{�,S�E[~)�{^�*i)��{�z\ >TV\�Ov�[gPv�s�ա����l�*���Jj���_t�|~���3��lm����59T��Hb
RT2E|�Ñjnr�������0����b(Q�X1�7�<��8�ٓ�A���t�LDj�y�MfK#�c�=�z^"���0Q6c�$ܦ�rbiz��"�j�@�4y�k�1
ʽy��>w:̀՟� �	�g޷��N�Cۋ��=���}�����J`��+i�AA6����!��6L5�u/��Γψrl���.�dv��0?����"Z`<>���ƏE�ҧ�E#z�����?�v	�kJD.��b�.�8�
!��%��~Ϳ��i�H<��ST�fJ��q�#�	����g�xM]�_5��3q.����v,UkCGKo�_t]b�R�.�8���}&T��J���,�4�9���g/K����
ȲEܴ3�����q�,�,]�B����";��P�����ZG�l�J�!uS�L�e�����e�E� Q�΄b6���)���oj�P�˗�s��BŢ���Kβ�]��
�^$�[�vX;F�5�I��?�����]��w����WE_U�<�`���%���@k��I@�&�):���Sd�	��M!�Ǯ��뷺�������du�<:�w @P{f�k��sV�!�c�	{� ��J
�AsQ�6���Wy:��ls-�������|M��J�����>�]I��%��M֐�
�Iӷ�Ʈ�D��`v���aS&��r@D���}�ð�U�=g�q�ď��7z���.q$K�CO���Hꅯ�V�����As��3e��׷�[?�9z		V�}dj�Q�Z�7rD��y��
��=��krY/x~����FBJ���q�a���7bQk����#wR�I|��]��S�)FH�x(��n�7��v�D\��!��?x���y�m�$,hY�	�x%�]�/R��ܙNAƉ���!���??���6��<ǿ�������!sꩩ)�:6��A��)���򩣯h���0���;yҤ�)ߪ���0�6۳4E��(d<uK���������9v���Oo�(��iX�������.�\˟o�@��?�v'2 ߅ܝ!��V0Ոm5��NzӐ��Zop+]�5yk=S���"	,YbP`hAl�!��;X�n��Wu��m``;�jg\֠od�!�5��F�ݠ��#)�tY���@/? ���R���N���[�sj�����8�iڧ�n]��D�T3k#�ᰞj�`�!_�S4�h��k����+�6�0SOA�8!�?6K����@�A2Q��q�sJp���(�M�-Yr�
�e�[����.��h�%]���2�:*��~�;�W�8�[J�t�L������*�~|ZȮ���i�٬K:+a�1΁Z�����"�&��X�*�P��iM�/��&����p��v�fi׸�+������������I��r�j�p���!7��	:r��SGL����3�㿪���1�&�~y�Uf���Ok��r,�[N���5߸���yM��1�Ǽ�g���'0�Q��U�_L���j�c��*�p߻� 1s]�b�K���r�fa,b���tS�_�cV&��6���̵���|�"�w|)�7&�=I^ѓ\�8uצ+�3���<��!K�QY��������Hy��O��=0��r�?�We�󸲫��E7t"r#U����n���i�8�|�߁9 =ķ4��EƝh�eaS���_�S���`��n,eZԡU(�@���>u
�TJy��/�PR}�r�h�������T��`�h'#U�p�-�m�")��!�}����W�:w�f�5?*��!��^�(q,��#:�唀?���~��޾ ^S�D^��J��u��1	w�]��_6�5��������{�?��f�4Mk䆱�k4�l�k�8�f��:|�
MsNm^py���Ÿ�.k�^��e� ��,�Ht�spMw�kj��}�`�Ӂ�vn|��Ɉ��'Yy��ch+�R���U�ٸx)G��Z�w�7�Z��ؚt�#���P4�y1��I�*�g�ǜX"�k��svv&\�V,}dNK3�G]��^E��L_�aͻ�'�FK�v������,��m�R�e&E�{9�s
����a���l��v���0HD|��D΀���!���QfX�c�%������c���؈�*����Q�Y��@� !�P|��.⥶�6��WN�R�8	\Wd<?.�����,8�٧�6����ՂO@��1c��֒��ߣ�aak��RO։93y�
ֶ��X&���A�@|�i$�TD���!��-�FN4���yq���I��2�oOu� K�� FI��ءJ��E�抍�XE(-c�и'3m��7���y�)�k�������)5oOHM�N2�O2����iI)K�Y]<��t$��o��)��S��Ҿ���ւ?��A��G�"L�Z�̽���_�W���Z��Z���������Q�ug�,j����0�<�zz�R����J�z��k��޷[p�&��ȵ/]��D���Ǣ`������ ������Td���z�lݕ�D^������8'���6;m�kk|
)=`��<��q.�L3}�ض��oP ����]�F�ګq��!�Z�U��5ј�* C���o1�?���vʇ�.��"���1��/�׺�L����ћC���被"�F�6���۫n�2a���XĖ^a�
�*���O.�o��uHC猞GR�ʝ��<�R/��fYލ8"aY�UOM|�L�Tv�P�5Ge2��#rD�q	�\d��l1Ug�YuP�rp���k}�$E�����hJ�u�Qգ����uc����`(cˋ��P^��J��~(v���g@�T��#ĊhŸJv��N`"{�-�\;.@��<d
{��q���f��V>����,���捃<.9S Š��/8_]�$��0z�Й�_�gvU&Cђ q��cp,��3�YE���]�Z���۠D#_u7��1o��e�秊OE��삟��6ݪ�Ŵi8�`��77�~ Ϲ%rN��d{��p�: �e#����9?@�����6��c�W�!��*�qt�<WI��}����"���������ͱH�Grlc�w�i^=E�!ƻ�}&���ۚϊ�t�`��OC�~}�F��U8V�S��R�u�����F�[ Z���N�>���@L��F{&;��7�$fXU�R��g�5�3l2�Mja�.�f�Wχ�i�;�M�?��4�J�tY����T�3;;��[�WD~2�/�h�?�1�I<��T����׬��Y\���ҭ�`�5JLTg��C}�)�N읎�@u1o`���۩�K2.=#�̣RU�Ϧ����������^s|,�<ën��F���pJ#��?�,-�}D6qw�V�eڵ���rR��L��*��DM����Rג��tQP��ӈtG]j��A�si�\���) �p���q�eW�U,��z���P�`�]�V�����l��*_Yś�q52\�l�r>���Kx�����K�ڼA����VT��q���Y�4����1^޹�w�r�Cq VO���&r��F,F�!��Q	b)ic���$ƿ���+�m欱Y�Dy_�"��N�b����}��,���*�b� }*����+چI�S��
�*r��ȤGXs?G��?�W��X��7J#DeZ��N��"� n0I
3�}M�=u�2�+Z�Y�'z����'�w@8>u%�;CMے��I(+Ĥ:��}XuZx�l��
���伕=�N|��>�L��@�ZJ=�wxs��"��2_>��S�F��	��b�	M�L�m���q��'@�|���;�d}<��Ь oN]G��j��E�B�.��zTv�"�3i���'����L���i�튯��&�%X�O�UӞ#���(9�&��������d�C�g��q�a/��`�^*N>�@֠Sg�]4�e�����rȽB�%5`�µ9�X����
ceq���e�7�-��3 �m�FyD�Wz�;��h�~Ҭe�$D�i�j�g7$b��2��P�)\���� ��]��"����IzR"��O�m�Lx��Y۬�nJ����wҮ���5���b]��]���줧�O��e$R�v[�r���<%<O�K�Zm3�y�q� �#�2f�t��r���wq)�����7����k�W��M"����K/\�^�Mv2-�ōIa��a^�;�Zf��!
���&~i�6����aŋv��W�mD5'��y�҅�԰
�̀�2J4s�A�����m�]�F��u��d���N=[������1j�Gw���(}/+��ؿ򨚤�M/����>Bi'�;[;dqN��`��NGmD�K�V��+��15�b��Wz$����y��`��m����[4��y 2�\��_�SOx��YU�OAQ[]��U��'����z��K�Xa�"�C)��h��V睂) �j�|jh=����F�O�:�~�;R5$�[�@^''��*ک��8�LHHBI+�4� ��"�;L��>�k�,|��)@�[S�c��Xt��xNb�gxj���}>9Ǣ�,�E�8S%[e�DR���2��"a66CG�N��]�#I�g�8��@�@>��,C����f�.�<�д9Z��_�P���U���(��/�C�qͻR�A`������uq�͹�-�SNGB�R����2��q�FJ���P�O�<p��Y�`U�9ŢJ��M"q�]��꼺���tw�n~���&WƑ�d>M��y��th�_I�ǯ�k�j,�"T�3���/)�V��ƲD�|N�5���I��L�	�>z��vα��`�ϙ�5�F��]c8v��j�ԗ�7�9i@(��/&V�#�K-���G�f7�	�[*�F<7����v�`���||����9 �(���R@�*r;s'.�z����E�I�/�.&K�k��͇ԛ�Q�Ŕ<��q^\���3�v��;˷�;*�M�L��I��R�
��Ss<i�/���6r5�Ś}J;c��f��L�#J�xUd�X�9�	Ƿ�����n_}>��w�Z�;�Lk����WI����|h�̓�5�sD�%��N��q�]�;lo#iB�$O�|S�K�I�Ί�{'�ZQ�쇪����+�X�Y��o#譓�b�L��}t����}����<b�y��P�Ld�G��N�*� (� ���R�Vlg��&p�,D1�ᅱ�M��bL ��V3�;F���Jq����w��ͦ]�)Cjƭ��Y�tH�=��R�=+`?Q��)(��S�Pn�������<ezᩕ�mYPa��o�I��pD����O�R"a�O�%};��9���ӷR8`�+�F���/���t�A�A��=�O���ZK���F����>��|VR?��P��B��o^e���_�� "׉��Fn���(H�Ө�9����COp�ht�q[�����V�Ө	E)'�}�M��+��qė!�r�8�j�L~&ݫ���r���f�G�ܼ�}W�d=NB��YM5l!_����o�]�ż��z�����/!\SIXl��h6/�B*'�`=��ᛞ�t�r�����?["C�|���V�&Ҭ.�h ��d�b�wԻ>�ؐ�5��5�-��2|�	�m{�������xfyL����>ȍE���:�EvwCj_#�������A�-t��g%�8�9����T�����|�h�a���)2�#�V�'�R�<p�/��ٶK"�ET��7��r����P�Y�s��c�a��4�/���٢���g�J�9&��6��g��`	�aXy쓾����=iGP��16��J��������uE���+�p�\�`��k�S��O�:KEѴ�!�vh��/.S�. �.�H���t0:�R��'ʬ-d#Z�(���ez�6TAH���i�)V&p��]��5����Dج/���r������w�!��h#����t�&�{�s�<��߸fs�E���Q�ٚK���rоt��@9�;��fP�%>S�y�_]"�5@~]����D��l���T����oD��Wlu�'6j��uR�����k櫼�"�n;��Q��\M�L����L�SN;���h��vn�G��K1H�k���(W�7�p\S h
��2�1M+>u�Y�v�3�SA���g+�4v���&��Պ-~����kw_J�B�ļ+�S':�����5ϗ�f"��ً�h~��c�v�b�{@�<�p�/e녦��z��c��.'I.ACsF"岱�I�h�CA���k�-P,� ����O��b��؝B�,��$���z�¿��܍A���!��1��.ğOoX,�A����|�UTKqs��|e�u�W��;T��o�����v2y���v�7�	�%��Q'�h��A���{�Q?������q@KkD/P�܇c��� =� >&C7w:%��@�ˮ�w�j]�M��t�#�J<�h{B�"�Ro�P
��s�%��?�a5N���~,趸���,��Ț��P�C,��w� u)��L8�3;�|�ҰX��qӌ�4S-zP#L���,�Gx`������N_,=��RU��(���pQ
G&c%Y�*'�6�Y6�<<?�!F����v���,���7��3�����' �Z�z���j}wA����I�\̺��g ��v��R!o���Pۻ�@M�o*�n��"[L��"̀)d�g��qtd(@�Vy��b��<==򰵑`�t��C
FV�t�Y�?_uE����(�����g��v�[0��li���j1�[^)��b>y��4P�j4�qjDzg�G���5�֋���{��CX$�^h/�ˇ�� 4(C"��Nz�Q�`Z�3�  \�xm5'J�=te*����p@^���gF0��>��,��yYO����O(g����0�d�G�C�e�Eo	�6��mJ�����p�3������6I�Ҁ-�'$)�P.�n�-���~�
ͷw�@j�w�M��
�M)�q�5����֐��@�]]���W(�SM��&!sݖ%���R�Ӌ��PMW��G�����W�\�>�I��W�oY����W��n��o�VL�p� {k��ADB���7�~�$>f"��� Зg�}Y�Bc#L���Y_�d�D_p���Z���>��W��gܯ���2����rFD#�n<������)-�o7�M:��T�A)>�c}�[_�멡���p�E�ާ_u��!��P��/3k�0?�#�g%2��y��m9�$_���ߪ�4+p(�ff�l~�g
���>˿7f�F\Q2G�U�=��bW�r��
n�=�qFY��3�©*؄����d��]ޯ;�R�b#��cHݝ+|hpGSI�G��s|��_1���<f׎5;{1S�C���!	�ƪIvc#�-�(Ҵ� )�+�P���<�TAjo�
b��g*���6"4��q���0u�9���/y��v��d�I���՚K,�0���e̸���O3�r6��ݤ��[蹬[�� Ϫ[����W-�(`��C�*!�]�{^�~%2Q�Ĩ@{)������ܧ*I@v>��sKz��#3���3Ņ�S��6�a�ʒv��A�D�� B�����~�*�fe��t��p&(H���.�_��������s��*��I�B� u3_[2lQq�<&:�C�$�%?lU���Z�y3� !������cf-����,0��o�7��������P?��Y0X�1Lw�`@��dF�F�7������r�Vw��(ů^ vE�聏�&�Ɲy!1
en����q�K$�n�Aĸ���Jm��j���Y��C%'V�:�Y}�����'ֳ�ѭ���au�f�q�:�7�`��s�Tr�Â�V��kKq�a����N?�Gf\��^��%��q�g���$��*	�,�Y\죆8W	��,y	�k,���-�D���V6�~�(L�(8<{0��m��U����A�[?��2��k� .õU�}��@H���B������&T!�2�M�}˗7�ۺ�����ZJhe�������M]&+{��7�Iy���>Xq���Q/�W�ve,(�0�p���,�j�+��˨�1���A�p��O&�ɺ�����$�߁ڔ�E�lqX�aO�>�B܇�:R[�٪l�e���#;inFe�==�"h���:�{]�:�K���c�a����Vi�9���F�I���ȏ��k���o�a�7O�/K��C��樨j�~�#.�&ɤk,�x5l�L7��%�����m��������R$�!ogF����a*�?���օF�SΑ�#���D���-J��CZJ��jH�u�2��Go� �3�m�&��d�ޗ��?<��d�&��
V��͙ ��p^673�H��g'l��)��l�����ZT<K&L�Z���2��fB!���J��� a;:�X�[)����J�����X5�Q9����|�d�u7�4ӗ�s�h��gvF��Â�p0*b4�o5��Ѝǰ��h�sL��>��G�KĐ1V���w�O�D@��IH�$&?��6�yX��ЪޒĨ �>�����>�b��I��"�,i�&�v��*���G>]&��U�r��z���E��o�/�	�GE���܍��θ�a�ǐ=�R���s��0���tY��˙�˃��.� <م���L�|����� �爻������6����D�$->��uEUUjfe�4��:BQ�ra�]5�r��z+B+<�K�Y���0-bk`�G���ǁ��s�8�v�<���1��G�O��7������2��N���%�ǋG%\���S��� ,1�O���Jq�.��
����`u-')@��C���"��sOmK��TW�����u��c������)����M�i-�^�6ύo�}��G���[*���?�W�?�p��BI�ft��`�d�SY�����������rK���u2�W~@fJ�������g�ZHb�:�sSC�%Fl�j�"2��7�&�p�t&�����~uN������k	�p�1̃��b�%�1��/�Q#tdm���Gm�uօ �Z���[�Y2�� �R�
n	2p?��M$6ξan,���E����I�]o��������5�	���gV��%��Ɏ]˫��n��L�Ʒk����"��{d_�Pd�� %K��'&�\-����YH� ��+���Ƃ�S��s!��D�7�G3��8��\�����D����p�aOq���gB>k U=�C���~V�S����46���P/G�p��b�t?%;�A�ne41��t-䰇��?-	$����&�O ����V�\�?�g2!4�&��x�&ft}H.n�����[?�Nʐ��J�N��m��~���7S�h)h}#TMD�%u��+߈���qb������XQҬ
$I���u�}�?uy����	�0VO�`o ��fS�l�=������j�_�Y��'W����',):7m�j�=���l��U�H�	��ۢac��@I�I!\������S_��D�_D�ਫ਼�_f����n[�'t��J�I����(����9g�%}�񅪹�rVN�LH��#���\��Q��[#ԟ@��-��]��A�E��Pl�Kp*O�^���"�L��8�|��~N <֪�����;��E��Hu}���S����A2�F 0���l_��2��L���_�X�`�Y<s�xծ� W���ڃج!����k�g����{��/`��G�"���¯���������}�{�'l˲�`�S�z��F'Y�ٞ0Js�z�/�z}��ΓǊ�O>< @�����"gW2������乇	�G�;���e�2�T|��󪃻R=c��@��s�j��=͌�X�죵�c�ڭv���n|)sxܘ�����p���$�������yS
��3�$�.��� �0��ʫ�,�Q#k�v�R�UD��f��#@N��YG.�AɊǣ��9�5��G3��-|�r��O�![ژ�k}2�x�7������1�:�\&	�c�ӛ��$�H�C��i�`�mU�V��X�o�{�R��'��^tV�	�v3����_i՗��$�4�i[vAz�s!(s̟�Cg0E�ȶz�CI��]~w�H��
��%Y�1��-�u�Nk����Jw�M��,������%{��9=&`�����N�㣰��k�����YI�v�����#�rb{k��4S���T�_�bc��>SZ'�5|�"�R�7瞕�R�1'���\�^yQm��6�u���T'@oh�)ْ�����d\d�GU.�a��}�"�[����������nI�(��i>��jC�!��_K�ǲ��ۧ�&2��w���V��+M�o��>���@vH8���vp�LA$���e�X���:�DX��O���L�_9_��Q�|���O�������ԣh�Mƺ��������/!�Ֆ&ϿPi�|��X���+�v���ǁb��v�����l���$r���N@m�,�ʐ�r���~�4Z���)�'BYq�]�c�4񾂾�_̢b�]ԧ9�w]�ƭ6['hA)+������;f���F�}@�Ӂ
��"�C;h���yR@��_C�>m�2����?��#�S7�x���0ɵgLkM���ќ:����o���W�ӏ��n]�n�_����0��f�C�CBѓ��M.��s}h^��'T<����l,8'j�G�d"�8T��;�v}����-��q��e��I@i �r�)�L��WV,�2��h�2�-f%[��:1,9���`���Xu1#��5�P1ݭnU�/���	`�e�f5�,`�����>�V��>&�1�Gn���p`;t9�y�u�xƥ��?<p5��Tҋ�k_>���q:��u}|�߷.-�b�"���������0��0q�:���Ac]�eû�G}'7��a)ye�OV�~@`k@��Х��b��@;Y�?���'$�"��u����zLO�Y
4�w��9E-塚�c'ֈ���l���"��$�q��5(�h cRg�E�D�461���"&�Pz������XE��)y�0��S��+��*:cԤ/k*��͉sI=PUn
c.=c�-n��w��b:��`��i<��]$:�����4?��Y��٨�נp���~L�3y��_I���H�@_�m�n��E��V���%0l�n0���'B��'+�dSX��T�q���=�Na�YI�>�z���sC��w#S"�q��:�J/��&�ѵvc~~?]��c֠��
��t������Yi���v�U�=��u��R��UEg<}��7C�
>���3��a)�s��)O�g�٘�}�IFzN1�A�1���۪B���?6�M��g�p|���2%�%s�ۂ��L5�M��QZeX�����b���ee�>��sN}�w%��/���6��J�4uǓ s	�|�LQ}��g9���VQ|�xK�V�V����_����0�Y������'x�i�y�1D�-럳��ꮄc��E	�ƙ��CK��Se�+��1��`�k~
X,���:ɇ*�xM��"�0��"�1��V��p?a_t��̮�M ܻ �aF$F4 �y��`��
2���G��t^"u���9]D���	ϰ׹8��a��!X���F����`<E_�߳�d�GZ�/ߍ���8��=��N)�0W㨭�c�Ї�08wmj�8+�<ֽ�U��0no�%Ns�g>�&�h�?�m��C�@d3T�f�7��l��˾'����#�?��a
���O�׾��X*���9ou1�p^:�-4 :��=�L�l�cm[AR�����)����#B�\���>��]�G��i��"]��MÌ�p����0�i�A�y��d�Z�|��rEF$�p��n����;q�[��s9��(����~��CL
 U�� ����Q��Ք?�+4��X�����Tٰ��ػ`X�uӏ���InH��q3�y-�6N��E6��`>�˛ϒ�
�4��k��<���;��yW���ڮ��Z�8[y�C��1-أ�p˗I{����H?нϭ��l��g�̉�D�'Wc���	
݅�<c�38�Nf����<��Vj�0�ѫ��<%�rs����9�9�OnI����Hp���m�� �7�߿W����WJu��_�4\ȹ��ɅVkfo?����];�@	#� ��6Iڀp!��ܬ?ӣ�Jlf��@k�A`��X��%�����̗���m:��<[�f�$� ?C���N�+a���/��ތ`L�-�k�:z�s]�m֐`�3$ؼ��<�W#H	v.�iCp\?D�hʸ�8i�I]�(���Ϸ�jt-�fA�2����ytŀP \p*����󐫏�*�)��b��0�:�+\������1��違2u#�v�i8V�FL�6ts���+oi9�ɡ>�IC���8'c�X3�[�_�E���T�2L��&Y�p-й�A~�SO#����b���&�� �}����9W��%l����Ζ�I;�Ċ`�dB��H��B
�����K3ta�o��v��;��.5M��]Q~s�G��66�7�#�y{�%��Ͼ|=��gS=��iD�Q�͇��I4��̤�2��ftQ�A+#���5+�?��{η7���a�p.aCL.��Q�d֦�ϗ9�-Yz	ܳ����d������21ocq�v��.g�.�U6�=����ZL�1���7y�5�c���k�K;4���y�f�� ؠ�G�H9aҎ�j�����S��I�@�f�XQ���Ś����r-8���<��G���	#m7f:!�S�
�S��U�*A������7�:$j��A^�WQ�N������̓-�����9t]�P��>#��<^=6>�e�d	�zg27@D^�%���� �V�v@�-#*�̥Ly�i�W�D����C����q���{_>�FH��7������Ml�V�Zn��(��b�_M��E�x��B��8��Ձ�c�-)�4����� ���=�z��V�K���~o�kn=P5!��������8q4l�OC���f^��Ӵ�۲w��)p��y9��Hɠ]�mK^�(W��M��ӻ���y��T6�=�n=-Na���CzGM�lm���I��X+�\�.�{�'�H(\P����^�%����S+���p�K��3pn=k��Ekv�f� �[af�9�ؕ'��	��I���0�is0�����D�=�a�����)������Z�課QHCz_�D�C�;����!��~�L�_����9�[��qb��=㫂�?��Z����`����(��ȇ��#�V���!��O`%�A�FO2�>��ǺI��@[(�UV��V�Tc���>oYȳ���\1x�Q�>-��Рns�EJ(o�O[}G�=Q6��������3���\;��
G�& �P�B�q�%s�r�Fu�ęp�Ո��.���gEff8G8S�|^��&wR�aA7JW�=�i��<��{y�#��D
;�O�:�4�kAr~�GL�X�?�^��;8�qPJ������5��7XK���,}G$AY�*���"aJ�b!�@e��t���碒��()�얈-C���R��0��G�鋌�h���a�D=m�8��-;����?S��������O�tly��'��Vkc��?k���rq� Bvj�.ː�5�/�c��ⵖf�86�L]�v��'�'۷k�F�h�^]{Hb�� ���ۛ*��^�XYZ��]m���rr,-�u�^��*�^^?Z�A=[j��;G�L��9*}`ڋ�u���d�s�^s�	�/7#-�I��A����t�v�%M%������1��� ]X"9c�٬��x_��xm�ǰ?ˡ.��=����H��@��&��nZj3ۛ�\R�Џ�diC :�uo�[�.pr)�S�747'��h%TIW���#4�:�9Y`��n���e�|7�!�Fm�OyTe\����Gs��ռ��50�Pz;���f��[c��\ُ�j�+-�Xj9�'b���4B��2�w�����֨ES�)v6�I����Ƃ�v�Ү�r?x��a��v��t�<�kO��F�g��MF�z�L����r� ��=�1�\"h��Ә5(R�j�C�Ͻc��4��3[CH�O�1�
�W����ĈB��ɣ�.����$���b�+�y��f%�5,60&le����3�7M�%{�Ұ�ZIH�w��0�'?�s��=ఘ mk�sM�b���pG(?�qK���H�.��i/�#_e�2�rL�t���w-[8��!l˶E���=�5wm��Cқ7�I��Y뇞�FϲG�EU��b`G$�� (��~k�E�,�0��f	ġ*N,snzK�į��2�M�	��bqK���+�mM6�P{̳���k�D�{_l��J�	�7�3�=��K�-�>x�<L���i&��F�!�0s�#�)j�ߢ���&6;X��[�|V��A�iӥ���vV� 'ai ���%���4O�8���t���ڄ��l�*`���VF��D:
�ms<���_�n|�' �����T
�`ҎeyW�K���(�Q?��H��^�=�}��?��{����窓����}�A`$���@���7�Q�5��H��Y?���t"�t�T`�Ӛd.۵a(�H�CO'�ʛ��'��^65X�j�W�e>���f���5�z��Rz;��)���݆���*��7�\��б�1�g�Z�h�AA��燗���d���%Q���0�-C�[�^��/*�������P��G��a,�Ș=7�A�ih���0 -�vDv��0�#�ܸ�("X+��f�Rc���*�?mf�������/r�Z�wA]�/����i,����mD�}9��FJ�tj�����8�^�t4�v�D�i�����yCBeKtoҵ�|`���3V��ȇq�_��YТ�iQ�W̘,��?��Jص�����i[��}��:�nN�"g��$��AYX��5�(��|p�5Q��ԕt���:�3ux�M�њ���ɩ=��|C%uŪ_o���'�����Lk�мN�׿�>G� �k%|�h�e4 {�4b�
, �|�����t�#�tp@�E�_#�tP����Zm��>�#����˜��8��7�Y��7�#�ah֣��� .���`T�C#f���֓�_
��b"@�J���.�m��������?��������wN��ѻf�6*pv ��6io���ޭ���d���hx7S:�k��67U8a���i���d|��ME�a �.�����u�3�4m�F�oϦ�^�X��Z�;*��[�yA���K�;zth �%E� R E���u��|���8������@(R? �w����d*���"�)�����N�E�Ɔ&�X��D�����SYh;^�����?���3A��R��8ٿC� �%9{�yC!�<�!�P<t���Et��K���������?��'���]7�[�q��UB⦬�]�\�S��<�o�|V����KIc-��qg)"���՝^��d.����w�S��h�0,#�ܱ���ڇQ�� ��dq6�]S�@�~��>�� ��['���5Sϳ>/�B1���Q�:�A9	l��7L����6�@�@,�4y�zG��V�B�X^��<�}908��q�j���0����MtJ�qe̶�!��Ocj�`C�w�xkIye�q� �n��ש���S�e|�q�w�:������5y5��:�)h�n��m��̢�Û1�"�m�������f�q^��GtLe�ޞH�Q��g�]1��ˡ'���v-��hȓ_���J���D��K�<�r�z���~���2>��u8�wR���/��+8T�Z���"���� t�c��9���ѫ�1��.�'U����VL�w�"f�@@�z�jrf�9��U�ta�yN$�N�h"�%=�GF&p�y�fb!@��+��o��
�~z��Ӕ���"\, e�r�ٗ!���7��>N�-j���ې)wc/\[��V׭R�YDf,�rl���e�_6�%���@N�X�T�O8$\��"N�L�ޖs��yq�gi��`ѣ�I�p���/�]�BYnԦcYF6ؖ� jW$��������l�*�y�$-���%	`ꋡ,�L��s��!�����c���E��O�O��WB5}��5��Z�m��N5Q�Y3|�ѧ�+���W�f���<���Bo�b.l9A����yk�}[�-�)@�+no	��<g��@H�=��,nܴ其U�PzaS�����+��Q����q����_��Q�37�2����;��)�}���n�����l�"+���9��{q�	"����Gm����=�;e%���g�&����*�ʽ�6�-�muz���-��������\��gyA������P��� �/���1�D4k$�K��/��{jn2��Х��<��Z!m �'4�1P)�L�-R��%�O��͌xʗߋ|X�}3��{���������3~m����yX��>gЊ[���\��=M�
Uv_�%V���f%Z\KA��Q\@�ܭ�p>;d֖���JH,�\/��b���#��}^�w��U()�g�|ڢ�A�!��P��~�_@���L�ZBf��]��fތ�8�΂-k*X���������
�]GY���HC��e�����"Ek�إ���!-��[��
��~|ܘ��� �W�j�ʿ�8{�}|�.���T\��y�ɇ��"�:B/8�V5�U�!�>BQ���|?v�;`��-o(o�(K�!Nz�p+Ƣz��e�bҝ���f�6���\^��ሂ?�p����u���[�ގ��^��3���T0&r;��#o��Ӂd��7���VxD�� ;�%|�/6z����)$�D>�$����m�g���䩓E��
\a��	�d&,��%+����(|p.�@��k̉$��̾X�ĳ�q�H�o��mM�q�w"��&��m�y[���{?P,ǃ
� 1���g��˷��!ܷ��3��Z�����f2)���xͦ=Ų�+.�H�LI�V�Z/g�\�W[���n�QH8���*?�t��K(V=h�z�8�v������_�`SPAT*�F�A��4s�1�p)�Hr�o/C0Ȣv�_��$�r< n�a�	]���=萑�_������z�cWp��@�~����n�'��m��,1�j�"Pv3?"��g���O���;
������@���
��a����9��\�ޓO�s�w�a����џ0��}y��~7Q��r�e"��������ۨ QwU���4s������.XY�?�O�_S;}R2Wm�  >,�	}�)"��x*��Xi��M!��\"��:�*ƭ�E�f����_�E:D�>���c�Q� �~]S�y�nٷ�����X�����փ���Է�>)���*Rr�3M��ȩ5A8%�Z�5��ج���cl�wo�\������g��+8��s�(�J�K�9F���d��0j�����Y�ķ�%a�-���.g��NH�{a�!өG�y<9�iz�����j��;f<��ŋGx�����R.x�(-{�Ȭ�F��"�y�D�P�t���00w��u�����6��d�We��43�z���?�z�ݑ,U\�:\/�$��
ѐ3�!��\�퓊׌T,.F����K>ɨ=	YUt|��Ҷ��Lw]Z11{�G˙M�p��5�n��mT�5�nb${R��X;�t��x�c��nQ�zu!��6g慳OM�VwM�(����wgx��fh��B�I��E"(����%�Ie�!�w�{���r`��=BM=&V]!��i��}NS$�����y��I0gE�P�5����o�GE�(0�J7oݺ����!��c���{�����?T}z��o���Ylg
��m��m�ȉ��i����ʅ' @Aݱ��hd�Zd��|;a
n��S���������� R`d&'�>�h��[��P�-�9� �
.ϾI ��B/�)�9e���b=Pn&Ҟ��͉�ѓ2-G��~���,����}��/�(�R`D�:�ؿ̄����q�ي�p���w$߭�N�a�83�*�Q7�A���$����~qΜh�C'�ժ�:�S���l_����=�Q���'��O&+0����ˈ5*��r�f%m,ط�VF
ZVM�*H	`dd��N�N�w�;�"�Ȉ�R�1�S;���!֛ȼ��7�gQ�L�X��1�t�xN�RwQ�ś�N�HY�端��a�_{�����34&��(�������Y}�Y�܇� م���a�X-_���>7h�.�?�%"����"�IA�N�\G��X=d�dUdh�z� �Z[��`g��9c����)�����>�(��W�?��,�Xg��l8����ҭV "�ӻ��MF9�u�d�
bQ��Au��Ϛf"h�J݉�è�ڹ'���t2�d�/����c�H%-���0㩀�k�^�e�Pc��n�4G&���;b$?��Em��" Գ�S@�{cu�rE�p��͒,�̭jA=-L�=�(�4Mk�Ku(���v@�\�Q��
D<v�U��v�-D��q_��Y��E��q<���5��Ȗ|@o�)1=j�*|���J��8ҏ ae�p���<�	�3���ۺJ�Mb
n�6eF�?[�8Q��p�~L��b/f#��]�����c�'��sZ��2���H����w8k���ڊ ��A���ˉ)���<ͼ�j��r��*�D���ԙy1��d�ftg�ؚv%q�+�<]�ڼ�RVT��mOvG�ۍ����!{���3g��S�X������(��,�����M��&�Ó6��a�Q��*A�9�z�s�iLw�����i���㝰fX]ִͬ?�Xn�s�0�׮ٶ�'Ź��ʹ	݉k{o�v��M�68��PIcH������#P#V�;� n]3E�^f⽞-ȶ�+qP�	��o˦9��H+stmm�P5z���G�f5*a7l\R��Q��b�}|����c����ǞX+՝�c��CTAe��Ə-��p!c�0�O?>��L܂��Jv��(+�������oWo����^�-P�C<`C�[�ad��6Z��C�;�����7�Z �G�9I���U��c�����5���m�@�@lSPbS']����G�U9ť\5��@=�x���skL��s�ڋ y%ٯ=��*4���f.�$�I(���&�#���ל¶!���p�qp�W�;w~w/F�S	[�9M�Y�0b���u�s����H���BG���*�*wqܓ�����V�."�a�n�/�ŦD{A���a-c��Q�#�m@o��A���a���yF�8�պ�Z��kY�/vo�0��(����^&��Tx���8@� ��RRz�E�C�)?��0�{9d�����`��
��8$�>����~�>w��:ف��x���ަ�FXJ֏�7Dδg��ҥʖ�fc{ʦ���r%������J�`vǱ{�K�{�Ϲ�������H��8��Z̺ �E��N�9m<�gC��XUT��,P�	h5�,�7`��ur����a��KAO]�
��j�9���f��J>���(�:��$}KL3K�A|���6�$�"޸u�5*���+݋!�#ZQA��2�i��?gObCI�����!D��6_�tr�׮X^��R�~Y��IQ����q�Q�Q�j��*�K3��9K>�==����Es���a<�`�o�{��A�UE����D��\�xq�/	�������v���F�|�xK���������V%=��a/2�n6{�:)5 �:e�٢���'��'�Fp�覦RK1���M'B*��_b��4�1 �[1^Y+}��o۝��S��-�v��Ҟu�F/�Nk'b[Hb\Ƽz�G�k�@��g�IR\��~��nG�9 �#�3,���Ѓ�������	����)HL-�����H%8��{�j�#F�h�=����S���W�3X���O\�0��˗�MBz�g��k���F�K[�dj>�8�M��Ȍ�}Q���$� 
/�l  ����Dec��ȯ^�ǐ�c=
 �
aC�>�%��=�S3����FfeC2�;
�a�{��c�z1~��6Kak�$T���Q���*{�
�-�=\6V�	�����A�l�I��b�X���������6�G�C��9�9P4�*� �J�T�Z��{�b �=n!z��8�`��	#��uk��J��FO�4�D�-�y��3�
cK�6��.F�����x��ؖ&�Ș
�L�,�n�Y+g||�7+6g��[@M���"�9G�1�P�~E��>B�#�A���ܼ��5A\�����[����+����?��V��w�A�E��.߫m����v/��ym���P8�)ƄJ�����H����eb���� �{�e��fo�7�]� ��ua�I�"���S�[�uQ{�R�����[E��9xJ��*ln�#oy�S���r�n�ďP��W���K�yr�f���6��8��F��ֲ�6��mw�����r�y@k*&��y��UrF����kE��*��$�08����"a�=Dnp4�~�n�� �|{?���Q��!���'��b	5W���c,�U(�����׾�/�|n��O�//B#�&R��Kq�Ih��޿��>~�
�# ��ĥ���Y�<E�2#rpv����Z�gş6�=��̷N$Y���1>�������|ad�j�bL��M�ˬ��� xL�1�7xV��6�)�w�\r��=��sy��Z��䳺����B0�k��/+�pվ�n)ϓ��1���3�7��vM������oTG����������"�ӊl�|�J<�q������;5�_YM�O[D^�a����u��ϊ(��#ϐ�;h��4�r�b:�ş4��Kކ-Ӳ�k�M6��oē$�Q���7�S 	�)^���ZT�Ja��t�?�<���Jj���IF�������pX�@(�����}��$��!� x��Z�6XL+Sp!�[�~��&���v�gû؟g5}Ϲ�nP��y��Ԏ}�7�ԏ�dZ����ɵJ{+�A�R}�o;���U1�G��x�����[��k~y�d�i����bg@
��j��U��-���������O�	LrC�N۲�B4 �~L�\����B`a���ht����
I�&��� ��|%?�߃��ރ���G��{:V�L��Լ/!6�t��~�M7_�ɕ�}m{������/�zU����;s�5e�S��@qc��k<�R�k�#���5�[A���H�����e�>$�;X1(i�Y���+I��osxg�u��F�:�Bq4圏 �u��_ƃb�+4�R�Gn�oV�s@�_n+}��@�-��	���#�%���9~;u|wY;�;uT�>�����͏ȕ�p��|��4�ڜ�J�Gh�׳d`�S&��2��S@�n �ho`��20�| =�t��t��N�e�� ˆ������G,V�����B����0$�~���˖���MLՀE��E�aLA�G9?�Ś�^�$}�GM�pv��L�A(�L�Q t��77���{R�=��������	xKg���\^j8m��ֆf��A��!,�^�Q�f�7�P��p^e��X���fK��P�M��m/���$�-m��ń�����;���{`z��;���`���u35�Os%(8��=-}�9�6�,t.���-%ةQm��Gl�ˑ��0��2Ź͚rbQ�e�G[��[�����?�l7� �Vg��[z7ԗ�J�=lE�6�o'�=���^:4P�V�Y�.]s2'=Fg�����I�$�%-H���,n��������k3������e�:��ȧ����H���/��{jPMurE�u��V^������X�'�I�ȿ�>>� %�\��U��Kd�1¢I6�O:��4Ya?��J�·�
�$¨��1�Y$�1�2�Cv<Oo��<�{�
�<Xj�y�(M�I��r\O�����l@<[�ĉ,�Uҏ��P9�[���k��fT�\:���t"��vQwoEÕ~*ke���3��x��&��F�dG����.A4�'^�ZB�,)��i,u"8��c��g[Q
�N�,�7����d�ٹ*d���e�4�����8+5C%x�/O�86�tSi��#'�|;��s �6|mSQ�A�Ԛ�6�����6!�P�AN	���>/����R�&�ԍ�e�����-~��S��G��|��Bv�e��uV�
�6Lnؾ�?0��0I��:��@W۹案p�k"��W�Lw�&>xّ���k��B�a�m��'=�ls9Q�`	5���M-m��h��@6�u�-{��>��d8O	���VZ���1�NK�A��\�V%p?��.�K��<�L�Y��ܪ��韉3>Y)��گ����J��� �Ps��-Eu��.�S�9�8�����w���R�[�Ng�����LVe��p#v�z��0���ե�� ho�����0Q:��|6��>��}P3����tI��+~|�O��&1Hx��NݟK݋:��@���2�ښd�+�n�T� +�X�"A�GS�[��z��km��E+���ƃ� �5����(�Nu�/�2(8NP�<-�����>A1	��	�7F~�oY��^-�b�0���&9;@x�ݣ#���n�1�oԣz`�Yfx: �ɨ�yȢsf�������s5adkI"A�0�R��R��4.n�}z��I�������t���r��h��d���h���\{��L�G 9B���r^.�yԊ	*������p�k��_����3��8��{��C���k�4=��8���Y\HB�\���wy���]�;H7,ɵN�&x�^� �6�{�N��a��b++����'��`Ơ~@�o��t,ܯ�t r�s'Ґ®���4��1N���"g�j~���&c�yq��MI���Yg��d�	2?V]��`"+����Vc�c��Y�,�`�|è�j^%�a�L2��c"phH��	���T�* ௿6����{�������6
 1U��R��m�59M$�	l_�n�b��ᷝ��t�]�e[b�D��G:�,�%��D$�����cd/��7��UB=ғ<{�_������Z�|U��lD�]�g:��?4�/�#J�����LTNP�a|�{���(S0������
r}�,�Te���=�q�є���Œ�6�)q�c�0YV6u{T)���.��0���ڦaF
SlgA
���料�I΃*g�x�ъ��5JR�7�}B�
�7�GIEN�p��xcsLPl]R1���i�%��U�%���{�}��g��ELWyҏ8��� �H�+,O�#�L�`k�-M��ZX��n�7(!v�w�h�<=?n����iʒao;Ꮕ�?��aD�P�X#�$t�4 �W���S�R
,Ȟ�)8� �R������`�-ӂD��ϣ�!6>?>Zg��\sǴa�eRE���.r2��߁�OA��~MV��o�
܃��|?���=�k�J8�>�b�eY�<O��*$��ߚ�X<6I��j\m����G�����=�/;�����ޙc\�����q���5��s�G��W"�)��O���B�\?ϴѥ���S���G�7�RzpA���s�8�B㽽��3��������AFx���*�u\Z�*"C
+�p9L��`o ՟��<�BRt�Fz��f���c���u�`j�_	�U�ٓ� �w{�}�H��c��/nhE��cұw)3���&�����m���HL]����U��?A�e	���Z>��C�S��5�&�ն29��3��hQ�,Ѯ|*��z��3Ր��˹�셂�7yv��� {���v�ٱ�L�z.�@��G�<�$�*��+a2tMr���w�2����Jn���X#����&p�=�AI�r��5�N�ZgT��wv�@t![�l���=���i�Me)��A�/ع�O<�;�
�~B<}��5��+�b������8)?1T-���x�_+ݩ�	��է:<���
$A;�}V�L�2����a���A��k7;k����!-���|�d~��Z���kt���W��ǀL2�N4)��� �L�,˘�I��q���'qe��)��c=L�,�?|]�g4"w��*�i&�ף��Lb���Xmҿ���k�J�س��䩚1�Yŧ���H�g���@	�~C<�υ��QFg�zq<����鲆��M�߲�}#x�|���D�>k����A��#��L����uH �-��ܿ����g�@��: �p{N��ro[�1��n����syd bL��x��x�_N$��?��ݾ���:o�, �	����",��´1�M�k��&�K����ś
�������^�$MS #2���@g쵓6�jv�>��|߽E-�\`��{^��:�ד���qU���ό�}ڦ,�X�5��B��Nnr�͟��;,�'�Ů�[��1��3;��W ̽�*�F��h�~������,�\^���3T�f���<��е�66�Q�!��)��_��~�W�F���c�U46Uhi�������(H0�|?4wa�Y�����0���8b�t6Xi���*ڭL�C�>�,ʾⅸ�D6�n^�J��7����i{�����-���F,�Ntԛ��wx�W��r�@�	��corY���˕X��Le��d:�C#Q*�Hc��};�gǀ����It�'T��"|�Ȕ��_J�<a.�E�,GM��^��������wgs#U�e�p��;U�?�&[�D��KT�$u ���m�/��Qֱ�g��
��*>� ��W�]%���E�I�������ve"T�vDL5�]���JP�ڷE��jKE	�L��T�V�乼T��8~d{�-Xc �X�aou"�!;iO���IYܱǜ˱KoP�:S�E�¢��qf��)���%�`^�T��ľ�4� ��9����%�y&��X�@����6JM�VG]/#w5��f����pa1���s�'�EL]�c��Sm� �&7|��'~�U_���f95�R�7)߼�k2:�Ë�A�����Pg�vc��&�k$.�݉C�n=�}�J�'A�/�K	�7/вҲf���e�1TzS`!����q� �HO=�{��"R���0�B&�9I��tc�#�L3p��V���x�v ��#3�˩�D��d0��F^=�թ����)h��/���}��D `��v���d�䉓�n����ՇV̒_�Ѐ�2'�r� R����I[�z���wlx��N�[MQ��_��w�]��_��R�7=�����o������ �*��I�J�f�0��ᅤ�3��&.|!��=��a���bo�K�	>9W2��s��>�zM+�W��&�l����	�`?�if�������`,�,*��".K��x������rb��1��zǤ�+��[ZVP4�%���v4�k�|�{b�����t���>�-U*`3��f��)BBt�`��/�~YJ`���G�]�*OCp��2�A	�4����*R�q��/`rF�O��L��؃���/� Ԍ�_?-W��(*RV�X��G�����i��؅��@����[�gM�� JrA^�<�m�I%Fv&6 �3����Pz�<7-i�Q���]��mc$+�.�Uj�3o1�5^~�.�A3��_#ɪ�|8o�+{���g�\ڹ$
�t	�ǳ}�0��	�ț�Kфpo�eO��&��ke���/+p�{�p@݂sp�(��A2�M��>�I��U> ��������)N�T��3���>�F�`t�󤭟��Hr�^�����4�'��_��Iс�� ��DK�s����(|������`GW�h%��4�� S����q�����Bd��v�1�X�S?��Q_����	޲찍���|��'�e�į�(�cU�`?�7��*�o5�B[�-ݠ�;DI̑)����L�!�C���M�Q{���b��B�2������)�o�h��h]�`vCh�������X{��ٞ
�Y����b�LGà>�5�a����QN�7�j9�3�Q�����7���96po��56�y^�mz�(҃���u9���:@5�| 5T��T��s#�B��͗��'Mq�SW~N�<�m�;�ŰO���>�]��#���0��$�B�>�|����	ȼ6��7�V�U~�$n��k��!_3YG����z���Ô�I'#K~�*XJ*�˄�o���¸�T���8����M�c*a\�D��i�2��fd�ꈔ	U";���4�؏sv�಑��i|�f��0�~K�JL; �n+/k'�0;_\����eu��3�l�p<���e$b��Yg!B��Pj��A�.'��rA��]pw�_b�N�X�����Z�mQ�t���ȝ�rY�F�d���7�5�4�;�Ot�/���u=��N�!�y��=j�~���e����n���po��<��#!�w8cC߾�K�v�����l$����ҦV�A�R����o�ܩ�!��ҏ+5WTM&v����U[��N$;��rr�N<noy=W(����k}�$%�,SW6$宠e7p������@~cdA�N���SY;3�F@:��=*�+G�y=�� `]�fNS޻7�S����F�q'V`d��J
I�*"�c
�4�V�/ʸb��6Fg�5)��Y�Ёce;I�`�[?����H2�Q�ҙV�&Q3�ۑ����C4�k�p�?��5�T�� :�F?g�D��`V23�!v��j����c�l�5}�/qg�Y�.&��Mo��(HT�ވ���/�iR��wQizn�8��#���Z��aZ��T!\�QZ�%+Z��1�����?�L8?���:���S�T�&�RO'�WB��"�$�	p�`o҇��S��J�p��1.��+���N>=��$,\�8��rV� Bm�6,U>/�W�P���:��$8���\"���9��{��%���:��\N�'}ey>/Q���2�V�͝	���0\U��@��vY�T��4�F�S8X� ��;���gs���Υ� &h�l1o(����#���h�-�u�<|�$f�u�E��Cw�%:�X��%o9fp¥z0�^ly�	[S�$�byw��w�g�rM���Fv��9s���q)K2���`Ln�wqks�"km���]�͕�w�����@1�̐�܄�3k2�e׮�+�k|�%��i���P���+.��2N�n &-�Ȑ�D�>4��H'�������&�P(������x���ޒS <����#"��:dD�b�_���z�c�Fi�?x7��"(5[r5-+���V��٨�y3
pjHX*$�%5;@w�F�� |����~H���+�Eػ��WL}��3e�d��߱�a�J�q�Z�2T�٘7��Ǎ�$�Rz�F�ӌ���3���Z]U�T��D0��nNMm�3�V~��W�0\��dqU���~�by�'Nx�j��h�wt���M���٭�r�o1<B�)�R�m�y8*g&��S%0���m-�{�������T��'�&�!8��I�0paa���)p6}d���\Ӵ�?��E�:;l�C���Ы�p���������?��&�ä��$�̼�8b6��#�^�]�Nt�ܻ�J��S�ϫ�GmO5J!u�H/�s�9	&;B�n���ɢ�"����J�h`~��G��*�11�G��B�(��J^����~M�a�����$Hrq�R9�y�␰����J�e�D_�S!�rrA{��t�<�[o ހ:��-��g6�Px�SOi����+�ن��y��pl��QMT>82{�!1���2W��g���c�{Y��o��R	�B�@�f�hg������%�d�G��b�<�/�h�A5�Npi��U����{��g�*]	`,1����br⳸�nb2�^�[�?���{w��Fw�nZr�
�@؉]���	{z�����穮���
n�R}�QK��nqٖyp1$Q����{t�{,<��V�L�=�X���ieuR��H�R�������%L&Vb`'��5|MEu�Io>��/�݆�����~N<P��qSH
��Pd�.LI���4���Z���|�[%��W���ڶ?"K�5���+����`U2��"=r��τ�u����)��K5I:x�E-.�d)0@I3wi'��K�u컾GB �0t���T�U�������t��|�4��%jd�됒��~*�"�M��j*���j���¥f�>(%Tz'#R/j���T1�����-��晿��vM�f�!�:K��44c����vk?������9��ư�΀�Ծ���\X����i�"�a�O�2�^����:j{�)�K��eIr7IG`�Ŕ�*~x�qV.>�hd��]M�m�Y�$��3���l�8|����Do�HTU���4���P2���Z wr�Wj�^��
o
��0���B�z#@����L�t9�=\����:��c2���c؍/-���NLc&��uL��E���jT?�׉�Ond4j��@q���Y�q+R�Ոޑ=���� =���z#�7�  ��^�v'َK�c�)b*j'�zع��Z���*�-&%l�kw�A�k���v2���(�XP,�A0Blh#�tecgcړt!蕊�W0�)�P/1
ybnutk��ԝ��mXcZ��٠��4���|>b��� p�7o�{E��,-l�L5�!E�/�Ɛ���p��L�����Sa��� �8ݎd<S`�z���p�lL1@^s`��/�;����d��9F7������zWCíP3���$1kS|����cI��,ļ7��'7a���~K��M�G�L�V��@���%��}^L�,+C��y��mqK	"k���#��+V<��D��&��[v�����7󆈲ǎ��j/\[�

��%���<�����fm�@�}1CNv,W7���`|�/#�r��L#�g�k�'5���׊,j�g0��2���F�*�S.��}�y*pP�{�^Z��}ɛ�����#�X@:r�ʁ��(Uט@K0o�e�/ �x�Q��U�U�<�&����+�*��1f�����)̪�n�C�FfC�p�j�푔5YFV�`n�+�?&Qe� (+���
c!�����!۹V$xf����{�Zp�@�ە�E��2�̯��|�p�b)9̴M��ձA�8i���sS|!��D�q����l �|H��x���Bs?<ـMq"&�%	,���\��s�Lu5����Q���,�r�xSN���%�|�Zt�cr_���ڿ=E	w��������)�|��l{몧�6�H��1�7%@,�j�����:#'�=q?����x,:웣�b�}�v�\�ϗ�����`�1Z�T��:l�Sw�ژ�Q����ᨺ�VC)9����'�S\�H�|���,��if���L�*��W퍆?c(��Aׅ4�oelZߦT")��,����_��^���KCݽl���6�^h�#�W�d��hh�c_�9��.���;��MD��i�c\�v����Y���.}Ců������;>���4��m��O#K!����b�v<<�fd�\�*W�"ի��u�X�������jE�l�O��K��KS�E��e�ZT.L�f-/���_������m�r�F�����Sc ���i����n"M�b��;��誰⊍�����DED�-��7�̌��\�}����#�s���##f���:����^����2B+]�M��=Pr;gl@wD������� �ڧ��͇�~A����o���aƐ=�]�S�!�m����s�%5	gg���т����aK��-m6/̄�����+�*�Y��Ԍ��� ���\�8X{_,�p��r_�v~���d,��j:�����2��pq�Q�(���!Wb���K�]c�Ӊ@|գ��G9����(���1:���F��NQ�bD뉾1�_����1��j���L?N�!��I<?��!���D�d�~GC�3Б�+���"��e��YL�(�d����f�vs�aNv)��H+O9��K�]��\JpG�3�J�Iv!��ȃ�����?�Ap��ð���S�1��Y�w��6K�T�u�v����n�s�2Vݩ���H�� �588��}v}����f���v���7Ub���
b#H�`�cml�w`�v���N����d�+)��ͳ�����-;���O�7wx �2�ҘÖ���:eo&�����2���f�[��/܆�"{���������ss*5�K_ `;#s\�����"��7��Լ}��$
�su!��}3�L��P����[0
i[��?���}Om���}m��3�C����:9���$m]/D���g�xU�� sj�g��h]q�T��cdO_~���3��˃��x����V�O�<Q���nA����K���O}�YWK5f��Ҷ���h�U���&+iRC{���N�A�Å��\�S;r�����植������f��l�Y&C�u�qx�#���c��i
�cjc��~�#���Z\$X,Ժ.��$�s�}u�z���<�����J]HV��9w�����F�*�c��i�k���q���F�G6sT�?`�[�*�E����_���ˈ]������P X\�+���(,�V�ǣ�#R8�}��<�ƀ5a�I�4\��;��� �.!��^3a��j����.��x�����V��EQ�%K�و�cŬ�C{�6h���2c��F����d�M�&)>�JGM���@�%�@J��\�$H��������L7Q�&��NHq�4����8��mF%k�dx���|9�Q�����F<@V�=�$n�/�c�F��J�<����˿O�4jz xf,���v?���f�ؕV�M_�<. H�q�ӥ�m����'�(S��C�3?�uz'yʸo������x�Ty�fL����;T����!x�5k�'i�V;�Hy�1g�"k�d�U���V�4H�`�F0�g�4�4l�.~��?�w�[��Y��4�:n�'�4;}����9B�7&�I"�N��^+z�BJ����H@Y�3�Mc1��ּs"%ǳ��'3_�8�9L�S]��`�zn ��G�\<�(Ç;��>P�㲂�6�_����',�jp�.�IK��(�����p�'�X�ZAU�ۻ��i���q��%#aX,Q#��5�^�$�}�gve�u.��܋�{`��.�y�)���˰�|ˎ�4�b���O�&-�BY���t�����4c���7�������||ݍ��vo�T����,^4�a�����I��-�� J�����'Z!�������D��ӄ�|�|x󨔙�	�N龤��\�/��]����=���f9R{V^�7��3:NN�f�Y!� �FR78�e߲_��#u��x��S��^'����K�Ⱥ���ؘ�tf�ѹ�4踴��5@�`�2�+���?j ����J����V�C���^���l�{ w�`�-����dc��F�¾e�#X��CU�6���t�OJ���*�R!�l�h������7��d��A�,k�b�,����,�T>�S��v���Kz
`��et�1�<B�K�*���6�@�vR$�g4�I�舗ܒ]�ڱ���x��M=HS�<M��`�(��3-:�K�u֚��k?�q!̒�U��9O4K��{���d�f���k����o��L�(+:�I�غ-�&��#%5�#!�>m��h��C�-��9��§*!�;��a�
�0��z�����&N,�"��$ 	wiZ��\����8i���܏?��9��{S�SJ���$~oi��IF��l�.�j{����E0WQa�:-����U;��@w��*D����<"��5I�Z�������(�yH�Dj��:� W5���9�0��Ŭ�0&Oؠ���'�DJBā�t�͘O�!U"/��mB���}@����9�-M��б]fS�÷��U|�%���5�G��T4P�>3徭��
�r1���C�{��F�'�*36�T�(��6,�r׺�Q)�o+���5�z2bd�6EAu�ċ��}�`sɪH��g�ʎ*_RS�!����jz���b��q='�|���.�.4�KS}luT;$jr''����B漳�t�y���e�Hx~�LV|ܻ���Pn���K���2�mT�w8V_Kkfض�(ߔXGK��/IsF���E8�
�{7�~?6�HZ��a��M�=A�dн}н�P��?��� Jj���������D&���O���������hD���q���q<�6S�X`b��g�VgP��#���˰�`P��4+7���z&8��9��ѤOW���TF��Ρ��v�_���5ɵ%l�B6��`�SD�ďs���	�8���F�n�8�qHo��01��ֵ�Ӥr �'X��h#0����3�����ץ�hBb�hf���3�.	�V�CI-wc�,�uì�q�P���\�e���Y-F>Ε�qwi�7 F�7�@����i_퍾Nq K� u��بH`3�U_��vn�j��2���*��:��M���['ssc<b�a�g��<�#�uS��p	��_��aK��ǉ����e���)8���5+c�Y�4�ʱi�ō#������~-�=���b3Z�|�hA��{/QS7B��"�f�0���O��G�i���%����9����$�SO�K�<e�A2��i�Ӿ��
;�t�u����zg9�O���[�-YT�|8)� ��x��@�ʺ�&�`l�ˎ�x}�0 ��V��o��=���+UЊ�� 
�np��=���/�Mї���?���^����DrO7�*O?����G���&�><a����~�`S\R�����j�&͈x�s���h��'��
�2#��NjL���i��R�L�9n� s����8��[�G��/:Qq3�H-�<��9��mOT4C/:�|��b!�U�0~��'��5�w�ׅ���١40�h6��V����8�������K�ce��H��^�eb�	/��1�B'A%�xŒ��m4��u�&�ɼ��]&l�N�׬��2Ӥ�\{�V�X��UMBېW�����x/���>�˲�Ƌ?6l�Ō�þ��GZ�O�XrEDe5}������	�}౻�\������t�f���?n�I����h$Fv��p����1ϰLlm�r.��а��@E׺�h�N.3�>>���]�\��I~�)��B����4�\�cbRi��5�g�uh$�/��/�}�c�բ�Ε^���32+dI�2�)P���M��UXݪ��6�|E}F=��Ջ���	�r�q��|0�$b�`{�C�ml��^�����nz۵���lǴ�ʽ����Ofm-�Ub�\�+�J
�	�Z��OG�]/_�I,$X���ү��Bn�"�.�������%+D�B�$�g�{n�&�	]�%V��V��g�[�3���I:\��Ԑ~P�J�M���?Cȗ�d��Ϣ�O�=�w]H������0�ͽW�)����1�Iy%��[*5��r�9/�/��Q
!�~/������ �i�C1��$�����I-4��I�!l�z�+u�cwO���f}3�<
 ���Fj�︝�]�dd:���{��F�t����a�Y��i~c���ݦE n�T3���ƣ��Y뇫�ъc&�=F�Z����ў7 #�W/�|�E����!L��u�E�cH_��襒tZ����x���ܞi��D��l�
VE=s�`l�!i�y�ɳmb6�8mߌ�෸����)"�V~"m�P{��Q��a7���Wys���@}��p���wQ����� �F�'��n��U��w����`�7*ܡ��x���O�Mp�����3��n�-�ڶ��}��K˰�E#�uH��a�*�nQ1N�������`�XW˝��Q e@���r�p�V���Φ��K#����_��f�Ty(�p����<�>��^��z��mRdK�uzˮ56�W���e����Mi�0�*�w4�S�ap<��� ,���A���d�)< ��"kL�=��X����������r\��-.&�㙆�KWn��:{���y7v�Yn��&U�ݍ�WY�C���)%�YA��~������~Y\�Ɲ��D*=Iʆ��7'4���1x[|��������=���c��'���w�h�b�R�0��(35+l:R�i�R��s�������.թ�L��)W�ۧ�Ψ���j�����>�c݀Ȯ~�3���� 7�D�ܵ 4bC�&��� �f� �ޣ����:��u�ǟ�/�c�,w�g>�_�p�ڜ���6D���I���3��D�;I�ywN���9���4��}�w��,o?-I5��ibX� ������ád�ﶵ�I�41�#�(:|�P;I.#YZR��B3ł -�
��:L.o��nK�_��I>~"Gj:�"1�*j���XH~8�X/��Z"w�#@:wp����'��m�\�3(���/��
oĥ����Be�����P���śLT��1����zG�E�V��T�t��t�9��R;Wh�~�И�A��'2Y��l�Q$$�k��������g��Y]o��lD9�r1���g��{��)�V��Bƒ���8�fk��W���tcz�7�/"zYXg�`��"�[���1�D�U�|0^N��zb`'�_�n_5�Cx��8�T��^ӂ �ȝr0c�w�+�89Z��ݟ=u%��	��z��3QjoC��/~w�~����@����k�JaR�D�~�#ک!R�qx��D���Z䀴&���H��K�۴Xf�8��ێ�#XnD^�H�_�x'���XŪWH�;�i�$�Q���~�l���vQ# �w�[�Hi:�`��j�x���P�f�*F�{��,�� ���-1`;p� ��<�-e���H5B��~�0��J�L�f��c��#��H��7�᝸v�x۔��b����{]r3M�Q3���FI�Q^9b�iJ����Kf]�/����e�yC�gR!��unsH��̑<b����Q׎!�l84f&�?ʆ��o.�&��\bۇ\j���PUe_5�n:�R�j����oj �e;H�a�ģX�T+rl����d�z�%q�?����B��U����&��~�-�Y���b �� !���8��%y��o҂�x���'�/�/�ϾS�@7G"�����'5��kpBZ�D�g�K�����i�65*����2cvk�V�ɩc����ELκ�"k졳��8�k>G�O5�ޓ�yD7iU�W+^e���ʘ9Y^��R�$G?RZ}��<Fh�����㌳M�!�v��5iI�5� �l$�.�ӧI{z��Y#A�^Uxֺ#�v(�>��FD��F��'������r���6_U���z��ΎaS<��������j�V����ɑ��?Z��N@I��������.ږ�Hq�kC���dsBc����
���F���0��,�a-��D[oA�;���JG|�h)I>�=�mƇ�M��b�4��FCz����+�u��%�֑K����d�����1T��6��].FR��#ٛ�X �hs�V$�6Q��@g��
55>��%�V��ch�T����ҥo���sWq|ݤ/�X�
Q�I�I!ݲPp�%=_�X0�6��X�H!c�<�@�+�J�%L �t�KH�~(������������-�t���%�}cl���U'��a ���+�~j��j��;ߨC�JP���N�������&w�hk��f@��������e0�B��:S��Y$	���5��s���Ș9��]����k��[��X3	�`h~�A(fT�z0��couy���F�e�)(5�^�W��\y��4���_��|눀87���|�/
���Y:� �h��������<�n+p6���P��$�A��ʃ��C<�����2;n[�"f�=�]�,W��8B�4O�Ǡr�[,l��6"��;"��.��j��V!U,%0n��?Z���ݠ����Z����*��[�2��������,�1��e�oZ�J��	"�V-<��mQ6�[m�w
#�̖Mh7B�"
"��{�\(���I+o|(-����ў}�yV9����0Q} |�E&�-=+A�{��<�&]��Jz|��'I���˪�Etң�RE�#�>(�
�0��Z�w�o&Bώb��B�Ef���3#��# 8�2"���4����j�K�� �P�k�ދl�?ށM�!��n�a7��_ּhj���K�۵񝶴68�5�	/��B�>H�P�ΰ��!#�0�����Yf��ܹ�c>�����A�yc�{w"�ˋ��jV�K`dj��m	�!�NMQ#����t��0ã����ע�=:#�S�p�W5� ,�C(m�=7��4���vS���}J��o�\�^��$.�T�
~O������a�C����t3um�"�S�DnO��6��q * [M�.�$���W� �8k���Ѵ���K&\�����EG��$�_3~�0�_ X�6�<k�����\�\���Q�A&���SA5)��QƊ�N6��r��eÛ���Ҹ��_�09��6���}0��n(P�t���g !bJ
����׫��m@�x�!}��PԴ$o`��c2��u�� �¿K9�aA�:������^?4+�|zL�l��M�by-za;�y�!���˛#4F\fO�Z��ܨH�{����l�@$�j��*��ɢ���OD��O2��m�J^���A@�G��y/V���)O��G�d���"�Լ�=�����o�����b���A���fL@�+B�_n��"!(XU����!�}��i��� f\�����]>u�6<�����-��	�˗0z���zSK@�8��8�z[:8m$8�C����/o��G6��o|G�aI�� 1a2)-�'FiƮYy�/��>�<��!G�&�#��%(9v�;
��OQ�7<�3�n��}��NDKvs��Pc��y�֫�5�V�ԧ�T̆�մ��HF?=�LON�C���8��?~13+8������H��7bjB�c� 킉n��:����@�(�I�~�ēC\�(���FR1�R��k�]Y��	��neOԀvsWm6Yu?�~��0f�c2� S���\�y�⛓�n\����ͯx�Y�y��vE������F�Lv�Gղ@�x�v��Ѿx�V�j��Y�~Z�?��������X��������k�s��ҰI���8�0����s	Q��t���Ѯu����i�|���H�5Ub�����A':8��#�w�b�A~O'���!NM�;1�I�Z���g#���=��p�
�\�^���`$0� ���}/hns:\�b�\_�0{
7N�*�]�I�����Z]7-�ei�ɔ�Y�ny%�4�@�J�Ԑ���D��4i��y�����<t�e�@u���iA��
Q�M5�hH����)<�R=���e�.r���W'�����mo�4�?`֠@^Q��x�ؑ����,��x��*�+�i# JV����v#�CQ0e̤�?Q{r<ߔ�`�c˯�՞u�����mT�Y�Z?��)Q�3�Rۖ�#�O�I_���3��|? 
u��d͏}��p���N�YV��y���\��$^2&c�C�f l9�B���`��t�3�%g�Q)@����¾��Og�O��� b֪�	"���M6�!�Y�?3�3�68СWZ{܌�ن�l����Sn��q]���s/f|�̵����(�ƗKD`C��q���Z:
��V�6�f �� +��H-0���J��9=�/��+�Ǘe9����k�I��h4��Dw�4�Q=m�� m}��.K�f1�(����p�Af���P�[�?���z��z(�і��׽����Ҩ����Z�Ϛ���Yu�K�E[�ᚗz����zq4	m�&��8 D����`
��6�-��X�{��P��Kz�$��{�I���Nb'��A��N� Z����vd�,	�<9+�=#�����lއ���nSkg'�r��9^_O]�[Y�I��~s��
�F�W�j�;�z�7��7��c�i�-����o���Э�l��������`�K����4y���Vbi����=�E;�bœh����W	�L�k��Y�(E�Y����ҡ|@A�y�N��=_K�V�9]�zsYRjߊ�
��zpg&8���3����n�	D] ��)2'��]Cd�䈎�b\�<u�D���e�>���WS��F�U[Irj�$�[A��Y%4G��Ԧ�	�Bj�G���HG1����0���/�Q ����vp�Gb��V\߱�� ��V� M;5D>�#�agQO��v�ڿ�4d؞�bQ�������k,�� ����ڱ2�r�ρ#*����AiL�]�ٺ"E�CO�O��
�n{�b�e��r�r�gg��CDLx��.��ɕ��4E�Tر����p�Lz�}�h�>�8�2�Cvnz9��f��t�8�����g�����eB!������Dn�sG}^$r���,K^Iv���4k��/��O8��`�%v�0��>�ȫ�A&�����+���1� d{���쯅�=}@��`?UU�jy�Z���2Ӻ1�8lK���k�S8�AW'Fy'"��O^��j$AI+��8��y?#�a
Y����Ґ3�ՉmNI��v ��&��"�';;�	��	��cf�����m�3@��8Gz�[�M�fH�>�O�������C����\��>ڍ����w��|�\f[WBf��j4��$r�&�����d\�u����ޥ@O�kDO�����r����lr� ����|�w'���k�l�?��$�����ΡL,��d�'��;#c���-Ng\T*W�gl�m�Mz3F����W���t�7'0*N�md�@T6�jC����aH�B��pmA�\"��K�9�3]m���8����P��Vt6��˖5K�G�x{w��7��H�c�CI]��
��n6z�?�XN��g�r�����������:�O�U���-$-1^�˲ۢ�f:N�*�πWV����iar$����xbA'k�o+��߶}{Jq��"f�&z���9�����_�!M������s3��[**����6e/q�&��)_��f��+������`�hY�N�t�AI��d�/�#2ǘ��P���Lp� ���~���,!a���P?��Yn�$?��A��J�9V0�;#m�\��>^:k��D� /LTG5UV�W��3�wl��sHrn�}'��̭����������G�'� B���P-G��Cjw�����yQE��D���F˾ ��r&cA^͏��F�y�ПЁ�,��d��;�Ϸ�gg��1�q���h��r�� �O~C>j^:����=p���d�/)�A�B�
���u[>�ۓC�P����>P"K��d0��AȜ~�b�i�)@�^����9�R�����IX�'���o`�[�J]):{cz�1�f=;�@*�ԙu���%f/e�C�۷�
���<�E���x�_�g����vJ�5� ��%�k���<�N�^�s�N,��&e���7�m9-��'�갲`�c�����FT���ɘ����~���.�$�SrI��Z}�K��L�%d@#֗#P���m�&� �T��N��n�IN��e��8�k�^�D]Nk����5�ӱK��{�é��$�c�����������kl�/�1x&��@�z;�d2��V�c+{욭�,�t�a���,̻Uе�:U���7OS1Y >좺�Pg�@[Qq�Be���8��� ^�����J�*��a�o�����}xp�����m�hB��ޣ(�S�̩O�8��:�y#��2�b��|֢�
�f��K�Nъ��@�8��?��2Z��4��K"؊6�-Q�9���	�C��DW)b"�ir}mf�,~��|{��O�{��:�L�7V��ΚH����[Oy��.zҳ�T��*�&��@17�Asy�GxЍ��ʧ`G2`E�\ٵ�l"S��f�
�_̳Y$���6���ۤ��wqh'M��y��fx���sdt�<Q&�ŉQ})牮(x6_r"���<x#�����O����d�a\����)�u��y�]�+���r�-�q�x���
��8����Mh��$O;k*�fM���%����x�KԻ�!������r5������R����|�q����"��o�Y1Ҩ�%�}m��Q�6ˬ�����`��Ì̓w3�������W�\@6�p�.��p������\oy ��֚�F�/s�{vFǛٛ�u�.���������Dg�@���Ҳ$��)��c�����A��ɳX�ݘª�M*/����'���E��FIq}��� �}����TiG����ᝃ͕`
#�������!D�{3+�K)@CF��'v2�n�`�7d�=w�CJ��~$�xUQ����'�:����X��Qg���!�]߭A����\���$�[H�8�Px�Ζ����\��b�]���cDV:��Y��AwKZ �t� ��+Ԩ�Z������<�X��.�єKN����l���G��w���t����"�b����[��d$DL��#r>O4��������1��,��3�̽M��!�--����ՍK��� �=�ȟpD���|��e� QX����
��J^]�$(�t�<T��;�m���e�>1�Im�j�8
�xi򽜻3<��n�c��M�Q��А��1 ��:!�?+(��N8�d���"m8^J������=����3J���',~<�5t���@�f,��*	fn���B��n$��\r���.�_R�u����bMK�V�I{�q�@JZ�.�j��6��F��rp%�BwJ���;c���yZ.b�G�?���5�=����-�e;��,�B��^��K$��0�2XXbUsj)e�͋�89�(�=0���I� z�_��] >.��K����_��Js�� ��YE����WB]؆�/��A7$A���3��4<v}v�~`I��>��E ��5�#�LZ�˥h]6w�α_��0�q��s�����?{���Ι�l|.ln�Y��|���z؅�I�f����J�5!'Κ�A)�>�gkG������Å4�6E�o�/�"��J�
A���u�>�B��	=1����K�X��lfn5i6��M��K9�D���W�%IZ�&��i�G�d[���)��bV��RKD�
��ySk��Q���hM��ڲQ��ބ<J�z�7�*���pSQ�&�&Q�Ѡ�P�����m� 
��XM?��;��#�)�S���=�|>z�W��^g�������[��j���+���ٱ1�eӷj�CI�v(�n�[x�f���*�J^���do�`ig ��K~Q����ýXX��(�S4K�#2W����D)�[MRtO�ci���5��{�.��@�6}dJ|H]������&�d����nt)o��r�+6
H�2�C���#$�Cw��G<���A^"�l��{دI�8�G���i�� �Jj��5�]I&^��;��+s�L�C�]�;�[��mA��A�=�V��P�}�8�9&�%s��fy��j�6
��Le"!C0s /z+�3����9����E��ӗu�)b,LK�g}*W�/���0�7���1�\��2�Z'�֋�ݰ���������P�2���0RԬ��}]V,����<K�lan�>ʖ���Lw���@6�H{��������i~��8��n���3x���������>���H!�:2���;Z�St">G�Մ8�<��x�k!&z,~�D��2\��r�tC��sSQ5�� �wP~j����q�,��ٺ����2��y�����e�+���S1C�Й챜���@�IQ�ߖ~t+2`<:搻�Q�������"�"3�z��al�+���D�[f�qo�1I$]�V��>O��3>���z���L���b�	I�!��1e~�c��R�����Բ�!��(D��SATv@�9�b��J��z�T��g�m���J����6�Dj����8H&m�mG�eHr��]��a��Il�Dd�L�]�r�TM�(��j�����#zJ�-�S���d��;�����t�^/.�!��f����s������i�z��췚�w;��>v!՛MR!ձѿGh�b��7Cb��9w���f��@�y�[4ڮ�C��(���J�3D�l���E=�N��B���JP�`e��vu�C���H���6��A0L�حkG�Ꭓ�/�RuB��a�Ӧ�����7�/���F^��Xb�9���\VQ訟z��&n- kN�V��-��`�#9 ��o�Ķ*<�H�j@k�jh6�4�#J���Q'u��Bn��|�{⡒���N���Ch�bP�^L����+���������+00}���ѐ��K�/�?ob^�FZM�f�i�
<���k���@3��
�7�N6v�8v�J��]��ק�°x� i�G�̂~;9�-<k��|��������A�9s����ɥF��8R�9��?k�4~5�^}a��:S�*W&�x�)lLڑUe�D���Þ��r�.^+y��m|(a�]���0�[�"$_�d�$@|:�g"mW��9%���:�i�wB�v���=A��Cͮ�L�R������۳�.\LG��-$	.����}�����\��r,į!��Z\�a_AD�X��Q	���2��pl�`oQ& 9wg��|ѣ@18��$��+���=K?Y����R�_HY*�H��7e�M�e�4^T~���0�v�.�F.�*�s�  �F�Y�l/_����2��|�{hrr:���\N|v¸�]M6+���Gv��T4�����x��'1k�# G7�h����h�>Δ8�������w�,�������dL[�
�H�o��)K|�M���m��^!?"t����X>����SD�'7�_'�-X�ӈ7�y˘:�}���y[�	�z��^��x�+>��0	�QY�'y}�%���9k�U�;���C
�@�%�?ն���'��iLY1Z�<����F��6_S�	^�<� ��d�Y��D��E�;�s^sJ��<�1�%g��L?����M*q�Ct��Tэ�ȇYkqN{q����_kzf�1�̴+~C�����������E[�� W��e'C�n4�}�i���:�͆�B�گ�X6���>4��0%��0l(Ih��0M�p�*)�Q�|$����Φ�OR���i�� ��>>� 0��CH���uϲ����ؠx�qV,��,D�*<1�Q<䮑l8�(	�9�8���cp�aͯ'G��Lg��Vy*u�]vH�pz�Xc��Γ��z����>��cO�x�s�ҵ�`��t�����������k�v)��)ͪhˑ�V��}���V��^�֕�dnv�!��;s{����1�B"�|fx�8���e�\�q���d�����|��Ua9A�5%�ؑ�=L���i���"]|��.8nf�)3�	�NG>�h8R����1���*"�9���vm��-�fiф\r��J��o{Z_��#7���#Y�1b�F��"���/�i(ob6-ٷݕh���z�b���Ȭ,���H���Q�%�R�zwjZ�DN	r�;M�H���^���J��X�C�'�bYNL�Y��M�TJ��ò�n�n���W>�I�9`64��L��{��Wk�[���ё���/d!����\��t���,(f{q���*�i�s�-AI[�?�eo�q�������"b_۲����e�60����]�h��l�d�Is:��brV�>�4}p%�a_�t�?I�Gf�π��{��*� =W�|�+�k�%k�-�J�#Rn����+>��0'�
�b�ko\R��iuͷ�ϲB�[N�f��r���`8�Kj�M2����Uu-���y �|����r��Ų$~�ί�t���8}p���
���¦x�@�>�:�ߚu��5��Y5��<�g Z-){�:����r~"�����x��sHJY�Ij^�I�U8C�b`��ȣ#km/G��i�̏QnA�A�h�W�����P�o��U���>e�J��VM+�G�d��Q�⇷��!4)����C�2*�`_-yi �U������9���7�G�h��F/��� P�@M��ψ���H�������7��d&i=֣x-~�	Hvl68	�\����kVTr���1
H��y�=エ�E�d]�Ԕ��;���bUɵ�ݞ�KEH�r`j�Z���+&(wȣ ��p�j��?��&��[���El��0\��~9
���8�Ap�����Ѡ���C���`�
��%��/����O�L�rΌ�_�f<!j[�QP6 	n�my�O�E(����{'�pCq�ך3���~��v}0�V�:Y�8
^\'�-��%��`�y�����;�*���Ǔ�}�����G_��(���t�K����C�E
T�ڙ\�͇vԺ��HFE�o�}xw&�H8��3sH�k0/e}�)Oۗ�Zy'��	j,v?�}Z��D��O::�K�p����p���b�n�ҜIk�_�	��K#�OO��6+��߀NuvR4?BG�A�4U����䄛xUP��`Œ�Q����D1��ߚ�wܘ�XUX�]��h�
E�#�'T|��c7�mP�&ݩ��N�n�1��^�+8���?�V��f�m-Sj���W�����Ϙ�a�Ds�~��^��;/���h ��w޸�c�æB���݆�К�o��C���tT���[Xl�R,�巊H�E���"��^��7�ם]�P�H�����w�k���}�.�b��p�*��;�q���s��ӟ�B�j����v`���|�p?�F=tJ�Mw�����0��Vb�"�?xM�'��#CȈڏ(-�:�
���pB<�cN8��y0��o�eq@p��n	���-��hd%fЊ�x�8����_3�+#��	n���UJ�%�/�$_�9�'5���5����y����n�T�2�C�.���Wy#��.{^�LT��"�ߘ�~����<��YK`V�0d�xK�!Qk�ؾV~,neU�׹�Q4ݷo�~�r(���	(eh�\a�as��l��V��V-x��
�7Q~֟H�~�4����&�B����+����̭|�z�fp���h�|�y`�1mJa�
7 ������-��[	�=>T`;?��ibp���Vn��y�[�1Z�y�.����i��P�@���	�菺[����CD���0�x���ζ���R>1�����7�1^�3j��,��j���b�����C�X�{-G]���ѓrO��ʔji���=���T2����ߘK��C�o��Q��WY�3�H����SP��Ho������!���Y\��t�U@2���4��Z�V��"��,o�`5�F�2�=|�j%4E��MK<U��6^����v�(�)�l�ApE��]�X��$UD�)(�5��v�Wㄠ����[�%�}`<�xb1�����"s�#��${<���������fk�h�Co$���G�&�׬̈́��{͕��;������\Q5��T�X�_x���M����E�� 0�z%ޝ��R ������A���jG1����/O~M�[^�v���;Ph�~W �������Ok/�l1W��N)A:�kj։�I���N�&���FOD��=�8aۧ�y��?.���ǈ��2|[Q�|�J� �����B�),�u���Y�	tؐ�]�iۆ�m3:蘊���h�!QHH�j�4Z `�����dԙ�1�t3C��nk�+DE�(�]�>����|Y��J�oN��tm�/���'+3K�W��')�f��L�0��M�;�����0��(�d}�%;M�1qR>A\`2�>�K��sq��:���|!4����ziY�@�3h��2�گJuXG�Zҿ�&�0F'��7�	�E�R��"n��:9�+�&I+/��s3Ȫ�����|X�����Ĉ��$J�MbX�+/:9E��{�ͼ¬B�NB�V-�S�I���k�D1���KEp"�]7�3�+*�B&�(��`��W��ÔG����~�,��]�����A��'���v0=!�Ae,���$���S��F�`�ix� �Q���#��h��le�,ԧ$"y�>9z�g��h7��J��W5�vO	A'P����B�-��
�t�}�?h@c����-*h�B�)h��&��?���+󀓂��ѫ��BЫD��:�b�-���\�=*�d�����i�J��2�󢷌�!p���U���qF'zP�%�!	�!ZM��I&R
t��z�8Ι��c�ف2���z�b1y+{��a;��-����٪���M��6�/{` q]3��X�	���.G���3"��!2�$5O��{�s��.���>��@��h�����3�˥���tՅ��Q��r��hT�*_�X��2��n����%��*Tf|݃&gO� ����4�JW��NԳG�Ղ�IJ��u`�v�6�r�r��f��"�s�O�"��?�d?n���� W�TCD����-Kë�W4��m	��v��sxuR��J`�o"�jU�/�]�n�!�
�D(��OT�__H�h8�|t�J5k�꣼��Z�CܽZ���v��]�z�d�q}ѡ�L�j<,Zœ��</��!��H �u�"|�!-�26��� �7y����!
��u�Y/\���<�;_p_U�Z����5���3�կS��C\����U7�����E�#�s+�֏	Ġ^�v���U���n++�n��� �ou���(���TKgl3HI�<T��J�\�DȢ���!�+ϰBﾵ��L���_l��� �P��WЏM�g,�MxY�1rz�K
TW��.�B޻��f@�*�{W��	X�S�eS�՚Y��z}�م�F�X1��?�F�cW��w+-�q�Vpyl�g��!�<�/��o?��.�n�"���x��Yd��>#9X*׉\V�j�=T�$V�X�T��W�:�����EŇ`W�!6�-��+�ꈌN�4�Z����ۗ�R!���_76��1�x������.�B$I+���_�}�3�my�I�>!$~x�h�@�,v^b�%�eK�2Y[�T�C*�K4�E�K�Um��f9��Q6���4Bz&9G6�f h��T��I1����8	�z��-��C��h��K�S��nf��Ph�t��ͮ���+Bi�V�Tq��rC�(����߬E����������b!��I:�Q�y�b��`\��R�{�������P拲 %��D��f�9�Q��U�����a�줶	��}&mQ��}9�������0x�~��N`��#���eU���.�c���:��f0�ĵB'��7f�} 174�Ka{��>��W1�h@'f�$�UV,����g�C�H8�B|<��4�%�i�}�G�����N�H�e�ؤM�A��j��u��$�7�2���}�n��j#�q*l�.� ����p��*/)EACM�P������8�R|�?�~��VP��Ŀ`ִǽ��c5ܧ��N5 �ȋqY=n��4�$��=J%�ܬ�yߙ0w�����=�1'-82tyq���}��*�T�I�	��!���S��q.�>�"E�۟�ɷc4A5�s`����<.O�,��<�[+ϸH��8(�,f.e ��$��lT�����%,x�4��n��Z,G�;N��|v♋�P��aWG�P5��R����uC����J�QD~������������=RӔ6��7�:P����yQ��_����P�x�:K�_Z%&���1�����л9q���8<��l���l�(�sѐ�ƽge�g����`3�]ʨ��_'�V'�|g��$y��w��d��➮��*\]J�9�5���G��J��	��ps� pyk�yU횇�_�@�Ss�bHd���<@���+�?�?b����^RÚ�\��x+ޕ���x���ˮ����kQe>CƘ�a��3W����� 7��pD���k����YUؑ��7��� ����/����4L�e�� q$�5ԏ�u�@��@�*�!M�l�|���e�^�ڒt�Ǽ&�5�,��mD���9��"����<��޲�0��W ��B��;V����sȖ'�ݽ�<Ϝz��vw#c���K�~Ύ|��'rB&,d����i)J��1�8M�G�`�dT�:�hKʴ��in��W���p�]O㳳&��og^ԭ�	l�U�$tw9�.�Iw�Ñ��$�kDLùe�f��R*D?Y=4P��\_�{��3D#�C��U1��[H�PE�i�t�HF���|]!�(}Im�]��u��a0�}p	m���;���M�0c5&=>�`z�>���y����Rs��Ӛ�3���"�Ϋ�M�jH�Ѣ��h����!�7ߋ15��c�Ć���o�b�m�'��(�WY�� �8�j�%>�O�/�* Rz�K��zc���ᷣR������x%i�����i����:�Z��k@ӎm44�=� �Bv�`�_�#���N�s�>�!���N�3�<l��2o���(��7N9�uM���3�ۅ����zT.�+�׋m#'����B�ԉ��ޞkƥ]!H���ؕhJ�ȉ�NjZF�z[:������vv|�(mk����u�F��y����L�O����j'�����i'3���s���=�ԯ0+<�,�a|8�֨y1�q��'t>�� ǖq�b�ֱR���f�|�F�s�Y�-��+�!�N��BA��sҮZ�r"��c�vtBaӝ���2�X�GةF9�!�ax��^�X�(_��f�-;��������\���$#@+��"����������ʥIL'̟�&�btm�b�'?f�;��t�8��-Ն���u��_V}�Z�gT�J5�|�Z�Qo�� ׌��6�3^'#jL^�H�1����jR���_���&ݱh������ �L��'��f�_�(���Ѩ��No� ��'Q_�[s�5UhZ6�s�F��Z��?��]�Nrs����1uE����*=���ml�~'n�A�a�*H�A�㌪Kt����71�b��a\�f��|�����m�q�R>aQ�O(�#>�+4I+��2���1 +z0~Mx8�MߎZc-�Pg�O����1x����@��8MqO�Mgv<.��j�-pHŎR��c1f���^��LQ�"��g)M��cv��K���4'emn m��FI��n+�n�h7&�o,W1�L9dy��Ǒp������d�q�6�iW�e���W�}�#6Nrȳ�~�[\���v����˔���3�s �X:ڽ|��1�ڤN�)�02�n�^E���Zh&��زQ����L'��׼�dF�r*��i��ᨯ���Pߋ����kl)@?Ch�w
��jm���%#F8���.�n��R�o/?�D��J�CdxeUY�<��d�m��	�sPX�b���%�BT��4�I�m�w�O�q�ƞ��B���y�����cm=�=��A�|��*@�<�Mő��W)϶��j���,�6>��ӏK�H�y�2|Z1��^/DK�.i�Q�1 �~��TD������A�O_&>�0�fIֳ��♎`Hr�YR��}(��A!���nb���+�"�ɤ�=�� �/5���4���ؠ��3�%5�]&����Y}:��s
v�2r��d3؀�����l?�(�����{Z�i+��vF�j�� +��_u�µ�3pW἟����CIE	f�e�5Pw�~���m]�,"�z�0������ҵ�/ڛ��Iq�@|���a�P(& /dV{Q�<P��T�6���P�w�]F�~��^��6�yC�K���[��:0E�,Mh�E�+�L�\@�l�qWRH�"U�bXۜ� ;&`p�Y���T  �ݍW6��6�&MV�ڧO��1v��m窀B�	����5,�E���؟��äXd"����4`�w)L<	�KC�]n��Ctv7�>u{��)�J?��i���䑭�=����x�n͓s]*��ߵ����ѿ�(7l���#}�yA\U�Ǳ� ZU���dP��!�YW�=�^ڛ�k_�����c��Ӥ�'X�ˉteUkCU���\�Y^��#صH���)Y��[�}aO�ZK@��}پs��q�����4+Ǥԯb*����$�>8��<�t`��6l�T�02YN߭�b���xB3��L�(٥B� ,ܛ�8w����8��Df����2��6�&!e
��"Z~�_��&*��җ��U�G2s��e�|��i8 �<j���<6�-:�u���X�5��(q
7Lg{t+d0������r�#���Q���-�*[z��
�%��ۣ���`iE�M�Dn��`=�
_ć����LO�6�I����?����?��9^z�4p���jLԋ�I4��;�~��h
=E�^��+�#e�	����U(a-[)��+*��F�����HD�~TO-��е��ތqd�n�N�(u�=J�DD=��N_Z���� ��Fڀss���M� ��+(٢�1�F�ֵ�TC.�e(�c9���0J��Az�$�ʔ8cpe�""'�6w:�|��fz�:ө	�����j9�Ok�Ƕ�8�� J�Z� {�z��d��R����a�����g`�`D-'��+�5wU���0s�x�����K+�|�z��D`�Er��� �]�d�T���?A���D��d�Ó~�(��o��{Z�^��+t�78l�(=��N��B��K�R�Dg��p[����/�`����~��pR��I��~H�M?�\��*����Ǟ�O�*�?����;����e���1��j
�G�"�a���������3[6�� p���`�{������d
�U��xX�O�r2���yL�A�Ɩ%�ps�`C�AC�d���Ffxk5hIj�t�c&������H�T9_w{�̿�V����XB8S�5-zC����	@���qܧ�ӏ`5cK��)����j�醗j���w\�UA�m����F+�~��I<܀�\��E��I8��I��Hp��VB�{`�($�(�,T��|R;ɰ�����ip5/Q�n9`'o�b�\#|5�&�8���j��e]�P���!���(���L=;�t�4��6��u����l" �oN�Y�B��F�'��P�r1�aw��(X9O�AG��^���'[�G�Zw�r�	���	Wa�V05����FƜP��_�c���w	|fW���Wo� :��n�<�� ��`{�3�ϰq�-n���)�c�"�ϧ/�����%��oi2�VF����	���j.�orq��rH!u7�ч�Q�f� ��b�3<Y3�h5�_� MX?��y� #��U��]��U��%̟���_��΂*!����B�~ �z 2>v���K�{#�Ő�����dTd��y�"����pv��	�>�x0x��{ �\m��v�����J���իw~Ȥ�7/�êԳ�2̻P^]�Ł����$�A�N��()'�N��%ߏ������S���ʮ�C7���*ɀ]�/R�©�k��~�5�F���2�Jp�A^&�2f�4���<";H�7�Ջ���3lq?�3Z�����x����1� ��]R�En�Lnt+-�<Qu_��tB�[-{.���bw)Xq��>
E~H�qY�pw-�
��à���lc�1�x&\fQ�.��_Q,�Q���І6��.Nz[dP�S���uʬ��h�έJS�*��Xa2��h�����)�m�]�;������[���  4N5r�!��72�_ !9>U�4�*^�F��H��
�_�$� P@Jٸo�2̀,���)�W�s��0��d,��טTT_�2�9���2�Yw̘���_���K�i��W�7��}?����fA����$oI��ݼ�ɍ�Ɉ������L���œ['//����V`h�T#$Vӂhh��QQO�̍�q �����u�����W�]B�h����l��*�C#y����޷�k-g��sF���\6/>C=:��r�8�'��l��UL��>�:HY���[(���[m��?��8Rq�Ϙ�WX
���>!�,ۿ�|�^�T�=�i����C��N��8������\$dP����
P�~�`��p�U�f��=��L�_��%{R���zP��
�?�xf��}�a��K*��1�+�Td/�:��y���C�z,CI�d_�>��.WU�/hG=���խR#Hn��Mכ���$� �s �pG�(���le��j�H�E�Ւ���EN���l�`4�|�v�n���o��v*�7v�`�e,ZSۂ	���j��i[�7�cՅ���^��@N�/�b��b��r�	�?d��Â�D��K8��*VN�U .`�x�d�d�8K+�3�"��9�b�	����K��u��v^ƕ��m�c��hqDO����%Yo,R��9r�	�0Y�ځ�
�#x�2�TŐe�ge[��^�`"�Z�W�	O�*ky��h��v��ŋ��bi��	7@wx@�^ ��;��?��uP�6�6�*����m�c0aTi����1�"܈���aR���J�"L���&�K�ە$��q�/�Fi��`р�{���(sO^ND���
5h9��R���c<iI�:��e���5�Z,��@iQ�~<�|����a6�ߖ�[�|A����eK��n�ڂ�N�O�c͟�hOŰ�������]PO�𼮚<x�wV��y�CƲ|�5�:G���X��|��	b�YU�z�+g	�;WJ̵�V��	[/�u��{.�^�H�'�0��AV���i
�}�d���RƥYn�=�Y$0?��0�_M6�k�;h;-V4�^�8f�����;9!� ��Ϋ���5dW��x���D�8��5J^�K��w���?om]/�M�	j6��� <ei~3�A����π�!�q1���$0Q�O۷Ʃ���28&�5ֿ���ޑ�����#���^K !��q4���x� )�X�����M�IxPֽ����B�	��R��}P^9��=au�/��|^�'��,���/�
8Ɋ�!�c�#�?1YV�*M~�/1�eJ��@�GFNeP�y������>
jƔ�$Z��i�pfG1�hL�W�H�wL����I z��ls���>�ޜ�1.�֙�^�!BTS�≀�d�=�[50Z@yp��N���� "��{�N_�_Q��5��(+��ݜ�Dx�`��Þ۞i��fm�;E���S#c���h%�ﺋ��}9�}��HMwB�����n�Sf��IfG֩��痑�4�?���E&��!�����椊�vG1���ʱ;\�T|������c��:�>�$��Q��__O�@�Z"���_a}�u�F1�6��3ܹW��%���uf�˔�K�����x�j�z���1:��uA2Y�㺺��2�ը��:�]��<{r�/�
����
q���0�%4ʎ
/��َy%l�"�䦽�t�G�l�%`�D �g�gd�Tm�+�������5s>�P;���&�ǁ��-+��G��z�*�$����-��^ψD�`'e��Qj��nǄ����I�?������P���"�MO��힌�VB���L5�
е]g~��R�[
�ר�

M�gq=>�����N�ӆ,T��H8:"{�a�ܢ�ɮ�w
=�0ئ����v%�?n{w���+�,t�	k����e �+�(�[}d�	��o�}(4x�j�B��w�R����i�L���U��~ |N<�S	��Y(*/�!����D|�&�DT�ĥ��H�Gǎ�8l=�6�Ov{Йsu���n�4]�V[u��J������$�|�U�r-��܈_�3���� ૻ-��=b&���E���Vr�S �m�%/M��W�Q�[LN�z'4/�?ӿ+�~?$�T��*��G\������Q��ԡ�: ��[-�������R��2��>�|V��{k�3k�JC�BH�>\����n`'�]n�VJ�V����@�+��f�=3���c^�2�vX櫱��u3��'�+&d5����&�1&��:3/�����Q��v�a;�~���_�ܢ��UEE�n����ȓa��z�!5`�f&�������+�Z)�X[^� 5/�Xѯ��Rٮ0>��#3�~��ob �`���U��g�p}��z�Ob$�F�kt�xCf�zsV�x���Ӕ#��QJ9�Ί�Mur��}�8�j($����9ma��� �!�#�D�03��NA�l/ĦH�Q�
�ΌlR�����LR]�Q$t�.�C��9��>�'� �|{C��7K�I���q�YИ�Tcq
|7��P����(~p2n���K+A+)F�'ϧ��*���ux����M��z���H[uA/[k����:������p$�aL�Sk�Ov�&/�=���'��y�7|��ܰ@'�Ud������� Ba"��覛j,,��bG�|I0M�[�۹}�\�9MQ��n6���#��Xn������
�R��bn�l�a��m�3&V��mZ<�|E�-E.��/�2|- ���d('�l�-�P�XE�{h23&͈�L
x*�ѧȲ�^���e�=.����hs�$�~�5~K����Ý�R�9玏ʎ�?)S��e�:��T�q��3��$(�;��F¥�u�;�.�o���4�e@N��~�1%���7چOZ鏄d�(Oj�ܤ�\�ʊ�W���/�-.kD�\�GH�ΟA�D�b#}fŎ������~zG䚘�$�4������|�>���VCc��G4K���h��-]Zխ�wLn�]Iq��0�*��5��:8��n7�K)\:�h����
�zϱm��X�Mt*@UgJ V��g�1�7d���q���x�BZZ�X&Z�w��&M�/�`U9Jf$S��(D"ס��Ш]�-!��M�o��MP0��5�E��]ڶeC��,��tn�
�7 �+���Cd��&�Y���7r����Έ�`�����[L�h_��S�x[��,�.�i����\��hEHWm�?�b������jF!Q���<�0b�E.�N��ˊ�M1�**q� �}t�@*�3���zKKÁq[!t�s ޛ�+���^"t���
%ь�'��~_[/�垷NT�e�ј'��C.*�>wSg�V}��Pǖ���!G��f��a�!Թ=Q!34�ɧ5�0�J� �L�õ��v�U�z4��C䖾\��#��s�B�.���'��q��� ��ȇ��g��d���	g�;�Dtϥ��a�����]"�pU���c��݀����#y���Q�	�Y�ITL�I����t�3"e��|�p_�@",�0ɁD}���4��<Iٲ��b��(�Vo�U)P��C�ט�i���T��R��D�G���u�}G\�3� ��\�Jr�p�E�����R�-���y;c�IN�'#��K�%��jN��+l�x��ZR9/�!L��ړS�D�E �#r���|�:D��
�����7ui���գr`@ �Al|���K�f?��k&��^��1�Y�ɘ�:��j,��0F�w
��Ve9Nx_�$��B䰙"�C �Ĥ�0��.$��DSr�K�֟���8�ۆԂ�1���b����i�M?� q���%_,);6�	��uk��8bl	�xB�'�q�,�o���t����g�\OZz��뺅x��Dz0�3�<�?u/���,�A���"��G�XY �{Ӯ���z��l;2D]OD�xo�F�������0���.:�J!)�%r
) ;U�f7[O�K����q��)��M�ψ�lHC.�X/��}�`[�s��.b�	Q�\�W�W)��/�V ��ϗn���s�H�.�q ��gh��9傛��'��3f����(
�ՠ	wk���Rv���|�5�o�>�9�&�-M'��'��o��$����or.I��|q��;:ʵMaQ�~Fq�����n	��=e�x�3ȢY�1M�،%�|��x��V!���uE~��y�j���<-y��v�y�OǚJ2���E;������(0x�d�+�3� <����4Zj�?���Ի.�6�V��}t�����U��m��O$7�2oC\Q:�j��)�<4�
!R%	|l�bC������΄�3q�Vm���2�s�6��p��):��<�Lq�|i��i��A1�.�b��(ѠEu�����i`��Rc��0m윩%�RX�8tiF8��v�`'�C�����F�9��JUcӡ�U�S��8��,9=�>X3x��EG_����ڞ5��mq%I��e�h�4��@d o5>��ٓ�b6�o�W��ٔ�v�t������؎����V�M:��\�l�6�׸����&C3H�Q|�'U�'�[>�f�2@O0�op���x�3K&dkh;w�=*��@�gU�H˭9��<���J
�Na�I���f�~?o��焼��M�}���!Ty��l�%w��Ф�&�}��Z��Fm�"G��I6��?Z�p ��CY����dl6$�`ȯ�r�:
J�R�˯�s?��{M�ܗ�= Al`+Yl�a���b��@jӸsx��Kc����ȕ9�� ��0S�n��BnE'_��K��EЌ��$Y}��W�.�Vؽ�A�$�łG8��ADe�N�� "3'"�|1b��ڗhʦ�!]�ɡ�b3�g��*���n렄��ҒyM���%%�H`�D�c2K���<@j�6����ٵ��������P���gI@DeW��&��Æ�u�3���W,tZtU��ϫ�M;}w�����镮|4u<X�IR@�Yj� 9�2�Ps3�nĚ"�����rm߂N�Ca=����s��:��Aǌ2���L���+efn�p�����;!~����*�89S8�-��T�#>1^a�a	J1O8���F.����n�Gj=�H���KR�\�����v#�+ɠ��yƪ�p�`L�2��G2t4��\���K�F&�凫CaX$�=��ů6p�%�-�U�*n�������of�E��k!��JQ?Qs)��g�z�0_��R%����.����7ޫ?��~�T��Gߊ�P~�/Ԉ���s9SONim��G�ho�C����h�K�� �W�݇�)�N���Q�ڣ��l}�笼	&ܙh0�i�w�&����XL��F$�} 	õ`z�'ZU��??f-�Ɛf����Z;N����v�u�2{y�����������L���Rz��Ab`8��R6�z�)��(x�:��7ޅ��9��M�b�,�w��~f�T��B���KE��øP�Qzp��{+�e�~5C/��8MC�� v	-DsUL�����ӭ �������=b�X�5��{v�7c)p�5\��ɟ�=-�x��{�B���i�|���Ҿǟ�EO�(a_R4Nl����a(�o���tl�(�I��d�<q�'EXܵ�8s(B�碖�i#Ȗ��nR��(��T����+��"9���v+�ᓿ���hy�L��B}���P�7�R�.^.�"�ӌ�Y���~le����,��;V.��&Wd?��x��JA���6cu�cf��\1��6v+��]�y����Y$�����`��9�������x�*�;�.27�����6����M��3<��V(�Z� �.U��_���g\3/ͫЛ���*)�^�EϷ�J�+d:���3�-�l^��!jgxM�����r "?��mBQcd��6��4�P#�с�vJ��������,Y�*DZ2����XϜsw���Bb�� `�[S����!��'n��)�k�|2�EB�P�m�� pa�KJϐsR꿺�+���f
�e��v����U�S��fyr;�:|��I���Æ�jV���^ѐ�����S-�x	<��v�*�$9:�U�M�T��0K�*�����WrC�"��^�L]i9:�� �� ]k�T��2��w��_�T��~��rD�^�7O�7��H9�\��*���N�B!�Q���Υ֨C=r����VkQ�v_����MB;�۔9up�^f�^�y��8�=v���&.�wH���}|�z|Tg�P��T&�ۤ����p�f_�.����-������,2��;�t��|̗�B���.�(=��l�,���:�ս��6���!C��U�鶪��O�ٓ1�b!�t�!{�ˍ�V��/Ô˪�q��MG��_b���#^�%3�wF��3z{ŉ��'� tY/�]qv���Qo�E���"�-��oZ�̾ۃ�����?d�!�R@Ҍ52Ԁ �֤���_�v	z+��o��C�τ��b�9ƹ���7�"���v��4�r7R��_ҭ^�܋�
�$$����ݖ"��Rdȶ��H.c_I�|]���wi�,������b�z<7�`"���f��у^�cq�N�0�v��"�O���^��)t�.�~S��W	_)�=J����QFo��!w��hVT��[����{v�g�i2#��2-�1�0>A�C�G� �̎��%��HP�U�Mu����0	-)�E�*e��ףQ����ē\����*�E!vg��ן�D+b-/�RW�������t�KLc#����³� ��"��T�&Z�J��sP���|g�?�z���^�#6�X#t�涀�#�:������=z'm���
�Fp�έz����=�� ���߾�F�+�똾5�Hæ����W��I:M�����֒�x�����ѳmM��� �)m͹Zb�5XM��}_�yذh�
�s�1$�)���&��2�Lj�"�~��b���b�������hx�*"`U�X�V`�0� ��5E!���%H�����!�}�Ԁg�a�%Iۏ��� �����i���x��0�YG�@�Vh���>�FDG+If��s*�ѭ�v͡4�J9����g�?���L�H]����@��N>�:-C���oٌ��s.X%,�7�(�?����fjU>MG�(:�Z����ͧ����%8��+d����3���35�"�3D��bK����4�,�����^��=&�-$� K�W���h湹o2>G����\�uj�[� x�.���]��24ͯrW��]���s�΃ϯ�T�	��Vگr���C	�^\Cf]#R>�8	�bp�6�Pမ����Amƽ����F��#�re��ɤ>�]:��t�m�2�3G�^���<���Fdɫ��u,��`X�%ϞːR[����SA.D�M�Rd)-?���.��.���'(䵭C���(�+&z��N��~rjbW~I�9��19�LQ�o��f|cQٲ��?���\&��Ob�wP�(s���]3y�q�뮍7�Y[[��\��&J���
J�gON	��RV��v*�FR�:{?<��Ε�uY�M�&[*zE:��%6�L/�.����
ȓFj1C׈��5X�7t���25l��~���ҹ]e��M��θ�%��(-�?��W\�����TP�Z^��*�l8������z�j�To,�3���^�%�v7R&�����r��`�K���V�c�T�!yX��!��)�P���,���1U��t��+~9��f)O����H��K�X��tY�;8�>�n�}U_  C���	1PLd<H2�4|��`A�cK�#�E9;b�-��t��yۮ.,�`���N�<R�� �	�(j<��ļ���eF4XJ�NN$�C��ɜHa�MU�w.��x;��O���Bt��O��9��  �{��\��8��/1ٵ#H�y�X���o7���� ��bV$�]-�|��K"�����L�_��.W�����7��XM쨖p��Ө�G���50��i���������^.�39KyR$�[}�^!S��=�T��6�j�:���ʈ
�ع��=�V��=��]���}~'��h�o��M)��
����HT
00U��m�I\�5���k�g��˝6��7��Q�uJ�ψG�omQ;hz[4�rf�Yߏ=�d��ٷ��0�$�Ø��rkaޓFR�>�u�}�A�)�DP���ݎt�m�m�]�y�,2�v���rI�6���DH��K�݈4y,�`��iZ�Hij�� ����iG�	ᮅ�S�%T~l]U�j���8��s R�p�������|�ҋ����ӂ@�´$8�U��@�.b��
1������n�-Q�Y�>�O�{��� ��(w�|j��w3�t3�;C�:>3�>
�;��j_��ʵ`�|:�9V(5H�-:�9��V�RT���vPc�N4�ndB��4T��8�y~�j���>p�X�`>r�ଐ.�:q!V�(�	��(�>ʄ�r(I�K��W8Q�)\H0ͨ�v-�઄���5�I�6�����:�隝��pi���A��;�I���m����T��������F�x����eh`�[~k(s`�* ���mE"�*�K2��sf|L�|�s�<�-�:�D�ki7Ԍ�-�?5��Ei�Dz'
��C!c�� �+�'��I�O�|Z�q�%9����x*�h�	0]�K��k���%�2��B�_8z��o�I�B3�+�P~�4#�B�r0PEk+�4M��&�|<Q����9���<��?���AZ�z0�>��#�����.���4���)�O5Q�n����t85�!��]�~��DQBg1u��?:�$�E��Ż��8
h�����K����\���x'�;��X�B���qx�+��@+�t�w�/��We��^YB	S�Uj��r~��T�6�g�];!�>`�]���`dB��J	��ǆ4��aZ�5xD ��oGV���5W��?�i�b%�ОP��a�*�k�#;Z-��h�@�K_"``�o�����9?K 2�j5���w�Z� �EvQH�rD��2���򾳒ޮ�.IyJ=H�9��Ū� �:�[��V��7�-ر
%��R%�������$�g���x%줁G���D����_�K�{x����޽be��H/҄i�zМA��\Ũ%Ơy����t����uc 6q�	ђ�D��
���P�v���ԗS+����,���W��-�Dӕ]v��g�a<a%��b�^.�c�m;���Cگ����U-�]�O�����d��q�W��^��g_t �#�tDN�fc�{V�/�.��jQ��R/�Hj�?S��"?V�펌�����R�>2+!�ԛ1��k7���=k�嶃��� ��l2:@�K:��}���)���I,��x�I�ky�m�"�w�xѧ�h��ƙT�#1�矏r'�^��o��o���t��V\��R_�M�=��7d0%^
:AJsPl� �y\���ϤU�kL`��sS�VZ�ge49<K!�Υ#3�m賀��#�(�lY���f�fp.���<����BN��3]-AIt�uc�gS��� L�ǃ���=��d"vr��\dwB��HѲ���!`�I߬o��>���r�[\�� 3����8��B(dR�B�_���9�����d�ɋų���3��p�,���W��8-�I�"�L$[���ׇj�?<�����|�&	Dxn]�'���I���삀ݓ�i��6�x{��%���^�il�2��B)�=�M���d?��� M"�N�e����ƥm�>���g�ͫ�ߓ7Z95�\��RNf-F������{j,�}����}H;�5�H�W�=W�mxިlf?Y��f�<���풬 .�ݩ��~ko��K�
���C�qz����͇�=a�c����^hh9R�����j�Zm͒�K&ˋ���#*Yhϣ�����9� �����d�B`> ��E�����ʀ�Qt���@�i`2�Ψ鐌�2����㢗T��yO��j�����rZ��5<T)8���X�L�#�馁c�z��QO�e�3K������tS��"s/��zLK5�蒻�"�� ��vt��n��^�Z&}ؗ�b�|��_��5b?�s ��x�Y�j ��P0�+vp�t�p_��Cr�P�!EV%�0��-(-���G6�~�_aԡ!ȧ�XUV��~:N`Z����mO�P���+n��`���FP@9���pgbQ��2R����h����~]hA6�!-��-sЎ�U,˞r��O�q3�,ħ��MG�(C8���9��ۘ=:�>��>���Ԗ��}�ML�*�W]�-�E=
��_�-Pu��y�ŶR����8ģޫJ�����4��a�?^h�X1-g;�0�0�(M����!��'��IO4�Z����"vƻg/�g�~ #��os����>�3�ur�r�Y�k6���� F�M/>�Ǩx֭m�ImB�y�2��Q�N%�W�7������wY��J��p��aa_c{�`V͑�b�9v�rΥ�;���@(#o~m���k���ZA���Z�OaRW���L�ݐ�8�	��X�&����RBv�=�xh��e�;+�HDSj����Í�S�6�6ٜ#��p�������%�P�שm����çY&%�W�Z�Y4Lp�UvP(��J|�e0m�Y�ᵺL���J��^���,"��^B�zrZhP��P겞���Mk�3��5P)M� �ˢ�݈�����b��i��?2�|�����ؐ	����#"e���v3��Bz���@x��� ��c�8�P3=y7Q���vS^��V��'�E�
����P��>f�5��������jU�v�{u�^H��DEF���O�H�g��M-��9�eapw�C�Z�zQ*p=IVF�=���1� �Cȑ���,4YuLP`�OcGco,��I��s����L�v��#���$0�(&u���x�7P@Q%97W�X�E���ֿ��h.Ȧ��;n5�hyw�⍒{>�K�RB&�9�kϹ�)e`�����!�|ʈ.��ݼ,�ir[=1�����Q?�ML{����5��T��L��k!ǯ!�m�kX�Q_t�<3[a̱I���!X^�#��S��t���v��)MxB��ģ��EY�;�Hd-���Q �&;� g�B���=�*�7�I��MOz���fr��a)�vG��!uU�<��$���?l�pd �� 2dz!	L@>{q�������yS[��m��iDk�k�[�T�K�L�^H�nᵧB�p�Ͱ��>tٓ�"n[$��h�7-ax��y3�Fw@y����=X�"��Q�K�lfv+���S�
ev/��k:kd��*Fm4Z{Ña�_@�s�:Ö9���Drord�� Q����<��k:�X�+���+&{�/�-��&�&1���>�)�pG�UM֍�d�+2G�<~ݐ5(9$��ȓY��.�/�w��:�x��Zb(�εKcp�������6�ǻ_�Ϳ����O�H��"�Z}�Z}���J!j��-����ȩ�_��z,<<�sU��79y���KYܞ�$��D�C�^�A't��9x*�4��c�O�����?���.dwHޤ���lT�%���f����T% ����RW�.�%Ƴ�yۻ9?X�
'�n�7\G#��ና�k�se����ڔ�#j�jI��X�"l�j5��r�����b�Zг�����@�qC7�֓�iM���N�z0�MNmkH�;�?�O-6P��/�D$��Hڮr
��#1��fNq%;MO���O����f|��ށ�[�&MÓ__���SQON�-�Y��SD\R�Y �ވ�T�Ov�u�#n
�L��$5%s�g v�7C�^|
��S�#+[!`�~]F1)}jS.~w[�y8 ��ꒊ�cĹ5
�_�(��)f�rw��{��H��^�O("���'g ��@�Jn��]A�'�|ki��P���S�S�%:�̹3np�������&e���5�a���	o���M�%V�Ȼ��l�\�_��+�_ߪi�Pe�ti�NTU� ���G�M�	�)Z�k�6!,oP�M7��7BY�����
e����58�������[��������,hq�:��c^/��Jƪm���	��μ(b;��4�9��]�y+0��kg��r��&������; 9ٸ��C���ϟ)E9r��2�Q��Ơ��sy"�z-a�.�]O~�_Ά��MnƉ�E�o�
;���lY���R��Ju,ԏ��J�T�Oa
��ƭ�ޒ�s�Aqf@Rҋ���f\[�$]���HWE"_ �?��6��x���z��è9����J}ޖr����\k�pg�/Yae���j�(T~�ִ����oeS�.~4�����{��!���/����ȧ^H�$�W@4�ci������A�=��w�q��|Wvw�M���L���ca/�&�@^Wʶ�'!��� ��+J?n�Zͷ��~��7qc���}�e(k	TD	��n��(����eAPT�~Z�D��g ��q�����iʢZ��On�릆��dk;%��-ms�m��g��|����U):�[x6�[�R/Q�}�`k�W�n3����A�W ���xpvx��X�Ֆ��W�?R���t��eG����dD�+_���J�-+�V�ݐH��_F�"S��e�̯���֤�uF�s|�C(|z�N�\t���e6-�9�4k]�_K97d��G��q����..�,�O�bwn�%"*`���}�xy�<�k}�D�Б�V�%���{#k0��&��ZM�m��FE���� A�|&&�| gb�����ei�?�NĲ�u���牧��c�Sl���/:���~}y��C�5;���y;�@�E\�vީ����pp�;ƕ_a7Df������Ρ�f�u4�dV:a k=�7���'�p���T�_��Saɭq��J��|S�O�A���2��M��f3��|����RE�L���{Tֺg��o��ȂW\r~��]�:�uw�M��M�ڔu4�7�J�V귴-5}��f	���ވ/�Ͱ#�G�'�d=���j�P���^�fM(/,�r5&�/� (9�AD��v��<�W��e[��;k��[6����$#�軯��[D���Y�-�45�o��E�Z�3�	�$��`����a5�����,b�h#x����8*DV��������d�p$/H�%�S2"�!�n�R��}�_���*��u9/0on3O�\�\���~�Q�"ˁ#�8��8�]���A+���ݴi>UJ�R6��ݸW��E��'R��I�j����E*�C��sm��u�Q(!@~�k�r�5�u��Ε���S�a��6�q<��E׎�FTȬҤ����)�.d�"�x�q�	���OqL�c
zZ\G#DS�K��D����ӂ���J\�
�OX�=�@Y���8���Qŧ�"��\喍�H1)���a�<V�݃Y,�`����q���������<�PȪ�g�A�4\�e[e] /�F ��e,�6�Le+�6��!{3��!�F����(��U)ߘ�8��<<�S�p��֮J�2�Y��84��p;�d�#��Î��j��c���9f#96��k��d�L��)R^�O!^��j'G�8Q�P��
�9�ҵ�)=�ģ�E��V$�����CF_�&�{m�i���a)%�|*�4��o	�)���� ϲ.��J��
�d]�>���e2m�*aQv{��ô�s��a�{�1v��P�$�\�Ū�x|�&�2�����D
��^�~��+r��eb� �-��,7]���o*7���Y��Nx��`b�ta��g:q�S�r�B�������H�vٳ��L���=!������Ѐ��1�ǨT�B���C���F�E}B}�N�B#����v��+�˝~�^��^�/+&��-}#��S�R�}��\�d��Բ#��:3�}�~�'�x���Q����,�Xѐ쎣�E�^��s���ڽ������tOfO(h,��=~�x�Y��X�
�X��+���,C�?w@J�fBuI������ ���9B{���ѻ㈛�Xv~�S�gXv砚�����`�X���+�o�z[��mr?�OB�@( �?@��)�����ap.Z7�Lr��uM�S�1f���ו�*��U�@���>S��EK0ؾ�^<��)W�����LN��mo)��m�����D�=u4�ĉU��B8#w.(D��e��h������[��D�'�~V�����){�!���6Ozx����2�k�|�J��_�b[�=��~���A�w�m�/9 xr�@P�UKS�Z��놬�AIM�����Z�i�L�Oz�n^��rCpI�V�8��q�R'UN��9��B���	�<���Ci#M�?C�DZ$u524PF�v�Aû�@�e�@#�A�:�DE5�~v3��w�-��:0�F��o�������q�9�*�ioV�𻠞�����'5ڂg��9���IK�}�f6�Pi�>���;�ZЗ��5HDnH�A��ruφd5��N�U3�Ÿ���?ͳ�.�}eӗ�:��[�:Vq��M�p��W�������f�J��N��/thj�!Ew.5�k��0�S�� m8]�C��!od^6Čf�	㱽��	� �>H���2?�gL:}�NYvA��l@'1eʰa��ǭ�%��SD��@/ �i��ǉ���ܳ7ٶ��v��t8���Vx	�݂Gw���eH���ͨH�T<Sh ��,>��>�@��y,=���R�"=Ƴ���^+Gl���:�U�fL �\�wI��C�	�x��g��*�w�A�*+֢a7m�{׀�'T�cy��?Jd��,�����<~�S�YpP�<S^|_yiCx���m^B�b�1q �^�+��e�qbB �Y�PP3A�Ol�t&R i�:Od�<`�r�n�jZ�><{3g	�B0vV�n=(0X�O�C͠�Gqd*+�8�xp���>x�C�o)��3�)���{���z\GN=���^x?"Ʈ�)�,�y���^eN����>�P���b����a�9�x ��[��3pm�䆸joƟ*!�"�L��g�tm��55#�H9V�u� �m��$�Y�_i�����_�h�2�bt�`�`3�������1���;��ж��#'JP?����mX���@B5�beI���%~�p��9�(�$RLh���Gk6r�;nS��ϲ��|1J�.��
��G�?�,��J��M4�\�7!��,]�_|��(R�E#{���=h��/�`�,dK}`Q��-?��P�>�C����f���,m�hus�|�JZ������NR��xB�S�p(��U�5`��\��&<� �H��|�m�GBV�~����9Xqljǈ�C>ɨ���O���N�ԓ@��^�T��z�s	�g��:ᾤt�)?H����Y�^���ǽ�J��:���f��D�U���Pc4Oϻ'���X/ʳ�A�Q�Hj4Y `�*��X`����8P��A�%1�?2ly�@�O��o,/�ytP�}u���\�&(��Ӯ�i��D8P��e�f��Z,�+�F��ϭ�C�v�T�m��m/'�C��Y0�0(���p�X�A����l*�-��B'*��|.[E��|����1��F�j�w8�r$3;�A��gp��;'NH\Cȷ۪~��dQl� �;�P���łb��W���i�\Gj�i�<pI��Rt�}�H� �s�7�b��xE��5�@1Z�P�I ���9tބ2��0����#.\u�@�6��A�vlb��~����`��y�̉#_[Sb�ߌ�ܕ+d �N�h��tw����uz�K��j�ufc>^��5C��<Z�gna٫��!O��C��~��B���(��p�LG^)u���~�L�ܩK�6��Pw�q�P��r8�rN*�:���X�q��#Iv�ՠ�����+����e�]d������/ٗ�í/,�M����"(�56s3�i/��L��rtD�&i{Y*
�`�&��.��z!Y��H��%pF*V��=t����](�d1ҜV?�<k�O��a�G��H��><-��a��u��ͪT5br�#�����bqTo��"����"�fs����5��uTs��d���h��G�5�z�?��u�V��TٻWDN�`��`G�yp�,?�����Z@`K��nF�)-�$V�6&e_��H�:��i�J�\
�\�B���GI��k$�c*s�S�O�><����*`�
F�������t+.��Ѭ��ވ5JKO����)��6�h=vDߟ�~T��}��jq�Ut�Ѐ�ԫ�@ŰOpV;E:�d����F��|^,,[��������@�ȒG4Yq�V-��p��iS��'�S�5��1�B��;�۝NcN�����O���Hh�d�E+�fW4Õ��,��m v�Ӣ4����q�A�t��qe-�D�[;��Ö�EF�HX5���-m�a�٫�μAP��Ry�tςcn�Y���Z���Y6N�p�������]�r�.be~�lk0���ȿ��M�zal��W�a0�oR�mƤ���х_�5U���kJ��UPJ�4�4�ϵ�Lg'�}�F���Ш��5Q{�0.mm�~�E��|��>�z}͖L�n��u��D�4j�]��g:$�ǅ��^]k!7y�g��&���L�=ą�<$GE�cu#�%�{����ҥ����tg�J&����o�u�]�Yx�,����LIA�s��,^t�zU�Y�>�0��I���\��x���I���a[SA�2��k���I㩋&tO""��m�7��ϓ��0Q@_zU,�8���R}��& T���4��a��W�D��aE�Il1{}.L�*ؒ�ϙRl��i%ģ�����R�u��
�m��B�x�i/�B��;��� ��L� ��@�p FT�Fua�����)�."�Cl�I�l=S}7�qĄ�(:X�;�Z�kD��¢�,>US���������#[e��Ӵ��j%ĂV������ ��6:��n�S�i��f٠ʤ�z��|V��n��5o��D�w1Ҟ�T&�U���՗ßH���5�5��V��<�ݥ���R�x#7�dGvQT�8������~�Ȥ�g�{��/ks���}N�z]A��ُ�G�7<�E��G������*�[pK�,�,�9����]L�E	c��@(ǆ���l@w�2�V�����&��\����p�yYY7�<ޔ�\uMB�X��)��hͣ`��zN��#\��og��jC�@��i��I>>��$��{5� ��Ў�y?���~D�V����z��K�wBv4�+R�q-L
�K���r���Ѿ�c.�w*�9��4�Q�'w�%�-?l%cv���t�GR��� ����X��>�SW�H�\�i{V��z���Џ|,䴙`����,��N��#${g~^�g��eB�W�����X;� ��C��-�SIt��R5-�ȩ!Z�L�;gz܏���ϸV���)���`��Yz�[�]��k�H��x��#�ؾU���α��}������+s2�gl0�r2�)˺3�ŵE���Wj7ڹ7 )䧠Z�E �����k<��X��+?u���>��� ND �=2JXSq��0�Z,2�6�q[4��E`�0�:v(�n~��	S�i�=�P����c���*Y�� =w��s�0�=is|�Vo�� *����H��Η��RTIP�{;-�F��2
��T�a��d��a�"�U��֟k�8���7]�Nܒ�YJ"�0Ƚ��@�&��+^������BrMϔb�y�>����>���拤�1==ע"�.U��LW�g���冩�����o���P���/�3Z���C%�0��4�	4
"�ig`ci5e���.u���,Cw3J�o��S4�bk��!7�⼷-�[��d6R�'B���±�Z���;n�k�:E�^M.*\�.20v�l���B���6pC �yZ�*�R?�Kf�!d�w#�#��|t�H^���RmԶ\ܑ��dlW�¿��h$i�\Uҿ���c���u8�AkR&9«,�ΐW#L-���KJ87h94q Ē�#O%)�]�Բ-@�g>�>�����K̵��b���"D3�>��դ�$#o��? X�B�&d��9�����_>*�cV��(�<�*�����9G���y7�oW��u�&�v��K����	m�!2c
&&�a��X���_��,�"X <�y-�^��Km��$a��f���l�Db���B?��J�"�ۢ��BP�G�@F����H3��$kآ%�]"�-ۛ �q������W���k��8�c��;��=��Dv���(�F�&4��Y�.�m=f�W�k�	^���`P���2¤��e��i>=�!s)���55ԆQ�*�0Y:�ߎuv��C3�!Z���-���#ɯq�Xb�+Z �9���,U�ǃ�&�%K�}�8r��l��S�#O������d���N�̂�� )�ƽ��SFafŲ�#sI�ݖ��]��{6:u�Q`&�pz��	P�G��_\QYZP耙=��c*18���T��|��pEx	-��ާ�����$&�
黥�e�=�u��A��&��G/���Q)��M���6h����l:7@�"Zd���L��@Bd[�~U��b�E#+ό�{3��x���n,iz�pwi)|����&j���BQ�����>��{�x��3�c�0���,i$�t�띄p��e�2EOVS�Z㉂pm�Xل�.����������K��CY^�ܥ���B���#��/L7(����}���k���{����@�O=FA�q�ظh=��<�<����V^��n�D=����K��s�(��j�����.q�B��\,�;.\a�O���;g�	��̂���f��\�[�Q���i�3�E�c���KI�g�4S�ލߥ5�2�Ɋ�T���?A�����v��w�(�L�G�G}f��
UJL��!.�ߨ$q�� }��F�v�1���ӈ��	z�-Y����u��&O��:bap
ă�R~?D�.R��\���=Q�j�W\�QQ���ű{ls��k�-��D�caw_��Lms44�x�{k�"cTU�jH��&�fZ�M��̝�n[×r�?��a�mCuىl�#h$���M�+�d;��܌:�Τ��X�Vurlb8m)0�*8Q�e�k��A�>��J ��+s����C>��w�bCYe�`�Y@�k����������FT �8��~�~q;Ӈ�SBH�-��|�C8j�|I��暋֎U�R>��t��.�>�C!� @��4]�Q#�c�B��Ps�X*�,$G�{�*��;��8���+������1N�� |���� b6�����l�
���S��8J�C���^�
�y����Ԗ���ޓ�}��ͳ�=�6�䌊�Dg8�`_��Ek4t�z����%=<IDݙ��y��t���O����wK�?��X@C�9.�Cs>�2�"�s��Ox�K@�2P�<C9��D%PA⃸+�n�ظ���Q�X��{g����^%�N:-h�!%��U˩XgX!G�UA��^�r0���7@#q3r�*����	$e	�5�-�c]���4�� ��/[�d�p�B[���ߝr��Ը�D�Ŕ?����T�r�����U�?y�!����%>�J��W���a��Q(��*�u��a����E�� �r9��<��:j�UP�A�U�%�=���!�%�?V�@sL/k0�E��l�.���O&L�_σ�]��A��
���22��	@ �ªG�C�f�b5�ؽd���N=���9NudS�
h�P��ɷ�	�Ii/��|Q��!�G-(�G-��~n-ɳ!��2�ԉu��J q�	X,��0\ �v4�Ɨ������6�r�C�Է2
��9����fzVd1�5�y��Gjh[����x���=���K�,���m	��r��v6n���g�8HA+�v<)I�󱥐EЩ��4>ܨ{tz�6�pضk���ʔ�X�di/������	^HFx���DI���rmy@a:��D�]���������3��
"G^*?�C�ŇA��������F�19;�Ue��%ے�|WU�y��(�d�l� rZ8έdh���1�'ըS�A��ɋMz�>U�¦.[�Px����8e�̯��@�@ɍ�������W�atx�;o˲��ʯ�X5O�h�����YŴ,��1��Gq,`~���q�O��F�߇��L�Y����p��Qb]WP��u���r�����s����+06�/Q&/N����	١cB _�y���߄^/���p �z�9cFi�@�<Be�'��Bk�&��\3P���S�~��H�8u�h�ܳw ���/�23���A�DP�b�43�ʍ�%/�ޡ�e�^3>�d�d�.���R���?!��I�ֈ�i�NN��UBR�NR/��=��C������d9|m�5v_@\��x&pA���k��­nE$zYt���}�24e��7Еݖ��
�=�b��o7��c�;<j�3�A�&��)1Aw8�Pk[��#&������;	Z~'�[�M?��z�}�6#z�r�
�1��9KU�����������Zw�(��'��!��J��#���!��*�Ck���� �}�,(&'*��vȻF����'����VFѸN�{O�����.�a���o)�i<i����N>u��~Ce�f�5��-��%�g�f�f�s�ã2��F��d���$�m�&�ok�A�B���K���
{D��Qn<*K8r��j0+�y�� S7X/�E�{#����a��ɟD\�S��a��P&
�>8%�;X>솁鍚m����[�8�����m渇8�
��Q0d>R4'!� �P�Q�#��3 P�7~yw�ߡ��G�n�e��@	::��g���mv� \�S�k�2M�i?w�Ǣ�̡�}��0�2heCN�^�����"ެ��w�*)@���@�& �w}4~��K�R�oV�9��@�~���r"�q�����?�u�"��!�?��U�H��4Cm�`��iR'�yY�PA����uJ� ���"�c������N��_;��V,C�H�a=\(�.���߷<��c�S2/�xkg	�b�O�����(��a�y���=�yC�%�r���[s�"ͺ�3(����s���?���gH�[:F�-J��&r/�:��B���ɭX�G�Y��*���Q�v"�>�W��8�Mh�Y��0A��	P�� ��\���꺅��Q��^F\��C�O�Z�#g�'�5Y�*r�I��.��-���K���rF	�6�ӿ�%���-�"�'�23Z�/i��!ΐ �$�.���UQFɝ~OIpk~r�$R���fGH��8"\�8�@���N����/�F���9!��������xת[�貢�W*�<Zy�ՆM��ս	�2O�&�����B����tc��Ç4��8��i� ^W���y(8��̚_����.��_R��E�%|�o��4�^]�!+���f�<خ �&�َ5xpk�W,�q�*D��6*o���qG�"�:�'�R�x�5�G�}��5l�@슛�ѢY��mk�OfK$K}|�0�)�G4�5~p������5�T�ʹU��l���
YcH��2n������	E��r�0ŉA+m���t��$Cq��"Q�;�^�B��;�aT�s�����x���
(��X���?ж���(��>%�r���}��R�������Eȇ���ǅI_Z�� �`|x��i%٥a���pJ�����&����L�.�������gL��G��?��z m�<��<�l���� �K?᬴��&W�L[t7�S�qM�*�aX�}��3IШε��c�����AL�+#awm)�Df����c�w�@v��4׊�楡þ�v���˩Go��_o68�����Ȣ�~�$������Zÿ�!��j��w'�dJ��u�.z�������L5J �5�]�r�����B��?1�qh�� Ŷ}S;�nDL����[
�Z%�G;f������d]��+��!��@�}�.�D��D�7n}��rWڸ��jX��z6�cA)�a�W)
<��&F�[V��S����s�/=?�֧M-@���M1�\���/Jv�=�V�wg��kв\���3vf�!<?�v��������{-p}%\+t�{HͩzZ�5?���Xq��)o6�I�-'��CP+��PLƁ���Gڏ^d*�3�=R)�0bj�]J4�WF�g���<�?iw}A湏�_Tn��_6�dGy���#��������i���G��7�|�K#wv���lN�^�n�[��[� ��v�)�[�[9�s��^�����)����Q8oұ�}����� �q��0��4���&FF[>g���������CV��O=(P���q ^�AR�[�T���O'[��pp<%@��3:�n:���q�ϖ��*�<�9���P9t��C�\�-�tg{?8m���o>�1x
�Z��(%�Dq����s"I:�tm�f��]���:yy	�2˺���<�Q�c�l��Z��GY��<@�vy��8Q��S���4}-�?�X��N���=�H��Dn�^�3~�$7�����Ҡv��0S�����BZ��f<l�Qlv�3dt�G%~Ϛ��ʣ<��#���O�iQ�~MW� Wۋ c�d�M	�cF��aG ��q|�9\٤�������� bُ���-�;�wq�����5��¨`x�J��K�~V��.LVF��_��VC��K�� �������.;0l��M�vtS�P(��$��延�I��J�
��=�S��d�N\�XH�Jp���P�Ӯ��0�C1�1�r�^èM�ð��\��ߐ�����wWd�F�_6>vz)������6Ü�9x�����m�֐���?e��DG��Fx�Ac�k��TY5%��wC���k���b�yv�]�u�Q�mWYR�T�J�]W��k�}�4�n	�iŤ��_�8^[�x��˭�/�D%�$�����&����ΞId��ZLN"R~睨�;�bp����1.�W)A'�[� ����_�wR�����>��!0F"���7�N��}�)�Q��퍻,�֫��E'm�u��*�}�@妋�e��
�ʖ�N���s���_\�n���~�΀Vmh4c=l�
x�%� ��#�uǆ�.����tLY�P?2T!�{59zH��,y'������
�"��|�!v���ߓ���Q����ߍ�E�Ķ�r�ma�&$6����L!r��+jf��R2��n��*��&���e�]�u�mJ��=B�@��ݨ�`�E֍0<����`�?�����1�+��%�CZ��/=���Y����6g�Ψ�����B���-2h9e�'����`]w���@���yM�0�-�u粨d�B�}��F��䎺��u�����-��͂��� e7[Io��};��TXm����Rr֍��O�Ƙu��-��Ϝ�9ݧ���!W�`�X�C�+�)��ga_��I%��KB����YT�Ze��ɤ�!�����;��(��/���K��̵���F����{֕��n��qEj�����?��R9�J����;���L=�`�����nͅe�{ĝ��Y1�,��!9�b��!�(�R8P�_~�w+)�s�)t&%�m9t���:ۃ�����𳸲�n��в\����r���`�W@=!u�H��L�6�O�n���P�ɯ��o9�. �rh� �:�o`��/%4x��c8��~�n�����N��ɶ��Y���,*�7��I�Y1��'�����t�Mj�Z:q���o|J�E�h��9.��Ŭ0�%�jM���t"o_'ӵ�� �6�j5$�}"��UM0`n:h�s�!�*�I�"Qһ��ϖ]*�dF���d>	pń.��9���
vڹj�R~��O��F���	^��snIUq0�O@�Ԟ�!�K=��F�jҰ��N>
u'�i�%�LV���a�l6h�:�LL��ZA?�H�Ԫ�v+�I��0�M�=�QH^}p�%\N���)xf{���%A]ϵݔ�� a���e���ۨ����ӗ�"Gp��B�O]'��t�g��"��E�afƢ���(��� �U�]�ި�3-[P�`s���ݫ'Kۧ����0�� ��I-=��ќ��o������OH�X-
��jfK��1���S=���Z(���'I��������Tcd���i�>6*wfg����)�w�W��).�9���;��u�������`Z��A�gn��},c <�����D�΀�-��"gav�QJ�����a�='TF��a1n��G�J���D1�=�K�!V��zks�c�U,�u�~ճcNP�uɩ�ʙ|�LۢX��9"=��g.O��zE��;�C�J:⻾H5w����=�a�m�����|�@=�Z"no�!s�r�|�x��zs�M��D���9�p�Cm�Y�9YX�cS�Ex�{�S�����߫;l{}Tƨ��щTn�U�P��t�7!|N����Hd��nL�cД��ޓ�a���xT-w���j�@�2 z�&ii����S8���yC��/�z8��h�I%��E��ʻ�:���)��Oݷ?�w��R�X���#��+���%�%8.��̘���{1ń��r1w��2awM�f�Z,����R���튻^�Z�������0l��t���_��&�7��b���̓����]���/5����ڧ�[�����Ǆ�[�Ţ��l���J��*�l��hW�)�� ��Xa�Mw-��O�NB�c�|M�[hD~���\r���~.H����<|��P�������}o�~�-�,�ua%*�h�_g_5�|�B�����.1���=J0Ī��ι�ɝ�\�NvNLQ��T�λ+��	�%�����L�}�A�X��\�]��ke���ɪ��V@���Yl(η��g>eM�͂C�!�s���a-�����vv�$�S ņ.C���Sb���������"��٫{y��?�'��L��+���B��}/{�qj�g�����ثb�H�I�げ��C�}�]���,t�*�`���X�3��-YN��ԛ��v�&�{���>�>�9� ��̹�ߣ��AtDm�b�0�9K�젦�z�1�T��y�*�V��˜]��n�i�"�� #���!�c�6�$��9I�aw��e�ƵD��\脯aR���� �FT��x`�'!@l\U��#�*�E��(p)�N���hѰU ���x�6�Z\5/� V}L�o�����q�÷���_��:Y����	�J(�����,/���%I�Q�KU�3��m�q���l|�A����&���ńu��a�1�_�6�d:�! ��'N�YBoNH�ǽ�24��mB�D[7-�J,�$)�
�4����3���S���ꊘ� ��-:�D�
͊��2��(��h4���M��c��H!�A�����MBʔ1.�is���}յ�O`�0�hL�ZU�׻�.$���?�1�%\I���V�~�r��K���TMJ_q� \�Z���F���7��p�~z��%�������H��͆� `���a6�2�"�P�
6u�&6.7l�"UU��[T3#2�9��E�}�>�wS�����b���!���|�K�
Jٺ]Ť"��_~A�!��~�<+Q���_��A�)Z���}��)�ڬ7�7�����6����12.�:���M�0t�I�?�!4�ebS�U�$;�ی׾~UCk֫�VV�щf^�G�D!l뤔	-��Yn�-�&Bxdʅ���>���41���Oa��&_���H;�/����p����`f+���'v��eF����#��r y�<TC����;���)���MOp1I�tx���������W�!R�T�D�[7Onn�6l���q���f� ���>�oL�Y��z^$	�_�~I�|�51\�r����4\�,�<Gz�X���k������t_��z��^�Wr�cgXt�y�i�S�8�Q��W��ִ7Y������_Ő,��Rm�~8V�7�E3�=��j7f6I�x\#N
���J�n���