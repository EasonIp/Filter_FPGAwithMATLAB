��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^���^�F�����b�}�<��S�����h\y�ӹ�+Y$�X5�%y�:�8�����;i�%G���oKp��5�3���=�l���ˊ΃�NA�|Gy�W�6;�E���f9<߄i�XTA�3vv�OW�x"��G���r�z�zʔ�t�A7��myOU�<U�2��qζ��'і��[�w�>\�����	�7�c78�o�N�𔃈�߅�P '[z3��j|��c|`���bo��O�%��ѶYɿO^�O�=-5X��4-; ���^ n2c�瞾����B��?|!�&y2�u|]�g,��|���*�)��}N�;+����'�'�p4�G������	����OR��Ɣ��?�^�<Y��~���`@ke	���+S .��a�5D���Pf[}M9"	�0��j��C�I��e�2v^a���s	��7+��w��[:b���٪�mϾ��H���3�{��H_q㝻�����Rݵ �̡*"��{i=�O���sS��U�^����V�)R'�)�v����Q� p��A���ӺQ�t�,��wR��j<Rl~(��.9")���\��Y�\"^̞��ǲa_>Q۔�<�v$ϣ���U�~kP{N�UZ�P��Ǯ�G�$A��_���]5~�*��b:��nNû�ɤ?���:�<ՠ��S!��Ɋ��&��V�!�Z�2AB�'��1=_y�y�M��4̘Wͼ�>V}���VԄ2w��T���r=恪��[��l�+���\�r�(� �`�p��@�)`���ܮ7g�3�5b���3�;��K�2�lPLνbg���Yi	%oSI�$�a�*<�gb�>k���m��_)-���A��r� ��V��W����#H�:'���ߑ8�T^�K%c~~x��g���l�m�a��x"������ץ�2) F�Ϥ܅@`,�����t�͑ö�w��W_<��bMH��J6+Ϥ�F�>�xx�A=��|b���A�O���brF�� ��@�O��!�"��u�|B�3xK���*.t��o!L���I�oV�~M�~����1�圆�8��7�"Y�ҷ���̞ͯ��a@�b�l��Q&����u��E�����7:2��d�օ�)�O+��;�x�:W"΀��y�I���a~�x�Ѓy�3�f�&[^/l��X�N�@�>��V0q�13��]�_���m��U=�)��� ,�ә<���C�4��'�1XĵeiW�d�4���yNP�����u-],�T���3ǭ8�t\N��t�;��c��VKdbL��Q���{����9W���k�׿e9fSM;�G��ھ��_'9����;%�nfgB�o��C��Bt�����(z�*�~oI�ޙ?N������V.��4��@��uq�9��%F����3��Xy
{X�؃)��J�k>�AϏ�9�$�X�7?-�Mb�z�?\���v��FUܖ�)�%��=b���y���,EJO��u WC����*�l,����:�i�p�ރΥ�TbA2B�ߖ��D/�U��sf/2�*������[h�z�n_n�R�ɺ�trT��׋U�fq��?w7w�ȑ����"�_��%I\��*�[B�2�\ؐ�9�����V�Nw2����WG�QJ��T����G�"U��mܻ���A���_��`�yޗ�'_�7H���qՏ�[��[��&��c��)ה�;	T6P.U�.�=�Hv>6{�y���BwD�~����ff�������(�(	l��h҂�Ư*2�A���V�aqa"E4�n׹�)I��_���@�=ϼ��s:>�M	ϿLg XIbfT�8g��HU�YP��M���E����
*��K&y�}�QEv�SA*Z��f��^p����q����p�eԚ^�qNȣ	�%��Ac��T�Bʃ+Iڵ�S ��
��1���:��YW��\�� @���,1����TŘ�]�"��n<�;P����{�+�����x��"I�OƇ��-�{W\��ez��]�����i�Ht ���G����z�]j%��)C9�v���v������Cۛ�X��0Q4Y�}��&
��-�=��F.Q1�idQ�
^��+��K�3(ׄ2�qDL$w���'-ڣ�GJ�4����~�ݏIk^w!�;Ɣ!��_́,�JR쐩vs�a`�W���q{�~���Y]Gے׮�Z�+�������ٲ��A�p$w�z�۔V�,� 5&�m���0��g/��BO�yom�i�ē�,?�a����(�Y�n�Z����C�BMG�|���N֕�Be����mã N�9�_���H�ۖUdu����'Zl;�@�����}�(�~�l���N�@ה�+D(+�F�U���ն�f1��V	dN7���Dv�� �!��S0(d��hF.�0�'�(��=��������rp�Z��i�c�0���'���qa�+��4��>0i���@^&�Po��g�Bv�K���4����c]�u�g/o�r];���fG��K��Ԁ�|�it6
C����Vn�(�j�k\��	(�#	ng+'ա��AP�7@y���mW��v�QN7m���=:��㒢�i�7t2����:'>|Ջ��q*�[���&��{|U��������6�G�قz�����������y��W��1��T����\ϱ W�5��eM��.���Ѿeu�^�.%P���L����4�k�3odR�1��@n���oє�z4��>�QM�Y�r��g`x5#�3�o:��L��9딍,(��S��}�*�t��C��nX�'�����}R��Hf�i��34��.(_�M��O�CdK�sv&�K
`L']��~TB� �D��)k>�֏x�N�����}7P~��=h�H������4���T������`� �Ƣ��pW�%L�����4 ^�j�^��ݩ
���K@�2���GO���	���Md�>�^�s;���]���>�`̝FrngH�����K]�h��H�&;�/)EN��Ðh�]�'�~lw0i������}��+����X�ᡀ�}F���Rd��`k��lF��CY�uc���	lX�r��r{�?��J�p����BCE�xp������E���$,���OC�����=�>��n��z�2�����Bq�%�w��Jl�w��/W��q�d��}������B�!!�fM�[��B&����݆�K/�4�t�@����+>]��"���3,I'k���*����^�wJ��I�3�-E/E��Ŋ�||U{lC�V�]�G-�p��^���/D�Y�ϗ��~4x;c-sz�q����R3��<ė�����[�^G�i��0����V�tp���0�E��N��3�oX��@��p��`��}L,qx����ߵ�%V���$ԍpݛ�I��uب���#�CN)�k8v�t:{�c'W�!Xz�
�������l�8�ج��X�T
 �6�,��i`��Br1����m��³�X;b}ހ����l+��u2�M��%߆6M�ט��q�C�����Zy�STUәJ�z⯽ď-��ߖ9�EW�s]�x`H[>�ZĖ^�*���Ą8��:))���+�:�@r^���������Q.S��Q�⨦�d;i`��Z�P�*cV0�g*�ٝ�Ṽ�016�;�~V���K*�V@����(�r��!�ӌ��a�L�U �NA
t����X�ؘ�U�j�2@B��+U������U�q�����~vjl�M	1?�'4�Z��r������)z�R���Bh��d1#�B�}j�҆nJ��T����&�C.=L�|�q_�����ۚ��դ��l���H��An�,�%�~���h3.)(+���T�;F���3�O��}0��.�QQPN�
ߊ�,Cz�0b���#j��a�Jx�uy�����t�%�T1/Ԥ��`��]j�\�c}��� �s��	�����(�[�x%˅5z�'�~ܘ�O�O��L��Ϡ�T��?��U��,<n��;Y�K��k���:?�,��~	%z���:L	��O���
��q)��ެOۙEAxpⱁ,U���,9q�}�uT	գ� ��f��������\QVk ���0t���w���r&t�eд9���5~eA����
�8�!Oᬤ�3�@(E���^�z�D�tZL�[�U���؆��2;?��q09A���rL�ƚ���Yԭ�����q+����w��^$����l�8c��H����N�S �Jx��2��I\:a�u�u)w ���$c�<K�cƓ^���W��q��D[�C�nQ���I��cO$-��W���D���B�V��t��*�C8mL�D���0��j_��=�Xw1Ņ6��8�"�j
W8 D�Y�!d�4M���UB�P���)��� �
����Gv��V�ߕ'���S�a����$- +wh=��5���	]�u廏V�F���3+��ȇ�?�o��'+@����w���P�6�����H�A!��u����W��́��$���Ob�АV��	 ,��&�OJ9�*1��q� �쫣§�(:�Po�Z�s�����[ب���/���J�&�B}�0V�r\�O�o5���<���I�Ĥ"+�:ADB�����@�H�.�JEOPò�>j���(�]B׆���G�'�q�e���p�����]*D���I�ѕ1��ޛ�"4@�7� bĻ×nӯ�p�?�ۙ�B/>tL�aR�5���U���8��Õ`/��;�%%�1ZaIi&���dѦ�l�h��}��.c,'��߽��¿�EG}q#噊 ��_��GÕ�s^ۯ"C-��X��ݍ�P2���x��ZTۃ��I1�KǗ�E�1҄mC�7�Jb���O�Q�9�^�e�Vѹ���Qҳy�{|�Wޓ귊����9�%PQp��TG_��7�C�2x?8�ܪƥ������� ��5��bԣ&є�x3#H�Ӗr��?sR&A�s�(��ͧ���c���Ba�LƊW���UX�j��&�/�Ȱ�ƒu��J��EABâL�Cc��$�!�eB������q0
K��Yׄ��2> �){�e���c����4���zx�ץ�Xv~�,���D��\�AH�(ĳ{v9�|?*e�y�o��(�����W�x{����i</��F�e������j�%�,ؐ����6�疃^d�<�'�ю��^����[ؿDx�m�G�V�=�}�*�O�cCb�uM7;���Bf�cP�LB�i폀��Ӳ34 ��	�{��Y��4�Y�J��\�2�S!��|C�u������%�}��ڀ��ӿ� ��gS8
�}��$�ժO5@8���Ǒ���m��F�656iA���[rD:X~�	�V��}�D�ET����4Ũ/�{��j������3�g����<  �y�_t�����-��?d��i҇��p �?����ސ:��z_��ѿ��#`��A�&&S�y�OGޠ�E�I�]��a͚��s��ؤ���d�/�}���=g����f�)�4Y�V6�h��[�w���(o�Wa*�1RLBg�'k�L_��`+٫Ɛ�r�c%�����慪*#���E�I��1X%-���]L��6��gv��@� ������S���>�5���ل�A�'�j;uIz�1;�3���X�R�y��I*�#�9�Ĺ\����7X�����SE�v���̅D�kf�c�-���:H�w�e?�@Pۻ���D����q�>:X�&5 !�ݷi��NFA9NOq~��z�82ѕ��{�>7��9�R���L�OS��ok-��͈��g]��\g����۱wĸN����N�QE@�rX��A�=^"��uzP3�kh9�zP�yU�m�i���m��l�����fW�uV=�p~1�9�7�c0�|�m������*����0������ơ�x� ��M�����?Z���h���]��ۼ'9qw�o��a|<�}wI%F,��Ÿq-	t݇k�kp����=7
�lpA��ʫ�Q�-'�pY��d?i�5���F��K��i)���<�c�r~1ӏ�b�u��v��\�ۨ���=�}oQ��H-?��5
�_y�}��uZ����<��T/��ɫ�l`f<�����s���������K�~;�HJR�{˺
�Z��u-��F5 �q�De��6Uy�J��Z ɓ�ﬥ	s��r<W��P�%��;�쿄�O�x|��Hۚ)ߤ�E��8�א>��K�~�����Bo|݊�iHBL��'��T���6�e�`�7?Lc2���C ��i��ׇ&��q��/��
��pþ=��@��"4��b2���;h`�U��a�U愉���7RɧwB-_�ɭ�Jo� �Fq=~���ˆ��5tk	��H.�m����t{Y���N��EN�x�d�����Ήy��څ_V
}�z�4 �n)�iV��Ըo�Pnh��Z�ɘ�zP�=T�f��+A��'m�7�#�E��q��`8����3����}ңC��-�2����=�{��$�&��5�amˋ��tX�U_�l�A{��b��>�YH�͑�m卣���p����נEZ��\��SC�zʮ��qX���K��}U�'�578�6|.&i)��0���)+ �#�ɩʊ�9����G4�S���'��M���y��N{���'�Z�b��{���T�0NE���Fg;1�7`�.7(-f���/d��8�g��6e`��4��J1}����Vt:��|�m`o��-/0���x�d�-��g`ɞ���R���V��E�˂������CS53����\):����Py��p��X		���$��K\����8�ο��N��ȥ}�1���c�y? :�S��Tj>�C�Pz:�� ����P7d��t���f���-�E�j�A7����{��]�y��`(�����ġ-{aKK<���5'�3X��<&�9(�Tؓl�=���g`F4Ҏo;�VF]����3���D�܅��m����3�Wr�h�&�<���A�hJ�C�,t"w}�	aN~Dlh Rnv7��)'��d��VۈW�5��@�R�Ug��H�y�f�b�G�yoY'}�ö�����Qۆ(l�zF��e���Sȭ���b��ZOo�W���?]�h=�v�i��C?��GYR�- �O\��dp�BrW����u��Ȩ�8�l��)��C�9ka�(�>�F�����Ѝ�/v����+֖��z�8�!���#8� ^�W_��P�������UD���O�~0o2���sc�\n��V%�r������[X�ɗ����Ю�TH��ȷ7�\�KSE���pd|S�<|���,����[�=���a��U�+ׯKv_��4;q���ᧂ\�B���n���Ņ���M}��3�;�^|h�h�Z|`j֣-����7K�����x���U�0��9<R2�������$k9�����{qX;��S���s?�K�%Y��d�5b�0�� Nᓘ�c���������ΐ��ſF���23��� V*u�q�{ݶ�DN�6P�XJJe��ꃰ���Kܸ�EM��>Ϸ�����M��ǅ��}��DT�8l@�ו"B��8	)�C�I��<v$�LƋ��R<�)��5�9�r�B[r�8���u����|/I/��^�Vw���5�yW�B(�޿��T�W�)�m���T�,�|�,1�A@K���x<��2�;Mr\�Q�n��T�73���?��=��3�p-0[T%19�F7`�MP^��f ��a��r$h��aVpLϮ�^�dM��U(E�m�E,��	5˨�m
cN�O�~q�pT������8�{���'t��
�LN�|K�ex���j����-�W8R0�S!�@~��f�����Cv
3��ON��ճ��3�j�˓�>�Uɓ�sY޺���2�QOŧ��A�6�.���rF�)M�R�5���epP�Ȃ���*�����1%�}���ڢx:��~��܃�a���I���Q�EW�U6bENH�o��dxS�k��#���f'e����o�8_���;�Jo^��c]5&]�����į��o�_?��u��F���@�8� ;R2��s0��MTB?zL���v�$���|�KF�)2��&�����R�jj�!�����x7���f�ɚ,�yI��~WOai��A����@���SY�$p����OhΈ�,���|�C|��D����oAJGc��u���H�Z�Y��#����_��#	b�˫���J90/Y�،�N�(��pe�TK5�=���3a����zPB� i�n��hx��	��������5#���zo�Vs�6E��.g|��c�p��W�Pz��	1�Ę��5]�������Ľ@����������E�L�G����78�s�� !�g�])�l8 �2MW��->������yK�R8�$�P�|��/";�O/��4����H��%�*����JB�k����VO496�c�R\�kz��w�\��U�Hh�b��h��ڎ�OH��B~iS��Ge<��Vڿ�~U}���w�<i9N�ߠL���(�v�M�R���i�ٲr�.K�k��A̰r�R��߂2����a
�#��s�LL�Ș�!��2�j�S�ue���Ь�m.�q�<0I&
c�幸�޺��e�Џ}�i�/���M#�9�g�'5P�S,��]n���U���kL��&g�6�.��6p^r{�a���b������8-os�6� "���ϸ�x��\���4�ɠ���V�[8�x��;58���b��O�M(9�f�,E���g!�|�x�wC�O:"}�\����XIT�yv8�)��t�Iq�e�^���E�<�L���V_�4p�g0V~K�1��.�O�W�\����%��^�S	�aI����t��Ӿ��S�� 1�&�PS/��˖����	r��UGbe��&-*��� ���旉��������h�����RJtyA������kR��WZH$Bರ(����4��>)p�.�&B*
��n�)����-A	gw5!'��d�*�i�q�PO�E�kx�Oc�9�ԋ

�^d^XÔ��ږ��[�NS��_)���l��D�B	��hXB�5��89����	���֌�}�
YAŽw��X2�?��)i���&��~�*9̐f��(�q��k����1g-�V/�Xr��T8�p��Z.i^rj�Go�Y�p���s �-ۏG׵3��?U��q>�����#|���f�-�`+֦��Y&���mUP�f�1�V��GdX�{�u��k)K�.K(#J�a��/�?win $G3��7-vDP@�t����C�@�ڀ��:Jq�p_���ͺ:�Ϛ�HJ��^P%�zt�t�De�Rxv%-�GMu�W���ɮ��回2_W�ld�N���1�
E�
�[_�fS�E�r�n���6
��e���qx�σ��o��!@�W6����[�|Q���0�q"���w:�vmVe'|��w�a��]�	�ک멨���vĉ��|0^�T�t�5�0j(���z�����*�@��u:_V�N�����p�L����X[X���ҠB)1>���"2 deM'K��H��80@���֓����|�^��=�,����d)'��ȭr�}|�2��f�-X)���;����۱��+�9�x����>��/�Y=�Gc^*��C0�������.o5�FPΐ���q��@U���M�M�D-�r�����z�b�V������[�H�9Ȭ�A�E�����Ӌ��+���c8rX,�ew{�Pz��^d��I_r���:�kvP�?Q���B0��� ��]WW�{+G�{��&j��;�*��}���|�$�^\��-JS��|���р9(�7�W`�eL�f�̵���M.2�4d��L�Ep���OB���)��j}$�zqI��e2�n��ǲ��D m�39���vy�B2,��B6��.#[���� /��"Ng���t�� U컉�ʚl�(r��@Ζ�}��}R��q�L����$	����Q�訤�Tk�5�C� ��!�pcs�̸��k72�������to�78�g0������gD�;�
�
��D�ܾ'��@��֦�qsI����N���bW�#r!O����t��^�=`BRF�k�߲b(���$���a��n~¨Xv�7�� H� -ۺv�eݡ^�
@�H��3f��`�������Q���k���J��ʷ���FG�&�+'��+j�&�Qg/���A���5n�=�V�i�5��'s�t�Q�b�z�V(�{�{��؊��3�md���8����c�Ya������3p����>KD��\��5D������o�4ͦ�Z�z��"�@z1�5�aR�*Ȩ���
�oƩh��>%q}wpE���q�݁wmQ[hN��3L��b�Db�Q� tp,&�U�!o�)�,�x�0�2l9�;@�)�-�m�>�|΍R�o�i,f�㔯B�Q@Vá'_�ɼf�!��*�AG4;�pb&�­������ި7y㧬���78Vᛊ�܉(�c:��G��� �8a���ň�d[�@�j��a7�=i �18R54��_6wYM%�N����d�F�k�<0���J��è9�T^�������z��S��[z�Z�φ	<�J�!A��J�\�<֘�4�2ģhi@�/Y�R`���z�����R�}k���]��5�B�{x 7��w|�jd�G4"~0rb>b��Yi {�9�����*�n�`�GB`��.݄�"#{�i��/��֚1J};а5}1� ��gu~�mA�E�i̽����w�iP>��>G�S���NY6���<v�f#��*?�"��=��m<�U�W,V�wZ���ҥ�T ��Wb�w��'���v�)�w��p�	�S�A�����Qw��
�O�d���V_ ��Tw_&^Ʀ�#R7U����m��.a�S���W������6 �1&;�O�O�]�wM�	�w[e w�dS�����k����4��\��x�����5�qh�gh_�&C�T����h�[��]i-�<�H�ŭ;�D�޻�u3݈��-�䢾�i��T�=�a���ܰ���av�uq-J2o\��"�(��������E����E3��4�̘��ם5��1	XjN`����hr�8PwS�8jC�	�l1�9�s����"�jm�d�s��+%s���b�����no��Ғgʞ�p�˷p����ϐ�z/Y�϶jFtȘ��׫�Q�޴'�@I�^�Xi~�0�=�}��h�j�Nx���	�gd��_���y�M��K��׌r���	�����;<jړw-��	���Q��Z�S�	b���H9x��s���͂�>S����BO=��;F_Qcn�q��!K2m�y&�w��΀g&��P=�q���A�H�1nj�9��M����(�땚���u��LJR;���&����J?5��1�sH6&/}b�[(��H�}�H���M���<�gP#4��+n8?i��}⢸�ㄥ��-[�8E�q�(C��<���!j'+N�KogR_q������h�����J�rF���9)&E��V"?��6A&�.�����	$��1�R���l�.���O��e��c�\g��k���OkB��]����4n=/sܳd]��"4�it��-̬+G�$kf�|lXR4y�f���\�r~{�h?f���>D~9�Kjnc����ݥ��i!�u���|�K����)ѻ��P-��q���+�.���ɓ�'������0��J���;fki~Pz˛��]=A���S�ks7���l��.��������n�q��tQΔ4�� J{����L��q޼z
�!D&zl�N9���{]��:*{�sC0s�f���#\�6{���uX�][>�;��[ ��[�v4\�ag���f�'����S�Ө� ��������Fz^��R ��^�����F7r#�_
�v�'��XM���T���6��\���ZCvb��t
ʳ��bJ%�,�Ց�����
:���x�8ۮ�F�3 \�zr�N
҄�C�w��o �ߟ������v*z@2��*�������U`��q<;9u��w��C�nl��t����?%�:����#rә٘�������1͘��C�p��)���� �f{��p��0E�1���A)5ĳ�h�ї��J1i����҅�5z��w�W��FeGȬ�cwlf�y���X/�P��:r��"4�D1�;.ڷ���K�_-<��nX��ozP��J�ŇxЮ�2�(U�s���xY���;��0y�2' ���nz��Dc-���?�̄����^5�*d)�ެ&��`��=�.7kr&��JTrhե�8t�\@�O1�4 �׆�Rn�S�@z�wm���M�o����1���O��zm��I:��t�_���Z}��v�Gʞ�P��T�V ��o�Y�N.Y�'e%�Iv��Z�y!p,����w��Թ*s$�aDH�;�3�,���� ~d�l�����rˊ����to�0iW�m����mgL@ c��nN;l	�Jٓ̓�~c�8��"��MKoۗꯄz<�Z���3<A�,D��~R�Zz�sG[5�7�S���Z^��$1�V~E�� ��]�2,�ªyS��Iaae�L�Ԑ�gd���a#,�B���Q
�'��4���'[;>^�G�r�sld���10��@��p&��Xވ4�2��V����������<P�����V�$��>/��q@)*K���[�t�}��(�\�|U��S�qfgk�St��|�=�
ݡ�a�j+5Q�[4&�m~�I�I��4�ȅ��Gva�6�=2�����Rp�x�fYG#X�{�qM$��/�� Y׵�*R��0	�u~!ӻU���UX�$Bd��Nyc����%Kd�W��t�� [Z�N�5�@%R��C4:n'�z�C[�ck5|TC�'7­Շy˴`�X���"�݋���5��U�>��Z��e5賈L���&�EA>�z���*̷���2(]qZ�Q�,(b����L��Zc�d�v�\��xj��5�=r�Ε���S6��\y>t�/F'���x�,F��-��u2���6I�mGNC���G����f/Xk)ܺ>>���7�7W�*���#��J,He��2Ž��t�(��X_�[��W�K�4���a�ob�oo�fB�����������~�:L�w �z��l(����T�q��j�V���7<5��~,�'�]�=�XǠu�p),�ƹ��Z�Wyu1�'��)�Qg��������JV�]�a�
�Ⴥ�K�0�BM-��$֛��\Ƕ���"���H��ИM����BB ַ_lAh$+��؂�E�(�r��p%��;���ʬj�N����E��q:�������un8۾��g�AC���zXO.e��_l���"Ӵ�`s��x+2qxƝ��=b��/j��U���	ae$��\���{���u2*�u���r����U
2�^�6iSB�@ϬU@��r%t��H��aPud�k%-8���1#�	���*V��/sO����w-��^ma��/R�1q�L��R�(���C����w�QTX����M�%�~�h4����r�I*f8����.�ژ.\���Wh�t��i\jʨb��3�E�}V@���.�x��f^�wP
��8�Z�BP~���/�S��H曉,�J�H]�P���0m���{��F�O�� D�̬F�
�ig�諨9OXD*F�����۵v~ ��2av�V[�'E��Ӈ]+]=�ϫv�vw�VEމ3����q��H	�/~W۰��|x�w�x��C�Ѻ���q��O�Or��������]�i�f郡��k�v[�I���	�˖�+�bP��d�t4���$tѕ�ґ��7�i��]k=e!V�'t ����3M^e.�]��~�R6�Q�u�-��R�'��9��c``���N�q��f؂U3��L��
��j������n�!<hԖ�O��\�a��ݖ��f2�Kl�bE��p�`I��:�9�b~ֻK��z˷�&O>���}�μ�T�g2 <$��$���IS��s�.ŨWEۇ�J���p4��t9��Xe�)8��}���hȕ+�B��&�4;���,�c1������B3�I�����f�����!%1M�?�h����>q�&,iE�r�����g����v�H;���M��&.�@j�k=����@+�lhYT ��dt�+��c���uݯ��"�^Xh�L�؎�ϰV�:�ٜ�y"�i)M0f�g������#/g��޺\zg�T�w�ҧhh�U]���I2�1��s��;�Y!ȧ�U���6?�i4_��́�����������]�||�P��z����|�n�f1j	b�r(4Jѯށ[DZ�)Uf;�z���
�8r�ڋOe�8{q�8��L���9C��!�HAӴ�S�:Fr2|X�Xpx���xv��6	��vS�v�8�j����-�-nF��-懒��g�Y�,��K�P�R��Qط�U��y�l��U���K�IN�E�"�ѯ��*��އ���x�?�	��JȊ���Lz۳���FL��{�ng,�`�	�HS������t���X�FK�'?I`�A��ʞŚkL�cc",B�<��_q�1�Z��^��zMͼL�c�z��kA
f���$�I�K0
ExQ���#�A�r�ȏ�dp�=}�_a�|�
<x�s2�w<2�F�@l��Bw	6�h�ڗ�n�R@��]�n���W�G[�Ԩ	�<Q��ܬ�����EFHN�N�>uK-��6�۵��Һ@��J��EuB0�-�k�2ug3��1$y��/��������K�����m�eq�	D���us�!	���ƮSe�ؠ+��<S�z)�4%��2"+Ú�R����Dk��]��E��Ѵ�\4�4>�͠��}"�c�X�P�BVR��Q9KV�6�9�c�O:���W��C�����@d����BB��"�P�XK��a �5UE�������c!Hj�J�"}���qM�S}b��e�ә�Yp�'�thGU=Kk\O�����C��N��E�Zz�� F�Ь�J�ցƂ�#��ա���S�wP2�a���\���7=�k�����>��,dWn��[#Yz�񷶩���D�(�B�&bZ�"M@��t�ó�[B�؍�0{��]=���Ԋ����$�ц/aҡ�������Z^�G�^�G�v*y1�q��^�-�H����'��`���zkNV�:��A�����]����`�Fr���|�]}�Q�;�~2�S�F
1%2`kI�Ш�HD�U<r����55�j��(�� Xke�w}j�sz~���S>�M1� ��RW7����3p�W���m�$Ѯ��8�kL�;1����QƳv%ȡ=��=�UU�<�g]�{��>�h^L����l��fXbgU�����:��:)�&ǐ	���K>��Y���z6<�/놧�����)*jF�����M��T+~�4̀;�pP����"m��-U��C���H�MW��rIC�_���kjKD�ȴUV//�P�.�}ۣ�F�7��c�a봇"[����ֺ'��-�\_�=���ゲ���Hd�;�k���+WKs�^��9ѱ����0�o�o���%ø�����m����pA��{��Mb�1I�*[��fnG��|���h�����&o�j���c0h�}�/("5��J^bOg��˝܂MI�e��/��K{�=��ZP5���EQi���A�+I��/$4��'���~ʦ9�UH��݂�j��T2m���4�p��(˽r��H%ǎl��@�6�1��)�V��� �g���D'o���k��O
B��P�<;N�`���{V������^�f!E.�5zo�Ag��A��{��[�==Ce.۱���;.� U<��8�Z��Bv�t�����W��p1*��1F��V_O� ��9g�ʗ�p����2	Ӯ8�h��#.����	{�th��,��,,� ��dT�W:�� ���l)m9�Q�T�û1�Gf溊-m��㉝��#ț�,O_�r��,A���
ɍn]Pup�|�&I�;=�_��e���`��&\�M0�U�!"V�����R�ac�9V
�D~��D��{�5�Ҵ�;�/J+���䙳4e�yk�-��^�]vuj��d�w�	v���Ӻ�+�/�Ϯ�ĪX.��iq\����D�x��?ո�Y��YI��*Fx���q�Cp����`@�.���+���ݝ���7[����3�KC���G�a�Iӯqkp�g�|��[�߸�1�ME�V�i�i���3�c�<�8�kG?�Ka�޻u�����D��Zs�SF��ۅ�����+�G�!�9��W�k��"���T�l��n}�mx��K�V��uF��~.�g_7/z!�B��t���z�)�)�Z��1�W�y�3w�G9�d�~�
&vYϡ����N�r^<ģ��h�1�J�RW�'�v�7���<��f�>p�Z�N�iW�hԵ�K���c�I�_FnU`ŝg�J����Zk�+a.~M�J��R��� ��"�������k���Ŝ��Є�3V7�����]�ۊ�QgZ9d���5�.����j�n���\�ʀ��L�K��_���L�4_	ވ��V�F�g�3���,vo,Ĕ��3��H=6��O5�r���Z����rZ05���qu���q�nMd��$�x��|]��Z�Ь�>OZ��{�,B��F��dj�����4Ɔ�Ԉ�}�bp�#Mj5�}�R�6\�����,Q3I��#�k�us��i@¬��FR*Od�y�����Z�͝{'wzT�hL;6l��'�	�-0 �ɺ�=��R�R(ǔr~�4��"؆.	��M,�1�Cv/�N��Ɍ���w��Ӑ9������ ����N.�G7�9�ZTdŚv��[��Q��8�?�^܀�`\૊	��'�L�{qa�)��G�B�P���Β���ʨ��i�.��i���4�(��G�� �E��C��z�����Tu���G�W�W߈E��Db�JT��v8��}nQ��P�/{�A���U�@��|��M�?�6Z�3�����$pɱk�CZHeh���q�A���rRQП	�B~�����3R�f<�!�j�0�?J�N;9b8,�י�f����+{U���H��A��B�3*K�U��!�c���՘��ٽ�c���F
�v����+l*��|Ό$m(��Ր5 ���̰�7�ֳ�c|g�s5��8`^���@B����y�g	v�6#�+-�SUN��8=��X��q�mY~�D�-�E���B�=J�Ǹ����Q)^�b����H'Gd�
Y�lԍU��9k08��)q�h����9�JMs���o���[�s�}I�C�{C������rQ���ak1�{�k�ヘ�S�
���\Bld/*�zqx��x��1��MQ�l�9�g�|Ih��VC�qאD���мƐ��*y�y���3�J�X�����븱���s�.�3?�>ٹt�?mگU�B�H��K�~�9�p��.���A���Ջj���㝼jD!\Uc�@��X�vK8�AIp�����\H5��3��f�VPY��[�`e0{$u�{�ugh�P����'���.p�[���l�'���XAY	����� �
���\�,��0l��%A�{A
���"��?�J�y�b���ggdl�V��yU^ͫ�cC�$S��z�{��3��{�<��J�.��{$?@`ؕVn�e�PO)���v����B����d<���C��]c�GV9��֨H�""��A��[M��|V/����Y8.t� ���~�M{�D���	*��P��=� ��M�rQ���cn�-����" c�0ۘeQ���qei`>������#���O%w4������c��
�q���J�ͷK���m�l�Z��>����0�q��I_y�Tv���2j"�H���z���ƪ��S|0��9�uk���B
�%?���2!݁��獕iێ'��DC;ݾ��3�q9د���I�����C����(��0?0QS��[8sVj>'q|�b��5�"ޱ^bHy���F0�C^���@/�S ���I��@��l�Ca�m|XgU�(�kj�ata�u.U��܇��H�U35�|�|��$�1��8���#�b�}�3�0��Y���ڱ݅cj��v,θJ��ǜ�
p=U�`�6�M/A(���z~���4�w�K�˧w^��s��&	��Ň�1E���Ζ�/��
=4���G�.���'+(O�����1:�c׉q��b��m����1���$q�p�q=='�5`���d`��2��d��_Q��eڨ���f��_pJ�R���폇i�8U*�ى�ta��7���e��&'\	���R[��JlA�jy������RG"�m���:wF�p%O�kb�W�J�������-_ˮb&56@�_�q:3=��CN!�t�/!l��!w~Sc a͓��X�%}�>0������ٿ��4/Ƭ�DE��7 �}�����f.8�)f�\��
���lR����~<��q% -#xÍ���a�������Z���SC)@N�D�
�-}��<J�z� ���n���Uf!��oiVt^8�\��r�A�t
,O�X��<�z�+ѻ���W�%��z���̂��s�[�)#chk�����͆j�5��v�p��h	ЫC���-��g73�{���췟2��la1J�1�+O�Z�,����z5�s�N��Ǘ6Äx{���l~51� ]b���nւQ%g��A̒��t(�"�z�
Ǒ�B8�b$���&���+�T�/
�Pha&������\e���ӽn�M��K�M�6anaLOɸǩ�*~x��~���F��k����|�����i�;�yy�;FrLv{�������������"��P~����g��Ld�^��Eg��`S&�:�l�r�9c1�\���ܦ�pu��Q�b��$�xA�5c'�p��'�	J5�?�����3�M��<�.	�x��w&�X�S��BCS�#@^��K
����t��L49I0��[4I|SO���Ϊ!Y�5^��y�Չ����
(B���
bb���m�g���ۗ�>��?5��%q�?L�ׄ`M�;������g;���*�\��Th�ϖ+�]È��nb�3��$���w%>T��.Q.ʹ�.%n wU_����Z���i���L2�
�iuI9�QBw��#I_�+�Pzy}�v�Z��Y�M�;�>��Dڞ�40����%K@�r��t�Ѝ?` �'13����l��4 [�>�1iY�Sx�:0@���9���q��SВ��$�(�G��'h��$��EXn\gp�VJ��p=h>,�i
�0q�i]�	xՖ���g�&���H2�|����"��U���ɸG�=?M���#���z?��UQۏS�/����^�B�Z�c��I��d���Ħ6��p�t'-o% ���.9��0��̃��ݒt�̗)��c6M�9V�x��u&-BB(�<WV�n5�S��u�//ﴓ�Ѕ�� ��aa�ӎ�^�����?5�z %�'(6G8)g����zP�)��7ª\������.��(�tN i��!��Q��k�{M5ݕZs�+"P*s����ʪZ�HL�ag�=��V̷R��A����E{:P?&�X����$@'���5����_;E��7g`�g��C�k�_`f���V�}��v�6T�u �q��{OCCJ#����G�$Sj��=��c����pBU�|��B���qH�q�F�R�z<q�q���jaa%����
���a���1#dOTo�aÌ�_� 	��5Հ�%�?����ɂh�E�Jg^F�醀y�]�8���ozF�f;�ˠ�I/3"E�T8��8�Z&[b�֕̢��V96�����[.���(	KFC� `"J;O_��� E���%m��(�q0�H;�\���&4Y�i��p�)���r��#�c��V��x�;�
��M��$ſ04�:Ո[CLa����/��Ж߅t6���m�Z�I=�v�6�h�n�e5�N��E@�°����i�<_��ڿ��+����r�7|4�[��0>m�
��x��MJ�4�E07!$�ml�08�"��akm�eU!*=0O2���6��`�ނ��~�I͙�t?�/�C�.rП��*��kIo����w?�H�9(����U��M�����d�E�{JP�܉����O��y i��'�K��oG;	�G�2[��/#� ��A`vF!�������T�e��*#�����@Vxp�NU:G���+g.8
C]0fQ\T��[U8�N@�W,�V�Rsg�o�~1����퐣O��m��)�?�����2�� c!������21*�B��#0��l��e"��� �W:*��� /�)C��q1�v��у�?���f�*J{���gW����3�'�f4��%h�[{�i��	w���]]~�p65��̽�т	��`pQ�ZИf�6��1��~�m�',��=wj�E�m��5vD:��Ԡ�!d�*A�:͜����s�q����L*B@�[��ve�{^"��A� gg�*B!z����Kğ�O4X/��c������@L�(��2r��R!οw&����3�~�Iy a�Z�*�\[���S����4WN��/.]s_ؓxֽ~�3��ň/�UC$����o͠� W���u��n� 