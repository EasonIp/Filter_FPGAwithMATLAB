��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�P��d�d�g����WG��򈣿ҫ�a���GZs�o��K˖"ƺ�ﺜ�e��$���NdS�L>����k+<7���bY�� �q0���\�aR'H��m�+�r�p��n�NT���,����h%���h+��Z���$�51f���'X�J�)��Uq�fM�PX��Tc��Xhǅ����'woV�cufz��U�o�L��@0�!+�bc������	�H���ɩ��n�m�q@Y�`�2s�{���.n�<��R�NF�?�p$�2�*qַ�����u��R�V��i�9IgX�pc���'<��jº����vV���:[>S��.��B$$���W���%1M(6IaaD�*-�||�z}���|�1������o����{7�?�F���0�4l|�L�Lw_~���6��&D_�E5B�\��<��@��w��>?o��p�%v�
���x$Ҋ�i�ũ9}i�+I��Vi��B@��x�V3���L�m��T$s%[P��`��@��p��}�g���L9�l��'�Uǻ􋮶�*�w21c
���N�S��<Ḃ����rZ\�
3]Du4�7P�l����_\�g�Q����84n�ߏ�á$�N�~=h��ztdȬ�����hp��P�e�k�J�p=��?��AO��L�)"�e���%������~W�����|���x j]���{�b��'�4�Vv -�h��+C�'�����幍Wо��ٸ/,� )�lAf�^q��/�������4���Ǫ+u(�+�c�\=�0"ڰ��2瓀BeU�S1{JcIS,����3~��0tЫ�?�7c=��"�zzJ�uH�'6��n�����=H��m�^p��œE��Oi��u�.=�B��SH	�nF^8��,���4��9c��lL��DO�9�C:���ם�Gd����
w���o���_�_��s�f�=S��S�SAB��r/�J�%@�'��!������fv���2^��#����2�����\��:t����?�ͥCTL=���G��w�j$M�J��M��Bv�ɇ?�i�<ZN��X�s��
�\�׭�����<mCIc03�fIl�s���]B�ì�C.���e]M�_'f�����-��fL}��Y,�&z�� h�	ZU�Z"��n��ѩכջ?�T�V>��8ޅZ��f`k��2����ȝ�~q�Gf���x��%��'��%XSĵ�o)�l7�h��r ����w.ۦ��iU|�>b�v>5*�Q������PA�:]**�lY4|Pa��A9j� ��|� �������NI��i7q�q�������^���6�a�1�S��ƀE�"�	�y��1FevCEY��Q,����b'dE��<<ۡ-��杰����P�֓�28q�y�Y�Z��_�˲�����t���4�~��+~�����-��p�u����Ab�n��,&�J�	����',�;Y2�Q93Y�tT�Z>�Eɟ/+��w�p��2®�gʷ��)�@8/���)x8�7�
4�����4�1. ���GO�,���ӌeL�4[�� \-q ���⺬M�,Nŝ�<=� {�+�c4�c����^����1$Yg�4��x"]L.�3�ߵ��z���e���%h2��r�nl�t��oߝ`��7�+j�X���"D�y>�]D�mŋ߭���G2�|�\�bg��G7i�l�����6}^~W�Q},���֜�n�g�n���8C�AUP�F��b2{���'E>^��6���%������o�{I,i_�
 (�g��[�����=��/�vp�d��FY�b��X�+���۝�b��rӆ눌-�f�ʒ�PE�-U��$T��l�%�oȳէ�>��;����@��e?�k���{��Oa�?7���\�b�
Qc.5��JK�ө\#r������s�0K��nl".�m�lV84��P�����V2-��z�-]�e��-O�OB��j� 
�x�w�P���Ie�D���|��	4���	���5�BgL�9�y��b2���Z�P�CXM`��*kf��?���z�;���l/�o/Z��al��;����U�L�^j$� ���9'���Z$!�U�r���H*�c��_������~5 )*$\W˘a�;"�IŝXT���;�!�0ȫ5�hp�Rs���_S�G3b�J�u���c`�ζj�l��+�0IbH���o�	�GԲ �Q�CA�h����fv�����-l�����$�6�k5� �#\+T�15��@��q���ΐy@��47Y�ɞ�r�u�2���e��y<
,�.�D�Ċ��MG�3e�Q7wsst����wq��w=�������-���9��ۀ���.Ԛx�J׊+����f�����\�'_�	�V�@2sC�{ځS���P�4Ur78���U�ja������r4J�=���>��s�QS5��z��D�3E�����IU����夃�Z9>J�O�n�º ��F�)5���O�eV ��W\��<�,(\�@Wi�{���=Gg�޶��5Ŏ8�pZ(��+�:�����܅�&vi�����"���cCӗ$$<�~|[��W@�e�z�H*�c�4_��[(�e�>Z���E~��P����&NӺ�b��xq�����d~9�<�)��AaZ�8��
�,Z����٪֕j΄�xn��}O�d�[�dZ��_.�%^�XN=�v\�����z�P��ag=?�oǐr�(��$ٍ�q6-�Pz��ҡ�:o?�5sVu�W�e}ߋ��E$;�ݒf�"5�^g3�/\r��s�a�Y G����k���;���\5[A�U��DX�3h�4��"2%�XZ�f�<q$�]�y̖C0�� k���A��+�>������$NjC���s"�|r�H�EU�J�����2���F����g]�l~�/
+��t�M�����c�8JHVm�:/�N%;��R�_�U����Y��ܳ ia'4��qXY�&+gPJ9i�~��n0�dZ+��6	|��ŉ���d�ִ�Eu0wq{|��d�k�/vD�Q��Y� ��m�M�U=b�E:yU���[��֮A�	��N?�}1��Q4󼭂��-�q�5�y9�/L�aG��^��[�\��S�E^5��ۃ��>ədv�O�\�E�˅��#@u�͏�<��>��Fk����T�
����`�E��eѾ˵!�2x��/</�F4Ɋ���v0�݈�K�#�Q:��
���^�z�����tAg�Z{����`O��ZU�q�K��؏]B+x�``w�^���9Y��[ �#�̏r*��<�?mu��];$���v��e�y�i��JMz��I�j��)bh9%ȭ�<�#ņ��#�t� {��Q�`ݍ���P�j���'�R�dn�@��z ap�f(�4��� ܂Q��pZm����;\� ��_:��<�;5X�~GV&�@T��ܖg�5E�[��<>��Ӳ��^�ҕd��v'm`I��0:�����3ރc���Չs`��Y���]@�Y�X
/��������K��-z�2N䁑�J�J��#��'����m���d6�o�l	W�Sa�:��_�����qZV|@���cF���o�c'Iy:R跋�?�#Fa�ސ�oL2�PiܳDʔ�f'��7�X���h
s�v���� �5�Z��'
4��ܘsw�d�E~*�F������_��������/����=�Y��Pg��O䠸����W�]��D�3�m�T��A(t���3�0:�%�N�F��/���ae@��; �����߇>)��T��U�^�z/B�,V$��V0�	:a嘆2&�f�>���a�!�޽ޡ��י��TU�y����/6�w�J�R�t>���o�bO	K�qB��mC�dS��X����r�Ks9�_��l�,����uEK\3���ڗr�Φ���`�PD}sr.�U�W�I�0�+�`2e�fR1a(� /+���v�܎"�ߛg�Au���3�W5%b/��Z�\yk�T,���%�+��٣̅/�
��**�=�H���1�r�|��:2rA�H	5w�@��e�}�0�6�{�Q��of�z*�D;����Z�m.�&�°V7�.�a���|��h%35�����:�����:�?�:�����
-Ѳ6?�3�+16�o�+��X&�u�sBX���K�=\��Jމ.�)�,��1�R�Eo�@6���l*��@��_� ��q���������1�e�����pc�O<�P��J��F��<p�])�ٽ�q��b�K�°|�k {q���!M&A�Нd��3�C�_��K����C�❒�Y[�D�)��J�N~3�ݙO�$\U�s�r�[\Ps���;�<yE�TX����P�;����3����Y�
��kx���x��<<�t�^�.�2�.\��E�(r@��!�!؍��n��#����]2��0�e��`���pN�JF.�H�uM��3��
U��2x���:?����(*���4��c�q��_1k��$ő��Y��������ЩD x�Y���'�wk���f�;x�d���<�A��ݔ�`N�k�Il��FN�����W����)�"B��8}���{n�I�ܺ��}3�|�����+�A���e_Xf]/ 3���;�(k�"�L��՟�^��bM;��3��M�z������Jc@����$U�l�}�/Ti�Egg,�j��8\
?F`�Q-�A័�Ϣ?�kC���;�z,�5��
����އf�Хgf;Sو<&���D�7����c�[��f'�j���@���}�4��'`�j�_���N��J�2?������*S��Ap�
���k\��ysV��c-�tN�h]�0�;?-V�����a3�q��}��%E�i�ȏ!<�.p�.?3��4N��#4�[0� \�5o���c��&B�}%��r6���jKX&�1�Q�Aa��Ɨ5��v��$i�x<��Ym���"�����a�m�0�ƹ���Dݖ�s# �s���2H]��UL�������J1���G5=��؞���=7��ɌA�@�����sgÙ��â0�e�8��oM�6���?H2�a�;�M��u���Ѷ�а�F�PO]w@S�t�_� *(�gA/:}?�T��!���M��`۽Q� HNǵ��G=��:�/<𑦵�n�o������r��	Z����6g�-w+�O#F�g�=Eh�<��@Sq���2��Q��/��5(�&��?��aN�������J>��h�N���/XK���؂�/>�(�LM��<��+�o���o�R��O6�����7 �H!\�4@}Ȩ������7���J�m-Nd�O�)N�5p�SG d�G,Q����<n}U9D[��]rv��+���Fz=
�Zk�������]���r1U)}������{�ŭ�Pe-5Q曝���l�U]����m����1�.��)�k�0^�-y��в��Ǚ�LiJ����+u7���e [r��~IR����6I����EQx��$r�յX��4/M�S�`j��W�ޏ��.k>TU���L�P3#zj��
���e<��jk�TL����@�����B#���$[��psx]�pGX�l۶�J0����p/��]�Ǿ�}쳩�nL#S���`�B�#�1�E���z�5'���7fO��c�	q�� �3J���ŀ�
�B�n���q�9�`	�C'T��4\O�d��h*����-?6��9æ}T��_�_=�
��Y��R]�sh|X��m��V�|��=��Y'�aܱ�/j���,��Q)��C���G��Q/���Njwl�5JB�P�Z����F�Uns?���
�����}S@0�� ٕ��:��H�zLn���R��>h��v!=��V��v����k������2K_��+t�o��$}L�X?���-[�a�)1�>+\f�-�4�I���$G�M~�0�~�*U���̱�=tu&]m�����PFz�Zslũ?�:�{u����MmBZ@gT���N�a>?�$�춫f
؈z�.Pe����	!�{�"*l�3&�(�����tv(�
/%���U��k��^mW��cKrw��gb9Mۂ�>Z.�¹�����6�a���B6�=j&��� �Z~4w�S%.����/|b=Y�u��;���=�B�l�l\w��H9�t�>e��i�&�yS��plb����'�D�6���j�R�T�<X,:�ii�PO6��8u
C{ӡ���H|^�K|ή��!�`J9(`g�L# ���{)΢ٳt
+\�~_Cu|S�=�Lg]�A�e��i���k���>d�L��q��� $�	��
4)��T��� �#��v�����V��Z����'���+���!;�Lf4X��ºk���]���a!��	