��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$��Q%���zY1�����3)i�P e��fy�n.ujvڞ�� �ab��b;�fW9��Z"�P̤�����_^�nx��]��-y�>7�Mټ�����mN�L�)3�v���f����4�̌"�cڹ� �j��~�Q��� �+n|�̕?W�
��
k�\d�"q��f�v(d��m�ES�]��o�[t����y���1��h@\6tN?B[4��z���;Q5��WN��ڸ�Rs�߈�E ���x���'wH��6��=�6������arti��x �m�P"<_�~�s�sW�j$���l�cT�0���4�g"�1T�/���Ƕk`&�מ�Be��Bt�C7�,3��1ɢ�9T��1e2��LI�����b5�ѕs�����~1�p1�C$��?�-���=������Jk`�8�<������r�Q�V7S�Ͼh�T>�+\<�6��O���xp���u�\~�g'�3Y��+�S�����c;��t�1�4���������u�C\��C�Z��Jhk� )0���K���f�L�c#�N/��IA?�/�P�#-7��-����| ���}���B���5�����o[b�����(d�f:��ߘS�T��g0�.�H���U���a ����fE�Yt/ʅ��<�3�y)TrZ�Wl�k�^�T<�̠�O�{�WP����ѧ�#�:A��t�Nh�o�yӖ]gQO8p19�(1�B��$�7�� �+�ԡ��`�掣<ё��elaߝT�x�^&�4�w2F%�l��|$�4����g�ye4��#?Y�]ƭq�J�JVK��ߠGw˨����V����U�=op�2����N}ٓ���˝��S�0��<de�{"l�E��7�n�����ֆ���iw���*x�3�����}�8n�c�>�GI%��
֪|�ޘy����w�����}��0$*��t;�Q�#��(A��`��h�E�����S���d�)�Y� o}��u�E��}E��j�j�ύ�7�sO(;UǕ��@�3���W&G��������؜=�u{J琹���9^L���ؒr��ď�I���H������y���ao��'���E`������J�]�r����;�K�8�%Xa;cU6��q��y���������q44�.�V�I�o;�C�0�=9�Iochy,
,)�³�kWu4,��S�<|���_�j	��7�]��������W.�{@��|m�' i-;��ց<".�>���):A_E���}Hw�y��}�*b�F�̩6�<`uc�`�`��D��fd�"��<j��"%���t��NQ6nn�SW��u�k`�M�tJD�#��4�~�:�]�~> �=����g� �K�{61@�j�� H��_g)���mݥbZh~�|��t|?6�{��Z�#}l�N������- �����FHLC�7��-�Ns�8��/�5cpM:��T�W�J���ۀ�}*OM���W���ǉ��|5|�S7z��twF��M�jSܤ���f�L��~ru�p	���M�]�a��+,����ػ)�W�?O��뜭;n?�*�WZV$����C!x�xE*��x\5TRm����V�t�4��Iy�`o�7Tln`��ܩ�M�N�<|�i��^����ѿ�2[6�Z��{P���.���|m��Y�c������;�+�n�J�;&m���#�@A0[wԁϦ�vU1l�s���!�Agk������-�O�A�]U��y� {�C!�B_���Ǎ�j�Mb�b��f�V�L�G	+|`i����)8�X�E�̌�gte4�C���C9܇�
)+�̴�4�˽s��dE,��8��RZ���ס0�WӜ���r�-�45\��??��1-�~��ܒ�7Sdev5��x3�J��FC�]�P=꼵��aN��vf��]Ձ��!�!��{�ˇ��݋�?`	�H&�u#��U�jٹ�h�^V!'=�b��xh�Ȑ|Z^jA��K��:�	��o��r[�Lp;Qӭų�C2���+�`�J�~�J������a�Rx����]�
BS* 2:<���N.����n�$�>��h3��m1��Ȫ��,<)���j�I�2�F�=j�/�=��R����B����iG�叕:?�4������p������H_��V$���3���/�jTv���WB�����v���(�$��m���ȕ��1P!H�z팔�ߟ����-�D?�+�a�m�I�t+�,p���T���L�@X��rnԠ
G9 �����h�}����8s� ����y���>
�*p���bc�o�M���{FT~ �;o�d���n��*�ܭ-:@�T7%�� &��r���jF��?2�G�$F�>jC�..���_��R������]�^J�"E~�_�~ ��r���$� M4)v�V�������	��<� ��RgK8�r���j�D��32�w�t�U^="��ޒu+g��V�t� �U@�}u��r��'��sz0hq|�?*
���j'lQO���0 ~3��ſ��w����tG5u/l�4��,�su$c1]1D$~:�뎆��=u��N���v`�ի�3��x�:��9�}G��br<� o9�4�N�e�|�y�N�Ѧ���������z��آ��H���їC�j��	�-p(��M`��ݼ������3�AG6�2��ܣ eeM{#��-Y��qR+g���3���'����$y`��[m9������L�<�������(���r�~���o�
f��
��恷cq�ۀ<��XdS.ޕȢ�\Zk�ࣂ=y�t��g��9�����h��S�hs���Y�����e�q.��T�h�-ؾ�c������O���H��C�<
�΍"4g)�Py�N����d�fO`�3Tzi�w�侌�U����y�ʒ�/YH%}ף�G�,�����U���2}6�XJ�'|�
:��<[�<�M�T��x�^b��I�kB+#DR��q��Nlr���.��ZP�ժa7)d!Z[ >6���`�/���>�^�m?���G�͈����E�֊%����!�{�|�4g+ó�ZEw
���X4ῠ�<0��a�e�o*&�Υ
+_���1W�uw
O�����m*?,��e��1]�� -�Ȍ(�r}��Jx.̖�':D�Lr���&��k���Ǜ��m��7W%�7H�\�Ϯ'���Q��x�� N�����`�������+�V��ι�zZNoDC.��3�{p�/b��/�Cq�e{���aש@~o��9k�c]y��	���q!t���WkК1�R�J+�8��
N!^u�R�ې���-�~�:LCN���ұw|A�
�~�]����hI�砋�<O!�/�|3��������SM���\�y����R�������[xB�{a�^:��%��}Kzm��w�+�A���� ���y��Z[��)I��b[�~�0$&��@x��퓄1��t�g!du2R��c~洿w�wfu��;�^-��[�'��,�f}�.����AwK��[��"xi&��ř��VpfVJq�B���u�Y;��C���#w��d�;$ ��6tN�eFg��K!����%����p���νs�Nz������z���3�|܄�Z��R��N��x���f��>�&`F�%ş�yh@w��b�ޜ5�gq��د���"���;�uv�ռ&�����׾-`̺+.��I/#����,ô,5)��Ē F���as���������4�(�E�=e>7f�p9;tiXNn}���}P9��� Mh�4!�Ү�2|L�]L�oX�h�s��>��9WU��%���=[�s
[���?7PA.ws=}���� !�4���.ǖי��$���
4�� �L����P$��F5O����a���Q~x���ҡ��L�v���R��=nX�^6����T9I�e'G��v�q�;cf�ӊԥ�*�x�J߱9s�)�$���,��|Jo���"��O���e�\����N2��I1e�m�B�ѣ���J��Q;J�7��(��H���ߺ�us�8����t޴�}q�Ȧ"
 �K�ӱ{a�ö`��n	r)+s�i������Ơ�2��B���=�φ�����U	fh��_!b�kF�<N��Ut��=�*0�Ҁ׀�H�EW��uXj��z���g^�ԁ������8��'vzl	YuG�E��	l�D��RqrO|<V�l6�5�ZGMp�H��7h�Ӓ�`��.
��꣭O��)k�v�
pFs�:zx�~]�����<N�z{9W�����L��z�^a�8��5>]D�T��7Jz d�`���6��]R4R,�u��4�xD:� ��{�LQ�9�i% Ԅ�۬v��|8�|X�B��Я|��F&X�G*�Y����zz�j{~SI�A�Vߜ���ȣp/b.��-���^Ǡ�I�ݯ;�2�����[�Ϯ͐�[���˦˯���y�q�>t<�L�<��1������{uF�<Z�����t��Ȓ�H鸖����;�����X�膕N�i�0�H�'�f�gV��V���jу[�[d	"&������G��_�_ ��ft&]k�i���2�NM���$�d�	?o8u�����1/I3�x��̀�g�W~(f|�W�K��VvH6���,�3ψg��U���?������J���R��l�^o;Ǜ�t�Y�U�{Fr Ɠb���˂�m3U�H�< p����y **�#6|��Ϩ�0k��O�#��9{N2b��#�s���'����p��o��s���)�ݗ���oC��W,���:��Q���,ti��WT��7�t6d�Z���0'?(���7���#��Ԙ�ƝK�3�8���C~z��=�eQ踠{7+�.����ޓxn"��^p�Z�M�>�v!�
c���ℸC����r�yI7���Cs��N��!���3���X��3W�Eؕ�����^�a,
�g�i�����isx�D�'ua