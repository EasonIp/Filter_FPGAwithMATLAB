��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0��`q�M�'���2&��Ȯ�W�4��д��|�6�K!b�'mY�`��L����TR���x*5���d6Z��B���I�aGDȩ�b4춙�J��P�K4Ī������ɩ_	F���D�}R��f�"�Q	8-��d�e�/h!��l�����][A��Y���b5�RL��k�&!�T�D �_eJ-1�3�f��<�#O�Y���RL_r2� ��[�.d�#(g��H���f`g~[�Eϱy~���nul�W��&S��e����׿�_�|x��p�1\y�D�ivM��\%���w�Z�$�E}�GS3�t���c�Adj�,rhv�i�񆖤��@	tsM�����b���(pC�ϐ-�"|{�����D ի�\U~<��7��0�/H[ܿ:w�o���,�O��Xʡ`�%�Ҫ�w��0!�7<1��)�M�t�#��r��.eLY��p����BH�E/����pFk���8y���/�֐���Żvv��n��[
���}����Ac,_ǅ�aoq̓B?G�V�~N����&��ܒ�	Ӂ!����!��x��jD�X����������9b_F$S-i���$�G��^�o�x���	�j��Đ�9�Se��Uy��U ��'�v��/��E��[��"����l��z �-l��w�
X�]L�+@��~��٫����V|o1���� 5=l[ف=�&\'� �*T�(d!Ȫ�+��:AY}�$���lnD'�d��`�l�,�;7��=2<�$�M��? &v��$ſ�1�1(-2��L�)/6O�	��j�n���E�c��92�sV���>�9K��m��r`���y}�Ӎ�R�����g���E
�
������⧚p�Ϋ%˖<}vb�R%N�QԎ6X����=5Ӏ7�S�ڲ��!�#AײV,]|-�KI�;�1��6��~��a�㪊!��o����P9�8�[.�%Pv7{�t�K����Pg}���̺x�����W��fffؗ�tE��7�U�]�SҚy�ИT��MK�+�3g�$/�44�!�~H�v���[��i�/�f��g��'p��p������a0���8�Q��zm����b%�~DVoIbyZe�J)v�Uz�JyՌcXn��v#~Sr�G ���R}]����]�`�Q�N�����˲���1�^�Ef�t�Ǡ�?�	F_�iS�<�pnr��ke4	��Ŕ>���<����� �Κ��5�m�|l?��K_�Ƣ�󾠒R?��@�i�B�?�Y����8J�@�k�UM(=�M��dl7�$�k�pw�)`�6Qwq����G�&��w���\1Ԟs f/~�f[�W�Ȓ��ۗ��8�:~,VO�����q�yhj]�j�t\B��U�(l���<K��㘽��mK�؆Ŏ�xM��}u+�F�5�0��NU���Ύ�� ��	Ӓ~B��;�~��5;"r"	{�t�|�XM3���`I��A��s����H_���<v�d�MWp?�S�!ØLe�,s��<�BD���%g��e�~[eeN'�Z!d���ifhS2�DnC�]Z�O��FV)�p��pm�iy]6"���Р9�tjC�W��8����q�Ƨ�wX�j��v=mKr��ml��̫�c$m�-$�(�Np��x��j�x�őNU�}����ޘ{���c���M���a4��4����n̼j��=�Q���~2�'V	.^��+.�Zۣ�w��
6�0A���^,.��U�`��(@L�k��
X1Ё���`���"p�1��#��{�qJ�Oc�~�w�5Mqg��vٹ\��@��ga_f6�"_�҄�1�*6����-�a���Nc���W	�v�_�a��p�J�S�t�~�v��a����n�?ǐȍ�������#,��y�y%5�Ǒ���1N���s��N��Q9aW͌�=�A��Ix�6SNc�̎����]��`)4k}Y"�M-��ۧ�eOPۃiRs%�pc�[|+�o�b�?QT2��r�h8L��T�b��n*� �j��~=�õ0�B�Eq3��ƚw���MN���R�^��ˀ�ӥ3e��w�^6�`��J�xN�%\`�>S�?\�鼦L�N��Y��`�d9���:�˚���,��hb��I!޾w��K�D�T�?=a1z�7ԣp�[R˸����9���]���ɱ��Y�Y�R�g�J�Ⱥ��k���	k1x���B\Hd^�\3�"�4���)'����2^V��9=n6�CTP�����<��-v ��3��R�T��vFduὑsR��v~SysQ�>�^L��Ql�9�5��'� Q����k��§����:0u�Y�v�_�Vn=�h+Oᠧf�1�.A��\���:	B��F9�����NG b�"�^���.e4���)�S3顮�I�`RϏ�/
>3�vk���8��Y?��������B�Q��,��Zb�1��w�n(E
�qs�O4�*��{ַ^H'e��w^V��7��V�Vj�M��S��*B�BL�У�5�y�1���+yWI�=���>(c}�]`;a�h�#�UV�r�'��I_i�K�V�Ǹx����Va+N<us��O�2�|׷]��k�02�{m���׼n�X*�}ԉ�Ǡ�LD���|aV�~G��w��W_�g1�\0}��Q�V|��ן�n�0�#k2mc�O䡤����טb�F}��ޗ~ܙ�)�dϞJ%���t���>!���}y�1W�hr�uLX���[�jl�f�R�o^65'�"�4�/�i�z���',�6p��8e��VP�9]j���鏇V����`�Q��F�tw� l���4j��q�$���l��� �8��F\��Z�6�\������WTU&�*u`d��д�Vh�Ft	�\�c�[��1l~���z/b�g[�u�^�bEa�N�̭�Ե�y�����\����3��/W��W&a�uL�J�zw4��V� ���,�n��P�>��U�h���Q�0��v��aPڍ���� �F�LJ�;�'\��d�<���-xj�W ; ��1E��/b��yv�K>9�W? ����HLx6��3g՝���I��B?�H�6O���+�񉶎m ڦlY�HH%j�Ub�B����q����b�^��|D�=@�i��3�+;�Wc�,3~�gq�zK��0
4x��,�X1 dW�*+��B���E��q�fE�&`k�I��v�of��g��GU�)���Yr*i^e�;���|b�?~�ʙ4x.��8�j�/t��[�#w��c?Ѱ��Tm4�4>�a��q$N���3ezo֖z;`���Y���-׫n*([ր�q��X�{��;� F�:3x|��O�G������܁�/�5��%������L�K�uVd��	p�[�.ׯ��O��af5�e�{��u`����9x[%
z�����u�A� ��vu��	}��ϰ�.����4��8T��;��Jo(�W^����}= ���z ��JLܑ�,�n]d;���T�0�� ����f�m��#`���5�}���	L�L88 ����b��$����;���Czu�c�O=^g�%��Mߐr�sL��;��&�Q/��u"�2Va5�V6c
�
���gD�u�6>��Ç`��J8N'��Fl��������`X:N*�u<����,�5���`[��´��-u(�J�TJ���?y���J��,'��;3n!t��7�S)�g�q�ǎ�C��D/fG��`��~�&_9r���y$��gg)�J?|�
1����<�"8R*In@�QZ��ɴ��^��M!���w�|��	5e�YA���*"�;�օt>���81�v�7���$��N�2�gK���;���ǽq�E&�H��q�q]ʩue������AVJX��x�J�v���s�_G��M�Q�%b����ȕL:־�D�8�$A�eaA��Z\4ͤ�(�'�ty���J�j7���W���8V����2E`Q�������5�i}x@W5�$�>���$A�;���08��@�^A]�,V�>��ӝo���P}t- ���'L�C+g���k�<k��>������+�2��q `��ˊ�ϭ��g�Y����I���(&$.~d�C筳G��@VX Vu$�bo����a��L�b��2ݛ��.�j�2��3�g��h�;"���=�dѫ5+�s��C(%�b��Q�l 'E`x/��i�Z�:���o�k�+����D����i�q�Cw=�ibƯ���g���	��B_�E`ā�01�>��������	�~��c�NSn&����n$I�_�lO&�{-Pq{
˄,���.a�3�5ሲ����)4x��U ��	:j�U�?��uo������9��)��;6vnx*�-��z*�F���Ě�l!��L�������6�h�qqJ�Ou- �*���Ok%g+���-���U�ȿ���a��qͨ��:Bٮ�)�
�*���0���e�9�����8�܈�� �LLp�{��=v�l��`�-�5���֘f��L�䱄)]2���OX�O�T���#�D*�J�Փ�r����`��L�vġkH
��br �W?0��K����e��{~�@V���ӫr��{+rYϤ�3��P�7`�לR�3k�P#_��i�<?l1O�I��"~��{:�6��$L�0�Q���&	�K��dK~yVx�ox�;���fRz�(dþ��Qi�����J�i����/U���`�Z~8I�� �#4ľx�&x�2]���o��Y.J�E�v޴ɤ.fQ�*��_~�B]Zkq�y�4�BS`J@{���&�Jށݲ�D
Oq����׏+=wv�T�u�N�|иv��(���&�f:�5��sN���9�Hԛ?���n�������Zp�a�T>h)�WJ�����VVlv	)_wZ�H�p����D	�a�<|�h��#&�ׂS�&l���4KˡS۲y�����������5�p��$�_��(��sy��q�`e��g vp 9.�i��6=��n�GQ>����{�kL��7	k3 (H�/���I��F��K6�<q{8���Ld�M�ĞtK����,@ɹ[���И�.l>�Ou��E�WǶ�_��"ڪ�Ӕ�����?'5�z
Ej4�@8��,�\��Á�2�R}��9�M���w�ygK���$�4|��$����fdn �s��.��?�Y�T�W�	�tq-S���*����բ9��je�lB�(�L����!��H|zZ�ysD
�.�MPi�U���������LB�19۸��pN �gCIy5ؔF[��9N�_�+�ż|Vh8�>��-�̾n>���<��]�	��֑*FA�O���gU�Dn?6�����h�8Hց TT"��3rM�YT�u�faV
k�U��GW����QH
��=3��Y�dmN�_ 9�)���n0�੨|�<���y�k���Y�F��/��$��Wz��(< 4��ç��&��ۉ���}�hBo	�$��[LO���,��n��N��L�pn�F�Uf�W&�/z������+�H���Z��<$����ѣ~�X('�6�+�=ӟ� �Pe��a(t�ż"�ۭa�
���=:8bb;^c\�<��Q�B�iͬ>/��E�tj%���`��!�q�=H���:+��@t��փ�h�Hh( Ca��u2t�E��g�H��Zׂ_��,ǧ8�x�A'|L�߬x&U	�S�h ��L���5�)��(�{��'�D�W��h�ڊ�K�\�e�۝%f����A幞�oe��#|d��/ёը�ɏ����׵i���%�~Y�D���Q�z���\W�� L����G�BD���u���أ��_�dL7<�fx�"�	[�X�+�(xi���44�AVY0������<v���;���\M�|��m k� ���;v���ά��<t���*f�yðc�J4a�����4���3��3���P$�$�,��Hu��K��ʚ�s^��vK �I��(� 
�� ��({�M_Xw�c+j��9�}�;5��i����X�jds�����ݕN���Ch�"�$f�ģ�gt�dv�o��#0��<�&V,�v�!���]�Be7;h�&��5.>|~�+e�6P�h�1U�j�2�ؔKwo|����Sp1?�.'Q�o��C{���.�#�&�_#�r��7���"�%�l�6� 95�S�깠fb�[�Dq�LP��]*��?��@!�3)�b}��I9��x��Gu%#�������%����=wǿ��;i�|��F�H:����P��z���d����l���Y|<jd��h���0䭔;��vt��GS��[ׂD�ց���5�E�9�/q8�����n'�	���7��=߸��ۉ�<�iq�J���Jc�~�W�q��!��ǰW7b9U��9Hv��n��)A`[;t�2$�6��%�.�|���%�n��}�s�u��`.9Ap#R��;��%Ԣ�u�f�d��!�]m�$�}������ށ�Q�� �͛ڞ{	TT�P�̆sB��+�v�_z��Ԋol#Ĳ���)�vK�d�;��*��|q�5ȡ�p\�%UwP!h���gx��u�%F�:^t�t ���z/I���iYϵa�C��r�a�x�R�|s��U}��~9$g�#ӌ7ui�ڀK�y��	�����UR���(68���^�m�`�L��{"#��*~�?v�2�ު�������#�<���5�7�q��JHK��o�v�Fp��TD5i^pőc�MsB��<s�������ZZ�������j� 6��jL�a#�Y��X�O�	��VWZ��a	�Q�;�U��9�a�/Y�ߑzo��f�o=���{����bV��9�vAO��vӚl�)�u�$=u���:�o��9'P�pT�ʁ$��)t��Y��L�������L��!��V�2��͇��)5c�e�Է%���<"V1E���~�S"�㐩#4zu�F��Lm��O��h�e����$�͟� N>2w���X"HX��G��?0���Ǳ}i51S�c�Zb��Wm
i�Sޕ	}S։1���j�$�
Qs.{"o�6A����2/O9��ʸw�~�V���`VY�;f׊^��~R���J��sÛ1���G���MIi�}���/� �*ꪷ�[ݺ2v&^�c*��9��؃.��Ry�<��D�Yc��G�Y	�����?J|-dv	ވ��"���1E+<9ґ��9�4k"