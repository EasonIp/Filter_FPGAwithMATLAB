��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~���"WYj����i� �N�7A!�@<e�]ң�;��5D�監p�.� ^+��Rk0;Õ\z�7PF���p�e��	��j�kdD/���1M���(���T�e+qr)zD���FWkV��������\���mk�*
`�R���	j�' �� m�cD���9:�DhT]�����۶�����i����ޙ%��d7ܷ��	�:���U��(�����#���wv�pFc�o�m?���<�δ�7P����( ��(�����1���o.O����BE�l�pSX�m����
'j�ߑ?�a\����3!���Dꁖ�0���?��AI�_$�nDJ�^I�i/p���Sw[���mF�AjCi�*q*j�+���ޘ�(�|������{���y'S�c���@s�S
'a�.ݐ�ȕ`k�5x�C.}��. [e�[���5��n8�+�Ķ�b:�)Z//�V�h��oĚi��~]W����{L��O�}�>�G�#��&���R���~����`e*�~�x����f$;Ԃ�u��d����{�7�"��^Rr���;���:,8���d�BqƖdd�'_�O������"no�%f�wD�x�	"�xP#�h萩
;k=
���T�������.bX���C2}i#i�\X�s��'��z4Bj�v6�q�! �*n���C(&�����v�ۍރe��mQN���(fc5w�s��n��4P.7^d���4_*���Z�&����t4("&S��G#�<1J��>�rۘ�((�ۨT�g"�M�����߼2o��!�_�#��k���-[5�q�J���ϠNQ���)����Qf���ЮC�\����ak�Ȱ���VOb�0S��z��US�~��0�,�h�4~�^��H���r�Y.r[�؝j-�e7jH���s�'���],4v�#0.�k�Ř��7;\�n3X�dl�pQ!uЎgAP��+h��J�|�.�U�t-^]����~�9�a�(�,�;'�:6"��^^�ha9x=w������n�I��Ǩ�y�n?44�5��{�΋u�D�yb!e�՗G�P��ݴ�toΛ���Øhu�v4���m��+'+��X��k��UWT�m1�����6t��('?��y�w�@��i &�cuZ��U��笡���$�O��"�r=�Kl�х/��󙪜���>p^u�� ����.�+�T�|�]�ʮ:�A�]��K����D|I����xP40�`7�tQ+6��%��NĚڋ"��F겵&�9"w�)f����mc��G��hڪ������ᢀ��0}}]@Jg�J���!3H��+�g���m{P�?�i����3� ��d�8�X'
�`���}~[�����������e.�C��n���<�`��[�~>j8(��w�v�UiXe��A�;S�W:���VM	�Žl+�^ �sx����K9>UN����� ���<ߑ:&���]f;ʹ�>���K+6����=���i�ٿ�z����7���&Neӷ[셼4����"��KT�tg�eֹz�� ��[2��T9&L2�gS`j��4�K���R�5�#�Q��8&��q�f�e|���6ݮ>�Ԝ���s>F����j���g�->rzKN�~R��"��Ru��X d��q�j��J~��;��@އv���|�DfIeLD>[�	?����������-O:���}�_��}�'�ړ�C���IkR͆��?���X�+d��>{�Я0��L�ސ�L���"���M�����ҩ�x/@#MN�fiȗt���W<"�KSF�A���*6qg�x�n!����R95�u4�m����AE4��Ò5���Ȇ������(� %��EZN@���5RQq�;a�NL��t��ō(�S=G���2�ٕ꒰�>5s�iX��
�8�
�v�K�ʲ��ՅLL��"�j)��2)rg(��z*�1v�Se~X��1~^��X4=Z�%���5GX�`;�f�K�	
)��Y	�E�F�e����'�Yy�wg�a�blIQFC^u/?�d��<��Ԗ�ln��P_Y]�5��x���C\��)�.�zD��sŕ8V�s�nw.�s�a�7K��ׁ65�ڌ��Ғ�@	����v����Ё
�H��Y|�
QIy֚I����u1�����GU���F�ܾ���L��"�I���W/���Fvh�\x�31u��Lݻ<@&}� ��L��_Ǐ$z0�e�Ԡ47[����c<X��c���:���4	�  p'�n��IR�:���u��f�V_��^�+</����v.Pإ�!��C�}���v��rT/|��B])�b�Ifu �O#��pEh[U����i5K����h`J�$���.!6�X�C lNo\�I��x�\F��qK2�Tr�):ٍn4�h{G��6뺯���y^{��p
�}Fm����|(�9 S��z�yi���#�0MZoV �J�~�K����]��B�?�4EF�6O�����AVذ=��`��5���������{�j����*����K��4c�ۈ�S�����:y0r{�/�3n��oac���WQ�����^i&��BLn��&�f^�=�)��]�M��D1iF���d/�r��-}6�h�4�-���p`�ZL-KU#��k��7�)�&+�N���r~W�	W@L�����w^� ���`�Li��Xw(����c���P�O*?M1�2�����?r�w��2�g9<@^|�]z�e�x��!�U�0��Xp��2�/?�v�<RO�j��rg<�=�u�ૄ�ce� �)�:�sJwo_&`�>쐊����b�+���O?0m{7�D=��}�.�!b�t'�Q�@�l�����[edIi<�:�Ϲ̽�=�p<{��_x=d�ty��E���S3��.�2��s�3���S&��o7V�j��+j�����i��l#�O1;_&A�3���$�2\; �����Z���b�Ua�}J�:�!���:&LT�����m�K8��\h=�jt����.5P�K�$3�4ە[=L�,�`%�M�_p����*4[�j9����u������O|aH��v�����x�8V_�>�š�������������5 �ƕ�ӄ��J���k���Y'�-*�UK3p7��D��2�qϛ���<�6b����|Ԭ{���֐��rS�4�̎xsT�6[T���Q��߅�?P�t,���R[d�e�#�gu=�,j��T4�|�`Y�B��_h��V�E+M����^�\�ҽּ|��6��g�]�>�T�W
槉�A�S�D�D�+�������z_�D� �P�ۇUfkث+��&���"�tm��lgZ�u?���IO%��=�b
��Z�E�~T��#�q�J�#)މ��o8,�*<Aa�+DɈ����lU�i������w��'�#���u�����N��T��G��g,H�]�S:��	����X 0Ef��mU�� ���M?����_B
n�S��ZRhx��F�d�)B�]w�B�oT6Ԭ���y��w��C S�l�<�(�Eu�|6 �LR�V�:z��W�X/1��H�⥵�	�k>= �/��F�?�- �r�d$ɦo�>���N���pkT6�&L_���T��ڭ�k�\ j|@��D�Ҥ�����z.��(8��ϤA^A�$kK{
����,�����F�n�,D@��Ɗ�Mi1��^���k	[>��ݱ��9>q�,T�p��5�X�f��2�Q{ӛ���za��#z�W��^D2{�����e	�"ݹ��b�_����*s���Q����!�캴�>vu������Ng6�?�nߪ��n��s*��◧��zo�j�I�'i�X�̂q��ɦ�f\j>x[�� LEb�TX-���6���M��Zs�qnX����
PLx�'�;�����/%����t�W�,��7�	��jS�6c1M�"٫�+	`p����r g��plc|��3^�1g/w賤�e�)�ۼJ�;nZ?ҕ&Y��J*{H��@#��+�d�y�)si �a�~���8��:�GK���,/��ǫ���� xXB���j���/���-�� P�ޟ[_��ERVQj��s�ZHP_�z��2\x)������D�LW�5�9H�c�B ۆ~��|L�����b`SF��,����w��@��7V]�;��Oh������Ah�
�~�ؒȧ�������_��qV��$ y	O �j_u�Fc,�ſ���-�b����9F<���p0��Ӝ��;���X�[�������:� �O�9l�������Gw^?>���5���P�/�O��2i�|�6:>7_\�a�+�աzpN, {a&�#���!�z5^4ۀ"4(�̥?��K}����(���L/�|`�Gyx�5�vQ��#c���4���i	���T���_]�ah����ΰ�v���|-2h�d.��v�o���������l;�Ksf���VB�Z$�-�B����Qn�h�qF�B�ٴ��k=~Eے���hnNb���@�c�gc�h��B�4y�z����}��1T�Þш����x�m��S�wuS�/�kf�)kӜW��ī��p�Puz��2�.X=r�����\l��wO��F�?�-�^g���^3tC�X��)Պ��{X���o�8x�Z�Wq<$Zu��-�U��aؔ�ɐQ'C�202�b�F��F��Yp�^'��=�����O�����,dG���[ $5z�������ۀ�s]�V����)�4�̕%j���si]A����k�X3��v�"s����M	S��s��Ѷ�Gk����,���b\J=�h?��z`�E�4�1����v�^
mb��F�ԓ�[��dT�:��� G��S���hP�G�(�N��z2�o0K$C��嚜Y���/�hUK�ȇUTaq"��5Z�[�G�� �$W�+�%��d��Q

��w|`�!#��0����n��!L��e���f���5��j�=�a�.�?� �vvq���.I�\�(��O�g,���֒zQFr�.J3�]M|�_��^&�!�	K���d�2O��d�!B����ҕ�b��V�"��_	;�~k�]�ƐL/(,@���N]sM�K��>�
N���8��(��}f���~V��_%Q%.׃�J�-�1���1�--_���E��|��V�Z���:���^���k�|]8w���&����~s��5�5���s���;�-��|S��~����i�]a�P�#��le��`0��`����D�N�:�;wzPAL��x�t"-"f��#7.]�m��Ye����c<7��aU���F��ZN?�
���ݻ@>�*Jg�������b\*\peӻͧ�! u�At`��ו8��RLY5 Ph�G�nq�\!"״%o�{�5ƴ�k6xx������)xt'6�'P��$$!FPTnj����M�	x˂�4����q�OjVL�M.]h\��Uѭ�/�k�%���}�e�P��ǔ`���G�CX 	�^��^�	�-/�2t.m����	�&N#�V����MDq[�)�`�c->�Ԛ�vU5��[n��d�E���z�?���.�<����FA��dͳ܉��:��	�e󼜖�$���|(�o!��Kp~�ju��mɟ"5[��#"�oI-a.��<��m�IV�g�m��yY�����G9�� owak�<�v�5?XG��� ��V[_{�&�I�A��]N?=A���31y���J�ɚv�����FH$��������Z�#G~gG�d�j��C��_��:4@&jA�hZ��'����]\�����6��gAm&�(V%�S��˂��k�k�4���ǫ���7�0l}x'l,�F{��v��)���Asf٭��Vw�]��T+V#r�Ӊ�t��M^J�zYh�Q�p�uN�a���� �t4����o{���/5�G�$�ɽ�ϫ��CSTV��h	g�����P�E�4�[����*�(��b�G�{�B2]���o2�>�"<X�%��G�W(�Ḋ9�48M��"�Z�*�t���@��#VA^����'��/�,9��a@� ��H�Y�A#oD͛m�� �H)4��X�=�*:�.Ч*�{��I#���(�f�d�O�$L��(nC��J��S'�AY��C���G��'�2�7-����X���v�}�T���:�Uh����8>�������{�+nFc���XIl�7�[o3_A�����:#/LS[5	���B]�n�&7]�}!F�k��&�P�v�6����uN��!��o������S��@UOl�,��?�y�W�N?�еfhf��S#Ц�s���G�#�"1���ݯu�\[�3�Kvq%ƱGe��BҦ�9A�Ab�`�+��k���1ߜ��~���7+x��4EI$���N�Q5�Cy{
ͽ!,��nN��x��lAB]K�
u�&�B�ۧ�v���Cհ�B@�Q�n$�?DL;�k�ݍ�o�����n�4
�T6�P�fuzA��#��)�C �ۯ��G�fa��]E�:b��@�7��9&��@[t�ٔ�	G����{����9l�Yv��#u�u�vތ'�l�������r ��%@W"#�3�C:V�U���o
o�~	�?`b�&��EqRC
dC��L/}&��+��61
������a��<](+Hɲ=�\OL����u��ZwR�]��g�����w�*��(W�F�z{脟�����e�;���%�ǧ���Ki`^}p��)��̩�I� S�g��#e3����$*��'Z���_Ff���õ���<2�Yt55)���+��X���`¼e;��!��A��:�t9/�NAoi��M��(g#%���^Z�e��l�Qyqγ���|p�9�c�����������+5�i�����X�d���I����+V_��e�6��@��)t��q�|��A�ϝ�r�R? �P�'�f�.��`��h2�0�4�n�ZQgo���h����_���6�s��)ܤ>��A���6`�3b���b
z�+�l��qF��LhC)�5HL~�3Z�ޛ�t�3���B[��B�= ��+�˧�k�Hk4�$����9�=pCs�����n`@; X���`�Qnc}xg&�z��ߢU�o0��a�~�Af+ ϫ�!�9w]�^����<��G`�ђ������	y�Ү�7
�ܑ�&���mu��1G���xں�3Q��_�l�r��8���@�0�o��e�_�fĩmW$p4�=�U��U�ơ�5T
��V��3�w��a�r��o�3g���uG�A[g����O@.�qH�DK�� '-���\uH`��Z;U�/
@�5���!rƗ����i/9��;n˒�t9B�k' 0��9�q�.,�}�/���VS����*7��J�c�g��[�6C�«�E�L8u�u3m��'����بKZ��D1�īs��Q�� HMbr�nl���<�PU?QJ���6����zG���.d 4j��!���i;��ĳ{�����k8��EA��r�*c�c(�|�y�$Af���P�z�q�/��h���:�3�5�� i���u�+d^J����� �Nf��m �,#��������m���.��q�u�R���*���YVĠ�Ց�DIV�b!O�YrVA�u%�7mQ����U����ע��f6a��)df�Pms��G�b�z$�${��]�ϥ�<�~c���)>+�͒ʟ"e�ͤ	���%�0��FU^��27i@��D���O
̪�������j��t����-���ܟ�)���w;���u����^�W�D\(�Q�� sɼ�m�������CF�}��`���6���񦦍V�Z9�
���D�	�a���$=�:��k)��<(A�'� 1���X���$Ls�͈�D�	���`�t��
�`��P�$�oh~�;�a�v.	��'L��W��rb� �]#�AL&��Q�����y���� �?����2Ԉ�\�>Aܡ��v-O�2cY���)���&h�VR9�}�>���=��G����'���w���5�S.Ѐ��Zս�h|�f�����#�<?%y@|垤I9��q?PBH"HM}���\	����vT�O:�Ť7l�y:8>|���2,�F��_p���
�VĂ^5�J+�e��6�+�o��L�K�u2���[/�=_����Oh��փŢNG*D���k��xѨ�o�:�>k 9R'��v�Z�']&�S�>��5��L�ۘ)U�+
jB�/>,�=����hK�u8�� ��Z�:�޹�ķRe�Kj4��'E�i���ǭy�ũ)��9��K�k������KQ7�y�Dg��1�`�7]d���¸(�$�DSA3��׻�Aw-�F��ңM��ˤ���=��ɶ�-ۺDB�}��Km���F"�n׆L��ه�����О[߱�FK@C���x>���*��LA�g������˴����j�x�B���O8I_�hIʗ]���~��4�(36��\�0~��(7.f������ֶ~>m�5i�js�~|��Z0����ܜ���-b�Q��̶�v��Ī�Q*t�6 ��VĺEǚ�/g��ǆ��T�^�oٞYW�u �������4M ��:�p簘鬷J�2�)����c`�v�8u�"���Ě���&��~%TU��-I���11�
�'@�,������֡/�~%�PvcC��!�ߦ�T�w�������Q'zr�p*=�����b�3��3�����Z>m, �������[7%i{��4����a'�I��,� ��t-B�S�q�WE��U�*^TŘs���'�Hag������z�u�.�#��J6􌮻u�]��Ŋup�Ɓ������VP���`@m��/�3����#P�n���Q����Ali�`v���{Fkk�!��=J����;�&��Eـ�}P�1nxɣ�����xd����j��P�k����ې�I��M�����I�i>���."��#�7�c3��,ԤAK=*��m�=o���i��y�=ʊ��Mv���e�n�\�&��E��ԁ�F�-�r�S���D�3���5�?S.N�ų ���=!t����Hs�K���Ĳ������'�JJ�V�2����H���ֈ����S�?���'�ͥ.\�)4u	�Cɤ{̞��Rc2�_���v����+?�����SA��W���0����|����B�Aɩ����ǂ�w���iY~�yH�ţ�o�o�̧�]��U��v^p������k�~�|��	�h�냰ګ��Z!@�&�pE3]D�J��ߠ7i��[e�)e	���q&?�X��W���������jA��*=�{ɢ�g��IleM� NF�ݨԔj�_ѽ�[����uE���0aw�D!#��?�v|B& ɚ��!���x�h��% &�U˩���j&�Ȋ�8����W��Վ�b�|,YRx���x��{˳OR|V9~�Z��Q�$g~?�\y�#w�	�6��+c�����6��`�GyM��V�7�\+h7>��j܌@Ņ����ت�2:��wg�p��>��z,���|��M�W@�qNź�
����H-�U_<�!�wY/�f�^��(*��~�pF�[|�(J�ɖ(��ڸ(Q�81o'ww������/�5�&���8	F)j@]��Qw�ȯ_f���1|��0��@��W�nK���Vo��`y�(d���2�.ೲ�)ܿ���ݯ��,��mTG��MY��e��� '��v�&�rH)F[i1�(�R�3�L�kJ/^ݭn^���8�gy����Hv8�����Դ��n�uY��6�-�_:��v�ӻ�3��Q�Qy�uO����U�p��B�t�{�%�xnŚ��	�q�Z����b��W:3w��ce�ӟ�gn�}2��G�e���CI�Z/@(j�k@�k�����_�V񢆾}?��MNʠ��7(J�B����U����U �7�Y�$����5�@��+�LG�P�#"�J7�͗"��]bĭ(��%H{�y��e�VIߤ�a0y�|��N�h��A�"�υ"�%�\�^�n�6�̽l9[;���҆�4�wk�R�����Ey�H�jj�f �ۂ��	T$Æ*��T�Q8���?�x˹�,��7�}��h��ɚ���t@���o!.�P#՘L�&�p�r�<���8�iۄP��}�>��E=*� ��p�^�qP��6�2���(�K�2�/�^��I�����ݗc� ���p��b����٧� jDp�e���q�IfyMѯ`S�jy�͓Rd�n0g�ե�� �1��hHU?�5�\�*��r���ɡ�\=r���Sf�jHn&�p�-G�lu��aז��Ƴ%�Io��c�_��ɐC�Mޏ�q���X�K�)$�}��d]����WP�ɡ�U�(r���J���X���o��0ze�=�A�|Ġ�t<��K�æ��5fF� ��-�r���Tw��j3uMmt�	�F�mp���Z��b��t�D�;��j�⽏f/wj�6+�F�w��P��\��f�{K��s���%������{�(RdZ}���a�E��R��4�jBiTYY�gX+�ʗ����>�
�L�U-{���R�p+��p��B$���*Ŷ�WX�=�PoN~���j��أ>���	'E��
�����#)r�*Z��}���Iۺ�^�,�����7zZp0i�����a�Xg������ΕE�Q�L�[<r_�����)\��T��EK[u���G(���N�|Req�7n�}yq%���/N�,��=��+�_�xlc�>�?����q��OW�M#	�����U5s�!�Ȥ�k�F���yϥ4�o'��AK���PL�a�ie�♊����c���9����ܨ��Z�G˝~c���Е���Ϩ�@&U��\�J�aM���r�×f.O��~�`�,������D�ejs�.�+��^�5�8�{f����;>@��(ۗ6E���e�?�1����^n6���ڂrрIyߧgZp&Ԕ��Ҹ���}2��&0��k	-�P�/��P;*մ�k�ORm��@��,�xA��N��	o�Ne�D���@�^	�ş��lx�H]rC ,w�i��v���M.�y$)���"�G��}�	���^{\}�����!#Sqr��
r<f��
Z��
u{iUhR�6� �!?j�Q�
f�*tj"�����oެfZYD�P����}S/o�hL�Dc(��o8r�G�8�3a䡦��"���8���3	�_�3�7FX����
�a���}����KO�N�	��ÚE���	�H��<�8��q]Duy�&���#���-bx��$|����2�H� �����Pj�����Ic�e���j�@�lf�szr$����� �ܐ٭����=�V�5��'V"�"$^_�mvqs�4T�)6d[am�<�CEp"�o��C�����#��/
{Ϩ�xun����
���߯���k���)^d�bL|��/,�v�!V���7�����Fk������l�l3�E��_80���]���ٰ�� Ҫ�y��̙}��o�u�E�=�	1_�����%�>��N�F=��L}6K%�����z-P@Ƅ��"6��/���k��ٽ�����E?[�_�"��Hߞ�^Q�`7H�-��X����Z��.����+�����	�&�;���d0������	F��������;�C����5��s�fR�5�)i�wƺ���H��08
�p�~Q�c�7��4���=j�ߴ�'�bJ��su�N�	7�@�Fn�J��Pۆ6>E���Iya�8��ۙa�G��@V�3'�D��PS���m:Z�[���$J_W���K�y=;��W[(ٵ�#mJ��H���<G�
�x�d���y)�|�mY�����.�0�0�9�]�C~���q��խ����O1�`
OZ,wVp����aJ�$�o�!F��5�a8���� ����������d��P-3��+���^�G�A�s����bF���n+1��?�C�}��7����
�Z��o`[�oۮR��|���\[��QMZ�����p~4=��js�c����:��0����OF{d�r� 8���^��Df�����~��|7����R�ݩy�sa�Na�\���ev��m��1�Xo��c������4��xwKH.�O�/�B��B����7s�ť�2���r�@bQ����w*K�	:)�u\H�j!�R���[�����Q����=T-�&tA�	Ӊ����o�wsp>����s� ������h���>�6�'�qx*&���,�x��������B@cvp�L�{T��b{ࣷ��sX�U�F�G�dFY��ߠ�Jg��Rb�v����i�<���g�zY������~g���p�H�-3���ԍ��Ka`WIz�^��>O��?]c���*1�Y�����> t�21�ȡ@u_D�7�=g��x]��j��T~*��1b�3,̆�Z����`H��� �]�.kA���ֱp�j�I�L)l��xKe�|E��R�|�aل�}����M���8��r��7�����;0�f�֌ջ�[�����
�E�U�U
_[6��[�ߺ�q���{�>��v���J"Ǳ2��tXf��򺊉�#@u�˄a ��F\+o� eW��Ȗ�V<�L�~��bgew�����,,A�5����$��*KAҸ��l�+^�����X�d:R��\[a�9hH�5Z�b�[~១U	g��g�߲ E��lXf�OU`��Eyr��3	�j�	E�}���vݭ{0� bT�R.��{��ɞ�ºL	�)�V�Hu]�@�)�r����_K�r��K���x��K�q=�
����X�.6,��-��$�ҍI���Te�`�����-�m��������֧��Ȼ����J�o�:��r_�P�W��5���|"�s.jt�K ���G�4EGN%�3U��T�P�Yo�(`J��H���_��o��M<?��!�GW.��Ԣ��`�1N!���8���l���ꖬ�{ؑ����J<,2d�e(�_�1Q>j��L<u������R�����ɣ}���c�I*@�a�~� 4V���!_��F�%[+h���x��}�A���A������(��)�n���hlLx^��6�1��m��?�-��<�WXZ:�=��ԝE�yZ�p��"�zZQ�ʭ�1�o���M棉,~���M�84T�Ӗ���NX��v?a�c�}����^w��3�d|Ч0�arx����=i��s��3�ŭ��Y�v��A��H+Ykk�[s��z>�d�W�s���5v9)���k�o{���p�ww��������th�$o�\u@�k����ݗ^��@M�R�	�;�����Co������/ؚ�����Cd�e{}f յ?��6m_���3!�ti'0=�#��Z�L=Ĩ��t{O%�w)��!��c���zL�8��b����:�ovS�I"�7V,:c�`Һ.�6Z��!�E<A�\��_pe>tH�a]Ʊ�l��uz���u�$�0m�<�>d�n%kڋ R�'yx�l�o���EM�*խ��-N�r%�~M�c�?RgkR]����w��.��>��K��MK���Մ�k8՛�4ht����IE����Ѕ��^�Kޏ8ٿ�P	)���Zo��Baq.���C�HCY��$TQ�!�9r���X0ޓ�L��AN�X��_���46v�l���3�#��Ë�+���e�K2����G�y�R�f�v�� ���F�Kp'�2R,S�8���]�(ex�D�+�8��|ڒs��H�z�ɻ�:x�joa��4�?���d����̞ti:DE�m�`4G ��ݳ���S��K�Tďy]�u�ROt����󉛳C�&bć�mD�J� *�! �%h�4����Op��AR3��Z#7t�����E���a��8_nj�^�'m�[K���Y��Jg��ё��^˜'V���X}�u���4En6�.�/a�F̹�+nj��l����g�mR�ŵ�_v4Uԯ��i6{�K�� :ĩYj%|լW�b
=*�0H�j�k ��\G�<kM�W�+& ��;H[{
����*0�8�E3�|�b��^AA�p+&<�=]�P�v_�N���M��Ǖ��V)�S���
��|���`�)v��lA� ���F;�fռ@Y����p��5�CM!�6U�X|�=���74&5�J�/�<ݼ����k0�~��V��ߙ�K�z��hy�,iǬ�����q?d�ǭ0fN����-�X!#�klS���m/;��Z�$;M�c=gmn�-�d��ƈ)�~ttӒ��xr׬U�����3�?%�U<�
�Ƕ
�1��g<�L�1����Y"��||�%���hs>gZ\�	*�&�ݐ0��҂����j�13���h��p�"�^���_1K$ͻ���5� x���
���) YD�}�5L����m­BH/���I���-�jv֝H�JA��%�y��ߠuJ1!-l,���Tn1W׃��P��Ony:�Q�Ev�u�T���lX��K���/���{��Nw>����eߖ賣���ά�5	@��]�g�acHJ��� ;��(r x�K+��`�'���o��z�`۶��)�%4�S���H�S�0�����?��i+�i�(@`����ȟ�ˈ������m�ݣ݄v��]<���� �2�Kt�I:����Ti���T".G�g�2@�I&�H�Zi�ED�M�����mT}��a��@c������D߬<⊗��-��ͣ�:�9&��w�I�I�	ʈ�o���.0�8͟4�1Am��)�n
e�':B��	A{������!aEp�s� �ֶ��5�8������B�}�*~]�VyB�uX xjh�ΖYq��\[�)6����?Tb��բ���ngČ��6+@.�X3�_2Q�e3�S",��'�x��F�����3	T7�Ŋ2�J:��[�+ ������R���Q�'�w�ӟ�4���;�D,bL"]��� C/�(�"x�'\}�I�K+HT�b�;
������IB�x��u�l�Eݕ+X�XGw���T�W`�׏>/`0��j�m���JPC�ўdƏ1�΁�e:UH�^�a��w�Iț"~�&!�`;�*���y=��agV�����n��=m�a��	���_:�+!��.<�Ii�P���=��ԁ\`�e���c�xb_PNz��jq�L؆������Ƙyh1���\����&<Tl�I��ǈ���Yx����[_�R/GSZ��t4�L�i�I �����o��?W^�B�z9 n�cVGZW�C�P�� a)����(Z(Ӊ@�)-(%�
Bz��Aq0�p� *x�`��k�j]��@�+��ñ�� bg����Z�~q���6|8N'f�[�*F�w{Sڞeh4��s��T�79Ś���fS
8�1f�2��	��0c˾�A
k��p1+��B�@|�I�U�;-�r5{��G�|�ȑ$;A����bqy�^��3w�T�K��X����Z�FI�L:9"lS ]�f0��XN�=��Dk/9��Y�C2�o�`�� ����/\�{f&M���FBx���Y�Nb��>/U'��t���W[~�U�����FG��k�A*���y�+5d��v+df����Լ�-��ay�랦&��1�8��Ow9���awS���J^)D#�g�n_Ir伷��:
Cw����|A�q��g'$a-L��g�gs����*��[p�(��
gT|e���>N��z�U7j ��Z��ONiH(�A9��E� �^J���tD�]�I�̬L�h�?�\�Q�H8���-"����n0lK���\���>3�k�/��~�Q�Q\E��� 1� �q��n��2��4�(ʹ��T���!>�b���~��v��$o����K���>ej�hĽ*��pc�wr]����~ a�p��ٞg��F�WVMwlx�]1��q������6b��l���	e�V��S��+$��`W+�y�@��扉�G\�U/<�G���Z�o��J��"�i���p�3\��
[[$0�<FG���S�Q�z.Әu�2K	���7�k�c"��@����N ��0��5 8x���?F��X��P�|H�=iu\����b�NS��Tr%{엹��Ňp�\�]��.+0��_��*��<���c��"o���|����u�q��B��Y�3V)@>��J\�tr�u��Q?u�����'�Pt�SM�c�l/��S{;�S��&{�B�_�;����� z���C�OUS�^�E���TY4?.�(3���Z�AS��U�����F����ټ�u�K����������>��ޚ��`g���:�a�>�����9�����/��c���ĕ��_ծ�hIG��)�������E�c^�!��A�ٯ������!�����T��,ei��>��s�������b?%鳁X`?�dF�e�T�V{0����U��f��,C��wޏ��_���u��}�z���c����i&�+G�,􍆨^�F)�}��Rk�#GF���d�T���ϱV�3�-����aZ^Ah*FU1�� $"�pq�9�Ͻ#�v�ݸp��Y� �&���c���ggP��C��1����}�=����(Ek+ҧ}>�&�e����>NeV�x�3��s魌��75Aҭ�Tr��<o�t��H���� ��`�ߚ-�4ʱԈ�XӲ̻�z¶�OT���������=��j)�1ui$�Ň�jDch�g�(D������ZE���{�5���݁�`�`��5�y�Sn.sf��&t����`C��zp�෇�j>Hqj�#�e�͊Y�^��#o�W��O/b�E� ��#VQ�_��U���x���¢�a�����sU�����{}�E�kd��$t�e��_�P#H7��j��G_*7�Z|Wjrߴ��b�^jj$�\�EF�z0��{����1}$%���|������Y��<݅�uUg=U�Kj����]��AA����K0bj`>��~��>���:;��M���My�ܓ��}L������B�.���B*��r��o��oe���nEf(Q{r�b�2p���K����2��>���-P�#ɶ8LD��\X��e�yY���P1��z�Ayٳ�a�����_���fVg�O�^,;e����d���O�m��ӹ2N�>�4��'蕞�8i�Rc>�)���N�e��֔���g=:�͇�Ĳ�=�ۣi�Z���F�<��!��#P���a����}�~�)K�"�S�����2�4ͪ��	{wɋ�{sv۴J�V���[��#�� �pđ��%����)������O�<y�o?�_�����ӯ8ml�n�]d��fhssL_��8>���:��"4H9��]I�`�Y:e�o� ��)��`�܋/9���^��Φ��@�H��	C���5��~rh���'��Ϊ��E�owv���M�m��N��Ի�v��-L�w����"x�dޱQ}*��y=Mզ�a7�!3D"�Z��f3������,ә���<�@8ۄm$�gʥv�X<�������%/�%z�H���e�]I?�CC�Q����������M�agAVׯ4Yk��O1��JF���ql"H��{����Uxȶ�j����:�[z�����i����O%�洓�F��Ye$٫����~��#d���Pu���ؼ0�g�Ov�"�X���:T�N\']��q��
����YB��:����[�#�Lu�I`�X��7�Â��@�'���,��
7K,>�?�7���>
� o�|�`�����P��8_۝�� c)
�6_$�3>"hˁ����Z�b�5B]�<�':�'����!8����Q��V�.QE8��n����L��#w���z�*s6���+кt����nBO��''Ў�Ou0Ĺ"����g(6E��Y��)N����?�{�:�������0XEv ��3��+�@�*��O5c�S?�|U�Hx�+���X�<]�

��M��&7�Tl�	O9 )��zϫ�h�4殬:>���,D�}�1M�����>`1Ȥ7l��@�;6e��d���p�:-e�,Aj8�
ȥ�4�����:�\�#̟oj�MUc�,���\L���]���JK)�8gq
�1����2�O�a3����V2L�y (m��߃�o���Yڤ��~�V�ʖ/�1��߁"��ʌ����N��x�3�!փ5�g�tG[a�O�)�x���S�f��{T��L����]�T���D�,Ez]�s��<���pH��i#��b7���!�r��Rץ��mQ�ȸ-`���� ?'9�������Zp�<P��@~��>�O�R��`$g��{tF ����[��aT�`*e�3�6��$P{�T��W�DJ C3��4���4����`�mX��0�S��{�dM�&����`��D���Xf<xP��ëp���{4�]�ֆb7��#��V��>�����0����'�˫H���[��FGK����{�g�kYGVe�J�=��7���B��%�-58Z���1aM�F��8��])!����4��Y	�:ӓR�#pp�cM O}H��k�(H<�(�I�l�5ElQ_�Q�X�ٶ/R�)�$��-�	�������k\R�ʐ�@�Դ#~h�~خ����}:�g%�T�r��JE��2/�q܈HK�Û�j�X$�A$X�Σ��+L��%4�߀:c��l��ȍ��?9}A�w��qJ�~{���Èd9o�V')ը$��3	�6��X��EJn��û�5�
�2��c�R��_>s)���'N�����Ra�۳�]L����2�B���aZ���W�y/m�k:���_����Sl��D����$�R%3�22����IV�h�B��퍾�"����x��{�F�h,wõ��C�����n��Ǉg^���<\��|D@!m4�S�ʢ�I��g���:��-_���p�)�rK����}_��
�,���BRc������l�u��tV����Ay�>�Tu��{��{��6,\����3Ğ�4l/`�'c��=�r[l=e����ɰOW�p�Ws�e�.+��3�,�o��Y���+[��:`l�H�5h�\��\F�Y�lgb���ɝ;�W�b�
�`/&Z�� l�k&Qa���`N����~݁D��t[���=�0Y�E�e(GY�.��R��M]b7����Ty��=ǳXmݒh�FȒ��`p��� ϿZ\<����zvT�͇����a�|�ǔ��?���:w�a�X��Q�/�q�h]Q�$��lr&�9�t��k5>��i2'��-�Qy�"�1�Ю5<�1t�w)���Ļ�?UM�~H@�|�|���?$�O�q6!K�~��%����k
_�_#����F"�ExHNraA������@���4��v����U��^����G�ߞ�2|��09j"�0сձK�����N���5�'On��	��1�y���j�%��髸ȓ2"�^�[���oU�i�o��޵�_�8���4�,"�C���@�k��N�K����<\���R��%_�^�V-\�[�,:N*��BYCg�j����0& `�*6���.T�\ʘ|T&����~�kY1���l�̏����0@z��-ք�R
 }�/f�vcU}M��鮌
0����>�������jX���M�6���p\nG�����̎
%n���*���$.��ş	Lw5���\��>�rG:���`����x5�4{�s�y�8��ޮ́���Nzq��st�T �#�V|�JR�T�.j�pS�����������8�!���eP�Q���3rd�9}8`���Ԥ��!Aa�ۋ;�Ͳ®��d�Xs=h�s����`h_�%N���O@l�Q����V���u"��7�̮��aQ�n pr��!8��)Z�)��t��Z� ��m�����ǻ/m��gk��V��[$�W��R_f���~��r�ɭj?2��gIF�K��O�x��K�ŭ!8m�-]G��S��c�	֧��܊���n����ɣ��U��0Yn�zu�&���YF�9oAL��з|���Q��|t�x/����vg���S�<��a�z�k�"�@^����*YD1�+�� �7%�6�D�C}��?lql�i@�CDM��)[�s�q?�֐�?�rȝ=h#o�]��|�Q�#Ny�<E5�{_`�)��T�~�~�����D�m_�e���̓x���Qg���n��8ԔRЪ��E��H�ҩ�c���s|VI����_�~I@���A-n�+�_x�� ؉?�ճ��H�9�����j��Xn�����f�aF������/�F~�ؑ�Ff$h@��AiN���%Y@-	��N�G�+�rXܘT�����u�7��C�Q�ؙ4�0����t�?�";w�^��pWy��X�ǻ�#���/��0�H�^m��dN���m� �������) ��n��a����<��a`�����b	m��P!)�!�������Q,�?������a��'����b�	��� p�E��c:���EC0�=u$��[/W
g�YJ�����G�D�Q����~�����~P�{�8ErR������ �O` !@8*�~Z�/�%�Y�X���gU��,X�5��|J�w�_z1G�]Yܨw�
:�"��v߼��JS!C)��nJ�n����]B�a��zZ4�2��>X�)�f#ׇ�M��0���^}�T�t�3:��y>Mf鴺z��آ����x
��#w5�)l ��V�E��Ø6��[��@z�řQZ�f�����I����g�;|�����	���L$ys>�����ݛ:�&��қ��'U�ƀ����M�X#gOw��z�ʟ���Du�ʇ%��6$�^�s��m��dN��A��c\RZf��''�9��uo��0U7�ᤨ8�凒ީk+�(Ҿ{�㲶|�	������;�b,zoW.����Cà�½�����}��o�M�0*b<"j6R�L�� 0��L,�}���b��⮕����M;����L���ǀA�`��<�*�k]��>zk���!�ʎE*�`=��&���k�XN`�%�1�V�en��&Ǚ��[%�uF���`Qv��@����*���/7�T)$�ߒRHz�o���%}z|�ܱ�!���W��ޘCT�<��R�O�u5����n��Hv1���¬�Q��&���N_���b;�|с��wVS�e��k��{�^�ꧥ��fi���JNA���j���x[��cE�	*Z�|�tZ�d�
����tir�F0��n���ڃ��T���f�D�"O�Y�6K�7��X���Ls����u�h/�1ֶ�����%��g��o_E���l��)��5�Z�����"�<_@�E�ޜF��Z�|��e|�l;�h�2G�S��t398�yƼ(��%��hZn�j�*�<�r��V�ɳ�Ǽ@���	�'�ٸ��9cW`s��t�*��E�u��M�����[B�E����TIo��W֪�TT'���6|>�G ����Ġ�*+)@E�)��bƆ��������_���*��6i��s/J��><�d�,�F���f�/`b�Y_�=��1�l�f'���C@��j��&�+��X���%�ޓ�	v�7�:���w%�xV(����Fȳ�4�Tp��0�	C���e���G��&d������� �v��u�7��k4�7uԄ����.dȐZ[��V�J�z�ꎈ$�]��@q�o�b��9����/{�@�2:��rަ�ǯ�;֜����K
y��Е;�%|s�D�t�H'�i`��[ҽ��N�6n�Pյ���Z.�q]�Z_�PU�	�˧������{�`���7�o&�BM=�o��� z������'h�z�O�s�A��/ďH���I���m���>�IC�)2q����?�B�@��k��q7�s�͢�ku��y��¯�UV�1����7���G;"HAӻ�,HR5��Q��Omo/�j���2&WĹ�Ti	�g��]���id!O��y������る�

C�R�'Ҷ@wP#f=S7,�Ic��}苩�^��n����m�Q��%O�@��p��?ssWXa)�J���d<�����}>l�*x"6beH%3Z�w4��m��,
��� ��hh\��A�xN͐!����I�Pe{���(Z���	�9>���S4vH�g9��4����A<8Z3Sش�~����y�Q<�A�]��<˨�ƻ]ۃ�'&��CI�x��/뉀ϐ'l���&K��% ���| O�