��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ���L����ѳJ���ף�6I	��7�"�D�}ے-��KpV��s�h�n]��[��;,��*��_�H1mTu�<'�M� ����Z�H�H�#����*ծ���p����*�R@�>���Vx�Cl/_G�b)�z)���e5��=")D9d��R�d0�� x��Ġ	\�{���> �Ueڼ{�g�_ˡ����T�x�\mB��޿8x][������v�	1)�X}� E�� �_ð[#�b�$Xt��C�
w��bGe���ʹ����UG٣�ɹ�~V��e"ѦΙo�ɱ���0�-�y�v��CPܼ�Fڀ�2@�E\1l�GN��Ϣ l�iRP'�ϙ����Y������ T�*�g���DO��� f1v�\�w������Z�2���8.�QV,���W��K��� *�,�J�6��jH�;�B�n]��CKxv���R�i-IJK�vC�?K$�Q�Ai�L�����I��L1�Cɂ��[�������x�9ئF��ty/Y��Tdto�	�^�S���/C'iy��^�,��)�:��K,϶>�e4��D��#��#�a��ÉB��� m2���pv �Ah���q�ݩ#��?-����A�1	�)W"�"Q�T�y��]�,�V��~���zZtˑE�qv��C������+	�i�����Kc����|���F���o�|B5Q�L�ν�!������q�"��?����z���AL8����B��<�x4|��<I�*��m�}��E�r{���K�B
�8� ��p�P�ĥ��X���@;;%lcKrʓE���Xȉ+A�|�7q���vI+@���dK�K���.B!xW�����4��P\�T"�8O��y��_�e�dY2ε��(y��O~�@�{�*�0�c T1s/���qtN_��E�.�p^z�����+��~���>j4�ф�����ا-P�,ӣGB#2�JY�N��ں�ő� �a;FX���̤���αMrd��$�6YQ1��IbX�gڻ��Y�c�~�R!���]��g�<#�)�jQ�_6�YΜ�@=8Ջ7+Gp?��WPb�{�Z�ף����Ȥ:�?�{�d��o��d. �c6�dTp��G�o��v�u}R��5j�h3ܚ�4'�Wn�O�� �8���%��������5dag5�g)G8*O>�=��/YO>n�,ɠwꩊ�Jx���!S��u�Ξ��gV�����o9%���sv�g��*8M�y��j�w��,�W컟�4��\u0�1S����*"�W�p�,=�V���qh�FX�a�����Kj׍�x�Н?Clz/[>��z���C��6�
1������BO��1�p�b���dO��y���*,�w�Nc���/�nH��ۍ�ώ�.���kNm��cx��Yf�u�@��c��O�O�7@� ����X��m�[%���@h�˼�����)E�Hڬb�pn(3cp��"T�i҂�B�ڍܯ�'�c�6GyWFy�V�.҄u8�D�5�b�:e�G�JV���᷏�e51�l���T�)��[1�[}�I ��gӨ5�w�զq��8k>�c�u�rT�Y�_��`���b�	x��M�5��e	����&�����i��k���1T���l�y�B�q��<۲qoV�4)v�^�B:��p��CY6�h�c���|4�2�j(��²?�$���t]�E��?�p��: �޹����Z_���`_�!:�=	� ��H 듞�Dc\���3Y끞����N�`e�|�u�?�i�����%���� >�����M��PE'���W���=F��i	��F{K�޾�w/@�Cw����'��0����|��Kh��ٙ/-�����}]�&΢�P��J�K�	1��`�W�������CtТ��4Z�֏^d�E��N�ޤ���� ���ٝ�(�>���~P�&H��^_��y���K|���J�b�?C��_������^)���<�G�.�k��G�D�����TNu=*��>�����W���NX��:^?���3e�2��[�.��$��@v��C��xb��J=}�.*E�6 r��S����<12���z���&�H����)�[��j6
r�'Ì���3�� �E���-a_�_&;���*I��,�G�����~͙M��pV7�\��rt�E;s�d����,���b<NgC�x$�Ud|���6�������h�#`H�?�X���+`u�O2�B��k~[��[����{�0u{�5@i����Ȫ>�׭�+\�d�)�������V3�5Sޏ�cpo��b�&}�f�IY�:K����uP���߃"����
�Ir��)�\�D���bOOQp�m��\������ߴ#�I����@�Jq��{�3H:ԩ�-E�lT��`U�|qV�J��!ج�R���u����ba/pu���B���N<e���tC��4r'V�؋7�1Ǐ�^Q3��٣��'܎
�g^�K�ݑ\.p񗵛����D���?�xh!-�"�'����+�3iD�p��ü��Ń~9�)�b�e3�kR�2�U^���{�������ۣ��u�[�����3��5�^�Co�;��SzL���*\�pV�l8�Pr��U�Gͫ������h�A%��L%�j� 5u3�˄S[0��ѓsAw�l���wc��O�odgr�e]��'$��#U�9���� ?x���o����xY�;��B�8��lպ*��Xq�;df	�$`�d��S����r���`�����)� �7u-�J��s�F���Ce��Rg�=�2�gE�A\BU����x4 ^��a���`��p3�C|ST�@�]})o|Dӕ�<+�#-�J������{���c�U��)*~�kw�a8���P#}��h9X�Ʀ�������Q�Ea��f&>����d��}���3����^�ԟ� �^+��O\�܍3A@|\r���՛�#��Ǩ����l��,K�#
a�	�X!(֋��.*T�����Em&Q��2~��!��M�"R�a��Vz!�=(Se(�b�n]F:���1N[�w�֭�e@2�;��
gR�UG�Ϳ�|\�W�mhIK�]��/�%����%�x�u]<���&�v��\F�cg��26�+&�'l!:5�Q�X��کM�~�bD���a��\�v/��~Oؼ?s*p�S�
+�e��GD�Ȉ`Uc�X��>��i/�u���dV���;�x�<[�6�+?y�s�cqC��&��Y��<���]��j����N����e<�?BԌL�?�7���?uMm9��:e�N�����	�	ƞ'������YΠ�z��;��w���A�L	����@dg\��Z�<k#���GRX�X����y�^�}�;Q�Dje�XB����xM�H}���c${Lߡ�0,�T�����'����`���F�x���䜓���}��O�t��Z@��B��¡��`7t*�&I�M��4.a����.��,hR׆K�h�os��'��@/�������������k4�0Ѕk^!R񷛑�FGJ��4��s��#(��扝q������fw�����H�5E�i6���k����*�`涶��Wh�����o۲چ�e?��D�@	���t�G&��\�
��<���ɕY�+���P[
ǭ�{$�{���9C��:i�^�9�1e<��=Q_f\�HIX���v
���2���P����g�]h��G�����+!�<?F����qTj�R!N�z�Qf���y�FL��9��?K�a�d�lͫ�xǱ��*c¾�<�k�����`H֨�S�P9�f���~Wg��lE�j�k	i{6���it�>�z�8Q�����Y��*�]�G�W:��=R�H��S��s�ɧVY�	����8У2���0W;q<��"I5��rx�*�..��n�шh�
qk��.�ՏK&p����6��Z"/�@�Ւ�˷]18�Em<$�"N�L���9E�Jv�4`o���G�f��i�am��`_<F�5��?�)x���R��BO��+<�`��޳�6Ȑ���7[�����ϓ�эT<0��.٤h��-��TI�leIQTjk2!�g���L�ɳm�k�����&B�h}A�ܱ��J��z'x�6�5�k���:�\�ћ�,�车`��BfA.�s��HY)����RJʴ�Z;��4�w�xa�'�V�H���.���|H����9
G��������q}������+�ڻ�m������]�_{SD���9��u��dx���XOQ���M�q�:n�lӕ^�w�GT�h����<R��ԉ�'MG�V�vZ�?8�Xw<�@~��=�O`��--���:?��(ܫSr��a@���vu,���%�E�lFﬔ/B�4�卐��(�w���U#�Hg��8
�)���;d9ߋ�5�kWm�Z��ڞ��\�d�P�3e��\�us0����Oh���k77�K8����(�%�W��El'�8��TM�����T�ܬ��=���@6yK�O""˾E�.YGP~�_>�i�ذ*�-5b^@{*�r �)P#�tO��G�\��	{��:��ݽ|O�Nʏ����E�!�h�w�g�� (�C�Z��;o�D��JK=�Qվ�������9����P$�.V����Ց��{T"9��j{61�+m����`0�(%�\U���<
�mC�~�g텡k����,��Ȇ0Y9EH����r��w�ls@^V��?��Q��]*��X�D�9�֚�Ʒd_ ���)8>8� T&q(��M0u�Ya�ƈ�ȁq�K�����&�V帞J��SR��)}�x>!Ʋ\��/�1�;J��L��E`�� 
lu��#�����i(�b[=:(��so��-�G%�V4����vf�K6���\Bÿ�v�����Mo�1��gsΜ�X�����軵��B�����ɣ���n��+�S�GU��
�ݭ�� aA�)�m}q8S���+7��Φ�G��C{���zO-2dj��"fƄD�<@ʗ��M��2-��XG@j�&���2F:�9_`PR핊��6@\�d��AX,��+ߠ�WZ9�f?��>���\v3�`�s��8���s}���#�cy�t�;�0����@ǿw�\Z���Hx����>asx�.SE�����ʋ�1�?��YT����r�)�˙�q��@@d���[ӥ��@A�dW[���B!�<�M�NI��dq�A���p�d:���|�a>�f��i��8��1�2e��E�Vc-�L�!8\��2���l�Q����ܡ��JW��-�":t��jx��D%��M��x֪n����W�Rri^{��G������V�w��X�	�9�G�o��浧�BBy0���D��fG`��;��[Q�ǉ�Į���C�{㊫�f��=7��%�栻���g�DI�$b�8EU�L�2��n��,��(ٰ)N�V���paQ�$I�*����z��Ѣ��~�+��YB��%�,hL]��!�q�����a�4 P�.$X�⢩rҧ�?�m<�μ�7Ls�s��q:G�9�^[��S���(����c��y�6���d��ſ��\9��w8��Ҋ�u���32Dȇuo�x��h��'���+%K��6��������f�&�\�(����C�}���}~�A��]R�<���̫y�C�Z1\w�ޅցS_aq7c��D�!��s
1�y��"���FN||���Z#D�E'�З��'��/����Dc�b�5��E�"A�K�S����ߥ3]õ�O���>�w��T��-��F�Fʫ��Bi�-��EVF�+�ϖ��F�.�W�97Fp�g+��� e5�y��2NN*$Wj��TpaG���S5ڸ��V߈�u���o������&��6|���)y������$�2��W�E+��>��[�G��+��7(�1���6a�Y��d�Ѵ�-�| ��ν�*8��P��3�̴����\�{9P�vC�Y��R����f�L��L.�Ś\�s��A�ѻ�67
��^}�����R?ʋ-�C ���j�+��:r.*�GN�hǩ��u��*ӪtE�����c��(ۍ�R|�r���?y�nV��+�3 #t������=7B�5uL�eZ���}l1E��{�K>ڜ��`�Y"�0nO��=�,O��yPe��
4�ꇹv���X�cHR����F�0���aݣ�i�+�G8f$\�N�D��5��>�$T{r�xy�Ģ���E�vt6����	ۼ��M��&z~�\�
�`��r��U��q7�"�{��1dh�Z����塢\���r!��ܢ����nv�
������7c4y���8�?��o:��Mϸ��h�+�iWN�%�� ��E�g���c�4��Qj3��Q}mc{i$;'��*���`y�5��xx�5I��գLw1n��Pv�Bр���;�}���,�0r\S�v��Kf��X=��Ƞ[���!�O#��.Z���}��;h$���ņ?�W�El��f��;�XU�&�
�����Ci�u�aƵ���$��ڔ�/X������3G����	�UDf+���i�z}���dI���W����,mO�
����$�)�kF�TS-�>�b-�7#Q'�Ab���(vGK @����'�|��%A.�(2 �W�a6
w�!rHF��F�gJ�f1+(�O$�L,��ɠW�EU�{���ʹF���w��[�>:�'��:V@�8H��n�O�K�q�݂Dr\"mu?�Y�\�-A`�In����変�Sl�Ôi���b���\�=#��!��V�t�����i�3|�M�����GiԶң�֝Mt�������cz!���s�%�}�����j����s��]��f������ Ė�İ�[zMS0�o�}y2JwJ�S=���1s�V�m�c|�.�}�-y�<���`��������p�|��jK}��w��;j�'�r�����Pu��D�UB��H���9��a�p9f�gڔ�꛰��W[��x/�� +,0�ޫ�kS�z�� d�
�k�Q��сI�~iR]s��,S&%���.cu1{-�b�~��t�0� �D^̜�ΐ��h��~F�'�Т>��`�������Lk	I��Qτ��)2e+5�R�L�x��n��h��'9Iw�=߰,6��w��������b��ԃr9q([E�
^ۛ/J��N��$������+0,6^H�2,i�}Xe]IpˢΚZ�	�)�h9%dN�a�l7n@�~;��,L�7QD��#n�zvx��^WiH���G���E͋˹V����V$�d�2��1��F�ѳ��5HXjzTKY�=[L_%�;�(T�(��"%'�ڧ(~�)r�p�괖�7�w9}��a0[[�eG�mЈ�;��^��]�Ժ���{Q��.i����z�=D���0�B�������1)KY��?�Ƹ���(�ma/�-��;�շ)�^�J��?Úi�)�e*��R��{j3h��V�����.b�oގɝ[��%z�g�#��qͿ�E��M)
f{�EA��-ky(,>�j4a���F�n��)bY����� Y�g�>�2��Q�~L�旒�[11Rt�@' ��H�Y��j'(����kҮp|�ӊ~;���m���M�:n>G`%������>:�
��~*���T��l>�;y
���}�4��a��Xtt��m�^��;+��!����w��+��Uږ�]�1r���B��e[�=��xQ�t�6��?o�ۀȯ��!�Ƙd}ݵ������h���&U�a+��N}�/rXm�Y���a���oX`p6oF��
��������s�����=tL��d
s���6�D�tw��T� ��X:�ک�@m���z�k1�+u�Z�?� ��ߖ+�kw�yzS$+�?���|PhuF�������~-ʟ���������%��Kj(������׀{[�?ۖ�у�z�&6� lC+�*��|U���M8�[48p0��pÊ��K�H��{�́�>���@����j�����8�-�]����i��@_����j�.�&`�$��7P6�r��ͽ�͘��' {�`��yp*��9��������l�{�{�!�H�Q`4���ڨ��@;���^�@�ކ�ʋټ%�!���w�a�џ���/X�n�#��N���%�'�7V��8����������Bo2Ԁ�_��Qs�6�#����or�g�ew������~9�埅 Km����i�7�^4�Jgo\���7?���d��"t'�NS1,T�GVJ[L�V2�$��Ym������_қu:�d�k�x���&9jC�C"JZ&'	��y�	�9�A�C��Ҏ����N�`Y�9іp��*S��
R�t����i�G����'�Z���\#��md��6��8c9 �=�[J�x�&�r�TI2z��V�����erm]w��=0�*���O}��0������+�tҚ��1{/����k�:��0~a'�Rj�bG�84���i�P���`��=J6��-�����+��ԧ3_��#�R@]���癛()���I����;i�1���,�����Ր������I� ��$���m� $��|�E ��Y�����r��Us��P+�v����ҷ.ЈrX�D&�����H�t�k�E��]9��t��&{Af��Z��UP>ĭM7�|��?X����;��Ԫ��S\!��#����w����X� ˷L���燱�p.l�lN,r����j$�B�-S�j�M�r|��=�-���0#�����%`�E�V2��¼;�Z���zR/�3|�M����?�%�Ы.���r��ލ)�=J�~��o��q���%��r�ԏ�
���&�_�N�{�<�e�����l��uo�M�����4��W��G{��wv��d�t�{��ߑ��t�\�ґ���+pKr�o5���	Z���D���sM&w悔��ā�%�? \
<@������/Y5}8⣟8k��T��d~^�`�٨����}��ʚ����ϸ��ڰ��=�C��QK=�޵)��z ��V�`^Q�,6��E��ۖvP�+��ֿ�@�MަU�Z��OY,�i�$���:9Z^�q4l��젙$�m��"��M�z*�L%��'b�1��NC�I�>�lR�@9BX�Ŀ�18L��B������=_S!��V�Y^3H�1�o�&▟QÄs�(U{���cI/�<�Zq.n��^�+��yE����(`Bc7�F%�k�8�e���_Yڮ��5�"09����B�O�c�p��i�u��鐓�m��ˠ"'�L�4�Ȣ�!(0	�)��x�m������Gd���> %��g$�`(���qU�m!G��F�_b�V*/%�.*�!� �C 1�K$H�nD��T���9l��-K[6�骵�t!���ْӑ��7sR~ q"3c��`��U�m[j��Vxj2)�j<uiv���YO�H��p+ke�$�f��
���D͈�=���һ+b9&���"KY��w��4��s�UO�*�4RH��<�0��٭���]Q�'ȽpRU���Ȟr�Hw{H�\����5���엹h���@R��L!��Ng���ܯy����1K��T6����k��\�q��nU!�STZS��T�@�G�}|g�b�#(\���`�_����������
�����Zo��C|$�S�3~h��	է��k�)�N�TF�pR�5��BYcH����I�w�]�>�G���[N6������XJĊb��Q׹[2,�@��㞘Ex���lq6����pm��N�SNXo����@�ye��u晣5�,&ԃv�?���Y���~�uģ���|��(�ՎR�)5�L𥐄�����Hd�K�m�#?�kO2R�qfm�k��c�]�,��ZD��K��d���h�l%�{�����ŢN���4�Ί{���P�Z����[ﲋv����nf�9^f$Jb{�	Sr d�&m_)�ɵL{R�M��~G�~eje�������a=��
����$����|S�.���Qw�ab&�ǣ��X���۾�F0�.,P�~o���1H������{z=���]Os������ꅥ�۷�f�;�uv��j����Wg6�����%J����K������f�P
����:�*Kͩ-��oWJ���C���z��/�Z]dt�u�y|�d���S���j�h�Tn�'�B��d��)����R��V���X�c���{=�Z!c�N\p��`�|x�A(�rbm����d	��;�ej" �^)���	W��� �u:��|���О�B$9zgN�>���9��+9���-W�����0�1�����Kʚı�2�垺�iKX�W`�Aj��^u�>���E:J1;��8V:�t�.���ä�ǈH�H�yV�m��u�99GM��<�I���ңM^�0�)� ��M�d���P�mPp4]+
�/t�����D�M���FV�2��Wp����lN(��J)�CQ+��7� ��|.a<`י�1Di��Ǧ�w��5?�*��^�T](�M����].��F�,�ubH�������}sK2�n	<�� '�QZ+���ի���9����!z�FዎM��Q��Z��,�ƃj�;��n;���Ԁ*�����Q)d;�r��o�3HS���Ґ֜���e�����4���;&�|�ʹ�9�-e�� �`�< /zl<��": 't�!�\����8UB�^c��4���P<I�f����m�"�7��j��[Db�Z����&'B{��S�۳Xg�PI�V�6?��as���t�W#�|���v���$v#��K8������~�����eP՘���c*����pf�o��׺����];tA}w�a)6K�gW�a�Z��|c��F�ۅ��"�
��նa�÷�a��G8��5ܷԼ�6���y�椕��s����6gz��C�+S��m����Y2թ���L�t16(9K��@a��|��vA���(�$��O�*[FӢ�t���v��6�E/�Ĩ����� ����I�-�F�èTۙܛH��`��FčBIX3��
�n,�˝O^�L� �z��`9]�����w^�Y?0��l(̎�uR	���h�z#YD��'�7���̛��q������܈����o���$�8a�q�`,;��Ɣ�%1�b"���2S��� 8��#z���
�΋���t&�v���K�F4�b���M�M��m��{��fb���߫z�yg/t��M���5m0��E 7Ӷ:�R�p�褁[���y��*�\��wks�h��8c��Kd���P�<�_�Z��,`�c=P=
�qwG�����&��}��&�	�5^sP�Jf�x�ui�;I���}����ϴ:�u��?]�!�%~ y��N��d��7a����Žg�{�z�����"���E͸*���"s�2�ܟx>J�N�Qgv�$*~n8��/0��AeT�%x,�_Y��AcJ)�t�*��>���>��C�aM�h����vϳ�uQnWW^Z&s��J0��bF��]B�\�Ǿ{��N��F�"� ���a��mx�^&I�e��������4�A��6�U֋��os�~��7
�!g�]��8�� h,�DJ%�kcvH9O�����a����+�[�G^�kV�r��Y�hύ���S*^*�D-���o�>`�>]b�	�f�,ű/�t���ěI_�!8%������e�nk�pN�����kAI�=!���*X�`�yp٭�
��%ْ�`�� ͒T\��(�u&u���t����i2O��џp���>�WO���Z��2���H�ཨ% �?�R��W �����2����v���7+s9$��@S�w
r���4n�ʅ|����Si&n��N�����?���jE�B���.Y������|C�8�Rw)����î�AJI���j_:[Ž٨{<���U1���yʖ���L�K��/ɓy�һ������V.Ӂk���
-�hF��*ֵ�y? �i�w@Ls����Q�ɖ�uv�/�r`�{���Fdn��g�	����)?͆H��`o{u�sph���J*e�o�ة�zW�Q��(���8/��^J�%M�&IO\�f�Z�8�@ǅ.��4�B��uR�N�$��1A{Q>�9�C�~%�$�IK��P�`%U67!:�,��|Y���N��e6
���Bk.̍D����8�V`i=��qn)ѱOB~�+e�l���l�r�v����l�cU��2��Xm��
�o��i�����C�&��nv?J���񀻻���@��X[�:-�4g*���G��g�P�Ej���P��`w|m�����)_�53o�(5��v�ioXL���<�5�9SaR����t�����y�H��pVQ+�oI��F�4�?d��J�Y@
(�'�w��LAPxrܜoHE��EMf����{� �z���8�xfi���d�b�ضǇ� ��?#i'~��`�b��Ӏx���5�^9�#��"�	����y�*�t_�q���-�����7O����
aē�����E��W�)fש�C��ǹ���nCcݢ�0�A�b�^���mPO/$ЃE�Ta7Z�� ���@�II=Rd�ʎ�\Z��wy���Z��dK�փ1P��G��ĳ:tI��ǟ���:�Ҫ����u�	����|�xW]v�!�%;���k�K ��HwwC�VHj�;�-�X�.n�j={���0��\~�P�E�qaٸs%j&�qaT���|���,
���?|��眱��ɢ�ڌ�"���e3���|\m6��fӤ�K��A0b�
F#TfP)��6<^�U5O��`,���?��	M��i'���eК�6���2�r����G�Ư�]���Q=��y���$��A08��yU��i���1�q�_䛨?��@ǟED��a:
�+9��U�䲹I�Q��wE���G;H�0c�s�(]�1�)�{m��o�BD��^���G@|1���D(~�՟��kB�o�JЎ��1x��`��W���G܊�,A���	�S��+L�tT!F&��s�/W��a�.��I}����7X�5Zm:�c�>��`��u��ۇZ�K���S��k�;a�l/$�K,ꞓ������3��+��ݿ:0�&XoA�(�M��\�O��>�>]�w�WX9ڤ�b�{v7����I��@k�H�F6��>���E&��q�q�ٍ�$Ì����\���i����.:u~٘uʇ2t�e�
�`�~�y�M�"8���e.���o�:�f�=9몄Y*���s��]�Ǐ+�Sz����2��̽0�����.����H-�q��Q��f�V:;;�u `D,v�^�c�\�%*K*��j�qSw�lDfB���v$WǥX>�����6Va��H���3W1��ZάH^D������ec̄���9�ʬ�V��aO�Z��ЂI�VT
xX��,+��Q��Bu�c�~����{���&^�F���0	,�﷤/	څ��{C�^N������q�2�E�Cy���"��ද/�9ZP q��IÏ}�iL�>�|������x�)�pl�;�#le���Kߐ��2��JZ��3�P#�j���{mq)z��W:��5e�L��܈�+��-�� "�%��A}r���A�(��:��]�������ZZ3���4��X��/C��2��B�<����P�p�����c~#$\HJ�5���L#
	��h�[���{�A����J����%�c���ӌ%��$�0�ۯxTGK5S�� u��QLI�(���ar6�Ѕ��dNM6Х孼K�N:2�w���\ޒ>�UO��<�]^�����m@���6�>7~t˭I�m-�vކ�A�G�Fq֢fR�7��{+]��x^�-��f ���Bp},��;J�����q$�Y2���;pm�_V�B'/�xc��c:{eV�B):3E�>��e��*`T'(j��Af1l�M�N/���QOy��zP���:Cؓ�E��b+���᳚���֩�=C�g;B��Z���YْC��؅	T,�����~�����/=�ߓ�� �V�k��"h���cIݤ�es���"�~ƃ��;�♽r�Ь�[�2�r�Ih���iÉ�����z'��1\
��z_i[��[�������e������v���~A��71�Q�g+���sq�_{u�+���@d�H�hכ��U�(�_㓺 jU̖u�G��<��y�9L�e��#���E��9��9�,l@�>�蒕A<y'
��U��_�*�y�Y���CS}�n!�����ʟ"�+�2��V���E_�=�k�֯b}9���'���*���C�Vy6��3�k����z�H���Vm��u#8/��"��S��t�)�7ܽ��Y}�ꕽ�t�/�Ɓ4 �ҁ�<�$(��,�ܔ M��*����^�*�A�����ߔx�vw�`ֿ�:���ue:M���CVb �N!�Y,���\�Yp�>>�浜\r��g$���BO<���z��Έqs4>4��%/&<�m'�^�ڋRV�}D�XT2�Ky��C�w�2+S����Q?_��V�a�θ�,�G��魷ic��[i��g��労�ނ���+�;2B`�n���[���+j����x'vs���r�R��k�6��.x��3śY�/�r��g�9��hTfuG6���/�|��������D�q��cL�'�@&/>u��Ft�ǉ��)ŪE����������ӽ�IXDe�ɩ�J#5��j��
�Q/l��w�*�/qTVU�Ίe͛�% R�>J?:FfO�JUVq�'��.rL��'y.�5��u��wҘy�|BE;ۇ
��Bw�Seg��1'�X�/�ע4s�*V*W�T� 0�5/��#���d��[\�i�	���fT55�T�tuU�]i;��!��.;���8X�ȩC�U�x���K�8�������,e��C���e��h������w�!|�VW�sY�����u�	�;9��KD��1%P \�[�n��y7�����a:7�I�'<���r��-�)�#P���p�v�2H�>m=�Iu�k��`L[�N���'�`i����lO2o���ob]@��p`�a.�����eըϖ�)#K@3;l�o4������R�$�}tK��L�i65�D��Mh�4����I���e���`S2n�`��^�a���_�^ஶG������sI�z�s�bem[�K���@�h'��`#ABy^B��̥V�~o[���j�k���$�z?>��I��U~9��˂��ip_��%��5��8�g��XO>�����7��������U��'P\�:�N��_�@Nb�a�R��E�J����B������Q�g~ڿz��&�!/cf*��/���|S��O痊��3�� �f�U�vm�m�����樖
x�Q?��Nۨs���=��n�v�䭭���!-��"��O ���3�Va�w�y��c�S84)X��KS�QT6Ϛچuɬ]�$��KХH��2�_q�}���t�5����k��4}�40�L<i�Rكv�&�i1�m񌖒�O�a�nT{ߛ�ύGV��>��NS2���M\}�qqC�T���f�ˈ��Ȼb�$�fS�(yS�)r�d#('NT2�h<E'����E%�5�RMy�"fci	�����#BQ���>p�M�t��\�Y����5���h��
	��pu�u��r��9l�D��ʞ�Xl!�P��ڂ`��֎�n>T4����\V)��`��������꾩�,/J̵O(��A��ɚ
pl,��$�!���{�x|��0g�� ~�x�\r��a)�3���d��I�U+Q��e�O��*��OQ�/���[:�uB�Z���!�8@��k����(79�!Q���E*P�0��Z��$C��� ����:<��HۥE�h!<�G��� ���nq-�q�� Uy�� ��G#
�{��+�C��O�-��O��Y�0D���	��R��'g����xb�m_z���v�g��ܿA2�!���t�\('1/ ��C�����%�y�&7z]���\��4��S�c� 0��v�ĘOA;�)�/F�}�z������I��9f�>WJ7���$�U�4�a(�����@��E�Z�n��=����S�	M�L�=��Q����#���{�:eruf���AJt!5�0�ù]�O�p~*�b���K��r�Ce^+��d>�-t9(p!����-�|9��@�l���0t9��%(Nkv���LBaf6�KAR�ꬉl��<?gZ��&W�E<������� �/(vA�����CB�6kTcs���%j*uD�F�wKn�)?��v��8K�ZėĔ���
	�B��cA����2�ANz�6�I����|	��"�F^�?#��{����6N6���z$\oq��/���C��\KĘ�714o���34A�R6]���"��:-W�
����p����RoA������tav4bhk��������#��C��4�{ͩ�T��nH��@�/�{��$ (���_~��[w��o�}HH�`��8U�#a�b��p�E�\�~��jٸ�k)v��ϐ�E5 u�/7ک$l@ �N�]dT��06M{���#d�
��6�ӕ���r)�K�p	�P,z�=_qFvD��m�x`���0���)f�&Lv��~�]��:���jx���slcO���V���]@�������7���u�p�7,��e��i�%��^������_������PH��}��;&Z�bi��"�6笓1�E�Ԕ`զ�3�B�Hr�T�6�ީ��yX�9
��l;:w�B'��v"|����g�Yb��b��w�%�*�����@�.�w�� �� ~*�o(�q,'�L1$ű�\�����r�f�Z��!���j��F�6��GQ�0$T����2�2���b��7�4�\����˄���}�Ľ� .n�/���'����7!�cd�./�F)�!��y,�ųcY(��.W�ݲ�vWu��V<+����w2��L_`� ��Nk"�u��R+	c��$y"UZ�y"�n}�Ė���Td��Br忠kj�&���	�� ��vs��B��o�X*޴�R�S	���Iv���a���˗�jJ�����J�����e�4I_��'W/.EO�3��1�@������#�Lst��R����p��M����ؚ1�Q�3��{Qi7�= ������3<�&}���z$�W+-A�6���[Kѽ������#����+��Y��0Bd�.}�ٯ��K�d&��{h?YլU��w¦X3���l�RBE奱��HXB�R'�ч������������� �Ht?���r����O���i�JCM�@��ϴ�]�2kg���-v:ǩAEg #`
ng�YLq�Vw��XLE�� �Ӎ�_v��X��M�kR��@C��T���֙�����S�<�ǙX�i2m��(���,%V3w��/�Z���b�����2�{�ȹ��.����]k��L�̍��}�ˮ{��GCL�֣�u& E��QK/�>���-�aD��sh�w��
��FHfH�K�.0R��mdES�_�E�7w�Yd�1��1�I�7m��#u�k^����L��n��8Mf�!������zu��Y�Z�&K��e�W���0�9���/���wa��BDDס�&P0�����w�\��E�'�6�j�-T�(ၭSpŘ���|yg����|�L`�6�D���Ƥ�/�������T�	��(���d2{����
wt<N�x��?#�����kg�V�~LM���R�ar�qc�6l�Z��!{�?�[�����A�J���ei�X+�<}Y����S)%zIvq94|�83���07?h�J��M����K�f��jY����e}=�c�h��CHJ]��-��	�����#&���=����βYh����Iz
w��TB�gc_]͎�>h+>��&��!Ņ� pxu%R��gwT6�e���:)ϥ>Qt�`�ҽ��lC�|��q*�&3n�nk}��g*d�����`)�­�����8n�s�J[[B�����"��G����K7Ă�]����ULI�,⥍�IƷ��oY��1�"3����4<�c�����ײ�R���<~s��R�$�.qM�jg�u��=�pEt�gV�C�C���ȧ�ZO�
ל�Q*O1�l����ё)иU΢ ~V;�HҤ� �hSY�|���ك[{|8ղ@��G��2�!_ b�:'�d�F��=b'�11UL�Db25��"����Q.e	��x�M���6>�d��\w\��,�x��g?�k$��Z���X���|��AK�}� �a2}���:2����D�~��h�݂΢��GY&�>���r<"Q?�- r��{]:o����r��5��_/�������H���Bx5F���T�݈x�<Tg�J����R��X�-�P_�k��e���D(��o�)D��p꜠
D�z����K���}��~ꖮ��i��J����K��%���tZ�P�~"�3s#�ŀ����D<�s�7��nЗy�O�nx����/�fS<y���A�&��S�O8���E*d!��Y�.�#ኜg� ��/\̖�3����H�1'y,�Py�����wYwa�m�q;C����U�.�!7@����L!B'�06t�
!������FÄ`i!
��T��0y_4�5��?(5����������u�b����1�&3"i��
�nB �1s�O���9$�k���^]#}��6�e�W Ū�HUE�4�h&��41$�8��ɕ������O�a&m��Q�߬eMG�p"ʂm�0�%�4V^e�t���R�l��9u��FC2ҳ�K���t�u���:<�a�{N��{_��Z�C�@8W��eB��gĬ�]ũ�j���ncƈ^�<.����E�C�r�7���k+p�3�H�����.Q��a\� f���t��^�2�鲴��u�.�|"��8=��5䇣J�9�l`��/�n|>�5�.6#i� ��Θ���-MВ\s��te������	  �6%5�A��!"���}W<�s(��Է���	��1;����$H��ēA-�uh����
�8�UX�VK:f(�qj(%��**m
Y[G�KE��>Y岩�+&�ci����K�wس�ϋ��=�p�ל�: e�%'�~}� ���(o�U�k]���O�����r�3������K�_EPL��nuB@�(a+O����0��G���4J���4�-��]��������&�����K���@E��͈�]B���c>�]�Š��*�ѓZ�!��	���4��;nFS��?6HY�Y��3���ݩT���br�fj�c��3E+@5���熠��l�U@)"%��S
t^�|��u�dA@CU�@���X�Q���-���{�_8i�x��LQ�!�	�8���nn�c���2��?�~,*l�"����2������TI0��~�2L��t�`��e_�m�탴\�'fE�=�V2�_�k��:�Z��^@��[�X��]9����i@��S9�*=a�xf��1�[e�efOu������Ѣ�>�q�2a�}M	��z�����K��	m$�.v9�`��H2��C����$��{�o&y̘�£ �gW:��E��&o	� #+����&ޔ��M��;��u�b=-&1��I&Ly����>�/}��}YJ���\̑����3��s�_��r^���=�Ϭ��s����>�	 �Y 8���9D�|�ZM=��	��LɾakD�VP����.Xc��7ȿ�^N�$��Gz�z`�����O�Q���/1C?����yOg	�5jF>�D���/�\�.�ٞ~�n���Ԭ��_-�i�]���?!.u�_�|'���~��_[u�e�ZaϸECF�5q<��S�qC-��X��}�)A���nb���SQ욅q��oeW �u��=��q��[����? _�a����tz;jK�Z�ܶv�R36�v�;M�ό�(,��Eiz���Ϫ��q;�� �s�썪�bFH�������ѹX|��P�mE�`崂��/��ЈA���_�,�˖��
sT�G ��'��21�|�s���s�Q�L��f�=�'�l6��v��g@��,���W7��o��kӡw0�}4v��|�y�%hGG��3V����#��r]ݎN�O5Uz��ƀ�V�)�eA��R��k�4�T�Li���K����F�Jb���7�wgL�wEi�,#O�t�M���(ȟV#�i�f�)���Q����b��j�R��"��Lq��(�ף��L���@l������r��;��g�Ld�_����9K��0N��14I��H��"������ ��ԺbО��au���I�3��ET�G�۫�:�㗁d� ��
G��������_!�ר\n��6pR�}��vTul���[�0��n�?ָo�?��̟ �&�7��ϙ���@�X�Ԫ�0����$0m6���%s��&[�>l[@��D,:�8�u�i�����{c�]��4yR��s�`J���V�(^�w�qR�?,�nԮ�Q���֥�����0Χ1z&���s������f�T�~��,��	��j��^�:-�\��mw	��M��t����eȼ�𷔛��>��/H�/M,NC)�sށc���0p
n'�8�S�.�A���4}�q55���tA�������L��&��h�S����e��VY�H���>P�O�k�����b��Vƶ�I����WS�\!��GX^`�>� ��M�@,�[�\Ɂ�)����(+3Q�;�=H�����?�P2G8A9���Pޛ�}s ���5c��
��+#�%�Lt���?�.>0�%���}�h�zʃ!�zv�Ǹ��3�X
7\��mB
�16�[&��WJ�=4���߯��t:����?�����-��߀�&��X�n�m��mϼ0̛RO�q�KK�ܥu�G����b��~��dx].�f>�+���S�����n�����1��LB�2�?��1%� 3�NC��}�N�Bb�V$wg��g�b���g�l�0�K�m9>n�ۀ(�8G�elF�[3JGb�,���H)����j[� PX�����2���H[�dR�iD/���]�-җ.9l��.*��}��)��>��v��ve�t�_�W��Y626xT�q�nM�f���y\pw�� s��p�� �#\`N����G�c[h�aI��w��[6� 3R�Q�ƨI47[?�N�?�4J�� ��w�(٧y$C)y5Z���D�u�d(��}pt�W'� !G5���e񌶤'
�(����XRE���Y�PP�e�-P%ç�W��7jf�p�O�b!\/l�����X���y��F�yX��dXvb�h�� Q[���o�&���(���b-I�=_�d���#��|���O�sv�z�Ls��):y~%1
B5!�����qO؍��%���9?���A� 3�`����WU�"�kƘ5`��D�m�k��;��;&tۇ�����CJ y���_]ɓ������/���� �:ĨC���:�8����ʓ���4�K]��0#�^��i��݉�찘)��@��uIj2�R�G,r�ɚ�r1\�T��HN�w���_��(����:WGm[�������c�� eN8��*`�'6�0U�$}�q�a�k�Յ�r�܊�)�v�"G��i?�-NBK�}��]�'=�CC���#�2�$/#gS����J8��8{S|$P�B�N, �8%�/�Ea�.������&�t��� w�a�0�\�����	 X��?s���P���@��
|Oi�ǰ�χXN)n��d��<T�ԯ�bE�ܸ]�i����"i��5lϭ��]>���>���$(4�qCR%L��qH ��x���.���P'MЂ�{}7�w�z7����0&��m�d�0�_�i�^���3�\D��(6�j�?�?�9u|̱i���Bh>?�Q�8aΓ���^�j�;�{�� ��:9*���=�f��;���ZwM9|`ağ�)�6�I��+��B�V�4g��Ǝ��d������H�b]��q�H}��YKc��m֧� ���gB}-L
e��H0Zla�_��i�O�i��� u%%�J۬�yqy�	,�-���סq)�ʫ4���uH����L��^��p����H6�Lz0�x>�����c;�]W�Ks�~����C��=�L
\{A�E7:�4v'���g�����[կ7�/>��x�@���-IFU�	ݨ��|���AX"��r������|��N��4�� L(9�h7$����3)�����$���*Ux9^�h7�����da#�Ee�%,�+{�qu�o��A��>{��%��<���NЧ�;E�5[t0{��,iaxq����)=��F�L��(���0Yמq �3��36�Xu"��>@�C�i
�F4�_�:�+�������"�N�?��&恒��8-��g���l`�]�6E�)X�T�u{����i�L�hc`�D�ӆ�z��֧F�3���|>:�/�Z�x�/'qL�ݐe�2B�B+Jd�ou�T΄IC/ewUȈ�"�u����-���^ŵ�l�e�#��LSX�j4ϖ�x�tl���36��S�~��������kcc>ݫ<��Ú�<����Zܙb^����?9�`n��ݧ��Z�CaY��u0��:Ƹs=8��k�U#]i��.2�[K3~0B�(ZF������h�j��/��9P��#�瞕C�I-n�ƃ��a�����vA�����e��]D�m��,��!�`�n,L
ҪW�>�!�p�)�#�ZCՆ���d��
��A�jI���χ�����i�����!iSK�)i�>�A�=��O��>mO�%x�=@7u�s�i��ʊݥJ%�I�3��C�{���mxm.I�k����\K:+~��\�1�ϰub`���*~��36�ճJ����N���]��>zB�:�n�,�������g��xʘ -&}٤�L}�&e}��ɇ�5D������h�@��1��ƃ�<��mb�2��c&�߲I��ԏ@�ѻ��##���s��� $�K�~�G������.���M��.<���6Y8#	ò��ӕ�CS����/����k�
Ʒv��w�H�xZ!���㭿3b>�sR�1����`��)q���{񋖑ڠ 	��c��� ��j����l��?z|h�/�|�R�x �4��L�~���>KP17#CC�-;W��A]@^����'�)5g+�!P�O��V�4)�����S���ŀ���?�2B=��c`3� ��'vb�������-/�&�w�S�,�:�mXttk��!�4�};�)(\E_<?��a�i���N����ĊYn���������\�v9�^��pj���$�֮�Y���r�"�O�`(tӴ!��.�Ism�v64�khL�T^B��9ϢJ��8;Ȝ�Q��	F���N�����D��J!��]�����P�n� |�aX[����,ډ�FD�DWClM�{��w.諫�Ŵ��h���.�O_��Xwe�[�I��Z0��׵���� �`;�)<\lZ�U��]�{}CCtOsj�t��[ (1dW%ӡ�<�ndm���i�~?h��</WxʦJ`��c��1�!rmz�Q��g8����"�K`��P�v���8���TЫ�E�ۣ��D��
��%��5�-p=��U`����g����M��S~�\�!��2�k�Y}��� ��n��}>\YEL�B�Gѭ� �P���p�p%���� �G� �� � �I�)��4J�CP�_r��i_8���o���D�kI�
m�π>�
@��䅧�5B*z.��T��1cGD��f���M$��MUAߩ�f���E�6��5Y��`HW�1f�,k%���3�8�n���0(Ir�J��|q��Wʵ�8a4�W�`F��j��1jhЃψƎ6� �v�T�q9�v��>�0����=_Uk#��&���.���B�i��4����{�sX�R-8���mљDTyp��@']�[�VEA�WH�U59��9nn�E0��Q�	�[�U]#���71�O�n�SL�!H�O�cX�j�����&p{�� �b^�qq]B>b[ˌCP]:3(�5@�LW�?�Ҳ�x����J|s�Wb
�xCy����TVd����Q�ɐ&(�
�["&#h� ��(Fʝ��5�e�cL�V�'J��
u����,��EyK&����g�΋O��L�ʧN`�0<ȳ!�w���9
�'���Oʴ������lqs�v�=F���R�W`N��}�<_%u��[]�KWS��<�͸P?a�.Ϸ[E�=��Wug+){���T�Lp����}in�c�9Z��������
��ߌ(%hEi�	�jg���Չ�\(�luv���۸��r0Kދ�oX��`�v���v�J@��7>追(��6N�J;MJ$R�[�-��l�s�@ve?��2�h��Kê�b�!�{���\B`B�q�2b�L�eB��]I���5d��g��7��ayE���1��&�$��5LJK����R0@�����2z���LY�S� B�c�׃|@�8����鹪��E�O�7D ��]�x(�oM�6���4����4�����3�ٍh_=��X��G��*oI�:b�\e�3�h�=R����0�v�n�O��PHO:��H�-4NO+�E����a�nË-�JGp�;i�����r�� f?5�6���`Hl������O_uX0��~��T�
�z�t9�<B�oP��,��K	Q�֏�`�ص�jJ��'I����d�w=�N��}i�=riwEG�|��O�?�o fU2��8K��1��|��a��?���W��չ�	IR�ԯ�d��� v�F���$�'�e:u�y�Q�7��i��t��c�Izg�w�^�q��d���>0�`,dCC���/�ؑKt��ȼ ��h�������s����o�������+w������>R���r��Fbp����U ,0�z)g\2�UϘ�H%SOtlɻZ'�ؕו5���N�zh��~���j�C8h�\��H�n�.��P56[s;�h^>nt��و���[�:��GĿu���$�Vի��q8�&
��ssؑ>L2Y)b63�;̌E-L�� ;p�!����E]���b�f�T�Ga���U�=4�,��"�p��I�ML�tH���
arP��.�n�4ڏs��)*Uӯ/�n^B�K��wq����<H�)�C�+P�1
}=��/����GU ƭ���;����ސIX{���:�y1�n�U��
��(�����4s�x�bIH<�g�`�E�l׭)�����u,E�[>�X�|�Ekm��~���]�L�D;������=F�'l�`�k�Oq�\ph�Q4�\b�����0��94�R�q+���ImJ!hgf�k�Z��s]T���ϴy�I~,)dNU�~��>j�^mOn} ��tJm8�M~N5��r�9v��Q��6�IT�!�������&!�c�9G)߁�\����CT�^�)m��*tR�ªX��I���VVL��r��
�@��tKï5�UL�A�}�N�D�m]م��H��:vIs��Y�pDϞ%ۀyW�0��p-����2� ,�7�Ӡo�aNdX���k���h���7�[=l�KD��Y�=��Su��V�²�F~GM4�����-�,�����5��J���Q�"�jÂ�-��9z����<�}�&e��7�q!�*h���qʰ���@��E��H�\�U�����N>�
_��1hûo~�3
��^&�fê��N���ë<�����b��s�s:!,s!��Be9����ak�wPGl���2��N!עS���o|�RPԁp�3���4����B�� �����h�p߸�̂�Ώ&�(X:��c��(��i�����Q.��Vk�%��۶�qf� s�#���/2��UФ�{�`�8���qU������.u�И��	&�͸q���ʺ��C"S�Ço{���QY}�Rw<���COQ,_���R g5,$�Z���l ���1��4�W�v�.i-;5�O��}�yj��J
����"��[C=�0G��|c��k\��U�p�A���f��E\�٦�q&��&��}�H~�,��A�W�� �����<3�̀�T�丸 u���Tty}DM,a�����q����$y�s��4���ZUi�no�;��]h��ɸ���@��fR�~�� |T0��?�kx��zM���A��貄����cx��]µp����Ru�l�[G�at� �t���t�#I0b���#��t�y���o�b39ajY�9=�EDd�x��!�SJ��bw{���l����y�E����읳���������hyh��3�+:�<�Wv�U��[(-
�u�?���K~�9pF�ڳ�����ǆk�!h����#�)R�9�Gב�X��$j1d��2����;��g����g����Y��	�$���V9+~%Ӛ]T�	a�Ұ�XR��Ə��?�<ٰ���t��x��������,=��u*�RmE{C���V��߭�d�gЄl�p\�c�(�1y��d�+����s0��FJo���ڄ�q ���)��+XGs�bK*#�>}[�(?�NƔ^�[?G݈A$�R!f%78�� 0pp���p:"�ZZO�GX�Q�>Z������<Wi��p[*9S�pE�2�롢�yL�6���|�bR{�zg���&q\W��е���Z�s����rRk�p��}̰C�����tEW��E��=�!��V�)���[u��V;.��d������xc,��}ێJ}��N�Kx�H���<��r�4��vB>���I�7T����ˢ6�u�?��V`t��#�lE诐���H�������]�o�Tʈ��.(�d��"�Ӓc��R��4���*�M���
�	p�U�[�+�n�[LDLo�֝�J�ߛ��x�fi[W���+�Q�+y@Ķ��yRL���h:V���S2��kۢG�[x��s4u� ��0�+��*]�#�0�,��H��(u`�WK[�'���E���qgǹ�Ǭ�Y>������lḱf��k����Wu����� _�,�>�����G��s�O�@�i�R[9��;	�n�[I_�q൧� ����x[��4ޗ��g"�|�N;�Av
e�1�B�z��e��#p�ĩY��V�
���S�V�f����88#� ۮeSsF-�t��PTG<�Ca$~S���� s^����sF{���y���|\ys0)^��.[���!����X�A����҆���pDcً��p�4DS��,�N���V��I�$l+��8�e3��������ȺO�~�_~���Uy���0���Z쏹B�f
{�q�K�Q��e���o�F�Å2)m�j�E�?85�,$8�]��xx��W��d}j�9E<��
�1{cԠ*��s-Ad�-�`СE��n��;�Z���v��>�����F%2�+{V>)�-��N���r���~��\��xg�j�@c�t�#1�1Б���֍;R[o�Gdyly�%��|Y�L�[�H<iH�*�z0�_������;R����Ӱr4��$1�j%|П/?��d=�K�2m�T�)ha�)^�V�Y��Z� $�����Eh��@����'���|��N	ӼX>�4�Ҽ8e�����L���
��h0�D�s��G�{��A�# �&�%����\n ��a�C|ߨFt��b7>z����&tEr��qx(<V4�IX�GBep�3��������;�K�\e�b~�c�c���5���k9k�h�Y���yGF	�k5��Bf�Ю��wY�Tf��q�u��R�+	Dd�����U`�_}1$@������^4,�Y�0+}�UKd]8C��� K��)	�a��"b���wʳ����o���.�N �;�c�P�^�h�"��U�U8��Mu�i�*�y���"}d�J|�}�O[��˂ş��(�t0a�C����oFsq]�X���5u������M�D�*��õ>�\�[Q��Ue}�������G��~e�Ѣ6���4��p��Gwi�����6��kK�J�-�%���\�U�<sԌx�'�O�ړJ�h:�/I�Ӽ?��i�h���+ ���ʴƋ���ft��!��-�s1�؞b�Μ �ڙ���=�E��Tni�_'N�)�6@�����V��9F�N����Rݝ�T#��L*)Ȫ��%�	�/{8t��!���b�k����1�:(�V9�\��AGv�����,�� ��������!��*�ks���Q�C��쯗�3)��[�"p��Bj%����R��/�|���ao���F�f��R#�E�^��u�����R"v��IEϵ��Dw��Vhp٦�	�:�6���V����k�і�lW��P)���BV�ڿ�%\E�X�'#:�����C�4�6�(Ra�k~S Iv��ca�
4�-^h���{h��]N�\�93�P��V�0�=��0YmR� a����jm�O�`�E�"�y���ez��@=	�+��N��P����k1Z��:qcBL�����yu��y 0�����H�_����K&h
����A�?Iv�U�S�ڮ��9m8�|HFq{L��aP�/j���svĩ̗�Rν���jF��ގa�*��S�2�'l]5I��d��o�����?bIˎ��Wp`M�Lቢ����"�pL��e�
Y�ۏuJ��O�Q�˭��Y:�>����-����bW@�$b����Fw�|��*���d�����'9�k����]�4�t��� um���A��Q��*���|��N`�P�m�U�o<�&�
p�Tp����8�o�!Z����"?&��+��0����"�Z�W��L��6�F�o�F����c��"�faa��*:䟫�(���aLE#}�a�&G�h�E^�+��+�1�Q���}�f}��usrL���Y*�祫�ޛ'�����P�o�����U��C��s�{*�9{K}DG�%�u�`�`.�j��oLmn�|L���oj�/�H� �3YGi�v'��o~�$+.c1k�=��WKt�_��]�dR0�`�F�R��v�fd�K3j'eFXJ��5�`v"����Ey;e��r�9���H�DK�S]�c�8��(�l�4j&nɋ&�P ��f&����g�ƥ�
,#.�@���lf���������bq��$��Ҽ2�@[�,�芾A�����#��B�� 2�Ǎ�Q��P����w]�0�c�K���IiCs��p���lCmq�e;*�U��dP�j�+�~n����~���'cb g�)6�I!�\�_3���iv����+w�D����cs��7Du�* '�7(�k��y���V�߭�>�ǣC6Q�	�{NQ����/5:�|���W���H� ��09s<��	R�<NSŧ�F.{E*q���|�h���p�%։���6O�I���I�T{�E��=�iC��x+]��MIr�?�>ӈ���d�ln{{}�h��[�!,�Z5o}F��{ݘ�����U�d�h�1�/��[���Zpr�
�L?�M�)��m,�.8��E�Kk u�S5�.��Z[�eȝD����JR}�JLm�F'�!K�@c�;=�:��f��Y
t?�{W���6����T�7e�W$?9�SHp����֯�8��I �&������#�tz���{��D�آYS��ߦ0+�,��X?����u)��eKi
T�ˍc��������樏���Wt��p��$�Z�蟪T-l/�r_`B�M`�p3^ry���-"3�IX�^b�wjO^���<Rq��
���꜈�`�<�����:=��7/2|��5p��އ��_�rt��CM�c���/�L�ƝG����|'�f�#	��;<J����X@�׹��9���MH�xH�
ģ�0ê���/x��nC�r��K� �E�( b�]��މ��p�B���ܙgc�2�szy���|��ڬC�������6�X緔��4N�t|�}|wn��p3��8v�W�Q�A��@���Ky;��� 1��HX�+�"��a�g�p�vҜ�#�(C3`;	|�{K���/$��uW>iD^����(��\��g����넥x�C<V�j�N"����tM�7@^�_	�w���C��X,��>Jkx�v��9�K�@
Y��Z��+-��C<Ϩ�>�vQh��WW�[�6)Oʇ�϶ov�Ʒ�է���?Lj�휙KJ��qv��u��3���q�aH�-��5;_��f΁����C�|ȥkFRȅI�|a,��
��i��GK.��W&�猒~���S$�\�ò`~� ��mM�i�	��� eqV1���{G:�a��`W���|َK�������,��Q��/�@��!e��|�<���4�����i!�x�d2�Q�JiH���t2~����t6��'�����J L	#:��y�R�L���7�ў��q^kH⃕��4k����=�qE��c�_q~���0=�x ���1��_��¥K#b�O������N�Z}�C��>9��=/IJC��YH�`�`-��y��	q���i�_��Meo{��Y�+@,��͍�Pͫ�:_�-�ᛒ@��d�4���t��\( �M�Z`�V��W��F���Deآ�BWT5����9��2:_w��c�J0�TA,lJ�C7��N�S�M}��� �1)��0)^���$ ̓ߍ"�Mtg������U�j�lrɢ�E�[1���	"��X��^��~��bI8���~���ٛS@��d���@^F���l�hU&�-���w��.�nPZ0O*�K��c������0��#�v� ��������5����S㎢ꄗ�D�z�RA4O�!��/�$0��lGN�HZ�J�b�U����u�P� ��4��a�Ni�k�!Ĝ�Ȭ���:�鸲V(4���=�~�
s�vE������*��N�]�aa�s2��F:�yO�m��#GL0����oe,n�5�V?���S��f1��"��>���J�� o�.M/���*��_���"(�����*i)W����o���E̻_)H��L��N�>gK]�f���ce��A�q�p�mCe1Ƹ��O�U��ϳ,�L����^J�z��ӄ�N�n���V{Emy�+�Wi9-�שH�{8�:�?IR����҅���l�Ti�*�)b��%�\�gW;*(R�u��9��P�ذ��63;y� *�+ �W*�?�Т骆�V"���[SkX0���k��Å�b��X���H�1p_V�!�m�oh��%�R]$�T���Ӯ��r�4*yQz�+��7�[-��0��[xx�UC[�ן�c�'�Q�����HsY���n���{�� �	�*�49�ۇ�Q�0��D3^�{��C�u���U%E�C}q�I�N�c��1��\�EwƗ1�m!2Zb����g3c�"`i.����>�w f|5Z
��jd�	����}����!�l����f9��:��k�M;�����������J[6�zD�o�R': �Z�pD�>��l�}v�|�S�Ksa�r�s�p�ɱc4�+�߻�A�H�ʿ��ct$�Rn����K���F�y��ٿ�!K�aj _�~�@�ޠ�t���u*��S�/��1��Q�i@Z*��י��3'�{�ٙe.�yqT
YE�${XWpDx<��A� �Y"ei�	˾�;R8�x���O�"c0�ݧ���m�Ƀ.�Sن\�S�0�a$�^|��D �F�';���Ê��r�o6��%�t $�d�ȉ�
����\I��a��&��S~kRn8'�%ܼ�p�1	D�~#�^4�F��!�`�8���
�s�rD�^�!�N�9!�4zTgl�9@��@|&����5-�z�GR^����p6��\�����B���vh/u=�WN�-������O�[��9ͱ,2(�m�񐰠�!gwش/�a�531��~rd╠\ n�Fz��W�jΑ�U�W�_{�͌�!3��5��Y��oc
 ��D��Tc�p���b��"�,!d~�p����Jq8�gqW@��D�;�c���+N���mP��9��kd�]e~d8���8|Oy���@�f;.����[J�2K��H�[A	�je&�V��o��e�;ɕ�s���]�+����Vù~)����l��03G���FFW�HԥL`�@����GW�8)�ea��%��&��O�������S�U�m�cx$ zΑ��<%_�����q�� ������=N�+���!;#�H�M�������+[��,$���)�^��9������=�YW��f�T6Y6��?(�U@pHް�1RT=��x��a?�L^t��ޫ�/��޽b��!iL�)U.XJ+����D���U�W���)����늄��j��8�ćt3�w!���ɴܲ��ѕ@F:ՓbЛ���9��;�<�E���[�7[����J����>��52[W�\Uw(9��]�M��O����������M��p��l�ĉ=�6����#�S?*OX�:���<�	�.}�*tP�P9��0<�OJ�pK�4�-f��`��ru�/��+�����v^|��'���ʼ��HY�ȝ�W��kY�Ҽ�#ح�K�5��D�<��pMOBn�>�πb>6��A�y��G�?DU�B��{|sh �+����b�`��|��-��^!οA܅�ޝ߰�Ae)f�����D�d#
V<JB�5�?2���p@�\F\����D&U`O�mY ������z;�R�!b͇,��T�^ɨk�*��j
���������ƚ`�"r�dRU�YY���+��O��3s��H�NIc����MD��ү|�n�2h�Y�@�Ġ���7��#;a��mu���81VUV�����7*A�Ch&�r�B[�Z;�g��V��W�s��^������P�mv�A$Z����&M��*��t��(�c�����̓vx_ƉI�`���3AJ5��[rK�,x��U�<�
r%�&���]=F�H����^����{��ڑq���|��;+����=K���E�uc�w�'
�>��q�)��AjZM͑H�Ho�L�h��36�gmCa�N�I�z��N�eˑB��4�[�@��W5d�v/MnO��2j�7#��p��ְNܓ{dqp�߮4D<�b�?����S�BlV��wnu�}Hd��咔ς���	+�/�\�G��m��Q:m6םv��^T:֊qj_�6�MO0�&5|��>�m$!`�踝�-��j�����!�1b���$y�_�+i�v�op헍5�*�0�*�SRz%���
:�~�T4"���A��NP��s�,)��[|�[[��ð��9gٖ1.Ç���������!Q���CX��w���S�`�4����7m��"��0+4>��]�	{����V�M�!�i |3� ���W�ݱ�t#�I����`�������{�U��O�#�$~����kb��T�8/c:��4��Ѳ��$��*�(�a��T�}$L*p�KTy�{C������\O��H�.�m�P}�c�Gw	qؚ�E{�)3_�USz���@�n?y����=�?��[�,��.io9� ��M���E�h�������jo�%|��ج�E�c[w�V{�py&��9�}�8޻.2i�M�����i����;кX�8-�k��>��2�<����s�:�C���h�J��@A���)Z\z��D��LL�����^ ��ߟ�cs0C>1�a�z`M��A�'�z�i��#9xt_*3ٽҍTGC>�s Y�vY_�8����6���5{ʪ����zE���u8-�3\��E&����0�v?Z"�%��@V���ۧn�� '$�n�伊��kĆ)��tu�9�f���D����u��(�bR�y��eZ�9���e���W��,5�d�P̘��P_�yI�bU	�JѪ%���	r.f,R�����8��:�Wk��k�b'<�pa�KAk�Q������&����&�'�rD��C��Dz5����Y�h/瞁:�������
��}�p�l(��>���^Kv�y�����[GWds.nյu��3���l����!�s�k�F�lm�&�c�|bE����$��1#j3���*<.A��[���IZ۟?��GEF2M�Ar4�5��RO\l�*�X�@C���53�}v�;L7/4��^��3�&�q��ZBW�|�����â�7K\��ԟp�tf۬y��FoR#u4��@�y�Ƭ�ZD�N��U���]nO]E�a_z�[������P~��#Y��^��)sT+nG�t�
{���)�;l�cS��$Go��łv�,���.F؜�Q��.�O�R��s�-#�]��1����Zà�y�P�F~-
���E���^d
ys*�Ȑ�k�;<[����0� F�΅��|��Á�HuiU��N��.\�;��I\�N`_�'+���@"�1Ӗ�]������ᯁ�*��LyI
��O@��js�>��,���QH�R����Ŏ� TX���&%2�	�����~�=����ME()" �?�������jwO�[}��&RU�>�����S��H$�^��Fů�8Ǥ���omUF�:8n�����f��,^�� .�1�]��\��W�o��CL�<2��P[a�"���O4���{R�M��t�Q4�bZ�^5J�*U�[���1���O��*4E$���ZT>��>�e;�n&�������r�� �R�+F{S7���Z �7�����!����|�XyE���(�_f��$`�0���M���;�����L�bx�2���{�1�KLQ�-csȐr�th�D�v7aD��u�~�L~�+�bC=��q��2U��w@^�M�C�����uA�y`�+]aa���Ջ����@��Dy�UMoq�,�l����|�z5�|�fX��4�5eL����-s8IX�^�Ԕ������+���n$�u��r��ـK�Cn~:�ZW���M`�F+ձ9m]�\�~>%ᒟ\a��DO��󵀸��-��`J�e	�<�e{j�Ec���i�V���	ܩ�"�2�۸N����z�\r���|6�;'���$����So猛p�����HY_��4���X����:�ȯ1��,�)y��j�a���E���XLO�,�m,��**k��n�U}z~ĸ�{5_{R$)pρf���S���Ymd[��Ԥa�e��{'v*��[ɐe��[v�V��I����6���8���W�e����'���3ѷ��x�KAƲ�J����R������d��g�֖�3�#�6P���G@���m��=[5�vp����b5�cIVX���#Q�{
�����f���P�,a��7�Ͻ��t�I�ܖ����L�=���;k ����P���m7����Gq	��;��9��^��j�8��0Y�C=�|��A�=ۃ�V����Ȉ~�:���`,wd-UiW�� ű�$�O��!$u>7�`C����P��@�B�uO����ʉ������g(M��o��������d҇�u��� �P�H�[���Y.��'����;�Il��U m��=�!���L�z�g�j{P2]59�{�?�S%��F�<G�p����3��<�k���AIoqpZ�gvo�(��-'eU��v�%5����TM6٪����n���2�?ϖm ���}A��6{� C�z�0�AO����o���">>J=LD���#_X�/#���t��iu�W���m�w�2��r��k��z��E�j��Ez7���X�o�܏@����

l��j$���:6'1T���e��������-��vU8�x���@+�}�n�C���&{ v����iɃ����jK��ޤ?g>ۜ�8�$��x϶�0�%O-�3�����#�7|�O5:�Ok?:�\�8*���-M�0�v�z�]�@���(v��d��_)n,4jh-J�j�8�������~�_���]�z�>;FHJ&ӈ�|�q�^؞-��Р1�?.��K�����Li؎�ޙ繑�i}��j����^�Ņ��ʤz}T�( v&�V��g�锿�g��s.����J�i>����懬(�D^;�,b�;����ب�	�*͉TTyh����k�V@5�ڄ��1Q G��1���q�k�@�~�|�8��ه5��@���oG?��ԯpS-F�M�osg?�.A����*�Z�8����iJ�[{�4Y�￴P�x��ȝ�I�d���&7�9�P���e;u���ܳGj�6����,��c$�E	&�'�J�(BQ��bH8 �a�=Ha��Ӗ@�Y���x>��&��F���7��$��u�F���I�s�c�I즱��|#ըD�ll�)��+1��z̔7�9���SO!�$����Ϡ|[6~dk��A��->���T� �B���o�TQ�J;��'�����\����/Kg���榁��/¾��׾�'y�:��>/R�e��[`R����֏E/u�x�r��qqd�->k�em75�"���`�6Aõ�� w5&����V{��P�v&魰���NאSՁ@:����&iq�n3��q���z�߈��W7����Έ���jU�b��IXa�B��]Y�ʝp4[ߨWpJjm0}ǺAQ鷑��E�k5�5&f���9ܕ�v������� �E�,pV�]>;��р��+�cl��/~�;��A�������*i�����IR�i!G?;Q�h?=��ʜ&�d�Nҋk�Y�a�wD'�p�]h�^��l�m����:;og���Yy��Z>��D8���7G�/"`�VG��8���ܳ���p�=y��/�c�P�e�i�u.(U})����Q%JBIq?RI��H�gZ�cE����I�x�U���� �5_V��oS-h��L��hh,��a ����{\��4�h�q�&N4��v(�w,&��}=P�c਺��#����jJ(��T�Ut\�8�����u=@��s�x��7i���!q>hٛ�3����{��H*�����r�_g]�wf�_���Dы�;C�g�K�e3�?R�ny|#çh�����ʠͤ�T:Ku�K�03���Py�h9�x.>��=L�]����0Ou|��&^����l��ne`��C,�>��CG�ҍEoB(��nh��˫�7p�/��?� F��7j���̲)���O����.LB�	�F�B�:�ˋ��<��T�k�X������"ϼ�߶�1�q�+�%�ȱ����m{(�ms������urs�^���v�U���6�0�}_���q�n�v��g/�O�����"� ����_f:T�ުh`8�4%�d�)�tj�3�`��aw��*��p�J���las�8�$�������M'�A4wu%�{��=��B>*?t�
+�J�M�z7���<N��y	�<���篹�ט�(ѹO*^�;�FT�>���餘e\�>�?��ala�+x�<��q͒_���Y�٨��U�Mb>ZN������9�yH�CD,w�D��Hm�0*�1���9Q���brvK��(�6k,^^:#�p�Y��D�֕=7������|C���1o��-�he��ɇ������H��Y�5�&Ԗ�;9(�LZw��)08�w��kԞ\�Gt|`���&�fP_4��]V�K�jr+	;�%g��-ϳ?�]�~��i1T �5�
��B�d�6_�;qG��@<�~�'a��8��F�n�-P�=
H���T��T29��U��#�(����p>5"�sd��/��.n�h�w�F��o7�O@�˭�W��3��oL�|�oaC�7s-}���Z�J���IY6<�g ��R�s�8�1:�E�����Rf�����,= 1$��k
I���
��%�V	�1��-8���c;Q��X�T���/�fCܕ+�I;��?��D\�_m��=?�s������L�����.҅�����
ļ�+-�������G�~ �[1��5 �Jb����sW�:䫷SC�(9Y��8��x/kwGz��b�`�Հx����j��r���Y��:���� .Bd���sP�^�:Q���i,�^5G�@�|9�%k��ώ�?�d�X�wq�/�[?'OHY��=7Uʃ���98�h�8�V�쎜E6����J-��Dj���.!<��,�K ?b�aǇ�i9"
���xؗV�B3���B�̜���o3<JǌY5�y�l�,�Q1y�XꚂ�2��
7 ����|�����#W�5�^��e���Z¦��{�x�o�T�X]�;p�\�Da�\2�~��P{�IE��,����S�5$V��:��
�D@�#�1��ϩ�x���p\�!և!̃(O��ϫ��.�])��#���P�7�ˈ�6�뉹�8Em�>}�L��u�=��X�����P�m��N2@�m+K��O3�R���-\���D`�\'Op}u����g�N��I��B/�"�w.���qɺ�vF��|�=�Zh�t�!���ќ��;�(�7�R#o7�sr2f����A|�Y��r��ߖi�RF#�rw���$�η�]�ۊ�Z���hI���y�:�1��q>dqϬ���F��9X�h\���
lb�r���o0�=�P�����S�S�eo+z7IL���Q9�X��?������ ��5��g�`�C�MK��!��b�ۉ��<�S�ۀRn�И`%36@��F(�r K�G�N7��Z�κĭ��Pbp`������)O	1]���W*�O�U���t'� ��Τ�Ǜ%u�#U�O��|�� d�Ia(E[D�H
_W���<0%�T1&.��X�ˑ�����T�*_��+8���=k�\���`~���"�r�m0�7:�j�]oP'AӠA �09�Q�q�Ҟ3B�Y�A�*9�k�̟�O�	�^���.�ȶ�W�P�&��  �2a%�8�ܔo������; �S1���
�c���g�׫|D�u�o/-�m���j�Z�L�/;���g��o�T�[C�_HRQ"�rw��R����0tg�(#{y���iV(S0)����mi�Xss��b�^�rrP��zd�P�L�E��$E�54��$N�Ӥ_+B�(h7�|7�"8���c�b(t�V,���g��"x���[�&V��Ƞ�pҤ����R-�O🕱�v�QOՄ���~˛c{�.��{i[�I���~)��ܽ#`��fx��74��Mo��Å�QT�C6�I`gQ������xI4�A�SI�v��ӫ�AT����4�SC|T��,�
�+��$Fej���@Iq�O*�o���#Ls�����}�����f���<�$��&��m�'�T�������Ù�Hb�ʥO��G�<.�@�c�g9��au�!,-����u�cK�/"�YC��PȂ����)�6g��|ccg%IA��(�����J��w0�� ƶ����8��J����j�f��5�z��{���fa�R�$�5M�d*��μ��HX��ܤ6�����ة9����B�ьp9Blqli�j��e�(�V�,yi���U����r�s��&��<g�'�r5�y��b�K``Y�2GC�P.T��W1��-�Cj9�J!>�#���R�)��G� Z���e77*r^�+��!��"w�˖"�'�w�a����^]�x��U�!w��i)y���e�ͥ?W��0_!%d/�u���6ou�$�Y��`~��z���7\�ķ*��B<�Dá��i�l�����	W?ی�쬥�/O6TjC�Y�N7�y;�ƶnK���in�ۖ�u?O�CK�6� Y�#�&H#H��mX�@�L8 64��$��̩���p�$B�T�T�|xi�]߼���l��u]���a�:��/��?�L�?�{��b�B%n+u��n��e��8ғA3�8����/�f�
9��_��ck.�0?���/i��V��To�� �bC z����FlzF3a��ҰXi��>)�m]����!���4%�Yc���,�V�Սg�	>�j�/Wo�*!oB���8��B�̒�_{��bM@0�zT�R�}�4�z�-�Լ����s����k����Ĉ�n��jF�Fz��X�h�t�X0d��H���t��ݿy�/mu���W�}�Zp��c��0sܟ���,1�Ѻlz�,�D��"<�`}�=BEEP����;隁���[��g.��x��i:0U��?9N{x8����
�@�Q�����	ؿ}�A��+\d��O�#�DWřܚs˷���/~m"i�I>���b�Cv¼�=}�@f����m�z�ҽԤg�_�l�����:�Xb�ɒX��[z�	��l{d�ߊ�A ��,V&�%�z��0e_�NV�X��t_4ұ�"���	r����@��ԥO�#��Ծv�w=$��J����Ǆ��B�x}iđ���'3�$���@��5�����7��-R�,	)�]O9/��U���m�ě*wu�j�4T�Qy�uQ��om�݀�U<f� %����+���d��&^�u�!3EL��vIB�c�m�dҜi�m��48�õ.�骧#�J��FX�J����Y'�'j.,�>�֜YxD3��s�A�y�KBS��_K�;��^x9{���)��+�e�\PX�y�@O�S��B����sgD�P�Ҳ	:�sɞ����`o�K�R�j\8�E\��]�B������Fb]�/16E�~�jm�7������e�5�=�*jḾHal�o�M��XԊ&��)�T�=�#&s�w��M��Q�Z��4�v�*��
�/��IN��5���Pm��}Am�@"�1�g�d�QCm����V8����u77�-���`�@�~�p��^4Gp���|�|˶��8wʍ���[��m_]+�܇M��gm�˜������t�a	ݯ��Qe� ���zkS�5 �cU�V�[��FI����@\1�+�+-�W\@�B.�R�,'?L�EiX�� ��P��8P4ޯi�?s5�[E�� ���%}�Ø�M��P�u�M�c��C����LU�
��Il*����،g��������5=ƪ7���~�da{	 h'/�~\�S�o���&�\[P��!Aҙ���0�ï� �~�X{]��,S�͹t���Ѱ߀v�Vz��e�ٰ�C$�p��m���o�yK�.�������[x~z)"q2�0M��@Z��:���N4c8�/�HZѧ�"Sq�w:̈́��U*�Qe�D���eU��t[���ځ��[��dF��I��~����'�h�bgi�=�J�T�z_:b�7�EL�1׻��(	��!x�mbJL��fo�d�Ĝ����p�m�BA��>�u��ޤ ,1��Bl��6dWX�-�-/�E��|���wH5^�ɍ��⽏?Q�lQa��~��g�� ����������2��V�zٌ.RX����H����[Sm�1���|4���X���3���?jut�fai�_=����38DmK�vdUYT�W��O��f���O��sfmJ<s`�.��]�N�̍J{��+���j��Kd�+8֞���z������fK�����߽��Y�Rݕ��K�� ����Y�t�t&~H@>�d��ɭbOh-˫�>V�����*��AQ��p1vm`Z���6W����}��r֞�����$x�y�Үap��=x ')�K�yy���r	*m��`��`�	ȳ����>\�2|�O��f�&^�h6�R�p:���>��Er`>��oq�N����=�K�H��O�]	�(=@%�-U���8=���ԵF��g=� 7�$�o�9���"}�6����K_ߊu�@���6�Au�f!5����6�ܛ�'i�u m��1C��o^U��u7���ů�G���6�9�B^�r?;-a�`�4t/�5����%�����S��ܾ�)C�qh��o��+����#�v�5�,��i��N�*^���H
� ��~�H1�RDI���/(����퍭�X�M�2���r��#3�#�4 �l%`Ҡ����/�U�h
<?�#��R�H�2�%۾z�r��%�W�Y$4|����"���_nC��� ���͒�T�0��-�C���b�{J<Z&�)���]�w�����^�ڽ��MԌ�m��JT�iAu���,e�L�zf��s-��+���(j��	�o��8���T��n���x;;iJI՝��Z<����T����6���ۿ�kC0t�F�@Y��1�7T ���"���\��(��\��\ħ����A+��{��UՀ�#A�,TI�)g�ĂG��o�'���J9��}ܫ�g
Ǉvs\�����41S}#t	�,G@-��O%[�ܬ�p	�?���B�qq6n
��në�R�hת�S]��v��C^�'8�)�՚�L����o"���b��M���v�B�._ޞ����齽�"��R���y|D��b�5�C���Ʈ�-گ�0�=
�����u�N1�O/\3���{����g�Q[&E��{]dt������E��,��?��`�,2Q��(d�ˈ�&��,�r&����Tw\�F��Q���wǂ=�olܐ��9�qjNY���@��*Dn�M���K�vi��x��� }iN?#/�����8'J0��zIe�����픂��x��oy�˔˴W����|�����(�3n��aσ6�.&`I���ܓ5�&�öiΐ���2��5���!���(���P�1��:Kpq��:OQ�3T�p^HR%{�~O����d�w�`�IԴb(̳v�gvR��q��nh�\���;6�7��
��>��{V���~+�ukB�"�(*)i�>������']NQBm\����'�w5�.�A+������ϼ��K�٬ì�
R�E�o�1� �Lgpoe��3����}�:��0�Y�{�$f�L�K�;���� �T�2�^n`�����U2��W}z,1�B��[�'Q�b��3^��IX������Gԃ��7�׉Y�3	���F���p?|���z��X�g<��/�Z�E�O�\([*�ɥ�8�	���M��"��#1��=��v��X�_��sSH^I��J�|���\Z'I9Җ���z�s� �c����fV�M��C	���R����ř�/���s�I��R�m�n����p*�`��9.�u�����w�Һ�]e�d�/��}������)�|ј��"3���73z��8�Z�i��f���l|@	B#"�+���(�K��&�Z�<�7�P�q�>���эG`*�0�Z��_q�lF���"��Kw��v��sY*���ȧE:��q{��K��:���B�-Ja.P�Ӗ݅T>�4c�r�0@�y�od�1����N�g�.�����p��,7�n��,�mP�e^A���If��[�	2Gc|P$O�nα�MP�u��+'`ͳ[e	�| İsQ}�{�?%Q������c��Ͷ���q~�q8;������#*)�=���g?G��Րb���[��%L��4g�?�������f��#[�;�����~��2�J{�����]V9(C�`��{�b�?~Q�%��	�ㅤ����"��xeRE�����z݌3h���k�`�	���0'��B1�@睙�L�$� ��&79����ۆ�9ą`�g�xXq���Ⳡ��}C9�����=>�dN�q��;��;�2�'� �w4��I�(e�d\3��so�4|5D�����`���U+H�4��4�2A��9d�Q��;g��˂��I���U�Ȧ��L���K��A�����A9L,Ӡ���,���GUM$�FJ��_��vܡ���U]�B����]H
��D(i&!H=�#bH��q��KW��xd.�6l��[��m�:[����\�s%�!"��|vu'lʙM�����(�j��2j!��R(,�j�⾶|`�e� ڌ�Hf�|��fb��0�q��W-��$�2�67OM}9IcӰ��T��:N����RT��e��q�9-�}�q�a"`p#O���PLȨ��x3|�W2�g�|vzG^��P�kg��=.	��~{�J��3�,~�S�nLlc�>��wvO��`Vq����^�?b�1
5�ر�R#(j��^�}�B�Ϟ[�kO�&b�{ېj����	7b�'U&R5V�u���j,�}��)���sb��l�l�X:
b+��0�Cd�i�q0���7|S�g-?�̂T�#�'�o��N~ך.�S�5=��b]�Ku�����8�U�v|6�m0�'D��:��2�%������F�2>�q`�I�c�!��݆ͩ�e��Ҝ�*��]�h��7�9W��x}m��{x=#�8�q�������u����n�G������'�#ay������;-���%Z��b�hɆ.n�>c/�KV��h�@��i	�I8D���1������&Ai�?X�%��q/ҥ�C�W�P�}�l�B��~����Ȁ�n�&�&��(6Ч�d������k�Fl�H��g��C���iG�?ܛ��)�uD�t����Jʕ�'P�̿��Ϻ<�+)��I.BR�1�}g�d��#��Q�t��@i���M�%F���^�����,.�Y�cu���f���)Х��G�
�<i�M6�R�RO�;s�	�x=����'s�^�S�݄���y��raʿ�
%m�Ͳ����a��<8T�N���8=�cηw�¥5�#��j��x�]�W�	L"mlKtPD�$i��㱞��F�	�`�5����u�isO�+��%_�5�ªa)po��]L _�譟��o֬���	�!���B=��ܪ婃��x�Ʃ3g"\uI��Zt��1y��0� p��{��`�d��4T���*�^
/��$�mL�v�|
�9�r���9,���7��쫠�}Q5�`}`�Sr<��A|c���CX��� �ָ�{��O.����q���R�W��ٮU��D5��D����V�$�L	@��@P�`��u�[�Za,OJ5sG��0@M%�dq8��[�9�}��r֔é\cXQ7ƥl����a��mWˤh{�m��r�O˲��nXkb��4��>p��T�l��N��9����>k���}��b��;��P^�fH[ �vq:��6����x�G���u�q>5 -d�`ؘ�.x�Xγy�1���;�����,f�dSO�O���FG���>��ezDL}B2yS�=���NkB�������.ǡ������qS�R`I��wS�� �(���5n�S�7���[㥓���3F�l�i��ή^��x8�� I���®�-c�q���lnex>ǜ��\���*4pAӯ�P=\�m%��۟���H������}}�^���!A��?���,|�%��?��� �aź+����`�S���5F�HSN
�� ���Hkb�^ ��	(���<)1_�ٔLBU8�� �`�;��m�j�l ���c{M��z�)>��t��&�J�������6s�͹;��rĶc�
�����A�S�j���<�9y\rz�7�/�͋�C��/�B��RG���z�j������mϫ�|�ޠ`��#{hm�bk��G�]qh�w�;�����P_+ɱ�4<����-�f�&����VP���q���Ie�&���Vs���	
�$�?��w=8��buI#jF����Fޣ��fIi��8|؟�)˟}tm���ߐAZFh�
@_b���C�UϿ	��T���i��BR2]>c����y�]�>��b��#�u�R�쉻����l��m G��>|���?x��y����؜�둾�����T6G�{L#���9��(�G��%�^�ֵ �v���VI�� �f�Ǻ��=]ɘ�:�h�(Pa�t{.�Ѭ`;��M�#�&w��Y٠g<K�����������J�!u]Q�:���!u5VC�1�ģ%�����RI9/�T�)r������kw������o��/"��kUm�B���> ��釟�P��"��%>���rn�d�ؔ[9o*$�\ e��kn��Œ��~Q�$�EiXb�cd/!O�3� V�8>|M� 3�+���g�ڠ�A�n����]b�1d0Т�@œ�hz�#8&�U�6�%��j���@D��v�l���.:��h�F��t������<8iO�y#i%�ώy~�
�U��%Y�%>�����[�Ǹ�Í�M����~saC���*�$���J�Z@�a?���&�5`�ax "�
�T�)��"av���X?M�Q�u�*���8|�XE�����bV�;�aU�k癤Ƨ|���r��y_="Ԓ?�ʈ=ha)��3�/�E�o�7椨q���c{�wZ?������^�`�s�Ɵ5�~�s)�D�s���9���|0��9CBf�q�<%cj�xwA�I�~��lp� !"}['��ts�h�$���W֯hp<�k��Ԥ���t�*_����� ����x�|�,塄�pD�`sN ~_�+}(AP���ͥ��TFž������*u����	��b��R,:��D0(P^␳%����(�(�� ;!s[��"=�ſ�x	D�U� ��C��dU1�y)��9��˚�W�k�K��n�V�̦#��N�����2Lh��iIw$8L�+��ф��r�Ҽ�ͮo=k�"cJ0��������P�ђ�
�{ �-Lv!HCG�l�0ߟt������;�
��U���S�ݖ��2���s�������%8���q�E�ێ7��ubO���T�XU���,��~�b}�u	�X�_-�<P�p��<M�o���|7��Z�~p7c����X��!�m�k�;a�*��ޙ�~�>ǿ�^f�}D-���V��٪�s&ÑqG��Y�
9����z6W�����Y 1�S�Q���e���a��%��[1��5�[��V؋�*�'Ld.� -E����E������pc�N!�a���w`j�7�����]	�D��0�sPu���`6�4��&TQ7/j�ő%���"�Fa��?�J��eP'^;�u載Xl|�x���{�r�8�	{.�7��U/Zfz�?��0T�,�.����k��&��~ Yf[�^	�6䛻uz+Z!�S��@�ٳ0&��h�;�-�{@z��1o
���Dl��D/��blɛ�F��f�й,)$9E�������#�-�U��wE%�EXI�t�W�uH����~v�W�_���|���N��Bz�("(��$V3��'�lT LuJ!���d�@r�F^��ٍ�ʢ� �[g��D����=�:Ze�G$�Jl�d)Һ��it\�׼O�	i�������nğ%������#d�<u�envH:��؛gYh�T����yy����wG�԰�;K���?�P�]�F��R��j�Ӹ����ʮ#�����
}&���3[� �W$F�.`�	m`b�+�< ����R_��h�1w��X�៿cԼ�i�K�l�����E�a�g߳g|U<q<���Llx��p6u��~V��C�
�]������sl�Ϫ�������i��(��{�1���|WH�6�9U�veܡݱ���kH�`N���e�+���h� . 3��Ȯ��ċ�Z����,����t�+.��������[GC|9`[�-�+��a3(�}JvXD��+SN������� �D%��`Ii_Z|�ϵt�_�d��R�8�%)D��+���<��:#av�����9R�`.E&���W3�������S�4A����+;y����� 5�hߺj8��65���s�e�	e��&��8������Kd���Ka����p
et��u��!�c�cOSFp�$	�o���'���P-T~Ck��_�؊]��מX
��tm�G� `[�П�����ɓ�(�,�"E+�h�� ���17�!�
)9��e�0�k�E�]L��g�̾7�u$���A�bxS�D��g�+�&�X�A�����(�ݿ%�v�yU,��|��?O�&��O5��]�(L?�_{g��Nn��)~�q�E�-�>�j���h���ʹ�!�j�	�h��~r�]5�2�D���U&M�ι�I��q�X@��i�:��°��_���&�2Fe|��8��֦�!#�uH�U��ᎢҎ�~_\���ь��� G���t�N�B H�I`G��y"+�����7�4�yD=�9�uq�^CTӖ�<ARQ������P�m8�7��-��4ܙ��<5�TE�ԾlX�|�o�'~K*B���$�싰�>>R�R���ۺ���޻7��S6C�o�,�$HrwaƟ�?T��>��@��$��B�d���-"��¿o@jR��w��D�ɓ}7���|f?U(�ǮY��j���)�m���Q!�z�5|�Zk	ڪ�� ?{&u��f4{a��j���|��"[UvKN�V��QD�:ӵL�<s�G��X�嶰eՉ�����\�!l	@�I ��-IA4�h*�9I���� �Tf��5�V���ԒYT&��"���)��I�Ȣ w/�<���y�}�b%�5h�Zg3َs�C;
�n�C5{|RG���C���67t�����[$q[7^ԈYP|��@A45�k#d� �����+�q�Q��:_�߾#�>F��5�q�ep߅9�*D�]w�y$��a%�;��PmP����W���Lm(J�^����]��r?���#��ɠ�,�3u�<�󀛪n�!s��������ǟ���cFD�T� �±�h>��@��A�3ŲCUE�3��3�~�͎���^�K��ت:'�JtladUR
'�m5����(�^K��['$'�X���9]���(�	#vs{	�t�� ��=6�u�Gx~�B��?�Qj�׏��Ƌ�0��̓^k˼��n�I���	�ݚ}�_��K���e&B�]%�JE0F��K�ZK�;@��t��#g�!�b+�ŝ�U��Qq���h'��񆨯���h>��+�߷;~#���=G�6��y�V�je�P��ʖ�+�/L�!Һ�F/;��;��F��U��=�X;0's�s`q����\�����0/g#�(��rc�V9���
��O�Y���D�="�b{���Đ�'Y&��l�n֒( .GI-�͇nBW��1˞뼅�_�N� �B�����6�0���M�=&���(����$54a�񑼳Bf��	#� b��X�:��J�f�@Q9)cS�meV崾�̚F�"�����ͤ+�ؗ�đ��ְ�C��Q�
B&�>�����T�3�-�x�1ܕ*o���'p�����E��}r�)Y#��zA�m�%�2��
ɱ�����������x"���� n����s��	qE�x���HB4C��Z��zg�Ӿ0�9/v_�r6>B��;h�c@?��h��ZbTȤ���9!&F����w�Ҹ��pX��V�!�\^��j˿fF���H�L����#,����*�L0�Ό���Y�;e��/N?$���9� TĠ�� �K�A9x �C}�E(iF%�#uz#�VW�.jU��0ۆ1ĺ�p�W8��#�r��^��F6R8e���mL�[�6h�c�w}����x��4�d��۝!͙G���Xb�r@��?�i+����5_L�NUKS��;��-Cǽhn�o$�jȂb��/�FtU�<7����J\�J��:� �r�^��Ҕ�ݍHJHa*�΄�V�� �uuİH�i���#�gʪ��i�]����<�\�(����O;v�_��Ϊ���[��u� S�*�����fh��#�.�UXuw\;t�DtuN�l�L%6s� ������*�(��͓�m�y�������%M��-Z�")_�֫�q��,!�jh C�G7}��nn�7����gM�G�fTb7cnj�$��
/���<��z�?�n�*g$wIEi����n��'���K���2���w�k;�Sۃ��|�T�S�:=��3� �\���ĺu�QhC�k˿���y��	26��ɔ�[���Q�s�T�����Wpr�U5�$�ń��l�?��3eI1�����ą̑KpƄ/	?'�%L��W�A��z(��di����ylL3Q�&��7�4޽�i��I�6]{i�
�	��$#�w���c e��rte��K)}ۡ������S��b�[�`��J�y�d��®��n]_�M�����|(w,��P/ƳZP#��(�������:oJ1�M4��L^��J3C�l��(�n���K�Q�l$�nA'iq�L�s_�f[�����{C?��4�Y }����	a��K�財�]v�d��\���"��bv-��?Dq���r>!y����Uz�3wA�?��[ ��fMI*� ~�'�@��t���a����CH>��`�=�#��Ƃ�9� ��4d�.��y�Ʈ}@.�7��/z�����&5"ѕAQ8�dw9{@�!Ϝ�����U��=�<
h����)�g���bIVs��K��ђO��ZH1Kɓ!�_|��3��M#2�ae��gy��SӟE�T�H���<���X�+/.��S㥉�|�=�.<�m�v�%��֍w<���yrx�e%�r��.8I�O>}�θ����7�6��N�����{��=��r��]�%���9��,g[p5+�?c���w:���: I[F7a(�Cmn'�q9$F|����u��QK�y��-���
ܥ���xc�%��'س���Q�(Q�7�����C��;p� �N��M�
����MnL���h??�r�E��7ys�5iY��K30˕����
k(;}Qec�����ɀSd��L�"�"j�,0��T�6@�ǰoƜ������~a� �,���[Q_��ł��\_�е��L�Yw��؟�͆�<Yf��{o��c�ف����-�g��<�{?�Gڕ��n;�J����`��o�ح-x}���@,9����y�;­����(I,���s-�a�+��H;�9ټ�o���d��;�|dQZx�s�qsqlљ��rKM���H����G���q�L9dP�8�!�eH#�#	�5)l��r	�b��LD���>@}yM�'Q�=u��tx�����{����_:֏�;!�4tQ%n ���޶g�]�����B�F�6p��y���8O���p�_��x�Eѧ�~GsO��Q��n�d�����r �=���˶�k�îy0�I���  w3���s�4`t��?�5VEm�r��}F����"��{ŷnsOt� �L�r�)Y�S�I?ob�`�����d#Z�I@՘g��]�\8�nk,�C�A*���Ou�N���]MU��"��8�o��ܲ�TQ�g7���z��
�6L���Ùx��vE/�� �/�aA�!�B�͐8�~�GX�O�?��*T{*A1K���)��X�g�4��X�p��/��P�z�F��S�z���4��E��G��m�!4|+>6�Ι�D� g�r��&��)�h������l�pQ�KY2S�����D�*`*ɛ�)��W���^tD�3�C������	3��E��6�	���#�$��e�tN��+�(�**�W��Mh����-~�x��A�p��TM��t:M��'��^{�L�0�!�?n�9���H�� ���u���W*���/���Im�8vZn���U�;Š�^~e�ā�,?ۺ�pkPv���O�M��X��7Q���0�O�65�?׭��F�D�`X_���`yU�M���D�7�z�Z�zΚ���,UhE�j?�O�>r�Xq�̗��B����Ra�A�Nd[�%�9���O4J�	����������ɦ_�b�
yۃu0��#�����V�CTW�U//$��9��>�x�)�GjX�T��!eE��ޓ�Ӗ[�Y�-�J��P& ���O{���S�`��U��J=̻1Bp2p����m���D} �)�gwk"��pB�Wq�#'M1�֧U����#F\�g`,o{�Z7ϡm�ހl��$�&��^��2���#dGmZ7|}���C?�JZ#����Ʉ|��vYUn�&Of�.wCQj�_��6e[L�"r0�H!�S����p��*��4����cCW�x�;�q1�?0���CϹ�X�y2�Q��ڢ��ƤK�`�J�f%P΍�	'�G<��d�c'|S��i��bG�����^@����>��N'�##eV}��~��S&���D&���Aa���Zsf?�,=3`��������
d��p��Q<��m8?q�ld�y���dO�K�����{�����<��<��� ��7$8��ٽ�Wmg��[e�u����ƹ9�oz�	���[:'��t����@�2�š�b����ɇ��@Qk��B�p�Q6|�e �n@"��e����,��#2F�Õ��ۮ�-�s	o�*a�:�Czj1e������s�ț�"������L.] ���𶈜^�U��1JZ�p��2�#Sa�P~K�j��O�&��z(�)�2Zt��>|���:R���q;a��$���=�~��e���{���9a��}���k�ޢ`�S�a�pO�E��~�l�l���w.6�{"W��k�g,q:����٤���C�fH�s�p��C�T�P��7��2W�9�т�d���p"�֣��*��q�p�&6��ߣ�Sb�g�>4žUp�v̚Mك��U���6I��6��)$���sq#�����FD���ܨ�� ��|lƇ��5�t�i��c}�ew輪�(Ou��ۭs�'��9�e�;fF7��E�P	��g�#OQ
!o�R���� P��|��s���p�X���H ����i��+#���Y��ۀׅ�?�]-�
K'�m���Yݿz���D�-Z6����l��kh�!��i
�
���,+N���+�@V��,���������8�D�\ɸ��1#�����V�6?� �yg3��<'?؆vر����c��8X?�`��f��r�lHu�����~��mm	+�K?2�?.[��������H|| Mɂ.m@XWl���{R"��f��wdr��I�3ľ`M��CƼ.��O�6�<_��S�	�9�;�y���ad�:��h�[J�߇JMȋ��u�k����B���r��V^�ٜcy'�_
y�M�o�޳�#bs���]�b ����<����"μ�6%��?L�����R��̔9��"˒}�`��������:"@��Gl_v8ے*M�։5������@)���
����[E���	6텦T���jP�����w�Ά��
��QƘw�	�Q��Y.���(���wE�R���p�nnw)x@�e'N���ϻŴ�~��~k!CK۹ӏ�^�d�Kfpj��>+_w��s!�[y�V��q2�o�m�**��6��$��k��ڊf�"����KG�s��� 
(Y��篓ܢ��.�K�W��|�NW��-�Ư�U�[�~��M���ܐ��@fX��/c�*`�_?�^�|�B�S��L�]�xnHe������M�\�u��ˍH��28O ��T;%�@wx�u�"�!�����-��ۻ]��/�y���F��U�����Bg���)�1���ȩ_����Z��|9ḣ/�$;I�J\�#��F��ì^���)����K,�&�D����E�x�kq�����h���-kr�-Th���g����03J��A�-�{����K.�e, �����k�H���D�.�4�������H���'�]����+�E|��#;n2ɿ91"G�]mtξD�)�G܇y]m�S�5(?h�JJq��o�e����&���Ƹ�����~�1��Q���[����H>��Y��>+PDB\�>���bꌻ���M��)'�����2���O�t71����t���VL3�<1��0��{�}0�],��'�C�x���ǭOs-��T���e��ܥ��s6���q�g�'�:蛩I��*[�wp�ޠ��Dfw�؊͵�S�"��r�	*�BD�h\f��2����8%VIe��L-5�N`�)p��Z`XljO���f1(��&�K�V=BG���
^.�� \�b���.y���i�yj�?@�+$��l~.��B8E勈s���eY
��֠`�\��
�x���:"����F�Q�����s�G����1�����xk�׫���p��zN���Ӯ5�����EF��0YS)��5S/�6�ri��(E��� �u&1$h��d���F�����NI<TPf�?)�yĎ�ͭp#��+�I��K�ROҎ�ߴ��OZ�����>���	��v���4��6�p�@-;�����w|�[;䫊��:�A�bz'��sF��;&2!��i/�,��/G���Hˬ��p�sm������ꅢWψ�c'�$��LRJ��E�	�C�]^�����"B�D�a�r����l0�0���b�����ts��	�~lޙ�ra&b���QÖj��PGT�Ł{:����֎6��6�&=� ��+�}I��xR:C�\�MN�ETG(�oc�gW��l�%n6�.��J�=^eA���;��,O��SH� ��N�L�ȷ�_h!2U	�x�\��GB�\�8�s�]��[N����A$�A*�Ҵc�u���-�<&�c�N�7���f&F;y�#�v�[K)��.ہ���v��������TŲ�'bG�e��oE3N�v%�O�&��؈\C�����K��	:��k��p$��H[�$����5>�������Q����]���3�9�r���pŭp�J,!�8<���(��ҿ*JE~*sB>�*	v���4�}R:�J��JEfif�@٣9����|�WL��pKUl���~�R���.�UM�-aJ"f>%|E�<|}Y��]�f�o�<H4>Yh�0����r8k�����Ƈ�I���8>��r�N���h��O�
W�U�*V'�{�>�wB�$��Z�8.���A���|g&��?M���+�p40��=��,!�6G��X%2VE�ܛٗm�(
/��jV�>����1Y/G�S\�MB�L,&��¾�N�y����<��*9��c�,$�A<����	�oFL�v3d��Y�����q{�k8�t)�IO����P����jx�A��U4�*l�6���&~(������Ld�� ��H�J��0�����P�0_��Ɩ�'�v�똨 D�~�X�W��<�XJ�j��GП �6�������٪r�� &��lP����[G	t�ǖ$ķF#U_�*~aP2�sa�eS.��C|ׁ��k���{�P�����L?��BD�MsI�0T�!�w���@,ا����'��уv�L��&}ϠEN_Y)/~m���T�V���W�wޥU��4jW���������F%�z��"��p,����V.a�ڿ�����V���2�kԢa*)�U}~΄�b��阛%�p�s"��[?m��H$$q%��'�	�f�39�����]r������)��A�loI���K�������D^n=��<�T��>�ϔ������_]�Y�T��sqb�8˩�ݮ�&�dW6Wm���ʝI�6��^Ud�gz׹]`�u������<��>�,H��~ym�g~h��R���=��>�g����Y�[��&���c��z����c�{�ۤVQS�т�)�}U��@݃�T<*�ұX��U��3��l�hTuK��m�)�?T2'G�e���7Wl�dy
RNn,j��ʽ�ȩ�.�	<���=��seօ�Op�?8=[�~�$ЭD��}�K _���ǓU��`61!U&MX�ZQ�xۼE����YTI}�iVŸA��F4_�e�A���WB%!��@������j���IH?�=�9oQ�R��c����Ys��`iun���:��E�O,3=���ֶ�Gr6?㩗�\��n�q6���<	o�@v��5�5����k,������:cկ�7�"p�3h�
r�eŻ������L/U�������w������������������u�w�!2�3耍�u�|��C��.�lu��
�\�'�V,�b��6��A��ثd9#GT�y!~ֆ3&��WP(v�
|b+����l�i�ij�Q �]�qW)�1��8��k��?k��]�Jx�3Ӹ�np�/�����-8u �W¡N���#��j�!�.�D@H�(��(�]���u��h^�t�/M[NZ��t4�%2)m�2�T%t��dG�������dadb��͘�
����]�Șk>�b��6�2�svhL���Hت�?���Ҡ���I����m,�=]�4�$�U��\[`W<Kޢl�{�7V�.����O���T����V�Z_����հԫ#1c��m:���a9׆u�s�W6Pr5�dΤ+;����\���>R�n��"f[�l�}3u�Z�\ y9��~g��5Tq#��A	 ��Fʩ�j)�m� �J5�f������w1�g2[b[yx��(ؚ��������AZ?�«1���x]�������K�0���z�;UhN�J��U�S�;p��g��DTS��K����:7�pWs���/����N	WPkR$Y�ن$.����~o�ɯ(�1�E��*Փi���8��oY��Kf�˷�N���S[�LJ��P�0�Wd�9=/�6X�P���g��;�j��s�B��v���q��/~��GEI�s���`>?X���~>D��t�$�&0��Ug����hIFz̯��0�<<�IN�x��yC.}	� ſ�	��Jk�`�u�W�%X�-2���*�sl�_�}��EE2��'�
O�j' �&c����y,#(��It��o�?/K�cSԏ�U���@����j0�v��_�᧖���9�_�)6S��;I�fDg��qu�i��b`��O�i�4ak����No��vuD�*�`�`:����nqzB܃#B. ��|�[UMC��Ls`��aA�9�֏Hwd)��4GHҢ��ӷ+o������/ݔV�y�pf�7L�aC4���K��cV�q�i ���lN4e��$̓+�.Ptd/�	NB�y.ʅ߽���w��:�
�W*L P� q���?�ίX�y ��5�r� ���W��+�a&'�'	ɔZk��t�#�A�&0����W�|�=Q�s�#��
�j���������{�� R)�
[����߱��;�y׾�v��!�;!ĉ64�ᬻ)���H�-E��ڥci�w �1{�����O$s�n����d��������:䎈\���)M�L7'�yL���ʻ��"�f��#�#L.���p9���6p+�:	�~�ftzZ��W�*���ɊDl�'�e�[�ᡆ,B���13��F���(���,s^K"���=���.�G��Źbdܿ���7�$��h�pT�t�s5�6���n�P�Z��+�?*�|�MI�S��uhť{gK{��dd���UȻ3�y����"	M��E�:p!�
��ˠ�{f8^o�$�Dm�_�aӾn�X�G���%{����!��;P�S�+�܁��V�z��!�f51!P~�kg]:�D+�@�]R��C
�.L؄ϣ�d������V�+]����7�챏��&��ت���S"��%�;�;�m��d� ��~y�H	�&�y�!́]�Db{X
��A��7�+��_g�l�j���R��<d�Cf�")F!��!�ڬ��1�Q���o�z8�b�*�]	?RZ0�}mωGhLC���D�e�fN�g`�\�M-@�R��UBP� ;˴ ���w��u�-F��&��%ۄ��Vȷ`�Ym���m��O�]S��(�Zo��``খS��k��$驹�3ֽ�M��ϲ(�$��)���|N�g��2�w���
�ߕ�]	�,}���u� FMI��?8�D�[�"�]K�A2�+&(����
��`�D�!��f��z��G��j������(��Z�k�e+3P-;
������\����3B���^�۱���]���*=_}��W)|��Y?��[��v�3�+�݁�(�:~�
�5��z����b0�N�t�
f�9<�맼�rM^hSz"���hGز1�?����wO$.M�Z��)�����0Z#�<���$)��AiO��sΖ8�N:F	ϭkR�&땺�,�!�Uj�,�  !B�VŃ{�^�����k;d��B���FP�-v����<�?+��̱њY����$��t�@W�˜���ٮ�a��iJ�F�9q9���K�v�KƁ�V쀅ũ%[���1������N�i�|=�9#�$%+|��X�<��w1[w�S��u�N�ɧ�&O#�Τjy2�^�h*|{w��4Ľ��f�\�"Ѹo��q��U��-	>�i_�$��Vwz^)��<�`����.F��v�N�uAL�XH�h� ޕ��6�ր(�I�r�S���%�<�D�}�=I��h��4>Rb�fmj���ZNM�Ym�!#o�왫�]7Kב������%JƆ���A`Gͬ߫4���6ۇC�Eӆ�m{�<_2��&Z�.��w�-Q�1���|F0��Ȩ �|c�L��щ����e�����ϏL+
�Sz��%,��!/��o�����fN�σ
=5a').�{�%�!+�����'�5s
��O@K�&�#e�B.���ߜb��V�&���7�K��������(y�[�Ce�"$���`xa%Q�Ï��\��E�-���!�.i�-�9�&=CNy&��m�.�-ۉhB*��������W֛�N���>6#!�e����������c�G���ۈa�y1���%��$r0��q���t����ӎ�����(ЗUr����VIa}	��*�B�u(ȭ����CUfϼ.��i������<�S�e�7տ����;/�i u��U	�+��p��P�)d�<�p��~.�<��]����+��]�|�mgO�{� ���h,M���ie�%��lusG��d�|ʁ�Mg�5�^Fs;���O
��ͽh[�A�m}X�ng�����S��Nt�F<�l_1�<�
3R�ۘpn]��s�{y�:1-κDT��|n���V�����Y���U�FXjx����|H2�d��X]�YC�*�&�I�N���lu��'�u~��d����K��C9
�"Ҩ� #U;"g[�YB�&�'š	>�%K��1gO����|Z��&�����[�N�	J�3O�/�N]#�Ĩ����VVek*"Qy�<��6�O6Os'BRpz��Dj����X0'�38Ciu�R>mH��
ʖ���W����m�sպh��l�>,tS9�EΈ�������	|_.������� �����%��_���g��1�I4n��=&�rg��o/д��ߧR��L���@����6���lsJ��ۍI��&��}��:�w�TZZ'���ڻSwm݁|�nx�J�e/��Is&�1�~��"|�7��F1���oU`�}	�����&'�M굮:̍�-���̆9I3�ƛ��Qn�<鮧hiM�s@�:�p� ��3�ŃH$͛w���e)��Y�Y���E�y����X<x1�G)���[d�����G����YEb��1V�h�g��S��Wu���o�U⫶L���kp���?2���S�P��%x�?K3�[ f�|�����j�o��i���|���I=2m� |�*��BË�MU�܀RҘ�}�V����|u�lO��Bq�r+rF}G�QD�HsҒc;Y?F��@�4�l�D4�s�q� V-~/�M��ϺY ��Y��/@�${���h"(@��Q�_�+���y�e29�,�}��!h����l�b�['�E]�Y~���)E�3��|�	k��(�e�C�3 � �ti�v�g`U��V'�߰�YJE;�:��u����w�ӭ1,STg�[�ɳ��٧�E�v�Y6�ݯ��A��p �{S�c�s�@�o\ƘW:U�T��0��+���+xB�2�k���[�xx*ZX,��itk3o���%ʉrL�`Q#�'��c�ߌG���d�0hqqaa|���� �upL_�$7���w"F�K{OhB|�ECu,��s���V�m��?]j�l���e�YpA,�*F'WCo,�h+L���[�{�X�c�~�.�� W�L]H��Gtǉ��H�f
?7J ��C��e���]�����O����|�S�(���.	�:u�+Q0�A�J<��/��Q�X?`x�f:f�h�
�s�j�%Q�'x��i'��xT$�>��O�$�U�Er�s�\��8��1,B��Y	�
�6U��<2v�*��_�{����t��J�[B��;a�M���$Ñ��<u��а̓��|F?˯9�#Go��W����Sug2kC���0L���C�Q�~@!���e�u܈&���p�V{�|O��{k�?�_M��0`r���o�jX|{?���d��/��t?M7&H%���W��bZ�cc�NRAY��e��H�+ք�Ȟsf��<oo��s��Mj#����,�*f4V����>�A?��R�TǢ�m+
q��}�S�]���)��ș�N�P�M?�lJ:�Y�~�o͕���~{�yv|
/*;]Sٞ�T\��[I�k˙�5���dt��!<�1W>!L�QH8Q�j��"�44Z�L�WJ4�%>�:�>��R�/y��M�G��c*GZ��N��w	([u��G4i9�s�m+�aU~���η�PJ�!�!BhIc�/+W����i춫�k7���	1� �@Gc fW`^	8�A�1�Z(,ca\�%;��H)��.&ey!3�w�Mco��GL f��6q3o��Ș5w�P����d��D�f�Q�x��)(]O��l�M���j#�w6pys�5�����O�� �G�V]�$6�h�'�N�q��D.Ly���$s���Ŗ�T��!��/{�rW��j�)��,Y5�IEe�}4C��Fa�N����4�"�a�Ģ�lk׋a�g��%y&\�s�(b��̧���Я�2ˀԉ���]`:����n��q6ꝺ8$��K��Y�ٹ<��ł#f�������G��2c��x���z���_1�7�+�x��lmo�akӯ=�M�~g'X@*a�x#�W����	I��X[�j9;�;�1@����ĵuIjM(�h��_��Ǔ�O����amE��۰��c a�Ih��pϛ�L�'�E�>U:(Fn<f�uO��sZg)�F����4����Xt���4����	Hq�nM����������~XP,^��$���_*���S�"�͉���4����,�$���K�Z9Ѡ��}�i@�±�tٿ�O �����{l�!�f~���-�qD��$��
�-������ukD� QN:p�w�$�X���}����iJ�*��j�>���4s�����\9~�!e��3#J�7��J�q��}���N���\����L��	�׎�+9^G%RTf�Y�Y@�9᳥���^� {�we��׉~YВYL1�X-
���� |nY�=���!m~�=��.8�P�q."ǂ��5;b�v���(�������9��bG'c6���7Lg8�ӎ?��u�ۗV����9�-�-��:X2rjF���G��\���Q��(��f��㧅6HO+��k�Y*6aP�d*��r`p�B�C�|�@�~l��B�n�f%�����;H��ԟ�du�H�����d�k���lS��j҄���K���2��iRF%᭪�8�>����_�*Py��]8}�l��_����y� ��DXK���#�ol\b�b7��٬wgH6��*�u��= ���L�M�޴�<<���J�<�����4D����1�wo��v��2M��_6ȱ�Do�[0P&��&�$���I�W	'ŵ�
��"l��i'#��`2� &�!4+�e���"�ⴓ��櫐�n��J���`���,�%����v/�Ƚ�$!;!�_�����9�=�?���}Xz�L�)�\�/���>�����-7sN��%�SL�M�Fri։��j�2���q�"
�`0xNu�F�ө~�U��N�^Ԓ��S+���]�FD$�$u�^D��H�!�P�j���|N|ռ���{��TL,tM,���mbEy��O��p�W:�����x��6���)%�".�H����n-fg�$�oSfv�.ä{���?4V�L���l��Od9ҤS�!�ܸ�K+e���1?���ݸ���F.4�P#!�>al��9��l蘜R������|��k�N�B_��1d^BEj��ĨѲ��ն9�ӽK�}q�(<�@�ǲ��5��蟙�5�?��.Ŷ���e�ʹ4��΃p���բ����r� ���]$ˆ)��Z(�J��칋�i���Ʉ<:>�B�J��R���w߁"������e��Ux$p��]Iֽ�*ET�V��烌#��0��H�?�뙂���3�}a
�黿�O`�q��F9�`�noU��O=aҐ�\����h�^��ێ��G�$Eq�d߮N�������E�ө��N�CU�<�R���n��� ى�����N���_���R�~��^لU��)�)�lR����w��"/&�`�cj��kj�\͌�m��u01�c���+KՌD �RI�?�=J�B"p3_�>��41HHq%��Q�W'��D � ~@~O��fI�Y꺹�9�0ԉđ(p�'���u���Eo��ঋ>Mv����ikH&*U�/T�f���^�3��t�;Y�)��d��l
q����z����ZL�'���d#{cS�ڧG%�	<~6Մ�R�?�;�(���
�@V�~k=�;*z9�N����Q^I�O� *�G�,|��yn4��j�t��0�Y�5['��#��!�!ɬ7��]pJ^p��:�.��c;���d8��n�\&[pB��n��P������ką>#T�)��	ͽ�G�O�%���$���,�Z�E~�@���o�v�-��sA5I/�`^ &TN��'RT�SGq<Q9� d�����I�`����]V�d�q��ʚ?�"Y��'}5r��Eb���ri�@�!��X87��~x/���������#z����N�k
����X���3���ɼ����,�3�c'�Ѹ���-6 �Z�B�E���7������9��u��ٴfX�S�M��O�Cfu\�(�1�V�rU��kf�3�i�q��D��@CY����r�rp�"�F-�>iW����&q�F��ާ�I��>��K�����r���N���Q��x�H��/_�l9q�S/y�����jQt��&C�>Q�UlwЋ<����k�)�u����WRE�Cq^�vK� ��:����g�U}԰zʓa���2�Ĭ�N:�R�'�q.�n�F�t$���ot���̞�Մ��4�W��u�+�RU�����D��Z{y��������*�@�UC��z����mKZ����eF���hG�&��3d?HPtQ`��(��}{]�![���Dj`�h��_:V81�K�l+��
ܢJ7�5ç]�H����	�[��/XZ��m����h�����uR�&�_<_� a
Ӳ-t��^��j/�$|��cb�����!�j�8�������u 6���.5%�Z�Ȃ��8Jh|0�+��H:������,f�O��,�Xm�F��q��R��}Hֲ�^���,���t�����'�\�a�u�E4Ʌ�P^\�n�ߗ�sS\c]!��ڪ�U�	}��g�6����5?% ���7V�eTx��h,����ΌZ��3�+�X�05�J�zl��lN�?f�^��c����;}�&<؅�d$&�1Ȃ[)]ld����iWQ~����.t�T�RG�;����cgB�;�M	Ӱ(ޟ���yܺ(���h��C��Z�ySyc;�ʟ���7ڏt�Gf�(���UpUO��NCQђ�ϖъ��W0�P?��iZ���0���&�.wޒ0��k:�R���h�.r��tlI�Pa�f��
��2���:>��4)e��2E2.�۽���VW��|����X ~�
C���f�����B�+Ǡ]��"�x�����ERg�Z�-)֯Ϭ�{/�$rp��9H�Ɏ��+��R��@��M�pU��d[��CӃ�(Sէ���Б��DgC!{y<���l�#�i.=�+��M���ҕ:�3���������KXN���N��"����[r��4�<-�4�̶X�pXAj�.�:�O=��^�>�� ���H[�G�����K����z7�?غ�J@�K������˜(A
��ɪ�F�j�В����'��Ҵ�J����pBU�TJ>�y�Z�����k�Ӭe,��'6^�]J[�v��muvt��V�jx�	zs��j],qU����;�T� >l�a�4����G*O��J�+��W�n]Ή<"j���ߒK���m�2����v�<��'P7x�7`yF��L0x�-�"�Bw�+���U�Z�S}��_y��ō��Ƥ���֜�4���.��eʟ5INe��1�c���3 D�yO�T��*�>��/�[�޽���G�O�Բ��唁?@�T����%�Ic��H�Q���e%O�ͳ���>维����D�*����S/s�o�+c�L�K���=!��K I�6A�Y�����i/���Oɶ%�M������"I[a�R�ڱ�rU;���\6�UwJ=�[/M��4��1n��#�Ώ��eA��M��3���_��X�E4�V"LT�&_cK�	S��|� m��c�t�QO:�4\�pR]�<�`�̳�з�� �����	^���9h�;�ߩc�b<>`4�X��`�����C�,���,�ŗ>6a]�_�<���j���Y�����R<=IL�Hv�Ży�PVj�M�j<w��h���o�fg���Nj��w,��x+}��S�M�a
�+�y�u�Y
��a�@�Φ���� 5XJ�/5Ũ1<� 
��i6%~x=��e䚳md=v���z(ǽBݙ���`�4B����s�y] �[�t�նv���n(��������K��g+|mW2i/�kD����{&�t;\���`����DXD&����J���:5N<.�Ih�$��k~�Kq䖳�߬��[�C6�2R�N�Ģ��H
�W2+����"z��{�0�����$P�¤.��h"���!��~Z�#�}a�]R�n@��I'KK��5��+>�����%NR���^aCg��x�M3��f¬~���Z�'8
�Ԋ�T��6~.G����+f��n����Ux'�XK�Bi�)p�)�g:[��>,i�ON�ɞ��̽��U]�k+��l�ܣ�|��� ��T(�{��in��X��~c|iH�g�Y��Ȁ�^�~�ݫy��nԶ�� �0�ThU��
�&�rF����/���N�q��
��]A�.T�"���'�M5�� �%�x-��l�Ʊ�C,y5jڔ+W���3�Wo��o���K�����}�Ħ׃1��.�2VD'�熻1g�]s�O�T�{|�JX'�$ۚz�m�����ο��n��P���g��!X��������.,'��t�sj�9��;��c	�po(q,�M��=����Hy��^vFw���=��|����� ���>��V��>�{��M�	��SM���6<I�D�B���V؉lʽ���7�[�;r��3�����a9��Y`�s/+d?`����1�)^��!�7r�ڎ��m1��H�6�2��!c{���Y�/Q�:�w�����IZ�1;���qܗ��B�܇����\���KOANՋ��u��Ϭ���('X�s=�dW�1�E�p���d\2����0�0bIP:<"+{��e�N0����o���+M�����^�2�&h��!H^�|�B��6��	�s��eV߷���ʦ#�g_#�s_�l�՘�M��3T�!�ځ�;��H��[$�5h�Xltl��[/ ��Q�9�P��<m~�t�!�E��Q�` ԶI��F_���ť	h41���V�&K2��D�~Zw�a�A�L��H�3wAKY|֮�W ��] �V勽�� åG%���
/@�f	NG���}�Gk4������L��v�?���j��|����j�� *��K:Pa�&C^�����;R�}- �Ú�+�Uy*FM�k½VR��)9�ZA�4�sl0���)�:��%�>�Dn����������OE��h�_�8�d�s�˄�[</!�ePP] �o���޺me��z6(���l�^~���k��ι��?��x������7��m���,=h��<�7�|:��@�Fi}U�U��"���Gg���.ݬ���GO0���{�;F���ۮ�A1����3�����׆{�b]x�Mu»�Fz<:[T	�L�t)���**��-����`�܏T:Z�w�^?�&#��K�L��^�[3�)RYi�����E�xOdaJID��*����ژ���FGCZ�ҽ�fl��j���� SG�!�0�0�{�̔�f)NҜ^�A���n>S���yiV	맭1��vd�5�H���p����ǛD:$c1J�� �tؒ<�=����Toa��,E���3�1;�3�V�[�!̡�%�fh��@+��&ݛ�����c��\h�"���PM�L����+��tU1\�c��<�_�+N��U��2�N<�WS�n;���]�׮��m��\����vB+!!�~+�>f�,�]���?�*4��|*4�kxd��ψ�Q�z�=���]U?�˭���s�h/�2`y8���$����<Rޙ��1��u�׈)�#�q�C�l���0�M��kf�Ւ�ZNz�!��I��4p"���`�ƢY
���'�"�#gQ֞()d��ܵ�(�a�\�����WD��c)^rH���k��o	�[iz��PӺg��&)NL~��,[V94o��>~%��-��e��:��"ɰ;g���]����ңKc/�p�Ɋ�ˡ���ϧ�!V[������Wy��|�m�N@Uv+M0e��%J2]�,s�,�׷�P�G�ԊI�N��U���{������GsP�sk�>��^��ַ�[�E�"�r�����ʊ���9gBJ]q�Ҥ��.�2Ss�7g{?=���^���͌�M�����qN��t�����;�/!��{��Oy!JU�&��E�⇡lU�k�Y�;��D0�m��%[3�����K�
�v���gWkn�D@�l2�[���	�;�u��`�������C�O	g��v���F�|�)��^�� �0D��5 �x I�'�_'�7��|����K�v�����iK[+��2�*�z�G�� #�\k	��v������M<4���lHҿ�	��Dq2����P@j��4CEN��C��t*}n�W��v����)x�;t�U�IxN���}��s��c��"��1��0�N����/�k�tN�T���O3,}���p��H�����rj�&�SIWҕ=
S�m�����'?��;?���g�b5�g|pBk�"�\������e�� 
��Ov�G��-6�{A dNؖ×Y�3`J�-�G��K�aK�b��D3ו���G��j5��4�x'Z6K�ȓ&tf��ڑoBy��^;yF-C`�����(�te�J�����#7�%�ЊiS��`��_�X9���B���>�jsh=+K��*��ft�h0ݥ��uht2�ɘ:8$��C�obP��D~��{���Q�4�^��*$H�|�S�j�}YJ�l���q��R�ɾ]��>�k�v�>���""�gB�}�z`�g�x`�Djy�^�4���us�a�#���B�a�d��b��0%�k�a�R����mb�Q�~*KF��5*ӏ�PD��"�`�8`����?����k�^ �)�?���%;PǪw� �Ѐ���&�ŮO�L�Н����ur��#U�J6a"޺�J?���w�����`��s��2�����՟�Le��}�#�4�k#B�48B���>!�=��G��O��V;��x8���l�s���gih��r��Q��1m�k�Pj-~}-扒�Y�Y꘨�����/Y���x�j��m���L�w����e0	%m�rG����ˁ�M�\����Y8��6��dï�,�+�,Nbb���a�{��%5�D�wˆUBIrr���X�C)����~��}�;�T��4d����+�,1`�a���S5T���
U��rt�Aj麽ّ�Xn��.�G��T G@a���B#"�$�����r��R�+��U��g����_�¬մ�0�R^�����U���ݥ:̝O�߰-s�O��鵮ck�}����耘#���t5�	�#Gi/I���������x���&^bX�|����Ѩ�������ё�	N�
h��&A�����H1���b;�"мJ��h��I�v���`�a�㜢G���X�%Ъ�*r��T�\�E��iGlU�p�lfs~z�@?��B7����O+?�c��	9�X=�p�	�g�CN�Mo��~\5�gj�1u��V��oݺ_���wI�)Y%d�Z�66N�#��;�@E��h�T*K��ȷ���ER����� R���C�O�ס��$�*U5+O@ה3m�L���I�w+����Z��m�ڂs\$���̖VQ��h]_��d���P�U�!��P h!�w���=�W�!�脭*�$�˛��7�u��G|�ȍ!ڃ�e�5�D{oO����st���9NCG��]cy i�4MI �a��~�Ov���`㸿My�y �3��m��6�& ؘ^���P@��!N7�~uw��1�v�,Du**+�q�C�*9�ӿ����K񇸌ԋ'�@x��J���l��TQΑ2]��=�}�� RL�I�h��'�3:o��^�/��7�u`G�=|�*vu«6j���$�5�a<��|̧���t���ƭ�@̏"�,)&uy���[쭲r-V��]dt��r�Ԫņ�E�/�|�m��w$�O(y�J��~ok���x	�0����p��/Ȉm�YYV�>lC��A+�����r|�%�&���Q <���æ�c��GayD��+L���0 /4*^�\�����m�F�o�i�B�4^�>G3Y��[q����5沦�W\�( 
���X�{i	�כ�g��f��͓�t#���7]!A�H��U��.wz&s1O�	�g��G�l-�����#�����ln�Z�c��68J��6��Z(�3i#	�!u��toH~�<
�	m�U�Ȥ���"�H�_�e�x��ʯ�ֽ8��Ta)[���M���Rx� ��d��О���q�k�f<C$h�EĚD���>o��&  ��/�P.2Ѿ��	��~�%~�D��P7#�tNS�O�|���[n-��|/���|z��pL���,Z�\�F�@x-_�.����9x!�% ���o|��2/<��b���Hc��XhB0�Jk�Ǆ2�v�w�/s����\��0�- �$SW>nX��j�	eF,�	I�\��x���f���2s�h�_b��;�ɤ'[�6�qH1P��̙�R�(�͎�=�P2��h�e&�G&�>Ս�D�*Q�e9���B$0�O�̏t�~\Uq��+G�-�=Z�:�uw��V����x}��;lO�Q���]�o����T��7�Rƻ��s"�W��{�g�-JFL7�3+�*��d�0r�Y嘐1�b]��e��R]�y�)t-g���$�_����ptT��|��M�_�����څ�9|
�鎑uؖ����RP
��G�����j��,cQ�d���6���>����i匁�n� ��������OUB"�?Kz@t8�]�h9���$��v����N!�3�ٚ6D�F����j����Ou�k��Y��lʞ�}E�n	��_;K�"E�*"]�<
����:�m�������(g]	@z�~�{s|9���TC�b��*�h���נ�:7����'�No�����S�6��-�׆�|�U��5_GY��|aP�m�����%52���቗'3kzYcHCŵ֢;���i\�������(*�t�B��w>�@-��~m �0�%/�F%w����"�F��#�<-n�˞�NS<��7�L�݂��(�@ϒ���⚩�,�U��>3��$�T����������HQ�m��J]z�@��8^�j/�}5<e�v��W��[y�־L`�=�Bb��u���Vc]�)���͸^=�K���[�~"���E`z(0�+�G�	64�Cq��p�eh���X�:*���Ϗ�!�o��p�C���G�Ӯ�p�⧂��%2��Fc�>�ps��oA%�~��:�����r\/ρI2���ФZZfg,8����nܓ$J�a�#��:�ә�x.����=Buy�u
�@W)��w'��C��(����F��=�B�f��(	�лjp�� !2�GO�j����b��?��l��sZ�<���M�(�?Y}��x$a�t;l�X/W���/�����b�
����^+<W�S�������/q���ëU��B��!Tyw]���Cyu�k\2��y9��+��� ��O#���r!4.Ud1���\�ڀ�_ξ�\�nCl+��T ��!b4�)ʢ��E�}s�j�:x�nXߵ���@�M�`֨��g���|d@`��@3�p�>�t~�o� ͋�kV_�X�#c�qF6�f�00����^HB��AC�-����j�S���:���r��Yw7s��<9�h� {� _�U���7���8/�0�s��S�ޚ@�vf�H'
tD��֡|��8�*C�sɱ�ǔ�"�,�I{L�{ݩ�i��㚵����]{���))����'�ƺ�螌a\�s��^]�M��`6�[�[{'7��t�w��}|NZ��  6SUK�Fvn=G�BA���谿1����ж�E�N�8�<� ��|t�J�:�K���#��`>	$z��>�Bc�ZO!Om1����5�N,��~�9�HdOss�	&J���!O���3a�%��*�|Z��^�:/V��y���D�cuQ�3T����QL?�)m3:L&e]@�#���¿)������a�����'P��`J�h�sy㾤��^���Ǝ�yF�qL�ͮ�3��IX@���8�W�����4^hX�8�U5�<��ܩ�ho"
��Y�9�x,.��2��Z_qi��ٔ8�I�><��8�6�����[�_���y}Ƈ�R����y�a�hY}}�A���}R
�[�+u�6�Rpi pb��&G�`�u5K��v|R�1�����ǳ*��I�QH��HM˞hC�JG9��?�*m�,���U!��i�q��9��zUr�ԌI���W	؂��p�:iF��IV�>L?��.���]/�j7郉�k��𻗍��1^����
���H�<��6��j�x�]w��)n�9�IE���胥�t�TJ�ѷ3�����G�r�$2�n����H��V���8���@t��ؿۥX�8�K��uO;^6@���zah��?:���d�.w':��yO��������{��I=�Tɨ�8��rd<�j�<96��+_366���- 6����gT�y��G���)L����b�H�찥`�p���S��^Vт�-�Ö�+lW�I-^��8Psp{zĔN�_�1am
��U�d/�2O�I���Ac�g0|�ږ�α�?+(&�c��%�||�ND��m}_��\���4u��o�-s��GX�E��7��6<#�H�"�$����8�*p
ǰKq��i�yQ.Ռ�=7�Q�6����q���$՝Fbb��kc�W�`� ��"@��x�Z*9d�9�B�A�qo`ή[�\�
���{,��|�P��N�Z��⍄�	1�8�b�M�]�D]��y?��q:,Sa�M�fm�JJ"v�a�� n��Ѥ��~H��F������"��J]}%'|mI����ޔD^![ )A����;Mmxƨ)��h��k��X��@��CHG����m�Lr�ԏ�J6����)���\:c�-;M�6שy����hŃ�\h�?ӅqUM. ћ]�٘Z����Pf�z���r�#��Zi]�:RV��K2g@��9I!輦���*5ϴ.=�� Y��Z�ge��^�3�"�JK�Y�q�38z���x�����]j�њ�\I���|����MMC��g$����>J,���8ٷ�2?,�e��=r��U��� �
���[��DE� �r%Nq#w�`��fVn����p���^/�/V�oh�	eF�W�t���R�&����PN1`�b��"L�`e��>�v��wj<��?��Y��|�?l�-��Ex̛<3����z��ߑ~h�G�W��v��wqN�) ���>w皬�ɴ�,�԰'�T��)��d���X󢛌Y�\)_(bnݰ��A\d����ϋS��%���kjyS�kUP����!�E3�/�!��Kir��a�C�J��\���kXm����z幘��]iHز)R���q
L6E8�L{G��j%$��Y��ީ&v�]mR�H:�LUMX��14=x�S�*�6ӧ5�A�Cm_x����g V��.M�Hl���u� �c�������q����B��qW~��kI���
/,SK�+�y@��X�ܽO�X%�*0�@䉚;��P���q���D��!n�Sot�5&-�'fPAX��"��Y����ޘ�:=�$��o�A{�u^�7�`�V��D�0�}Ku��S���G�{��@]5_���s��\��c"�K�[$u`�Hʄcd�l62�r��H�qj`����w��O�����)��̨l����ӧ���/N�1��h�!��ыY�7c� 4j�R�+9��d,�jA��-�@ E�n�Dɡiki�����:��.;B)� �Rk�R.n�M�žP�2�����S��RtI��R��A_�6�_qu��o�_�r��3ܠ:�����B��&S���=�� Dx �ǹ�m��G���X|x��7����e� �-.� ǚͮ.����܄�r7��ּ�-�!	�u���ĞT/E����e��h�ld�:���A���w���p>s�Q���ba�G�"�8w�9�}����L�N8�FN�x�n�Jy���)����^3�3�Q���{|��[�j�Ι������1&�� ��KB�M��پ&���h����K���]]�Cx�̙���C�(+�����;�xڬ���G� x��~�P)l�����⼐D�UP�y-��K��l5�3��1��^J��h�R'��c���Ə��q�)�!���Q9����9�L�ZC�g��zFATh�״���<�Dv.�7�7����z���~��Iɹ�=�������]��~CxbKl}�O�
�g�#;	�W�m�����Ή@���To�F��� ��hC�b�D����̯4���5������4J]����*���_#���J��C�vbCz�GW�[V38�Q��̷p�������Y~��-E"C�}f��}�~�t'C����޳�E
j�҉�#�`O���'�r`:ESQ�eR8�9�D��.�a,@�I��a�U�����X�M:����a�;TecV {(f��;��l���/�*a�q<�FB�s�5{���vf�r%s�""&]-I�p\���yS�ˆ��G�g7n�<�]��R��~�?��}c�<QڌZ4���V=k���rk�\w���2�i'�P����ٓ���p��A��bR�ۻ� ��i�3�X]NH�jk7�Za1�&S[ԏrP��d�G��.Q���l�X�',~��iU�F�(Z��8~���z�F��h���F�w5ۊc��� G�]�v#��+��Ӈ���ķUϸS�Vo�̘���:����v1��л��u+�%<��y�-Z5!����2&8�闸���S�'�Z�Ł�?AϘ�2u~b3!x ��{��LE4�P�Tf�=7z8�h/T���
�J�F�G�F�u��3�i m��wڷ��^�O)j��U?�K&0L�C���A� �}�	4�bQI^�S����k��9���)�;���L^�i͓��@	��Ӗ�4�+�Y�m	�48�!����qE���e*(t�,���T	���gX��\�GRgch�u�ā�Þ;�����n~���3r]&R�W��/˞�}���B�9\�aD�aϑ{��hx�����KO{6�nKY��}��%θ�d+�	
#�pL�A\On�z�763t�능׺kz��>�k ����c�=	�SJ2�qӲn��u5TF1���~B�H�8��[em7HƗ�7	�_�����������Ѱ�Y���A�~#9�X���ֳ����Mm6n�8�0��޼���x�� S)���"h!��C�'-��v�����Jp��h�Gө�[���դUd���x��u�m���B8������!rea	�m�����r�,#Mx��u^���8��W�Y���1��Ȫ�����p�k(~E�w��"g1�3<�o��9v1�H�s(���@+{��{Q�1��(ҫ �n�1��Cf��o����( 6d:گ��4�[��"��0�_��;'S��
���o�A�
\]�v} 9Ϫ�Eۅ>�T�7��Q�v]�H�x����Ţ�Q�ǧ�:F���)��M�w⧗��*�V{Ոc
�bG3�4��j�����\������&�V$.O�.���0z3Ӣ9������������&����N�(5��P�s�����R��K�ẈN�+Ŧ���а�h��(�2;�amn�	0�� ���$���݄ R�L�z}pt ���g����'��v���F�!EH�/%�R�����Vr0�ѷ��۱w�)Ō:G̖�h��:�"�'�f�c�nQ���\�!n�������)L���|�rtAr��Ĺ�	���b�\5�V (���y�pv�)2�)9R�T[I$xi�GjO��_�6I`�i�9�$�:�`��E�,�@2��K�:�!�x`=%�IX�ܚn!]Wps�� �O�p�&t��b�%���,zH!Q��->HM��(g~h5��'����)��z�:�B���[����]�ѰG;Nj�,yK �ʎ�P�OxO�f*���3�EG�6	�Ц"ٵJ]�� :�v�#�q�����	jV�<Q:�\悑�[�0��)UbǢ��R�w�>��A��>�A�wP22���mx1w���vW�7?�#/���.�8M��G��62ds�I`�ۂ�T��Q��#�=i?X�,���u�)
�q��۶+�BI��؂?Z���L�StnDo'��Pl�7d���:�&jJ��<6*�ͱ�HkH�X�#���q�QJ�#E��ӄ��=�ү���Q�o�ԇ����O4q���P%_��i�&�@�b�mX�{��y��<��N��7��K<���
���v��Y�w����޲�d1�YVv��Q&�硏��U�����	�p+ĵ����*'���h։�P����w 3����uq\$Rw����d�d����A��ye��+u|L���͵��G���M����(e�߯�S?9&��;'ԠɌP�y���$���~��d=K�t��i���`���W���L
�1�r\kxO�!K�y�h\�	�*Y�S7x�R��E\�\:t!��Ն����;m��=��^8�*P/�nɤ���qz�]=q�]|��mfs���[�8���M��/F��ȣwW�]]o~	 lHl&`�d�ymb�15����
�e+�|�7��h5�$I�kv�G��N�9��{�C -�� �`7֓���.��D���И���\R�-3x����|,?���w�ߟrNR?���sXƽ˲�Kc��S�bHɛ>P���iu�l�D�dkcnt�vwr�Cl����fp���V
C�+V.�pv�ܛIN�CG�5͗߰��E0l-Գ{�	�� qN����m�S�(V���o��{Y�+���Ȩ�S������qm~J[ۍ�x��%�� ��B?H���[|!��"���ʯv���@tΙ{u�"�!���e��#S ���H~��?�@ ��BPE�?�?��U����QtU����b�!�[�2��Z��ER=��M����S?�f[I7��"lH��1ɡ��\���V�j�v��W�Ý@��������o��P�C����2�;d�2���d����p����	X랩�v�Ө/ap��d���9
<ѳ[�Z�:�=�mz���!�d~C����-�uq��*��:_sr-����Oa�M+uJ���/��m��U�� -�ʞ+�)�6�"�3������oX`�m�Y˂cך&����n�x����E0>Z6N*8���I�,��Z=S�+���aG�ȏ�q4E-g����z[���=j����b̨MN�Vf�j]l��+a(^�C��������?�>����W���z�.��@l35֝!�����%�X��H|������.��:�Dw��J4 ?��r$cAJ-�fQ��zJ@`���pc�.f�Jb�gerq����"w�е��n��V^�8�Ӣ~!�R,�П;L\>Q�+�~Bo��4�0�-1�"
H��XC�