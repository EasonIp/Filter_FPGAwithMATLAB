��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�J��"4�=�7(�T�JѺ�ő��,\��s���ӣ�F�؏B�v1�fR�Q0���(�>�//�y�-��S\��n0��!�a}��T�Fk9����������3�^��T|��] dl�M>���+L�nf��F��j��X�%�R�c��@���/���t���(�xι�Zr<�L��DN�3�T��{w�WYDmhgrQdK0( �׌gc�t<,,����� ��DQ_=��ێB6��˞��;���+���%4����� �����$F8���D�U��/� �ׅ$��p:��=%s/�ǀ����{
R*n����uLz�WC�*���hG�A�%�*,<��Z�ry����t���$��ǊGS`������T�z�`�["�r"-H��W�%�vy���%����>o��+!���z/����M�0j��d?���Y�:$��_3��;��/�%�c$p�Xj�y����vO����_��u�ќ(��vӆ��$=���<g���l��g����-`�/��=�2 ��֤&�@�J�vM3V����k�\��ۀ���!�5?�V���_��c7�9eSA�55�i�;I������}3��m!��o>�yI��!�+��՜�4�K�~_M�"��Ml>���(qd��@�X��*�?l�|C�1�:HCT&�F��v7�^���Ҽ���:�[��,��@iKnin�1�ϰ�{G�\B��#�ಐ;ks�w��s}�H���Z<	�k��z(�+���:p�fO����^�5�n�X	�;�5���u�(ʹ�;!@���T���A,s?�%�� �}��ˑgm����'^`/�N �+5�u���j�7_��s
!��g���%ٮ�D���	~���;���dU��f9��:u0{�o�����O���_-c��n;�Q�9[5���t�j����������-b���p	�^PKC-��Q��˒4�2�$DcUD���E���P�~Cؽ���������g**�4���뎲�8��1�U�n!}�ɨ�)CR�^
�u�6E��>������	�^�S'���1·ds�Tл{��6xM,w�x|N��S�����w��쨪J�����2Iy8K�p�]�o� ���nV_�C����%�OYw��xĚ�X�\�m��g�(��)�{��qW*���y+@�Rۍ��u8�G� ʯ�÷D����Z�U]�uX{SAWlX)%�6=xN	h��D�1�Ep�&���WXfC5[e��7E,�Q�A�T�~z=KE��	�h��J6�z���!U]�!k�2�`�J����c\��d��4 ^Y)���9�fj�Y��f�����M��&�pZ�/5������Q��{��@�g�v�2%�pP�!������g�5#u�d=i��(;Gk08���������	5q"�z.�l�Z
3�K�����0
��gJw�%���m��?:��=��j%|4V�(D!��JӪJ�l��<���s�ܚyy��n����_7@}�7�<[��qY2}�6]ۃWȊ�>��*���{����4��4���	�}m���[>NvA�T_����acaĮ6�42���Py�Q����nk{}6�zzw���8�&w�D�&��D/$#%�%~�P��P8Tӻ�:jp>;��Bzy ����
Mq<�?�Z�t��A:���sr�	]�r9�E���5Jb������P����iP&��c1t��5�G�7~IwpfYìCM�/ȫh��q�7��DX���ՄxZ�Ǡ�k��[2��D����l�JK�Ԙ+�	U#9�?�򕫛�������$�EDc(�C<m24��]�p�#�|j,7�����n�����i<ܳ�#*�����| ^w!}��v��U[���K�ɯA��8g߹Z׉M��	���d3b"V���k� pL��ߺ�奪-�E?�-�L��-�D�&�G�7&�b��"m�n",�s7J���|�"����s��<�)�(�R����fXT4s�[���`8��^g$�`��8)���+���?�x����Q�q�Ë��"�����Q��&X' �>=���(L*Ám`~�����bW�o�T-������<��%�vS��Vr�6-�U+��AID��J��\�����Tc�x�Ry;�,(r�Q�E�N�Tٔ$�O�f�X�@Z�j�D�G�]�uP%3�+x�iсO�|��kV��a(ۏ����D�_��#@ �m2�����&u,3ׅ�?�� 9+fI�G@����:��7��5Ѹ�݋z�+O?�g���m}Į�}K��A�c���¼��dnx4�2g�w`z��ۃ1��;���L�ӎ<� ߎ����+�'�����V��3��Za�#�?����+O��	��M���N���Nh������~����S�
E����̃.%��[G�.M+_�<e!{hs��B�7��c��r	��6~w`��rŪNxv���`@��i��l!� �����(�
���{�:O��cKw���Ef�����$ȭJLh���[���uO1��cKx��FD�yr���׫dY'":u�����K[E%wE6��[ڰHh,����sn+��hc��:Ea�F�������Z�IO($)v�_��PQ>���p��2ok\3�F�j��<Ý����ض���d���8U�"��m�O��8�KRO���N��vIƦ6��y5ڄ:��B6UQ�{d�K-%@�J���i�8�fR�[����h��C��;�z�7p��;��9��G�����\?�SD����H��H��ֆ.�����%o8��pެ�
���	�G%PՄI��p[K�B�i>�����$¾�ަG_B]�[�\�"�"�~M����N��[���$>X1�\l.IB�V��Xb�ңao�k�l��m�ed�k�� ��_Q}�����Y[n���V��,i�'�C��9���&w���'2��4:�c��(��h����5�D���ɋ�u�	~k�֜�ְmbY���=�;@�B컆}39�|���y1���ļ86Ϙ����S��>���Ս�́m���%I�v��Y�/t@���ir�t������J[�ۤL�L����VB�F��d�4b$���]pq4��.��O�����Whu^�
gjrQ ?vK������M�T� ��N�%Er/~��[�g?:����g%���\�'���m�ct&�h����d�|�->��8;�$o�^dOhB�$_���|����V����B�4�Z��bÐ��b��\zʻ����3	(U�_"L����C�KC7���n���]`�Af�="m��Fm��G.rV{��5���̇�{4ڄ^ä�d�R��z�L(h6��\�RQ~M�1��՝Y�(��\>��?
Iǃ�h�(��%܌尺�)um,!/9-1��'���o���0e�b�(�����q�f�!	e�GO"��
�WN�|��Iѻ�e�y"�o����u~��������UP!�:��SR�(��ej|��#(Ww5s���2��7�0���`��m���+prc#������}�"�6|�cd,�y���*��o�p�{׭b�I)��ERf��Z�p��A
����
�y�W����r�+`�,�Č�'F}ppZ��H��p�pP\feǣ�:-H7�
0�&.�ۅU�2A~�YT�>��g�+]$lے��qu�+�W���5"_���>&e��)	�w�d����~5���H�]��N�>zU�
ޥy'B�4=���2~�*�z�_5nZ�Ku��iܩB�Wn�p�����F�1��Ә����	'�˒�B��W�F{`!�N��&�ګ:��a��7�`k�����9=2�d��묷,���O������.�Y���/D�I�fZ���x�|n����(�iK���ԥШ�N�:珋&4�{���>�<Hn8�DǾ�A/��xg��rB��e�O���P�<,3��.��~ �T�I�Ϗ�D��>t'�U���/ҷ��%|���RY����vs�������M��f�T�1�}����e ��>nW]K�����˻����	ZC��A�3�T�?��vx����H5yX��n��z��Os�E��6�xw�K)����!���^v�&z�����K�N��t�[A��N�7�iE2�h~��֩x��0oZ�J����� ����d"��A�v�߾�Ӿ��IzGr��c
�
��4�Cd/ ����0b"j+Ԡ�i�~�2�1�o�T��L��ϟ�����U��.M�l0����!R���T�����A�;]�G����a0�����ya��T΅�k�cgUN/R5_E1����Nxsk�kKf�_�:\֨ן/%-#����kV
�����y����X���`�
�ſ�x��[����|��Ķ=�.U��q�p�Գ��![�Ĕ�U�	״�E�{�|&q��y�:I3#�b���qܶ��Kg[�Q���t�(GM��/�n�$��{J���S����x[�)ތ�E�J��D@8s2�������2��U��ӽ���*����,��f�l�qW$_+��;��R��T�h�64��l�YÕU �`$����C�
߱u��c�-��-����0���iq~����Lsc���\ڳ���c���ę;L<�e�[ά�ՠEK�~;C��~��dJ��<�4E ?)�,�j8(<�"$^�]�q]�N����=B���r�tE9��[��fMv����ӣĞ���y�B�����(��H]�^�ɴ����@E�Fr�.$�Ԥ�9���oy�Uط�\R'�Ƒ�l����4 D�Π�-��Sy5E�uٝ�+h�)C=��� �MCN�D�w���Ϛdj�L�K˴����|�1M��/�cs���W�y*���>���R)�]y�c�yP�}�*��߯l�S] PzN����m*�y����mP�|l t�]�E$h�^Rk�^�4W���u5��m�؝�<�%Q�fo:k��3t|g�((���FRc,wo�f�=x]��$Ɛ�I��`�9 Cb�-p�'P ����3\G���-A�ua>5Z�#��;`'������Ǔ�`�n�c����B-Rwo�}N�� �KR�z��Q���5-XKeE��������I���m̒�F;{ip�<���Þ�ͩ�e���zmK����ML�ާ�x5�Y�Q!bM�<��ȈvQ߱�R�����^X���*5��.뒥pH�W�`���г��O�t�� jSMy>r�G-��B4�<@߻@3�Z\.�m�8p��T��U�?���=qT�G'�<jF�NA���0�q*�̒�AȚ�@�tk�0 �z�L��P�Vp�R��w��ܨM7�����-�C3,M�<2�Y��|�(/�tp}H36P�29�*?�(oR$$��I�L��g��Q��-! ��=W�cC�0v�,;��>�%�Y��=ܑf��-v��$�ѣ@�q5㣠��*9�;���zw�}�����%r��eqI�.��X���j�;�m�Α��������K(ۄ�ጋ����l��u&drAiC!܂z� �}��&e�S�Y�xj3~U��]�P����kZ�|�2�Ⱦ>��sK�D�˂���-E}D�:��9��T���0�6�8����y������)[��Yў}I��QVP�7V	_V߈�Wm�l!�&�C��%ȸ(Ig������u��2�DPM����<b�Ƥg��FV�g���2�b��}S)��K��t��Ṡ(�)M0 �QN:�U7G��z��kP���L��׿�ո܃����rCտ���Ƅ�XkrMeBbu��`lA &�.�� ��]�=<���%�������mOG����bS��XT��')��+�@������Y��S)i
g ���;
�2�'����y�|�ϮC�l��ڌ7�	w��B�Ms�c2�;�E�8ֵ�:���P�	�4�zmb�v��¨5�,�Ϋ�f�,�
�(fsѹb1"�� ���h�����!�U8��7I�ٓ��E�M���z�M������.��>�7��W_�黚x4�[�1��J�V&qܯV�����$�
�A��[Y��q8�'
o�8`�s�ca��HN֧j�1�.(���9� �����4T���cQ_�0Mw߀w9���gՊ���d����N�tR��e���9!5�����
&��3Xx��L��Yg���՘>[^0��D��k�R��f����r��k��3������ؽ�:>k)��yW���E��_Fw#�=u�"��J5j*����9ȫ�Zx�T��%�h�1�
/���-9�|�'����M7��>R���B�b3�eK>����O��e����an���}�:�0�\��~Ic�$�/�&�V/�Y]�s���o|��E��\��D�q;8���R��K��$��*i�p����\�a��U�t�CfZ����쑺��([��,�e�?�g/�H�R���0���+�؍s.�+�7�I��Xk��j?��=?	�$&�b��]up�� \S�:M�y J���8n��h �Y�Pwl@����@}� C ��ر�[ǓH!�h)ag؃�uY	��w_N���d���.�%k�B�)r�v�/�@��q��������D܉Q�ö�I��,k�?��	�3\��Y�Z^,]�Vv:V��j�g��^�;���y�8�C�q�]5k�)�����3�z���;�TW�U���X�J�&��o����x�z�_{��b4N~�D1c��z	�J���Ό|Xb2�����,�&j��<�v�A��fyü�:l�����-��0����D{����Ң3OX�`a����f�2�ߜо��x�#�H�u�-�2�t����}��I�S��n 3�h�d�''�	TI'r��H�g�nMI!���=�,��nܚLģ�R�l��#��H�C$o��ɅW���������l�wM�tw���Ӡ	g���B��P�o�e���Eȧ��tr�j �����$�6�~{A��\"�ǹ���mwxB_.�z�CwQ_BDǖB��]�Z��h'��D��窥F	�1��Bs��u��G|��]��%�/�aJ	ȋɈ�v�/�yc��	J �+���	�x[	w��=#�LL,���2�	3/�B��q��Itꍈ@�/����A�T0#m�`�0��/F�^ĉ��NZ��{M���$�I������ ����ґq�u�Ǫ;�ʧ6e��S���cfy��njS,���WFH�p�H�j��Ճ�Q�c��2�8v�ȫ��g؏�x����c�b��M	�8��t*����M��� &�z3{bk�({T֫�Gt(r��tL ��i�ke#2�!;S��+.q���T_��&�� �"�{�a�s��D�H+���4C��M2�eW�s���d�y��K0���W.΢^��
�B�k�nڰI�;n	iR�*����ey$�ΟBb/�)��W(�;k���U�B�[9�30�"�����hd5,�1�L�v����rVd���Sˤ��0�u��o ��ǛY�,nD���F5{b�(�X%��j:ו&7��A�7�; �������#���t8���)gH��\Q{�}�Zc�"�ϴ��Y�`��q����# �W�;�w�+r������µiC�w�o����G�9F�I��7o�jV�<���HD�b�Y�d�1l�9<��X:bK�/oHdnt�VH��I)��H��1=�\8� T�}%�H�#C1c�`��_҄��!v;��_�:�۲ g~m [vZ�s�>"�Bg"ʬG���h�C>��e��h<����A��Ɩ�z�'}�(Ɏ15�X�I�8녶�u3&Kb��r��Feo����F�e�̾���C������$��[����:�� '�T�@�]&,���R�����:��2pC��{��7�����]�9���t��|��.Wz������}���,�Q��d'�=z_�:����:�$̞p�<G}�T��V�x��u���mCI4�J� ��s/v�*����0T���z����IJ����-����l���Ty='1�`��3fgUp2?a�4�����k�<oP�UO�2ъ���<+���t^�ZS���GJ��Mq�<Ui���H�x��J���H�$��1ʔNS�UZ�C�O���<$ �V3����C��n�'��
�s�GX�H+ᔔ/�(4� ��?��� O��I�"h��������W����-������,�i��2̇�4�K8�}�{���vÒe�0��0�?���`�a�������&
b��Xq�jebT��L��V�*����6 j�Qχ'"4�
o�E峳޲C#�"��Δ�+��@4�kS�S��|q��2N��)�ɘ����٪pd�#ˤF�x��?=�gȄ	�[>m5��K�)���
"-���Ͽ���k��һ-�74&�,� �H�Y���$e��8������v1��|h�I��V\�34ք��O�Dae���'\<3Oǯ�6��\m\ѺO5(� �0E��Fh�����-!���^Fs2���ܤWX���U�b��R��6�U3�嬑n�}�%��U��^8�="�bՠ�t��&���3c��]@{��R��L�*���Hѩϭ�!T���Z�T�r@��C�kq� ��9�Г4�5�n�c�U�x"�.���A���#OKa|K��<R1[�����O�&�xI���O�SOoc�
s.�Ȋ)�1%����?z���7vk	��Y�U�T� v�s����L����Pb�������;zعV���P�Z����jM�;�{�&�i�f���b���ZX��C��ᬣ�!L+�`������;��i�\1���G])�T4x�-��i�N�H�Y$Hj�ںk=O�ejm�Z��8�c	<��P{ʊ�
 Xq�Y]Qsd��vt~.C:�S�W
�ǳ?���B�D*r%�� ���{���9On�D?/�+Y�\�5�B��l�l������g�+�b+UqkG-���z�w��;�cK{
�� ����E���_6mQ�6L��&k�tN��Ԣ"սZ����_�=���&����_��?�+��a��)����x/N�V�����KbX�̮���I�E�v)���d��&]������e��}�d���X'Kzewސ�_ �BǕ�!{Ŋ�@�& FʌASv�{� d��N��Ś �J
�fp´�:ȏ���G���J]rtf��PR�x�P��J �H��&R��]$Մ
���W�MP8z%�J�H�U���U+��+rֶ�D�ʠZu֔eA�Y홈����zSMf���o���w�?������t�&&��Т����K��0qhd�qT���VX�=�xb[��:y�P1Q��2�=fX�L�r1�>;o´�+V�+������М�蟕��p�� �6x��
��$M����*4��#~DG�~�p���	���[�r��#O�Ȯ���v�^��54]4�6jZ��p�/[�u\{�'�2��ʝ��������g�Tʼsy�Yh���{b����杕�|����k#��;	�H%G� ��G	`�a��fd��8$o�t*�R�K��h�l����A�Y�9ê�q���1��9�M`H��5�2W���/ ߺ җ`��רW)��ך�Td�gXB>�г�h�(]!f:��_�`ɮ���>�o�9�a�\ l0*u����y�]v<�E�5F;"�������7�C��L�pQ��u:�.��g���l§�t3����1kP�Y���h�a�o����D(��.&�@$��3KhAX���;�dJ	,�Y`9
6�g�vh@:t�l8؜��7CA�<\H�AB��@R���t��Oir3��T?t���5�VM��:�.w:؀��>X�5˘��a��5�>���4� ��|VJ�@�����C����\_�L��ev6mN��]ѥ��B\�Y�5������@m�dZC5+s2Ѻqx�?��|���!��QEf��	�C��z�M�G��vF
�5H
�ǅ�W���^�&����9��	�$��tH�Ww���1�7hY`%���]�w"�-3�o� ���(q���v�ķ*�&�ݞ�
2�z��&8X�b�q,W�q��T���3K;�2�țឧܚ�"[��D������4xO��u:������8�TJ�\J���{E( =G]��c۴�8'd�9{���c`��%:D��3,k����D�����"�7{�?)��܁>s��d�HA�c������v'o�j�(AR�0\s�)9cz�D��g�#t5�ڬ��)�:$v,6@�d��(����Rl7��n`�Ky���׉���(�m�We%g���|	�!k]�fX�O[ .�g<���:�|4ܒ`����D">��H�����+(#�p��i"n
a���D��9���������Kh�B��D���G�cМ���8E2�*�G�6/N���}b����
��"t��<�{�ߎ�?K&D�SB��p��2���z�u��V����m]��x_�v�%4��j}�B��?���#��\����5�� �S��{�(�Z�v.N�ᮨ�~Mԟȿ�|�(����vz�hHv>)ZU
�[��I��8E�Q�B_y�_�REu���33![-�J+4S�i,� ��Rb@b��n2<�S.r9�Gٻ��eY�-����-��R��a��6,�); M�Oo��<��v�5���v2�i
�|�"��K8�R�a��px��x�7�!?1�dُ�*��3Q�������#�ۡ���G��Ϡ�!�v����-9�9�H��g� �#�GNB�<D��I��H����j�_���M�0�SUi�l��2:�{RN�8���lA�lѵ�/�Hd����8��-�4h\���Њy,�����Yy5�.��xՖ�5�����4E]ဲKW�in�$��i#��E^�/��B��u��Z��;^YuR���[��6HD�����K�����L�n�	"���M�4l,=����������Z=3r����� �~��j������r}`q�y^E>w�w�{�"�7�8;7Y����'���[��/�8�.�l�	.��0�1>�.�j|�/7߇��LS��\pWc�5vl�.y�~�r/�2o�$J��wAM��*���S5�&r��3�l��<w� �|t-�Cs���5�U���UT����k�f��ϓ9�p��6�m�M+*e��<����ū�q��4�;�7]����W������S�k½^�@���B	���͡Z�0�����Y|�ޙ���W9?5$�"<�4�6⚀����ښq-��"��4�t*��ػ?�|u�J��\��Jy]��z!�\�D~e����ztC�j��/4|��W���;��K왙x6K��	sz��oM��/���n`W�IfӔ�</���@��7�x��ْ����SA��[PD�+�a��=���ՒC�$�|��Y�Ï�`��2��A�~3��=�8��" ��F\R(�/�6;&؅5<z$�@S1)Ӎ�M��mw��K���T�wlɿ���g9g�dM�s�}�:rMQP!�OU'yO��J�][��>M�-�4���G��;C-bc��5 �!���r[b�����ҍ�U`�Ҳ&��ɄKc��PM�ɻ���׮c
���(h��U*�ў�$� ,���.\+X��G�[�8K��H�D\�A�}�A�G�?�k$��%E`һ���d�������� �.��J�<_ڄ�rꝝ��~�֣�]�_f�(�ڶ�ns\�G5?�И���b&�C�8��(������i���A�����ų�����i��š�U�~�(=$|�����T���B:�Qt&�eN�I�ͦ���
o4q��ћ�^w,|���>���C-
�4��J"���C�AbRm�'���e;���Po>^���E<}Y���'Ӱ�o��a�/�|*GE]x�b�ى���:�$_�moNg4>3m�/���z�R��h��u��5r� ���J^ϣd6�ټ���r���$@0.o�7��-((��2���r�C����i�
�k���pu�A�$^�����cM�.��#i,���JX�*�P�¤�{����C��KG/w�U*S���?��8W<���F�7�*ׇqKp�}$�'�����Q���z��
'�c�qqzt�ZAR�GIC�6c���6��R �+f�s,���8��ir�`d>e"s=����(�=�=�0�'�O�U9e:�S� �H��>�A�.����f���F���i6I�9���n�&� 0��Y��=��2Ұ��o-�?yJ �S���Ԋ�|!��ï�X�h{7Ԗ0�������M埚�X����+,T"�ϚX�����<K[�娞��z�49(O*EYe�;�o��=�qqh���)
ު;�=e�X�t�����,��;49���q�>TC��S�	�?Z@�~�zK�涬x6�lR��{���)�GE��\�������� �e�fIa�|ťk	^�3�2��2�Z;GU��<�oū�����m��z��Ow�M �$AXt�D�����>[z���h��e�
@�{E�
�q��/�6Z�I�y+���W�~c"�o��[�t^�܊��pJxħC�O�(�2��"X�.XmR���1f>��U�P��n�*�9)�&X.E���|r"~�h�Sʣ�~�=�� ��Y�$��a-�7bFp%`f>l=]�:�'%�ԯ�.���P��<�>�\����	mY`-�����^`�,�.����[u4��{�s��k�말U��`5�सBfM�&�S���fMw֔o}z���AiF�Հ�b�*�o�ZCY����l&� �}�KejMsB|?��K�~A� ��0�dШ1Ѧb�*.$v�s�j�IOM����V޿�)5��ډ,{r��F���������B�5�G����.�|���	E�)�L~��t�����_���}\��^�%�!p��>g} ��@'�ᑸ���cOM�#����;E�0Mɞ���v����V*��4ܓE�E�bR�`�v>�,��������O���&�@�M�{M�ى��{5G��ř��}���X�3[�<,��s�{^&qMz�C�&���)'P��Q.,0���Sb�Ì�PJ0򡖒jH`�!�#6<j"wL��S}�Fb#��H�G���~�(w4~�A�q3F�2��zϫ�+�6��S�4�R�B,�`BA)"tݫ���^��	٨���c`$n��iNL��Mcj+m�D�W���	E8�f�J� ��?�5�e8��Y�P+���ȒG';\=����1VJ�+sE&�e�TrוH��:�����eB�/  S�&��'�g~�����et������$��OXL��&��%��R+��`�1���V�1��ļ�<9���
�i���4�$w	B��8y<�m�'�{����R1:�P<�;�ط�>��h������zGT��������d#ه��v'cg�9��
tA��V�)�#v��e���,�$���#7ټ�=�
R�u����Žq�bI���۪̂�6L��e�O�o<����7�����Π��y��n�T|�� XY�#��̂6�����T����
���(���-()�V��'����qK��K�(��9��$
�VA���Y��ڞ���������-K7�I=����A�������pY�Uy�w�<�M�䩮D���|d(�{9)���m��>��!�1"λ��f�_PF?��zX��1���" �d@V���2�s��w>cz������`��c.��G+�8Ή�N:~R�X�m���16}$�c��U�*�����3�d=@�:�����/1�%e5�P���τ��/T��SB3r@�&�!h�pl�{^��h���ZZ�?8v�B��0{�*i����� q\���@|�
�1�v�2i���"�%��yO��Wyx��V�pBSm�N)'2�'')ȿ�����%T�@h����#��Ix�+z�K�*��Ⱥ�k�������'�W$�n1k��W*�qPh����Iq�$�Px�(�!��;�\���Ě�f��s�V���I�]����,Q��@�4�/�Ğ&N��mt
v����z���E�a��5�O�0�-*/��� �ӊ-k�4�FI8\��(d�],z�
'y]�J@I�+h����Ldu�����U�@�_/Db��k�5f�dg�Ao��B�V+�	��=C8�"��
�����64|D��[T%!��b�0.|��Iq�q��J��t�'K��V�t����a?�)4r��}`̱M�2F3�p���@l@��Q+x�sb�RO���U&����)aCY_��Y�tjq<*`�
.~$+sʐ�W&Yp:�n"�	��lXx@�R�Y������!�w�B�����i{�!��j��_����5&���6|���+�4N�����꛲�w��ձ�N|\)��Bb�]:�ܮ������l��2};S��$���f̿���{*'����e�s�j�5Z�8���6ih���[�/V@BN/Ǎ'M
	��4 n�⦆QX�Ǒ����U��C�Y*`O���:��$=�z�vW���y���95�67hb��>[ej���?�����*"b�~|蒯��$Yѱ ރb�AoH߬�?Z��_������КP��΁�Ա�>r�Sh~��ж���%�Đ�z�yR�\��v�x��&3��e��})��n4,��:��E3\�'ee�f".�5�h�ڀ
~��U��C�Y B�6�j��y��l/Ya!}��z2��0�@���e/�(OW�z
g���<�#^�̈́9	s�������� y��@񌍞�?|.*�9�>��%�2)}�G�ɤ��
5�i�IĞ�d����a+�CL�s�]5���_�p���G�UjC�i*�����n-t$����S�����x��O>}�Z�!Q�:i���'��w�[��o�b'H+���_�Z-�,&��T�hxk���X�mT_�۴aO,��W��%�� $���d���h)Je:�����s�&��8T#�*��$T!C��t݌;�_x�~H�h,���P��,���Do?�\����*�y�&�c;���a�e�Z
u~��V	�����y
ߖ���#�}��1TѦ}՜�	�q;��=+T�N�Q��"ûS�p5�ziCi�P�?	�e�ȟ��]���D-�Vw)�e��{G��*�'�D�G����_��֔��p8�m��IbӴN�E�b�N�5�/�(0�4�G5]c�Y��H�����?�@-���@	+	�����$�#��qOd�v
�C�Ea6�H�۪;�&g`��@Kk�p�JJ%�S�9�E���s|��8O$�+��D ���2U8�ѯ�A~V�%àϠ��W�d��"�B�AXdfܦ���̓�}a�s�!W���'ea%���me�,��\n���#��bP.�"��#n$G�k�4��`�qZr	|L.����b�DFK�]�&X+ xSM��2<��b^�����L�
h��-���Ќ����7�u�&x�]��O��(���3Hby�<�1�ʪ����~R�bZs��VA�,�|�:�<�@�RB�r	��}'������ m��Q�l*��!_H�*�����`ò�ȱj�N�*$C�����ǿ4��ڧ�j����s��QcB[j���Σ�:�Ss<Gz��|���'�P���$S�an��V}�8lulw0ʵL0u���[[���2b�|�����U���I�J��]��,"����Vƾ���d�!�r^��
v6�3<��,�d���.x�������YT�W�Ê8�X�����K6��+PE��3T_���!��/�у|N�O���p�����/��%�t���c?F���JV�hiʷ���_]�Τ�bG ��3v��D�-����m�˹�K�y׳�6�M��r'��JH��9����Q����#S'Xx��[��7��5�.�w;9�g�	k��E�f��ReVe�̩,��a��,aUO�.�����W��;�z�'8��ׁP�����v����]��I�����h��t�GO�M��ڦL>��lv7[3�כ����ź��K��5hU5�<�:7�iVce�h�!���1�
��O|��	�A�{|���'O�&W0C���t�Z?��x%�D)���p�]# 1�ݿ����Y.*�<AKZ�vC�Ƀ����_�
8i�H�z؂��@CR���9��h5U��nM`rE��%�tc1V�O)��$@��fKZO�r�e۶��Q2�ň�_��h�l�ig�ߐ[3��t�J�I�1�Vumľ�x��8����B!���o{h����܃ܫ�����!��,o�-��C4��{?u�i%%����nҟ,��Z��rs،O��?o�<�LE8�A��#��|���8UϜR����joLj�/����� �d뵹�I�j�ҕ���YQd����%O�/��*�{����(�i�Zd�#nb{�o=R)0�M=�a����ٖJ�X���t�qm�5��3kE�1�d�� ���O5Ơ�Xr��CZ��M���J���t�b^�aЫ�W�����t�����5�bC�T>��B�
�ݍ��C�FY���W�*������y���W{<d�}��2��R0��3�@��*	��W���s�VG�t{��aD&�y�K��(�v��d���������^�� �6������!y����&��j���Q���O�Mr�z\����c�I"J\��Xmoh˓׍z�0��(EѰ�-���RGP�9�u�����+�_��4�n�(�(/�e6��!��$���Q�����iS��bSHH��#Z��q�w�0����/
�
�.��ʖf� �#.�W\����I�U�"Wh�ǻ������%=;��v�ݬ���|G�C��}����\�>�/{_V9���Ķ�����E|���1]{�M���I%T�Ŋ~/�m oH�XaT~��R�T��Lv��D9��ư���.:z��Rݬ�ם�d�L7�����T����J��6��kP�L�.��B�tG�Y��dC��>\�۝���ow�s,����.���ծ���r�LB����˅[�[��T��eQ���_�OP<�I��v�t���΀Z�����˛v�c�E�
+m�6�!�#�_���K[ ��T�����2J�?���㐆��30	u�)���$Acu<̗**�4��`MП�C��3M@M�$d˿��P�`7݅���d�dV6�bc�zS�}V��|̿�(C��0�:��n?'��"�w	�e-^I�}/ �fGS&\`��X��+�g�xz�4 ��2�GҷknR;#�:�>G���P�T�Lˬ���'})޺��O���;b�0C����|�Q*��E�Q�?���*���}��-�%x������7��lڹq���""z�E�hG���.�bUB�-Ы�.t��lyHH�I������x� ��ij�m(�#�'�������f�$RV�`Db�81�����&�����77���޸�퇳�[pƍbr��@ղ�PUx>��h�������/+fް�n�����c�so��:�g�W3�1ѐ�;����&єƺ��E���=sf����e][{�x m�����X��?E�H"�i�$��ت��)���^�wPYb��*4��3<߬x���;���2�䪆��M@4�ao$ ���	k|��1@��'��	l쒐�I��p]�r���p��{Ӑ�z��a�`}|U�G�,M��9�׻���aY�=hT(a�-#J$3"�y�t�p��?j��WplT��ZFŠ�l O������PxW����Q����)�(ߵX�m�6K�6�A�Ȇ ���<~�w4�B��{�D�'0`�
�P�e��9"t���*"�~ݨ#r@m��Q��pf�e�8��N�Crs[��v�1ώ�FP��|�K�vY'�^Kl�w�J��0Y�i��`�����[b��Ea��7�q�5*��F�d�+ԕ�E�ڔג�8���&_ii煠�לٮy�.��L�֝1�4��'���' �c6}�$é|�$G>\�d��#U���)��L�ƌ��=���C�6md���u��u��ur�8U�+��hww��j:i����+*���?�>��(��5�YO��Y� ʭ	�ъ�'�s?���&[Ї��GàWJ�n�oc�@����U��3��Ĉ�(&�ܒ��}ߙ��D� &�|�����5��rOj�.X�����,��������$��B%��W��}�Bqk��%��l��c���nܫ�B�B���:/��y���
��8�����ݥ��M�4����P\l���Y�Y�X���s���.�]��Vg�e����=a|�e
fk1�U�ʽ<߹H�\+� �2ql�(�W�Ui�jz�;�Ԡ :�oㆍ�8�i
ȑ	��ϻS�x%N��&j�������'�H�f��͠eFL��|�\R��Ux�_Ntz��/��n7���C�P�q	M����ɮnfV���Vb	�?/ڎp�fRR��I��"2y�.*�?�D_j�`�s���r�o�[؝Y�߫3�
�/d�>���t�Ϸ:�٠�S))%��O�}�`-�/�i�q	��Y�'��BJ(0��ta,t�����(�`A>\�%U����fW�k�mL*�^��z8.��6��0��_���7Q�M�1Hi�
`n�M�c���c�G?�Glr��������}�E�s�5�{>^�s�T�x53�ޡ�_��5�:��%N�A��/\��D=��#�n���C�lXVX���w��g�ײ={�@����l
��S�ՠ��o0�)�s;>ܻ$�vN'�;c��R�U.��q+�=A޶^���C$(�i����(Dm�:�'�'X��?H��0���S�� D�K����&��=��P1ǲ@e�\�{
�q���4�ʨ����g}VV�;�AV��+(������~уn4�r����S��BZ���,��/��RCh��,������c�z�:>CW��D�uZB�v�Ju5I���^a>C[X��X��7��ZBu�����#���iYZT�2'�ّ�)d%3'�-�gTJ�5��3"G��!��zsM���{h��}Y�]b�Oz�q��Y��u
���ѳ�b-�V�j�V�y������9�}�E�����>�&��a�8ZKn*�C;0�#����O�լ���OɪanX����ܳ�#0,��?�V���
V�P/�BP��b��f�Q�:��bi�j�7���y���Ⱥ�ū�X(��b����w�Z;n��m<��L�����̚�~�ju�yܛ-�I���_���!bBКN������0��Q�����6 ⼓T���	s+.��Tj��1��#� �d�c�1���U��qZl���,����d������~eO`i(��Z�5�_���w�,߬����QemxL��;���v�D�v,I��g��Z�0[����e��D1�q[��3�%���6LUk-c�x����<򉱼"}��
�p*\�>�I��l_�u9��Q��M��X�8!�mm����m�]����x��ܴW�f��c��BKQ
:G"�q�@	�j�--�����*o��̝���'�jt0�̺>(��ِ�z�z�!�!���\���C�OxX��/�}�P�ot¥E�͔gO��1{�y����e-ewc�G��v-���Z=�R��݊�r̬�?�$��ea�H�_|����3A7����W	K��f�0,tWe3�tQO"���n�<��~@�Z'S��͕�Y�^3�P^�~���Z��߿3;�qu��hh���l�s����/G��f�_=��u�������
��bM��F>�����vCio��>�N�mÈa0t7��t����Y(ˎC&�q/�g���ٖGb�Z@�Z�95!Y��&Z*椉ē��_�+��h���y�xg��8���d�vn�����(����	yc�ǒ Yx�b�>'��=D���b�j"�l8O��[4J�wI����j�>�;��>�X��Lc�:��_��A����j�0c����{���z��*�3����{nK8��e��z�HE�&��d<�Q�5U3�pR�tlӝM̈́��7��4
r��7#%ds^�]Q&���r�`a%�j�h s�r�3�3g1q��u{��^nX�nb��:���b|�SH�?�M>4���~�����~��ΙM&���E�H֙�Ҟ���B���."GjP��1�,���طC�l�����c���E����LF:~�ai	[7ݸ�w��x�}�vuj��m7i�l�0V��/�ok�Q&������?�5�2[�����➍��I���
�9�Z��X+���%�D���	� ����ԏ����i7�"�?P��b61��
L��m��6	��Z��CR�AUCcI U��g8�i=֠V�Y��0���6�<ť<�v���%~$Ѝ=�ѝq��3}�_�2v���w��Ã�Y�y�&[�{���P�<�Z"#��D��^���ʬz)�T�����7��XM-�4���AI�	Z(v�y�*!$,#j�V9�3G��%k��c�⯳H%Cqe�����tZ��S(���D��]��sKTSXM�-l�c���|�f+D���{$	�.� �O��v|�0Ү� 棯�p����`���l0�r����`�<;zȅ��xd����`�J^(wףּ�@�3��YaNK?z;�{����%��&Hcu;��@���}�`� \ ���w..�Z�3Z�Ϡ�)��T&sލ 哨p�?Af�:��%'�`gPy��Z�Zk6��X�Ƥ>ϕ0��;Lo{B�I�T9�/��3AK|�u�..�9�@�Pt
���G�=&5���c� ��e~�����C�	~��� ��q��@��c�ǥ��J��L�\5���}�V�x(A�3WĤN�M�"��N��&=�S�M?�<�6Hs��Nኝ��h��$��Y�(�Lx���HP1���~���k V�Q� B2����;��lۯ8��%9�ޮȀ}t�+d�"14լ	p������	0U�@��ay���C8v%�|�i�D��4��䵛L~�p�0�x��`8g�)X��9�S9`x \���*̟8Z������1H�::��xGst�T�%nH���2r�P.ߟ�!2��
J�8e]ĕ\�z=tP7E{�|�A�����[�t�k7dՈ"��T���r"X3H~�����n��#}�ԕP������zUa��XՅ�c�2P�Խ�Ŋ'���/�o%x�_�uR7�����	��!��yǃ-T��)JGk�����lj��]��.�<H:
�J	���K2�%����?cT�&�."�^W����s�b�Z2�̼�lv4����ӈE~���ِ�`�K!�#j������S>Ьl�1����:��D�t�"���n*�=\�8^�)����KNLMU[��-���b2oq�^\�'���<���l�<y��G CW
��`س�O�2�)�T�(��n�St�eeri�/s��Y�K]IuRHK�����ʡ�;]�����j��oY�5?�u0���si�C��U`l��Nn���ޅ�q�H�w��E��@)*�.���� ˽�4j,�����������T���6�)��:��]��3��1��"o���~<&�K�$K���� ��j�K$L�ԙT�ݨ�5_�NT,:��X����m�G0�vn�XIf��D�3q�Ri�^���*����5L@H&���F.%�_�i����9șn��� .�T�}�1j��G����$)�V�F5<1��
�DK!K�O>��Ih(� �[�Ck-G�O<�'�k��49��x��e@�.ǩ*��%Ѫn��Kqf�tS��vқq����m��bYb��6l�B��8����mI�>)��A�7�Y����E.�hu��M�E<���6-qnq�8썛������\�:�L���c��:�N�1F	ïK�i�|r�(Mj�� XQ��W���6p45��)~��B?<�Aë2�XlHݢ�;2�zD6�@NQ�cм�O��av@���i���-0/����^))�π��?�2";]�=��{��8{YR{�3�m]�d�x@��].���3����-�h�V�H ]�8Uv'����[�dCks�x]%M�/Y�Դq�tT�!.:)�#Ҫ���[�+������D\�m=l�j�η���;ꜿ�yT��T�K�2���E��.Ex�EHAQ�H�ˡS��S��p�Z�_�#ɥj��pHe�(h@*�*I��3--
��r����x��oY�<j�S_�0dztu�C0�p�G7�*���G�"�iSB_�ۢ��F}[��O��e��3��ۈ�K;2XzB�r��i��I+�v���p5���6P��H���au���D��*���[S�+�g�{n5ej��ͫ����a{��)�w�?���`s���y�lh"l��|忁ġ�6�Y-�p�VG��¾lL�`؂�A� �oV�
+b���:D��cs�b,�D�Ly����#`V��� {:����*Y���F)�$j:�v����4i�6?x���i[P��v&��ܺSA��Ӽ0��!{�L{x,�N��dQcTO���Wl���I;��Z'żP�>�`nGrT�&��,V1 J��y�
��m�ok1�҂o=�g3�H��j!�e���~_l��t��S/��\r�e��A1�D�Ng#"KeT.�<OQ�.d@��t�]*z�R��RR,@'8��Y`=����ٚ8%߇m~��*I���n0q��R�A1�}�
 9��-2��N�2����Pt��L0a�1`@�M�3�.�k������OL�~����77�Ơ@@�=�1�����z������x�c�Zv#����zP:�Ҡ��7\�����)�ŭ`.�F��;����L	�8���(A)g�IN{��~�)~-���� �c�,�dQh�[��X:2����z��ص-�#�59SF���JN�?���&�2�������[��r�w>���c?�*zl�	Џ���tGPv%��R��|�):&x�k)�S1��Ocwv/����6��O&���e.r�F�;�j��{��3S�o#�F��,�+�ת(���saq�ڱ�K��X��CY#�W�C�,7�ЦZ�iT#���F	�y�@�ѱP�ȑ�.3dE�w�u8���;U'�}k��%��xJmIN�6�4�OSX��
�Û�� ]{@>���JkI��8�*/�^���q�Nhn�F�yR� yPK4(�nj���3�������S����F�]c ����j����-�}�^���?�.�����"s[���i�(�f�Fkӭ��M�6�a�,Gy%u
�U�LOH#gϿ·bT7R�؊�c�E�,�@���_2SI��R�x.��,�]	����7�N���2�;�J=<���(��h�����;��,�� `�%�� ,[].��re�1�&?�:Â2#���㳻�N��*OV��<J����^�ߔ�QOi��ӳά��t��m�xu+AV�B<����qO��FL��$�H�>��u�Q��_�.I�*���8(��Y��Pކf%/b^z�#H�[�|)� �	��������I��ai�z���e��=L,��w���~n
i)IH��z+�E�rg[�R����뉜��y�K�)����A'j�Poq��⯷-"�LH�S=�^d����%D��D����#]�75�A���svdP��=�$h(E�����|),h��x���݂<7�G�9���YG`|kU���yw����m��c�d�L�H��a	V拮��L����~��u��cDyz�'X�0V�b*xK��n�U�y��ʑ;�/�B�#�h�%�J�[zc��r梄��{@��t&-��ت����xǘ:�q�N$S�x����v-y���E�J�%J����݄�=͍���m�zK��]Y�i�Eo�a˲��Y�t�E3��0��D�ˑx�K�'�4=J+��	d=���#�	Be^�`�1��{S�h�ږƗa;B���aI����	�Fs�����j�~+4�2=�j��\�'��8H����>-�=�N$�¹��7&*��W��^��dZy�+zk��=z���(&y��\���͠v7�!�F���-*5�����������S�t��m��Ǎ�TP�J�㙄'�vb�=��P�(��zaB�KԾt��m���&]WD4g��eE�i�A/�B��Ms�T[>���������Q�)x��v��61�LCl�4��!�O	\��a�����a�C��f��Qy)�-�K,��3�r�2n#���$���7�.�r���\'?���Ыa$'H�'����7��ϝ98�"�|)K��;� ����z	�h��!��7`	/QV_֕���
h$�ț]�6'�+Qk���h`8���_��-'ʝ�c��u��竽	���CI�����TwF"p:����n"���$�}�6{�㢕e�,g�Q��\��<^�ø`�����nosu���<�]��� 8�}\��M���|-%k�m��/:w��<^6�|�	�fX��x�ޟK*2m�O]�h,	C)�x�R+������Ȉ�w�a8
ɩ�t ��!��"��FtC�wC���)�Ӱ^0�V��5x���]ͅ�v��N���-�ܨC�-1����ȶ���9��6g`,�YT��=�r��ͻ�hݠ��]}�L�6F�O��RRi���7�&kp�����)�."�0ZAЛ��Prγ���/�B�K�n�3vMD9�|�e��z5����~$�B��^!�xϊNB�[Tj7�)����׏YV;Q;�_6�����T�O��M�0�
2~� e��8�@�ςH	�k�>�Z���r�ƭ����Sݖ��,�p��v��4�CrjFpS!�c�?���Lk��_ �q>�XFI�"C�ǿ�]>G#�Ù������:G
��*��=s�3>���ל�X.[�����_��H-iE�*#V��n�U�66+f_�a[m].����c�O�I.�ʨ(�~i��/��![�$�0N�~#��w־1$�v����Xʆt�h�H�r۱�E�0�^�ؑ)�9.Pà��P�,I#"Lop\/j��R] �`D�T87��H�*�Tw�6��D3�0�1LlZ�@�'����[ikT��ҠB��w�U�`��,��e)��A쀥�N���8�^�A�cV�n�,:"︇��q�� ��cˌ���vcZ�'r�50x�~�P�������\����Lٕ<��?�xTH8#�52�Y�� �߭0�@i�2���~cn�+��T0���~5��b=��. ĕ���U�z�?�kAL4=wz��T�̷���BEK��f���*�Nd��*��3�ˡ�Dob&������F+`�w�Q��=簚������b|��1j������2ޓc�Q�\�fy��N�Z�&���P�}�"��� *����b"�)d�w�{�(��v���ֱ�Ŭ蕙DØ�D)��@K���sYlk�XVx�g��xJzM����醤������h�-� �2�����؜��@A�ƕB�;t\�fS۾�kI�:?�с��Y�z/)̃GZ��^!���"��	�iw������s����L��|�'q ��2�d�k-�X�k�l[�:��;yG�'쪗�K�*��Gj!G~�6�Nm���N>q�QaO%)S�c[�By8��t�T��4 �4�EZ�e�$��6Kқ���C�g��GCC��6(Θe�����F��23,�����#%�`~8�y�Eo��i�c���?�G�&6�"���4�C��c�"��_��#�t.2:���fR~�  ����B���w���I�ZF#H������J�b۔s���}�U��[VS��MX둎nő�pj8�G�L����Q�$�$TSZ�ccd��c>Y���ݓ~R]��s�5=n��?�5��%�S�uB����e�Z�6֝�mkm8�4�J�f��I88�qS���j_�Ϛ"RR�Y�p���jrl�.�\ 7|iO�ʅ��_.B9�_���j��ȍ�"뀈��(v���;.*��"����Ba�GB��`HJ��?����%��ڹQ���GEntU�����h�	��;i��:9��J��2��Xoxzz<�[}w7i���koSh�#ƾ�*Dj ł��x�<U`,���i`Ӷ��Ġ:
^`IՅd��n@&��+�m�����#���uڞ���t���ź��|��(p��j����By!���Ms
�&S���т��2�����
*#8�y��%gK%E� �Íif���tX�QQ9������W� J��G���>Ȱ'����͐ճr�!35�Q���+�a�]�c�y�ƙ�q>�`�2���ʉ�Ue���NZ:�Cm�)h����6R�E
?�g5*;*����
��4�e�p��=�H��c����3�5�����W�
c3��c�FQ�9�!\�g����Xgg�W:ժP�<$!�M��#q.Д�ґ
\3�\�t?Θ�L��%f�Y���u��ⴧu��ޘb1_�7$yΦN|���yo>̗��t�)1��f@�W�ή@]��?>���e��{V(p���6)4��)8�n����B(of<�U���s���FR�7[ԢC�u���E�M��pʟ����
7ņj�H5C[ �j�H&T�ɒ�)E&D0N\��V�����=u�v0^P@�	���\g�'T�stU�uR��I=.����+���Ñ?�v]����n�
)�=F���]�[g}��P"���t9uAa����9�W����������)8�=�-�� �-��ޒ���q��G&�����(�lC7�kU�K�Ә��YD᫠[o4���+�9��"�6'1��;�� O~�`X��r_��9~,c�Pa��?�\��h�#p��U��x�Q�_�>��Tx�-����Q�3_]D�`�J�U���t�%� J�B��)�_��e7/6�7�g����W�1�V�?��ĉ���+Wܵ�"���q>\t���{� y���$���d��R�3o�l&�bĳ�`�F����8���Q҂#��6Ʃi�٢�r	.5���߾����\����I
g���~�0�3iG����K�=� �U ��B{�N��H�W���ix^��G���@�=��m����Wn�}����c:�OR��2��y%������Ũ���e.���)�R\V4r�Y�%��zEuR!��'��q��ça��:���H'I#5��$��׽_�i�p�|{K�X�`t�hlI�C5uA��W��iH<v�*��4����j�P��%v`h���8����Q[�����c�@���X�Me�5���c]������6�7���H�����8oM-}���cG�" *M�O��r}�!�x��ޮz����5u��̤<ꄲXj�M��	��`:��/;���=HK�Y(�?5��/�;�$��`a`������']�Z������1���7���?��^���I�:�=��qQ��!�ɮ���6���i=���o�ǳ��Z$�{�F�C�q[�������I��<�e�7���Q�楳~U\k!�!ٲ�-�.���m�5��H�}�PC�P.�2�hxo�����a���(n�G%���#�v��-1Q��b���'�$�*J{�t���%�U[���滔ż�/��-�V_m:4PZ�q*�^Y3f��_����>���ȪPvNv#p���E��Jw�4�����S���'py�,D�ج�^ �,�Eܾ�Z���i5��Ę;�h�ʦw	���S�:Z�)3�r�UbMu�K��mˌE�������;9�x^h�����ap�0���;�l��cVg�r�'���pt�?ޟ���,q�硋�J"���������C�9%�y������$�8J�Ay��D���,S��&�����l�� %�'Z��1;~K!��T��K];�峣�NI�Tf�%�E��҈�٤,��9Фk���b5_���֧�.Fq�g��W]��xbw����&j��+ls|!�W@h��߻Իd���������uU>�������<�]�>�#���-��p�)p�.$�|�=q���P��I�����JZ�q���C�����>}]k���;.�%��|�_\�.�]OGx�>�V�N�;����%g� ��wV����F� �P"�.�6�ㅀ+H7a��%��?<؂b-��C�p�������=������7>Ha��2�a
�f�GE�ǣ��'�F��_���|E����M2����Lӝ-�-a����ѯ�-|�<��D
Q�k�ҡ�J���hdYj���݂�mV���!Z�^�cb[אּU�iw��q��#�i��h��4}B�����!�����T�!�f.�6p,���j����J������c&�r��2��ٻ��}`(s��h���D�>-�ɬg�F4�gS�s*fQ��ꇽ�0������l��L�7յ94�]�NYj#��=~���%)I� P�g��pRt/9m��$]��S?�п;.�1��&��<r#y)a���萗�0���o��c|���1�JT�П����ӫ���ߊk���<g�P�� �e�n�b�7o�}�YP�Ώ�p�"jֹ�4���$ix�s�Gx_$��f��ʐ�?!��czNd��b�j`h�΢3�\���V�SCu�ƼG��EB��휄�s�9qE|��C�I�l��NqIleOY�(���\�T'�Չ��Cӏ�߉���Tž�K��ZA���۔0���7�|>x�yH�;!�\�|���&���C���L-� ��.2(im��y81�{+��:D�i���$����Sj*#���x�am���uf�?�7�*޴S��(��4��g���զ�2�	�*�Z����w<���>C9yk�J��!�OG��m�,�>4F���p�+lB�y�yL�Ni�<%�fb޼�!B,={<x<�Y�1��9�/�VE��L@�H�T�O�����Bf�@��mS�o(^�2�V���r��>>@�yfG��;m��)KXek|c�[b�Ƈg�|��/�'��/�������/ѝ��hKS�M@���'P��
e���~�ΎA� 4��*;���K�����j���'�0|��O�8�_,.�!��i�+����EP�&t��]����3�_�V��8�ʏզ�0���]�VH�rV�p���:5l+A�#m�׾C 5x6�_�#E��J����c����.��8 ������ǥ��J����qA6pkp��֙+|\K�Oó�Q�r7��'p�ݴ������F�k"���ϕV[S�A�j$��
$U���6Ua[ʜ�01m�KCBOhz*'��V��rl��TӾ�)]��-c�h]��2��xth�^�e=�����m+l�������a�$8:*��rtЁ��+v|��1sO+Yכ�A~w�|R�&�����1X�q��"��4/��k�{��"�W�V���ǫ��Z�}���0�I.��W�[D"�w�w�� �m:����	����E�9�7�k9��>X�{���D!h6�����NW�s�s���ξ�@)�QI��g�Iԓ-�~�+�l����6h�7V��Z�·�
�㢀��8Y�lT(t���}�P�g u˰�lN^�F�ɛ�Dō�LE�Ӭ'�H�1.� �u3��3@2p|�w�P�-ݛ�(t�����4�$U8I)S�r?���>ƍ��qF*�m�ށE�M*{3�3(����'#��lɽ�F��d@+�Kq\Ec	d%�������|�2Λ�]��+�ﹿ��n�����l���%�x�7�O�p�a>�h��#�<[���CJ���<`F��2h����	�D�O:����
t���R���5l�W��+�E��x.�n�Oү�zl���6�uzn=%���w�9G��P~��`c����fA�vP|����}a6�H@9$��u)F���Q��X�c���qT���g�߄el���D{� �=���6n�򄑦�ѳ����W~v��x0��B�%h ��XQ�O��C�-�zX���/4�Q���*t��v6R,�m���p���!u"PQ&���*�( D�J��:��cҺĒ�_�'��]���y2��OV��R���M6�
t�Pf��4	�st�����9{Mʈ���^6Ħ��!�ɴY#����U6�)���?�z��Y~��rIѝ��&W�(^��\bzZ��o��!�e.`g6j+C�}O��0%�GY�$Sښ�J���?��E�qu ��a���~�}5
��*�&o��y/q}�P�ANPK̩Ƹ��ôA���?������������`��Z����|�ȩa�J`XN���иis��K�(���P$�)�iU
��P�U5��&��j��:�en4&����O�%O������%m�=ͥ����p�A=\NL��j,:��f'��?�4Ǡ�qћ@�X3��Nj0T��3�p���P}
��r���ڒ���R%HW<9��P��M�pT��xB��E�!>'s�@Oh���Fg��8��V��~�cQ�O���¸إw$(hW��\'�z�:c�,�E��ɡ���m�0���y���R|��+-x�?%��1�5{hOIfx��?��ә���Bk��!���Z���X,�~��O:���!5]��&fH�w���=�9���n��hbK+!!���~\~��&W[f碤��\_�!%8��y��<%�@܈��a6����K�8M$[9���� ���e#�c��#�Ԁ������JZt�T��;���`��\޲�>��T��,J{X�p�
����B���.�3RP�W�A�ܨf	�(o^X�BS���Ѕ�4�^�RIw[c�FlOH>��&�2ɚ�{��e��;ٳ��(�����|�?䪖�똑�[���S[���d���|(fĈL1GX"�%>����j��q6���4H!��G���8δ�9���@��4ׂy�Fɩ�Θ+��?�}u��+���*\H�(Vg��Y�sa�~�����#wuk�Z#�G�Y#~h>���;�.��� �@��f�e���r���[�l���m�ă����}�Ӂ��iR��p}��Ղ��o&A���'fT��?ek���n��B�������t=�C����â'Һi����v�[vk�D��U������R���3�5��D�VO�,Q⭘��Gq�]��}~��dJ�Uƚ��f��EK��,��Y_E08���>����9�>�޵< �~��!��F��r�as��7�R���j��W���{�k����g��J�ƣs�Z�YD#׋��-o��X\3���gUx7�-4��N���l�,5Ҙ�u�G������Omb)����$�;7S�w����m��T���1�������;V��b�yH�6L1�ʝ�)����O���Jp�|YѼ��_�u��&A�����f;�&#�#������3a��ʥԶ&,,$��/���殕���X�V�f�b	��6`�1�j�S�Ogҏ�  �:j������_�%_�9�[�w6lҁ����̒����>_+�E�J�0���/JF�H�� �#�ri�1�#��+�~1 �9���li#�Kv�c�>Dtq7��_\�c��&�XZ�G�/\Js��gޙ]0Y�1��<���Bt�&�,>W��~��|������M��b�{�*9����a^���B�gӀ��W�~�`}��EP�u�뉊���褵���u��G�[{�������jS�Z�aVz�N�2�������ÿ���%5��$c�&��'E��?�*�X'�$j	�ӑ��Am��8P��{4:%bҾ���_�t�.a$K���s�#��}�s�s�,��J�Y7���u�_J�/������p��X9��edڳ����|��9��ɢݬ�YbH�#�"�ZB^����ki���	� {�p�����-��Ę���x�n�;��jG]����s��M��ͮ_|(e�R�SU'�~w��&�HJj&���PV�l>�v�Q�[Q�-��Or*��nk�(�sM�}Z��v�UIe{��D�`�B�t�L�3iydٗ�(��m5�8���W�ߑ��[/a�����_��;QI�8�L���)�
]�˚��]�A�U����{�ݺ��~PmH�����U1y��v��a���+�733�e��d��E��J����'��Y�E�o��K��;R��fUe(�$׳Ɏ�BǪ��h��߿��r�����Sǆ3~�������B"���Q�*�³bzG�o M�D���d�J(��◮:�Ǫ�#�Fki�Jx��e�����4
nxw�Q�-R��m�Q����d`F@��t\ՠ�i�.R��K���=j��ܞ����l�mJ�k[��Tܘi�\�M�֍�t�қL����8ȹu�Lq���n�H#0��ΩT�h��{�*��X����G�?`tve�$�0�E�2!���ב����T���b�,$k�ë����k���&N�eKOZ:(i&���,�o�[^�����H~R�Y�΅���8�������]e��A���oHB�_\6�KwV��]�}���R�i�7|�=�� �4��)
~:�]�3`V��O���ʵaG�F_0�b���N���Z�7�R�.��\�w��}�?�2$6��&�ɵ�jf�4{0Ej0�s�0  ˞���{uF��.�nqq^��K�����5��:k��lq�KWyp$t[nH��iC;Mv��&�+S��6���W���"%u3�3O��e����hZ��$�O�[�r��R>���G�:� �ͯ�bt��0!P���Њ������<`�M�8?;A�t�*B���5�#8�A�L��a��P樮�+<|�0�8���(��8%�N>@��m!���eqQK�Ha� ���b�D����"�l?G�����x��=��E��y;��Y�=G�$N��l����� �7}*��rHm��=T
�X֥��v#��**?�1�i�XcSm2�h�Z�E;�4���w���<��Ɩ�5�/I@mN|���a �Y����Bb��G!�7�0��EN�T������ڍ�%��ٜ$�X�J_�2��1 �Z٘�K���Z�[���ٕ&#��a�X*�������h�^�mK�K��}i[uO�C&l:U>��v�ӧu�����GIr�'CD�1���*�D�.R�!��h�T0��%k�� T�� ���y6�YLz$_#�@I9mE��T�fhh�߲��.mهw�UF�|C������  ���F����P ���n|:p[��Q9�a�z���$!i	4��s�!������#Ŭ��������S��,3�8n�ϼ�BŴ�|y����⋡��=hѶw���0KU�YV~Y��*ϥ��)>�>�H�u���t���@��vfk��^�_@�ek����{��sĲʷ��i��Q�T*Z
�z���J���eg�A޿b�����՜'�n�MG�j��l���dꑳ����(����E��3Z��U�����g�M��B�dll%�<�?���ؑ`�^��/j�g�,�G���'!�-�nT��@�ѭ�2�4��op\�����f˳W�M���r�d{��Xc��5h��ҫ�&`�\�N�C���J���t׳Ԣf��a�g�����j�?�����S|ci�Z��ғ�K��H��~���g���Kh7�+;J(����2��������b�d��;۔w�[�T���_���֣_ǒ����>��-�]C����o�vt�f�c���e��LS���w
����Į��>�u/��*9,��������� M��{��z�0���+���rYBiꭻ��Ϭ���[9>�����Ȝ�!�mI���8�w=�Ɇ���b�K^��y����	�%��t^��!�?�pcuʅ�F�d ������RM>�~��>®�[���?�R�����Z�T%w�Ïè�gK� |3����CI�)��h�2fHT�,gN�K9�Hg���s���8��GG�����V��u�h�*()�$�wB���Ի�6�XF^�Y�Q���#�q�E�7��N�~��؇��D��)"s{-
1�zdv,*��^ۤ%�!����ܿ��T��ꄸ�i����TP�E?�zs��[(����M/膝�kQ��VU�����Ӽa�>��j�v8�����]'��ߘ"b��B����u��[���ib�K6�JH{�,�Aur�9��EۛY��M)#��ұ�JQ�aM|�i��Vx�׭�z�a��}�h��N�+X#�Tr��Ȱ�ПCa\x��zZ��}0��N�������H+x�0HuHv#�e7^Sr�h�<�y�tP�M��sgo����������#B�<����F�9����蔜�s��+��v��}U��(2��6�:t��P�0�X�s9���腇��)���]S,����# >�Gm�{yB�qJ$:N���W��4��-�G�������9yO	e=��WL]�3{H��ыA��Q]�(d�Vok��Л�xG��7F��w5%�Ce7|�X! �S�G�_p��JQ<���?���}ߗ���sv�����B0���P�om䍞x�eA�6�a�D�!����R�	2ba� �{6�;�&蒒3�R����%Y��޻{_b�n��9z�/�J��1H}�"�=z[��͓���A�����K�_j������$��c���H�D��ƕcv���]�����zz��@C�T�C�ֶ��Q|�|k%��W�W����%8��`Ų�/���>�R�e'b�M�:yAEm��`���T�t��>
�*�I��i�]������ �4O����T�b`l�MM�m4����{�� F������6uϔ(�[������E��A��n�IA�q���4|�"��ԜRV�sEӶ�DxM���:��)p��-�xyb���`9q�-v�m��,��0���'�Z����Z<\�C�a?�^փ�8=a����1���� ���&i]��o�&�ޱ���̥� *,oDj�L��ŉN��
~��C��yp$}3U�⢌Ee\����g������Xy
�A��]kD��>��?���83'm,է�J�+�Q�x�En�G���o5+;�s�&��6���d�yu�g�H��D4Z���dU�3�x��;��j@��j����^(h��g��-NSD^h�'��m�F�2��]��9<�>((�!c:�m�6OO��d��bz��#��/��+�QO�p�3�j�{���|�"��B����4�*f�`�'(0B�̒�h�D���`�>��LW#ɹ|�c,>��g�YUK5g�T�������I�/8�H���ܯ��)��朗sNX��&��1�y�Y�l@���a�ĝ?-6@�6Y%��U$:�ȍ�����h	��z�Oh�
�#��9lo�5�������^8 �n��0p�i/����(N/H���l��y��-�Ϥ�E�H9�W�3X�2`�yZ�V�R|�k3gy�҃{{.���2�:��@���k`�Ra&���qػ�a��� r�V7Ue|>��
����/��iC:s._�ϰ<�� ϡd�:q-c>ٶϵ�Rve38�_:�~���j�bh���G��5�S@��b+�po�����A�hCv��!Q��$0�U4��|̝����҄6$��V_r��3{T �V����q5Wϙ�A�x:�7z;e\���	
T���9�.qVB��G�<���� �%K�C�#6<bm>���Zw�*�~�@�'����څss���@ހ���z�S��s�yӮ��7ʣ]��&������,<��WWC��;+&��/�֡��h�N��
��BW0�QH��ɵē3T5|���}W�6u�����L�*��J��=�;ȼ{�	h@�VN�6m�/��칠j�8��g�r�{�h�̷-�)ߺ��[��nJ�*������S�!�?�h(�\#�Кq���-�N�����8����NXTQ�5մ�Y8n�񛾇�Y[��&:c��6�NQg0�z�^E���|�r_8x���q'�w)�A���L%`t��\�Ro�\^�*���/�SA�k����ܼ�%���f�c��tx�F�۔\>G�X���q)�f�����c�����jdZ��;��F�ɘZ��/0f��t��!�2�5%��jG|aT��e|�mU��dĝ�ma�F������ٺ[��*Meg�E�.�<2�q��/�&��j�U��w����S�o�J��<�
DܸL��G���z|�,�S.�ؑb8:V����k��ޘ��T�*;.�"E�kw��%��T�Y��ґ���z�l�u���yͫ1�2'�e��sCyK�����G�: F)K�E�o��v�M{
�HT�|�,2��<0t*�6�V��B�8Y��߆%�3n��%k��~�{n7�麟H���.��M��c:��"�S�G�N.F��&����D"�;�~�9��K@�Bk����_�\c�[����Xm{�fX�_�b|���.ͦ0%�d�uCW���8Ԟ��tomU��T��;���>:!L^����~\�	Uf��	���J��^���I\px�E]�#%��ӫ����{-pM�� e��Hnp��LT��J6���MB��А;,���ƠCsfs�b�/[�=A��׊K��x�{8{���]�ȶ����{W��nQ�̮�-��"��'c3���Qi�2�[�&�P-6ds�Q�`���.zr��z���XO���?�X"�rti����N��ʺ�	 }�Eh��tN !>���,`*�#�N�z��*b`q�P��ǆc��!K��Y��'':@9Gߍ�h���8p.��&��$�������!<��
�-�v_��h~F0\���<��dT��U�~
��Ӂ e�[^�/��'~�5�<��{�k��f�����RJ^e �`
ۙ�ӷ�N��PDFc�8����lu��MŜZ��������(�� *eY ���*�Kllw(c�E\���ˣ�;B"�ʆ����~ɋ3�c�����e�ĦvA"n��u��7�����iq��h��D�b�*�]����I��ȉu��5�O�>����I4�6��l�}��}����6�Uh�JH�<B^�!��E�G�:k/趐-8`�;�Y��?���k����Eb'�rץ 'w�Q���R��s:�9�)\K�%k��ɨoڝf�.��~1��G1E0C8	��4�R4��>�4c�P�>���Z"G��x�I�|NY��|狢�(r�c%]*� V�JS�տ�8��E���b�
D~o%:�7��Rꅓh{����=s6��q	X�2�A�\u5� =�pB�)��+���P�E�)c��\vw4�N�^ګ�I�pܐ)��Ȳ�U&<Yeêxs�3{QC�؍z�N$�H�}@�h��[^�&\�x��W���Ĕ� ��|���?���Ƃ�^+�ꔸ��SY�!t(eV�m,����?�3Q2��CC׎С��% L����p#VW�Qno4h1r7��@���2Vk��s�4)��{3���غM��h�ԧ�r���;K�\\�`�(�f2��+��~�ؐ�=vaJd��J�D��1�&"�������^�s"��<��q����Gk��>ow�7����=KX5us;5�t�-���W��)��G6� ���+վ2����l%����JQƺ<M�M�w$�K�+�x�~7������V����n�� JUl��{ٽr2�7cf/|�}�n��\VU��ӹ�T���+j����h�I��ry	�8�HPGF� ��M�����;`b�$�p�R���'��Je�Xu��s�ؼ��K�0�rj��M�g��]��*�Zx���	ʙ*zU�e^����}��*'�h�q>=f�-�A��� �Ϧ4�]�a��������4��n�4at�R�)zܤ�n�3n�m�#�ځ�"U���A���O���k�:������	tJN����w��P6b%�)=F�/ħ%z��M�q鼝@d�v&�^���O����?r�["��ïY.ț�� V�`�U^�;z�i�	!�\�H�.J��w��c���-���ҭ������+ק�^�<4p�>^���w �+F��3��/1�VT͕$o���ܸ��\��`v�`9~�sگy��i����-�wQ�;"Aj��ڇ!���������<���M�C�������nkj�xEx��ís��%ꫧ[`{�����د���5vil"������-�Up�]m>n�K:��_b�( 1��˻���~�*���XkE(��0Ҿ�����2<�+w��8#���j��M�)V�7$��<7B�X�Ȇ�1�ᩘ��/	�-Om\ז$�LH�=`�d���4%��$�L��ӐT�3/�eӦ��DA#���'`�ݘ|p�n��tI6����\N�_�d�+Ʀd�mH�fi�i�"��;*�֐nE/glR$v���P7�;��������zLtJɎ���eáƨH("�2"3o{��%Ӿ����lA0��"�8)�;��)w��{PP5U��e��եE㥺�WY������ϝ��{]��U��vra�J����W��k���9@q׺�g8�/�;�*Ķ�#=C��B��nɒ/�����h���U���~K�\��[�t_��念Bq{�ɲ�L?�����9V7�^R�}�H�`���]1����G�<������`�ʾ��&�M��ocv?$Z�H=�v��I�m��4	���p!���F�	o�I7%&!�Az].�@��l�!����s�\d�5��7i����t����� �s�Yꔠ
�p���4̟OV��i�x_fǞB�����T�����*x�}���s\	�iC���j�c�H�
�s�І(�;�r���!�����%��-3 f@��e�<�'��S��7�����w{�`�*m���Bq�^�Ŝ�Fo���t����
��#ќU3�D�<m�ʣd T���tR![�/���c��y��ݨ�ȴ��g<�2��O)����0��jnѨo��}UcG���ng+EIZ~�~㏔(@a)��Noy��'��	ڊ����[J���$�9���S���b��,��^�ΎQ�ByxﬅS�l>&�غx�qamr�AL;?�� �Fփ�H/ž
�oSQs�]�ͯ�P��"W��4�W��vx�H�l8��UK�聆p�`ဈ��J'՟�#��ha���\�����)
�{��X�-�A�����U8ar2�
�,�G�L6j�s��r�x�	�՞��, (��i��_��di�'t�7��
n�$���|:�hB�[�	0Cڼ���Vi#�?�̙�����<�ڞ��(��`w^CK(���B�`B�S�����2>��&�� ոpZ!U*W Iބ6m]op�`kM5#ꃜÕ��|��V[��ꦻ�����'ߖ*�\�;� C�г
c����iÅ)KfS����S>��� �Րu�>�͹I��
.��%t�n	6�%H��m#W4!�=���Pa��O= ���P o�a�h����9�=�@Ί�k��{��Q�9�f�1./�;�n(V���%�����P2	��uϝ={%(��<�g��Z�+څtؖۼS��K��;��E�h���!A���b�H��g�BW�P��J����;��qs¸���C���[
�^~���Ǎ%��Bu�9'�4)'���#���{�����N���0(�5��X��hڎѨ�k!���A��������!�R�x�g]���V�9$M!�M'��u�
�I�﫶f���X�= R��lҩ��ϰ;dKֻ�tH���۠X��|`y���@b��V�`��	>�B�*X��O�ݾ�(߀{2�ڞ?�~��r�Y�d@*,\}�1X�'~�f�v�֮���[���V?��q���j�X�Uk<��q�r����;�n٢YS����Hz�u�y�sWvk$�-ȷpo��<&K�t���6�Ӽf�����#ls�p8C�[��r�Bh�ʞ���kΈnt[X�6p��MRs���%�z�"������cNMY�i�D����� i_�)CMbj[IfO�}�NH��F��U}�%�x���p)�
>.-���oh��`�=g/�&W�V�
� ��q����S#͟roc%�HLeyJ�:uv�D~nB��G}���e��M��E���̫���{HJ�?TpD�	�PRP�J&��^d1��H�X_��B�%�cqV���=���ˤV��m4(�.V`�D.���#���DP�>4l���ݠSw5�#H���ZG���|I蝞A��;�ܰl���C��|���gu���8
�"u(�
[�.E�|��M���C�qG��>�n����V"��S�X��YQ��kS���F�RH/�΋�1�m�mE"��(6��5�p� s@b��!��y����d�4˻v��Y�;x[�,��$<[��c�Gm{cF4��������)I��m��"S�x5/��%Ny&~�&Np��{1��G�3�G��nK�r�ej��8ڣ�����_;d�?��jHv��᠙��,*AY�r�D_?�/�t���^ xZ�[���V'�@���G~��L����Ʀuu�YxjJ&�����iQ�z�G��^��Չ
?���"0�,$��vυ"����ŵ~�Þ��N��,ŋH�s�˜�wgI��!_@���0*H�a#jc����T��,3���#)��>>C.���!z���� xTQUݕ�|��;J��4J�5ѕ(�����@����+GP�Lk	���R�i٦���Z^i�JM�g����v�\/�8�ڃ�gg6�0���T���/�%�X�\����K;>��s�!����|�Ƶ��������.�3	�6��U��{��8�`�#"��p�1<��2�j�*�B���(T�v����������		�h���� ���8hL����H\�Y�R}��9Vhb��B�~�+����7�.�Hx#��J���s?>�=��{Ul��5±��t80�YW����`��$�_@8v�̢�R�������D(��"n(2D:x�l�8�8��^��r% M�+W�	��XN�Ԇ�p�Q��&Q�M� 20(��O#�4���tE�1'��bjᢪ�jUiKS��)�h������r�qoK�	g�I��˾u���Y9����=��6�~޻,bߞ�1�0zѰD+m{CC [�����HEiQ	S5��c ��G��
�l�j����H�X}dq>���� "�F9�r�!��$Ki����A���b����u�-iIb��k�S������vc��ұ`�����J�S���m�?���%�O�#��	��\K�;�ғw�i)��s��?M�f����?1SS/��6�U��;�ok�]���{X��x��T�O�I��`��������=cĂ��m.�����꿳M�=��/��Ȗ�m����)Z�6pd�a�wB2�˓�H����@�������ݺ����Lܝ)i�E�?l�4n@��&ܮ��,,���u��6-^F���cJ
[b����t�Y�����8���ƫEw��
P܈f�򆀳�+>��Qt2��Eگ������\{�X�4}�&��G9T���zW8��2m=ݷb�4���)_n��'�� dg����_U��k)�|��'	�M�&`�}Zk=��xY�n����a��S!�uO�=G��l]��%�����M�U������sOHp�#'��h�egI��;�B�5��B�����L[��]ݿ��Q� p*|[P�HZN�Y����H�����|g�o�Nw��3\�f��Qt������z�4{p`S�,�'�v�D@&������B�M�`��<{�q��D�jF�!��Ĺ����Ն�*�Z�f��/
#`����k{Tzq �+9&���ِj� �%��}���W]�:���#p��e���*٨)���լ�["�qU���#p�ս{�N�l�X�W��<`1�\���aS�*{���>�*_�-�:�ƒԃ��<��h*���a�l\��M~�\�N�H�*���/��>}��s����]ą9�?�]/%����e�	�9��w�jg�n(債�C�}��Z�
�e���ԥ6�1Qu�U�>�>©�u� x�+>sZ9�_�Q����o��l��fg��REN�n�;zj����o���-b���o~�4k\i�����2��0d���T��T�	_b���.Z�)I�J����̴a#Qo�op&��X���!Wt���I̲�"���A�$ߚ�c_����.Ua���y�@�mQ*�ڲ��yj5�R��>:�<y�zj��#o�l�s�&���͑,�8r0�A�aA���`}�X{?�}�MR�z1(�>�ۙ��DL�B�ĩ����$)��׉4[t���0��,�h�d��2��
�J�``q��i�-s�eyp`��$jЁ@I�ai-ߝ�x8�r�}ݮ�~!q�$��,Ռ�pq�t ð�f�����9,Al���� �)ᮉ�Ri(�Q�{���j;j8�}����:�	�����q�0�����)�e�a�-�O�}��c���u~ ߒ�D`3Z��.q�M4���a,��w<�[7~���+�D�r���,UN6�UI�d��v�����$b��7�d1�!Ŝ�(13��U�g�s-%%^[�{"`�-1�g�Я��4U݊I�v8X$��H2|ɖz�#Z8b����#0!�����X�%�j�R���jg�Z`HaP:g��GXw)���R��}<�Lp2��P}��x݌ 逍߂������כ��:�h��	Cw�.�l����W�$)�^��l��1��j��#<�<ۺ*wU��I~�tHU����T��P7m:K=eK�0Ƿz{��E����&l�˃�)|�7&�c߫Q��s�
��K��O�G6�g33]���	�9ڡL�2x9g8��"2[���@����f�!\�l4_`�?X�*|������
�f���n�k��+�(s]K�:� �������� ��Pgಊ�Kv�X<��i��0۱� ��o��>B6�/?)���x�`����o��/��a"�T'�Ż5���y�=_ڤ yo�T��m�g�W���#JM��As)�O����"o�o�[��`	�t�����/��,<���D讎�l�	3�Hʜ|�Fc�4,|td�	9H��\	��ώ$��-�_�ψƈ��l�~<�������l�P�"E=���*�
�e$�Di�d�����'ܠo�6̸�thFv:i3s�Z�>�D���4�
8Ơh�c����O+���l �ґ	�/��ķ��P
�S�.$�{쐂�����[�_7Ll~1����o|�9�q�V�y��Z�(,C*S�)yg�%� ��g�%.sc|�B@ۛ�׌�Kb��⾔eu�BeK1W�W�Wt�P��Sm ��A㻐��-3��{��+Ek�p�7��M>� �q<��0�(�ײ�wZ���?b"Z���MzK�u'-�?;����)�mz�U����u2KHD��2"�>q����,ˊ�c�b�gI-	�o�����������9Ⱥ��wyh�_�q�����8?�!s���)fx�JȬye�J���Ti���{�mM�w��b�a&���_DO��wQ?ןa2���$��j8���un���
~��zF��iS�N��6 ��w��j&g�
��Cޓ��Wi�:�:(�� �܄��_I�����τ `�c%v� N�;�8��}Wmu*�y{%P�q���q�Z�MɩKA`�I��wh[ Jn����	4�n�M&���\���s0�.�&4jh��%A�	���=�/�6��5���Z�1l�Ҟ�f��ǀ���;�^��$���n`JU��h��{�����)߈"D��)CDz�J���]/w`���9���n�j�-�\:�l�2��V}[�e2�zNݘ=����͜��p8��4R�4~�rJ�.�u��o٥(�}O�s���4T���g:�1GS
?ߐ��[j����.�=ʽٜm�?CA=�A�A�G�5p�"¨�?�I���R�UJ����T�
ȼ���7����b<�V6�w"�%Vz4�;�w��L�ͦ�+d��{��̷݋CB���|�O9X]�u����j6,eI��3\���<�]˃�ȏ^���h�X�t�	������ q�q+C��ֳ�'bzB���Pt�P�NءWA[]�z������;.�+���z����ĳ��;q�1��,�+�ɛ�cE����ګ����/�g�s��[�`��"��ͩ��֠�B`��?�Y����M�l�b%�U|]x��Ί�nP;�+�!4�E�g����A��V�1(ss"\�i5x��%ep�Udl<Գ�i�����Hֲ
�>���)�K\���;�+�"iV��f�E3X��M�5����nL_��U����0m�,�4�`�(5�t�V�SE�W/h�Ř�vݫ 4��ڽ!�F�����:�:ı�\��G7^[�M��r�)��K2߫4���Q�"ҍ�JiYe��Ӿ7;J�65��S;Eq�x� �~^B�_������kۄ�#@Q��5j�f�f'q�ja�'��C���T��5���.a��������7��b2fm������`�MiF��|x�#�@;������D�t�Xy�6��������J����_֪H�����w>�̋>=��$�Ҋn�I�{�R�=G�{k�i�ߘ��W���q�E
E:ݿ#٬S.���gl��REtx���E�c��B ��%�YB�b[~�UϿ���ap���@2܉���
-4��������E~$k����7hk��x2��g�l6'm�
�Q�	�{�6CB�<|O��y����p�fk'R@c��;I�:�(���CܧЯ�Hj7Ke[w|�=�(5vӽhʺ�<�;���xn���%��h�@������~�҇�#�M;RzO�~�5����+A"�{0szūQ���S�RU�Lv+����Q�B�f��c*�Pr��E�L$�2�r*��A�R���3�d�&��`�?N��(�|+b���
L[��ܯ�]�S,��:���z�:���j�Ƹ����Ay�z{f�/�@{��L��"U�"��S,��@>������rT��uI7���)ї�Hf��箄������I��ۿ~{�s��O�l\?���2nd�«��
��(��z&��fC��~�g�!J~!��KX��|)�D����sg;�H�Uu)���(�~��,&�wxO�8�w"s��G��J�m��tR�bt�r�qt��P9V�C�#�	���x���p��*&jB��(�P)�,r�y���X�Dk�4�1�M\B�C��qP1uj��r��*q��ȫ V���C�~%�1t+�O�Z�ҳ���v�,����Z�7��ʬ���'�j��-�I���)f}q��)�O��*S����H=��!���Ł\� Z���b��\IBO���\AuY�^�F�v�9"k^*(�}J�C|�3Σ��8���2iI���A�kݶA�^>A0s܀�l���`��옅d�c�����ْZ~�2��-�!��A�-:�����4$��D I@��.��cz�/<K|��hT8qa J.�����Vj��۰���k�R})$� �/S+���*��=�G�_�L��W�Q� ��p��36�,��I�:�����C�VG:p�W����3��@I�ukHi�`$��M=��Տ'p����Ms�$'�MN{��K��x�Z�4buvѼ��/I<�ag���ŭ����_�2���m3����z�o_-C��؃�2��zD���=�벐�jHD��]4����s����t��i)uR��X�ۺ��W)�~G��0��1n��i�����C�DrH�+D3*�ײ�l�<g�%7�.&,Q�D��r����I�N�2z^�=�յ��<@�^Upk#�sU�o��A/qnY����J��}��E7��n�5-{a=C�4N1��{$��ޢ;�|��(�=�X �Z)"J�wv����H)�K��q�X�{���"�#x��
�-<�EE��������+d��A���o��6Yh�/h���!�و��f�nfm%75�ݩ�黎c�\>��1oa@�7/p��`Y��儹E��-�2;��+2#v�:�M�A�B�m�o���aQ$v5|޴���f�Q2c��zI�Ut1O\y��N���oH2#�?��ܼ�dAkd0��$��x�{�<0��b�ep���0}O�PLK��5�QDh{H.��sD��+d/k*��!�q3l���r�������}y��QNsޔF�z����h����G���n�x����<��%����ɨ�)�T�+�Uubc�$.�\G2�
x��������An���&ʛ`��x�#�	h�/j-������m�J{Z-eN~�l�a�����c痞��k��YZ�F3/^�b��0Dt�.*s?.޴f�4`���36�E;6a�n�`�X8q����7T�慈�s��@�2;N��o���6��2���dh煗����~1���(р���#�����Ie ������nF�
�Dd�d�}�����Eؔ�����,�Q�av��ҕ�jA�%�l�*9m+��s�߀�*7��:�@ ����:��.�i�.��[g��$���1��/P�/&�UG�X��.��g��o,7��u+II��'�yD��<���ExOu'-�f�^c�]���Hۦ�z�J�Z�x9.���{-�6p�6̟͇̓��S�p�K� ���5��m�n~���ȥ�:'�3x����dg��k�`Nﴪ!<���BHĀZ�_���+
������)$�J��vב*� �z��W�r}z��b�[������l���40�@�h�?5q�B�W�����|ĩ��t����:��o$��I�i@�du�ԜG�}��+� �
�Ͱ��f	���zj�X�B��{��*�D"�%�^r��A�Z9��a|<d"���w�1�����7'ɳN`�&h�K���ly�W�nA}�h\$�R�����pk���(n�3�>��+����� j��;����2R���e���9�/��;8�e�KBҬ+W~�0�odϓ!�oւ ;�4�NRa{��JL]�_������_M���h��=W��s���DK�vqo��)e�g��f��^>��>��UB��*�^si>�:{�Tc�۠Q^�wSJy�*@=��qH�|+gc���%C 㝻��l֒�VЙց>��(�8;�)�Q�y˕������Sm�N�k�+	���u�4��u�->�9.�6�q�����^x
"��v�N�9���c�^eK9���S�(|�n�%^��)�,�^��p��*���tk�lJ�l���-�^� �gqk���L6%Cf���fO��?��:Ė���;��mV��O)��)>�:�ݦ�Y������!r���YM�F�.�YB��Rڷ�_�sI�vCj��T��}�.��ؙ[Z��Lua9�]�ً)���NZ�[+,�e�Z��ȧm��S�J�!X�U�E��Qh=vD�!a�T <�JV��)���,�o�`��/H �D�$M�[(l �C2a�Α���� x����yI�z�cN��*Q��M�y�N�-�X7A,��yց���N<Q~�R���"ܳ���n�T|w;�1kx���X�Ggi���Ly}�[�GP��"bT�Ҡ����i��
td`��4�w����ѫ���ot!!6�m�#g%�ݓ#@����V�8�Ū�6o�g�n�����j�� \��V{���y����v2ZA��,g �9���G�q㺁��lJ�E����@63�'	�K��A+[r^E45�)6Du���Vxu��/d$�Ԛ���zK�qb�4SYP:���6&�(S8�ؚ����֤�'��d!:��b�XT"Xc�t�co���_�W׹.�⚻�����tJJ�I��م� ����=�uk�Ń�w)��cOi�i���j��������(���ϩd��9d[�o[iDBS�������do�a�y�W7e� ��+ �=!��(G�5��@������̰�D���r�ǽ��Y*��+���ן~�yw���#S�٪z��*��̧vf>%|^� ��Nw�N4Pݓ�{ �C m3��鋆������w��̑��-@r��{E���n���"<¹j4���N%��
�����=�L|�|rM������8�g�n��l�RB�qwx�o��,9�
1��t.�8i ��{:iz����*Φ����\�51-ڡ	k���IG#A��B5��d�$Y�%��:܍Ztg�lBN0H��µ��ӕ]͏$���W�dk{��f���'�<�\>������l�`yᅨ��*�v�H^@|�߮5epBa��7O��L��O�9ū�`��?�e�n�n.Ը��Ͳ�������a�)P��O�� VM���w��S.�� �-
����]`�X�@�R(9��R+����%6�G,Fch����*1K�-�L-3$�DUɱ@��X�ᴨBR��c;�����yy�4h��eBg���ޭ�u4��̉qZ5�4����N	�!  �D)e��},m7l9��!���p�K1m/i.�o0��ZfB�<�/g�$h�4�Y옑e]���M{~�56�̿i@�`HFn��iD,{��͏a g��.	<��/1[���m{,��V��i����'anZPo%(�2��}ǖ)��}�Q��_A����)�s��6��*`�O�](�E�"�!�'�"�OJ���uWaҞh���?�eSݡ&�xx"r�T�N&�����~���W�����z��K��h��n~�n"�lS�g�|�rM'�F4s�!�~К5<��e����8fN�GJY\����j�D�E-��uZb�#|�R���qX)�+�B���V��q��$�s1�a-r'r.@܆�*�ZZ��4~�o���H���H*��-�P��d�V�����ːYդ���p�}�w�ꋑ O�[�p�F!����3��,J��s98|�r7���H�vLʶ�]�YrE]S#�(c«y����h HDE.�n�_�ͯ�oz�o�ӌ�����dm�d�����3ՒLS>Bta�P:_�F\z 2t S��d L͚����h�H�'b�J<�����z����c��w���Z<׆�����X/͟
2�<���V!�9+�6ڌ�7�K���>d�.�!��g�A���J�z@�*�9��X_h~
���8�2%�TU�
2N9,��Ǎ�D�#(�S��GI0d�~�b�Rvu�%�ɶeT[I�!��O�T�u�]���~#�t&4��M����Z����Y�����梻Ө���m�f��ƞ���C��/�qXM!{�fd��)�:�P$��!�m%v�fZ��su��=���9��ڻ`4Sl��<�0s���?Y�YtvF[�T[���$��w���%�
���N�k;���1�o��\t�O���պ��h'0����~t�r0��kd����O�iJp�b �ڴګ�Z�����%_�
��f�aC?%�D�צ@��ĳp\k.H��j&������r����7?.90�vVw'KZ�}D��N2�5Z��J�3�:�p�	����'Ixy�����c�dA�d�����@�3�B����<��#��}�>7P���x)`�?�'S��obƷbc���(��s &���+"*�2";�1�7-�&���GQ��}�� ��n���+5�R9�0na�M�my@�ÂF`T|̓�%����J�(E'yB��f��~nP�9���^����u���/�����&��3r�G�l��1��`:����|w��k	�Q��W�DM��o��2m7<:�,2`�㘸T� Ð�r��K� ��xk7�;��g��7�2Qr>�DG]Y�W8����E��˂�]o�� �3�+ȅF�=��IG���K��b_��q����~�sn��P\$��M��F����'�e��_lVJ*��bc�+�=#�s�����S-��]��Ԅ��,�g�4���V��ud�d��}'Ȗ��.�wT�(H��H�����,p����l�W+��^�p�1�k�%�FޖM%�e��V�6�\ ��gٰ:�Nb�82��}rC@9�N!�ǂ�h�@g_a�.��!\�{j�_w6UǌL8�8T��C:�M5�x^��7��࣒�����d/��opn�SA�"�{D�0��)�n���Q߮����� �U��	���F6Q������X��!��S�����yQp�1a���ƍ[��y7��MZ�dI<K3���5�PtF"�����<\v�>��&7a"�:zS�%\�Ð\9�[����U�	;�ڢ��̓���,�'�����)�g7"	���ЮQOmu�?��w��U�\�����y����-�Q�C����<A�ι�dU��5O�@m�T9�p>Y�#F���jQU�hӸ7�W�z
��X��a�� ,��om��	�^1����k�K>C��eN%6> Q���(��S��<���k(�V�;������PL�9�,���<�M��MB��AE3��F	C[����|Ҏj9���=�J&�M�>��2F�N^��?�N� ��J:��-�5�O��>���c��߷0�q�(e��Ū�Ec>�Fd)0��l.�C<�������Z) |�3a�I4Q&=��9lD��o�gO�%\�`d�7�yh�+��K³Lh]5w'+�BE�soOz��ɑ�Z�~�#��!$���,�؅����.��s�׽mr���n�qV�՟\������%��O��0�,�j�v;s@���T��w�������-��=�i�okS��Չ������[���T~��p.�Ҏsy�����L������}�BV�'���i����g��
U�5�1 n��)Ƌ���'?�CDa*��ρ)ʟ�^T]�Ռk$Dd�1)�q^uO�{[lA�)*S �yP��H��V���8{9J�j��?�8g�c�1Vn#�ob�Rnhȭt|���iq�2]�1+ݝ�`K�a��DG�	��Y'��Mz�]�f���9���G��`�m���[�����޵��������(+M�8�v�����ڡL�+�S��������w��0�Ӿ�>��a�@�1��f�ʅ���EU?�u�كg���e�cמo,ӡ�ҭ��rU"��ݷ�T�DHZ�� �쯣�(g������y�)IKm`9�F{�r\������2E��ԗ֋f����C����]7aS����Ntժ�R��g8W��*��Mw����9��e�d�3�cwg7�T ��"(}�B
�l�(��8ʻ-���5J�b��P�5t�N��	�M�K�%� J�v-���H"�o��b���8��6���z:��ݥOOm���=Ѷ5�tcSB�x]��w^��� x �+�ÚA_M�����.�NoP`���b�u�ik,8>�OzV�]��;V𑁍�`L)�#и������,�'{d#ȩ���4��,-@Β΅f�H��ۄ���y����HYm�����N@z	s�X���d��Z��,�o
ן��V=����xL1{讳���>n��r�h�K	�}r���v�,S�<��P��ͦ��<���T��J4,[ �P��&��c[�����e��lYV�C���(L��Vj�)��Y�P�B#;_�آ�m,!�E^
�L��_�����������3kF�b����@��$ơc�c�Dtu-`^��9�*�A�V��U�<�6�Cy��o�8ZA�P��4lj�d��A2s��Y��`�ͼ�Y#�H�3�i�@�<���Y�|��nǥC��EĢ�})��v��)]Z��m�z�̕�)��2��wE`�X(�(u{�BY�DR\��ՙJ�"a"s��=�;�k�t�� 9��i��3�5f��ud.�f��X�N6�w���?�*�0;"t������=�Zx��Z�[���qm[����o��}���'9t�o�]5�^�#�_���SW�.D�'���ׯ��j�^*����(ƶs�~ة�&�=�WK��ZN���3?3�B+��!�d��oR��7Q)*W������MqUk�H��>$�xu�3��Y YT��o�b�7x�AK5yr@d>�i�2ѵ�@c��d�@���)Ƈ���C�r�pO��~.ѾH�5�@���J���#4�+�O�Ի�)0z�3f�oջ76�_n6���ǒQ�]ȩ8ؤ=Pý� [M|���!��Ť!��;	<ȃS�am��n��o��bȏU!�{�a��c?�S�v4���cq�^���3wCj�I˫��dAg|�X�r��c�/և�4-5��l�p^v���~���V�(���\�� f���f�HuK].����̈����<c4q���In���4^��)�s�J���W��"u{�.�p���A�6-�a�c����Tu��h"e����\l!�y}�kQ��G���5�/��~�d�rT��"����.t��;�o��so�>�z	�ਕZ��w{5`uY�AAXG`��W8�A������n�b�]�eb��<���w~�%��1����_�B 6���Ih�CB�GZ���';v�6~s����s;��A��U�ӟj�g&��}�k���xl��鹍p�Z+#6^��~35�RH�2N����X��@<ң6�i�9��S��i�`�&�;��+��7<	��3�rZ����P��$[��$�&������-�B����0M�R���֧k���9�"0�Ό{h�+�_�B.��|�_qnBk���!Ҳ7��U0y����[���`mI�P�S���&��d�@i�$�V��D,�T�b����RF�$�@���������͊Iʱn$������R6���f������ �
%��w�c�W�j�O  񲼌چF��lgC���E��q$� ����g��&a��\��W�v(�S����<�3�i�<�Yu=o�RU���f�\"�r�]3���(Pͦ��Ps6����<a���I���M��K�E5�*��k�|
�������D1�-���M{�m�#��#Z�O�wƦ��u��\�a�r������U0?fg�=��
�:!\�X	�C=E�)�(������2�s�U�st�le�pq�W����-����<T��iͦ:Z�Ph,��4�M���׍�*�Oƽ+ފ��D��y��RK�b�5
�꙲���K8ű�]jX����WVL�N����4K�ʣ�AXy	��A���ݡ��'����TV� �Ë��af��h
d���7E}̨���oj�9F��;�w�7(���C˭C-%�gm����Tt*T^HPc�Tט�72b��&L�3���.	�L�O��_���������z`�<�Pe�z�"����1+W)0�漈��� ���_�HW�C�����J�.���𭴰�2]���"*�x@��U�m{��C'3~C��4s�y! �ުnkj�=�>]4�*���]��፾�J"wCT[Za%K���3��������3�bc�q"���*�dJsfQ��{$�5�t��E�Q�!��r'�0I�垝�ě�udu��d�}^�.�&"�J0�I�rCX�L���k�핿t^��Ci��;]k�5>[�)�)�c]� �R4��ns�X���a�t�z���+�P�:�z�.$�iNF)��wgӆ_F�Ъ*]g�G�Ab7��1+����w�����2��I>��{c��3M̤�B����,�v�Ho�;���[�Y��|tvV��QOW{�o&�t�|��ǎ%!Y�F6�f?��<l@�VShŲ����X�QRY�7,nJ��=�3W��`�y9�{��jC��ȟH�7�#	��k�z۴�j>n�V&��$������
_ɞ{��f��M>H4�oʱe���$��X[t#K��S�k�oّ_�~w]{��-I�q��}���D�k�G���æEB;W;�F�Y����G��N���de��l���$�D{g��"@,�w[��oU��zj3'2��岃ߨ�P�������ˣT�eD�3[����߁.l+`�3�P�0���_��9b������<��62���[P�C"��@AV��� �]OƎ��#ѨdҪ��L;ItOIc�S1�z�0��I�J�d3Tol��9�xUI�*y^���ՍNCu9d��I�z��QR���ٽZo�*c�>�o=��`�2������8�ƓB��r������=�O�#%�ȑL��FX�
�܌rx�T�8���;FT;O<.���2���9\M�V��f�AG�M�y�+F��]<G���UC�F��m������Ѡ?��L���񔜞� \L�0�\m�y=B�����A�� �z�CQ�j�*?�0������H��?C��
�LS�ř�����#���(�_7�q���L�*��yt]�Q[%���]j�Ku/BuɁB�Z��4
��{$����ͤ<���)=��=\�Y�1:�	��~@��_eN&����!�6]Ԃ�S�J� �������`I�Ҙ�)İ�Z�u��U�b��>&h�^�õ�/k�,���
�x�j'*m��뒭M۾���	��t�.>:-�t!d�(�]�RDy��{��Q8*)R���m��m�Q�)�s'�?�c\}��vJܱ� 9�gc�b���¢Z����v����s%y{U<[����H�#�x��'��U����C�k���^�� d�̂i��E���ܙ�=r�*ux֏,��Mu�y���t
ҚO�I��K����$�,b���*D��[�J��"���&��oVZ�BV+�8V���ƅ���R��|���z�i����-��Fػ�x���8��%횒�&-��tDe~���  �^T�����M��+de��:����=�(���+�Y�V�z=��rm��_��'R��|lY4� #�ݮ\(;Q��B ���\w
>�����m�d:�f���s9@������e>Y���"�x��*�̪���/�('��9?y�6飖6��%��g��"5�(�ֻay9��qIJ8�6��\��-xDH1��Xb)�L����o�����_+����4�yd{R1^z+ya:��)�'JpC������?"⌲8�:����E�0QCR}oCI�Y΁{����>�k����r$E�%�y�2�~pǿ��w�J�yo�q�qvmA�m_V`:�GY�}�j!���+93�A�(jp�#u�o��~u��ǧ�շ����hq�H�";��P��&M�ٸ�P�>(y2L�[�9\�p���

*^n�x�� ���@Z���]o��MX���g�v�(�=',v����H��Vj]K��ܯ��Mi	{[m�v��X�ڳ��W0��C����h:2aT�!�E�m4�C��Eq�v���ܚY��)m��t��DmV������V����·���0"� `�8���r-��v|^�;7s�Bn໪���4�vS0���E���/��4Oe��ٓ�`�0��O��MPڠ�qy�U�sg�%J$�`��h�}X,��=����&�Y 5�
��F�����@�!+7 ���2� m�M' OR�m�n�3w����E#9=H,�vipC�PhHr_餆3�(�]��P�ŕ��*K��Z��Qڙ��$���b9�/���G~~L�m��k��P�.CY� 5?�@:�-_��t;=����$�8E7���|Y��'�B
IN���q �$^s�q/�hԗ��m�'�T����f����'t� g��$m㔾u$�^d�
����rY�� �e[Ӿw��
��gJ��F�[��c �=�_��Ģ�k��G���V���"C��L�l�+ETʯ��0�C')�3�۳����^����܄�&�'�P���̭Kf��&��I(��eh�Ϙ�c��x=g"p�152��Y�B�1��Hd4����gDY:,�7�X�����X��z]{iMJz�&Z�6z�eLT�۪C���n����?��ܨ�_��VqL��K\�"N=��GpATѽ@��	a��7�QЅL�M�`��1'�0H+�g�3�!R�߬�E�ܶ�0�$;'#���+� (�$�5��fd7I�*28��������e|8	�4�Fx6R���=ι��� P�C~o���T,��ّ�j;2D&��W~�n��5UE~��v8������`L�3�Ϩ�f�B��Ǚ�#!�j�V��p$4���.�x&t8�˰�*C
xk��M�����O���3���M�\��YY�cn͙�H�&�6D�E�g˲ύ� G�o|M��@�j��2s@�����?ɝtpnV%v�9��=�����kI���(�(U�6޶'���n(ȉ<��mt�Ft/2Jc�O��މ�-�W��~�|a`�栦�W��x|��*�I����X
��:�C��:������
�a?*��q��d=�B�-čU#�x�*�c�Ҷ��e���m�`0ܒ��䞱� ����>T4=D����0@�����
jh�5!ʀyU�Sэ^��?}J�Eim�y^���Btx�'����+l"[�.a�����.���@׍NoWNC�!W���e�X�ݸ2����Ԩ0��@8ov2����:��R�V��	[@ �x�R�`��%P� wH;_Ǜ���Wٵu�4Ѧ��˷x�����T�f�G*�n.�j;;���w���c�vC;�hce�/m������sc�k��L���-x�;�#{ӖK7�PA}��r�V��gh'J��'��Zq/�,3)O0�OtʡT;�2��qu��(S�M�!�0�W�u��~��L�2n���z=�ޕd_lF�q�+�1�v9�S����X�8ש�0�|��.���b�e�]Z�# ,b�[١��ã�1_6W>��t�>�
���[��q@ql����)N@�n���b�? ڴ�%�FD.�-[���R'�|��#�!/�v�j��%)�b���֯���ll/���W�"�� �D(�ٶ��~���<�x�˫��/����~��X���%�����Gd��/�k֑���Ȫ�"��~����X]������Qe�}�ȍQ�e�
���i$tWȳ,!k��k?}C�F{�.��Ί�T옞��(+���!�J�I��`�Y�K��R�� ��Gq�f?�TO���*���
��x~�P�DPǿ�a�ď�dE�����/�׋�!�$/V%3�mVW�" �5c�p��w��Pi9�Ѯ�C��j�Z�W��U�Ad|kBⵅ�	�(�����p2-.Db��n��e_vv��9�_
QQ��LIf���q���J�D=c.l�w/w��a����t���xt�TЭ��^�B-[3-�#@E�/X ���E*�5�3�C�T>]@6~ �V��#���,oT=����4H2P%��v����/�Fe��}b�q;�"�=�C���|���N9y�j��lߟ�oe�c_S�����ɩ()*F�>��ϳ�r����o��_��ܷ���.{�$v�{������
8+A�H��U
�����M���J!�5�r�R8�r���ZR@�)��F��J�%��~%Y��6�vX�J>G��G�s�e�����{H}-�UH6�s���� ���yAI�;b��L��E{e���e�u(���"�o~d��Yg�5(�RS�0�&����e$v�>��2� ��;��	f[:ǫX���*1�P�$�<f���P*��5;�+�W؋W�3=���B�.���Ļe>�fI�2?7�_�����H��� UnF�.�&�\$�}u�r���Jf����| 9Ƶ_����sJ���3��C%�7�l��>wO�M��GAy���pN�_G��ҭحb!t�L{`������z�n��~�s�$V���4�3?�o�q��%t�.x'Q��T��~�B����}���ݥ�k 9������Y�TXA��Q�V�����}(��+�0q��J���[���o�pV۞?��`�:,��^}9���E�w���.�UR_�1�m^d��1�gFC�
9�^ґ�̿�U��&�	aX������fY��_�x�s}�f	%����ɻ��q6"/$wl�F��F#[!?s�qT��avrĞ�`��edQ�B�,J6�zگ'���l*.cS}�l�	������Z�}}
�ǯ?Sn��h���L	�9!�:�!zϴ���� _�m={#Ew �Ҁar
���?�
�����!Gn���xD�{Au3E�fRq�w�%?�5u��UK�qK ��t��֜�oD��wTz-�Aq�s+ 2Y�������aHv��e�,�h#+ٽZ�s�g��4A�� .P/C��������:�����������.�P�O�H�����I�(8掽5�>���1�>d[	g��AO��n6�'y�A�Ou�+]um�%���!�e���0��Iϧz��n/k\�j�����Xx�:�C��<�!U����$kq�fH��Ap 3Y���>\j)[@�No�H݌g�7�F�� �C�́ث��i�ʢ���J��K��ꡞ Ps'C�� s���x$��Uc=~|���c �^/[�,Z�Թ@�#������f�ΧȾƓi�Xtf��4���\��nW����
���Fa6+>��ڌo`賐r�� }�},e4~�M�K<k�{��4����m�`	y���0��<K�a�I#Ӗ�D(���[�$�z����8kY�ZtoI����I�>Ǘ}��!�V�槢�]��i��w�5�,�'���) FzU�ٱr�/��cZ5U��'F�Dj�S����ah��	)�S���'�� G�DtL%�(J����,���4pw��zf1|��ҙ�B�Z����8yzy��_)v��Oa�����������~��RXL�\\�f�Ƹj��!�>�-�C���'{P�?��8�L���a��x̀�� �&��y6w�Ͷ��dH�;�m����B�:�-�� ��jf�>&����y��j�}E��s8�J�Џd{�V��ʬ��k�x7)%1g�Y��w�es����6��a��K�2B�����3�s�����gm�]��ۜ�W��ܩNdN\�>�&-j��B�{�����������0.�	K�]*����Vu�ڪ�њwn�W�`~�f�hn`qyb:PPe��ܲ�Q)c�5
^�7
�O���|'<�2^H4����ji(r[L��Y�Y!���|���Y>��`q����,M��W���9�y+�?���,��m+��F�fM����5�����/"���H'��懻�)x���ʅ�r=��i�N�071RAZ�l% ��Gt'?Ab����SќY�ա�MҒ�N��M�������Q`W�Q>z�47�D��H�B�K�	:���ߡЮ�g�?�H� ��yu����L�V5�_Lv�t9"��Y�����F�{ٹ	.�v�%�a�%�XN2� �^o����XDEH����<e��M��rJ��K���P,+�c��6����/�	�h����S�ꘇ�#D,_�܈��W��u~��Y��qu#����0N�o8e]���ߩ�r�b�a���`�f��A�W�|U�5'���CU����p�O�t�OK�%jA��|l'���e?�y�bmRs蚝��fy��J~��F-��_��?G�]XQ9ۑ�1;Σ�ؔ'A�4��ջ{�jv��K��5	,����Lj��N�p����gn��Q��@�6NcyS�(����-�z�D��KFc1�Z:i�s;�1��(��}�ˈ�]�ʂ��T5�{
�R��9巛D�V��=�@�1��,V)�cK׮�D~���O��Z�ޱ�ee/�����ׯ?&�Q�]7V�D��=�H4ʤ���n`��[�� H�>�Y�l�4!6d�����b���i�o;]�#��&��Vx��5����M����!wO���ခ2>�m���K ǄOf�vG���d��rD�1I�p��,�t��a���Mo�Ey��em��azU�?��>������'�hA~?����E�������V�������m�[@f��L��x�A��X��tUv��5�s�c��u���Ri^O� s2RZ�HZ�FJ����͢f~�����b{-�3��Bc�l�k?ۜ���hJ�W�49� �,|u��p�,nG#�؆,�K����в�ըNaB��P��j8 ��U��o1Q/��%�%=�E��*{O�a��B��ߩʼ 9-�**��������v'5�(��e�sW�����9�6�.KpVn���ԭ`���z����>�ܱ�R,�[�q9��{�x�`�O�Ͷ� �:�[�a��G���T�������{ƘxX;��o�펰3fJە��)���G�튊��~�x��_&�x՗*�ר��=8�Pd=G�RVs���w��i,rz�,3J�����*��ә`�-ޮ&6�B�0�^M�Ĕ4�	#ZP�]�����2k�w���q|(��B����n����������Χ��Q� �TN��Ҭ������#�-�� _7�zCoor��o�74�u���ᆌ��Ƿ(�Nfc�i��jD[|�,���7�|�4�k�^-e�J&e$�&����m���_^�[�ib*)��m�5�4aeH�}�Muq�Qڡ�r����h�d�kE���P>-�s�����J���D�f��,�-�
������TưUD����m~ç�d�X<�AV�N׉H���Bq���hw4����N %��?YQݗ&��r}ImPEM�YP'J���q�Vnm&�&{9P��eߓ�q��"lM1yM��)�9)4�$��x���U���w����_KtՆ����ݹ8zn��}���C�_���~)i��{L�.-H@(K�+Hr�c���$�����3G~E�@�P����[�\����B�=�p�a�f�f�Jt����f/��$Q�/(�z"ݔh���E��A�OJ����ߌ5��Ն�;Rsc'�!8Fq���%�'��'�TK/}�����زJ\�B�`�t����P��yGq�6�+�v��fJ�v8M1eȂ�1�x��C��@��{���8D`X�۩���i�{�����AT��@��$�d�!n�-5;Q�F>ȃ)E�*�aX����gѭ@�/��:	'҃]����3k{��(M���P��_��a�i8~?���&u�~GwMw�k���%�1�q��krIb���iO04�,�"%#�@��m,�w���N���O�	V�ϊ����lP�L<�?��<{C�P4m�̩�m���54�Z'�?��m�ǅDM���Zc�iSa��$��c�/�I���\̦�;�U�j�{�ɻ��s�	 6E%Z��Ҧ�B��E�L���N�ʒH�^B�) j���d�r��OV)����V�)Ϻ"��VJ�j�#lH�e�a�q���]2�p�b�UJ|U�2������D�5�y[�:�U�?�������q�m��:C�{$H���D�Z�!=K�M�4�;}��X���`
���ց�g�N���p*�0G�v�d��� px�xY7��򲢂P��NA(0NVF�@h|5k�T7�0p�ԃG�\{!�Q8F|�o2t.�T��B�卙��8;�dI!����sK�x�����&��H^���Ĩg@
�j��=����!�i�M�m����̢�L�CQ�r)5#`e��
0FvQ�e�U21�v/�5�l��_��I"���V������\HϘ��P����%\�1���X�2���S(��5���c�z��ԍ�����Nzԯ13��׫.�I���<Z*�1�ϖ�"u+���`=yk��=�����7�����������O����b�j����R=�����h`�A�Җ�XW�Sґb�#�� �� �W�������n� B(|���q�S�¯{��Ni�[e��$J�5�n����B��|�o���3�<ޑ܎��W�)_��BY$�{��Ӥ�ǎP�#�^��0�����@�I���#[��o�,~�Z� 0|���%���A�$����";����oL�[������˛�,b���yV�$�w��to���p�i��~�y]~�ŢsQ��daU�����U���q:�+y��/"�J1W�+��1�1�d���?���K;P��n�C�o��n�#�/M� &jմ��1�^&jk�a�k���U����� ��S���5��.l�.�4�f��<>�JQ4�nN_�o��q���k%�S��8��DҊ>Z�^=�)"����}�bi��d� M*wn�+����	9ڷ��ˈK�ڙ_+���T!���pv��e�%�6��\ͮښ�ߊ�����/���*̽q�h�+~6�)�pb�8��ؠwɜ�c�y��]EAaEv,��^(S��iek831fع�O�Ôc��XL��@����;����Y4���nj
�B���(`�A���
�jHi]
~����f@�y/��*�Z,��Ps���V�b��Gn�f���� [�)'�>
_�Ѿd�$7��ˎ���Z���J��6ª�ij�|F��T�����=?<7��W5���1�N���Gr`e�K�K攎z�ED��w��7��Ɯ9��{�"��,�y��+��qߙ*fg|l�X�[9�����Y$ �ǽ�k��3�|�����K͍S��hm�mN��1��P0W�-�u�y���x��?����Sc�r+f���eX`O���3����*Xl�Zt�c:�r�w��|����EN��*ߌ:��5���e6��z�.&�ߡe�ż��r<� v��ޢ�-kM�
�ϐĂ��Z�������fw+�ؾ�c"}�*B�h���Ec�Z�ۼBE�f��G�($$��P�˭�=�Hb0��1�+V�W�G��\���G���	k��̼^���
=~���٪��ʻ�?�r^�_���CB<�o �z&��Y(�Lsc�(����_�rD;ɘ%t���B�~0�3l�"���n�/���e���7�55VL����Q$��L�g��h�Xb�h2�|ƨԯ]AR�A�P�?�n��P��"��T@w��)DӪ#�;��-��x�?^�Fo��lQ�xW�!�m${�����k݇�Ȝz��y�V���3�ʻo��RD���025���%��J[9B�{Y��6T�Z�05V����PLO3]�GHMD�'΄eȨ��{�`~'N gsCja�Wv�x?��*S��jH���"��R�,�F�\y�>�X�}��"*[�� �#�3��=`mi�s�j,��r�Hʨ���[ܠ����\�A�I�j6�m�d<�LtE=|I�ni ����V����~Ǘ��iU����d�O`ڐ�~�J0������8B0˵�k�w �|Wywtg.ם ��um�>k*S��k1z�̆��)%UL<H�|{)�7�4\o���{P7jl�<�{nL���U�ȧ�}��m@��8%Ђk����N= �������z�1�����w|�]�@��I3����ݦlq��X&�y�`?�%��_is�(�����d�ȹc���q�,XS��>8�w���'f)\��A��8� �rM6��Ė��H����+r7_�D�z��),pb�w�)y]2��԰4��ջF^�m#��(Z��Zr�������3�_F��ܗʙc>�g�ƏmO����Hfd�fi�-f�u�!���ޖ4���
�r.3��p�}d�#��5����<��O�iP݇6ƒ[J3t�Α�%��-�=�@<_X��IqLT�HA~#*��5�ބ�i��{[Lv��=�p*B$"'ggq�Rs� x3c�?t�}(l-ih��#�����;K���L�C:Ձ�b��G*>��Nu�$�)���ڢWi�����7�H��v�j6�D:����c:���mzQ&��Q��H��J d�a��\8ț�!�#�+��NAs�,���-���iڿ�-%��&�Q�c�}g��6]beZAI���{OG%�2����[`��������y���TK�v�E�Ra2b��F� ���!gqU��kvi�U��Ύ=
	�s$�5�4>~+�*o6R��E'!���YJs�aS2� 82/��=K���>�#ł!�rz�ٞ([�n��	�!gV��,��/,��?��"s�2�#���˨�Mi�Z��q�z~<�\�6Z~��P��1����oܾ�=;)�Di��L
Ln�b����;������M��iC����H�PwXX�%�1�`�3�m ��!��Jy�b�R��Փ��yN6Ǡ:��n�N|��И�Uz�et�����<�Ȁ�j0f
8��?-�8�����qa����y��-��?��,�	?L������;���jwFx�:����d��g\�l_?��W%���-�9�Q������0��M��
���\d7]�^����6���8�\�Ae��X��ugv1h�q��K���%1_��I�9�pmj���*�=OUd�Øvp(BFϾ�]�H�T�N���Dʬ䀙j��
��ss��p.��|�k�>.��uU�(���Lt-��4�x�N	JW��Xq[kLUa豮�)Or���1��?<��*���fg��S5��iƐl@Ck����v��</f���	 f��</G���G�CoC���@��Jp�!�����!O�aUz��� kR�i״�:���V�Y���s��x~��C:���L�sMd�Xݾ�qL���YW�!Y��y�C��+���u�:�����:����'ۨSg����2��b	u�*����~�T�P5�$��*�;w��F����Q�Z�^�`�kn���e� \J0�I��P��+#{` awRJ�D���6�+s�|�V���H8���m�sQ�P���׌�[���]�>-Y���}����R 7��T�0��	p뾰��S7(xƐ{��\� ��*��ϣ���ވ�@K۔+����-B�������"�t1�JQ�N!ٛ�ynpM=�%X��~g=��n�9ފ͂�q�<�S�劗 +�d#J�����2h��^��j:��a �)���J����9��Jeي�b>�pb�����U�dp�| :{'�:��c���=���ۉ�g�T��LEd�/V���k�ezK��-��[?��F�����$�
C9m��O�A�j]P�����q�ZF_�)X\��&%xV�\��`,�rrܡ[`�Nܲ�����/ݠ���On�CH���~]���:'!�7Z%�zP����qV��d| L��?���~`�8�Ou	H�/ju�+�c�_�U�L
�H�P<HH�
?���)�>�i �x�A3>��ݤ����r�5�*�m;	��$ɴ��ESn���`��U�HO:�la<S\�b���6ѧT�Z��s�:)¿��g��Iʽ��N���o~Q��8���P7QeF������Xeyss#&��t�,i���P/���̱@Kc�ڴ�п1�&2P�H�II�k���趝� �6�N�����E�\��j��g��Ze��P�.mW��pZDsf��T�ыG����Y=)jҧ=Sh+~�s$��p�i����òH��fkM�e���u��O9��I!r�"�2��Q$k1oK	�&�7��|t��-��L��,LHI~���M8c�A?�P]=�C����mw����EW��E�_�D�O��&��}
`����+�v�Lk�Ѩ�壗���M��J�x����T�~�����3P5>#�h'P�:����e���ij+R���R3�� c�냙�f1~�.&��h�;���n�ހ��)"%�/A���[.J�C�)�6w��_N��I����F�HJu8�M�E0~��^�dD?@�J�y0g�6Ƣ+)K`%��_���N6q��J��eq�D����٫t���N��_�P҇"R���}����ZEU�?9�	;�Gƽ�bJˬ�|�._���Z�I��c���9�ر[ii��Kl B/�û��lw����M���d��m�T
0�`q��ɼP�,%�7<ُ�I�a���%?_�8K�j�sV�
�ODXJ5��[���j�.V�v��攅ג;*�&���.��g�@�̭�5�r'�⻫T��`Zo>X��i��0R���ab�������M���̊��ݘ�HJu#"?WM���>uZֻ��C�-�_�]Q��k�\�l��t_vvpw�3tI��A�Gj�Ŏ��-����`%{�w,M��x�2����9�}�.䝩�\�siǂ��:}6Dh�W4�J�F�5�zXe������°~]��]���RC ����l]Q�(�L<��gI�i� �J޵���?i�*P�����k���#����~�6�z?%�D���3M�S&��� $Ǚ�xbL�@�@�B�;�ȕ� _���n��3�ř�u�>Z�'�Q�
a����*7�	B�Ej?X�a�vx��C�������C�����]�wڽ]�	���\)?�ա+���݂ɷ����W�f��Xר
7a6��9F����z�L�CS�>�N
������
�3�F;���0.D;5����cb�����BA����*N�@��E0��04��5�}��p���%a��o$�2M�j�y��Z�z��	\�g�P�#2� ��m9�x��Ũ|�@�ռ@�T�c�Y:�|9(�HR�Z���q�j�#ūw�:�ź�0Q�<:����J�4��s">8Ũ�f��>a�B���]�o������ϦX�7����� T�ü���'n�l�-����f5�4�YFq|�\ojA�W?�q���v�;�(1+�nE��${ޭ]̬��� ���<c�#l��i�ˢoU��hؑuS��؜�%���ZK�����PD.l�[W��E�م�Gy�yF�P����ל�]��b4~��^'����`P51?t�>.NQE�]Aɧ�9��+��q��1�O��B�Yu�h=����k���e���jS���*�wf��&�I!ATS�W5��ҁB�B;<����q��|�n��}���+0���1�f�$mBߞ╪�0��A&������̞�OztbgRl3�؜eiS8�Ȅ��*[�S]#4�5b�Y�L]�ȱñ�u����3 ���r�����@�BdE"��Kr���z���y��$���ci?�37N� .F�G�Q!p��`
�#z��qw��Wl����4.� ���"$�*���x������o@9U�m�w�a�[`��%�A���6�H¤�dR?z?�T,���B�P���9kP=�q�����C���1I<o�^����a��7y��d�R3��Xdz'�g��Ԅ�(F
Vg�+��\ԛ"^P{��|2}�b�t�O�HC�L#�p������v����o#�����<��%�Ŭy�o���UdJLf��.��#��]o���[-X(��9X��k�܆Q���Ю��:F�5��&-i�V�@z
�m�u���Mؑ�t@�i��uJ�D��O���Ƚ�9��%Z�|+��3�@�|R��j��}ݮ6��	���B(��N��i��2|����~�΁�`����#���C,�|!	���q�hcM��gw��b���{4�zC^���L����o����_������+�v`��'G���{f�1�1�Z<P�<��~��]�2��o�za��[C�ɸ!���VwL�����)�'R�a��?\�`��7��U�7������Bq}&�Z<`3������\0?NKb�n�L�֥����eM�˝��c�����=�ĥ&n?>�	�;�r��|�R���Y=�,Z!��&|S?�F�U�noI6��bQ��5�����O��TP��\�2�B ܍$��Y�G��8��Z��-��g�����Qڣ�|�q�/<7��/��ZA�}8	��e�� ?]%�F�w@���d�G$��\gr"e�W������#Y�vO��=m��i��6s�z(��Ǳ,����TB�15)�BAS�y��ݵl��-���=�Dm�d�U�kJ�V��;��HKH#�֊��Dh�+0�;���ˠoE\F�����Y��?N2����\�J�o�:ˑ�[d�~��D���ٱ�\�lӪ�E�9�<�R�3�7�Eā<������˹�2�G)݁U��c&"au��L��:ne���ew*/Fb�ߛ���l4���1�q<S���ɍ��,��e5KL�^8�P��ω����P�T=+G3f�N	�yMc��sE��ʈ�a��hjMݼ`��K9��c���9����tE�Ywg�-�B_��f=a<B���'惡�����9+\�B����aԤ}�h��ΞR(�lBN�&�;���y\����w���}��	n�F��9��3��[��������l�$R�
{��.R�FdY_\���]d��w$��bnQ8�=H�'Ϧ��H$�j&�CH6�笀=�荧��b��)��#����@;v{	�A�p�����W(RvV?.�..9X��	��&oU:>*��ʺkd���l�:#�)v]�_������cćYZ��*z><����\Ȧ(��@���H��\��[ΐ��!a��?L�+lH>�GK�4�6:��'�2� E�]c�_�U��˟�+`i�LIb�!��;�����z��a�8�l�O^_;i_�����R��j�w���6�iu_��^ۉ%24%�|�a���1E�B��`#��_��C�z)r�L�2	���u3l^��[39���a��=BE�Դ����9�?���P����}
��ӥ_�
�C?�����j�'QpÏbo
�lD+d�`>��ֺ5�E ް?%P���i�&2'�D�)X�-k�������\#���	��`����H��T���q�����@_v����E;P.��>�r/1�@[���*�_d8��Xo)@�� ��g����̼�L��c̲}t$ے��+�g�.�{�]iv���s����=HZp�	G>��������x˲��P� �`��y����w��8��zy�͎��E�jB�ۚ��x�e
�.��Ċּ����p�Phrm�ћ��k#;�"�{�v��M�g���gX}5M�}�s�k��$-*R#�IȲ��R�����>��t�7�}e�����B�3���x�/�
�M�fE�xʐ-,`k҂l����;��n��<=�R6(`H��X��.�i��Cl���݀֗I� S�%+r���m%0��`�'�a�U1j�<I:c������^5e�`�NnB/2�S��+���.O���C�ҏ~�L�E�!Ԕ�����%L����]�؉͎_�n�m)�m2�@����ռ{5{��h��D��N"
�������%!'���F��")g���v���}��$�0ȃ���3�cq5Ϫ.�g����V
���H慪G���f���
�n�/m�Hyh��9 `��'�ɽ����oy$a�@�4��$��AT�b��f;��	��j�0�s���ht�t�߉�� a-����Q~Z� ���`�JB�Up"t���`�i�EU����/��F&��]~lv-�h��L��&S@�v�nX7��?Z
��f�����ﾺf�|P�Y0b��a��3�H�Ν��Cg㶎��!K{�t�'#�L�2.�7+��}i|N���o�\�P[qRKM^!B�)^h𱙂�O���-�Vx�D�+��^�%ؽ���I�ϲ�,w�Z�����3�z�m�e�p.�k�9��_Q�O�GQ�p c���3��y�:*`�>���b�7�ǳq8��)����.�{�U/bS�܉��ؔՍ�]CexD}��.��.�$�\%�u�`d�F�4Hʬ��^G3����}Z�������^,/s�����.�c꨽�Ny�!�������T�^�����&��d��dR���އEK\2?&�8/���'�hCv%d�P�Pـ�ʂ�������7ɦ:ެǒ�<�b�y�F��J�"�,�AG�O)J�����{ƩY��!�Ѧ��P�GI+m��?���k���y��B[�a�)ۓEBD���#�/߅AP��a��rX���{v��%Un�F�!�b�@�Tte�՘�S�t����Y��Xޘ��񻲩K�y��}��´:�h�c`�3��<v�X� ���u��;�.!�H���8믿!
��:�k��aR��yB#c0˖Ն1�%��F��'�`��:j4b�k���F
�C j%��H�v��#��3�[�&]�Iu�Ч��B �nsHA84�ߗ�K���� v�@J�^��NpC�������{��Z̳;~�>j�6��C����2���g�条�л����\�A���9�>V3��$Xk��?<Y��/�� �Mvq�;�I[Fs$[%�����5��ӺO�2����biy�tXܩcR���~U LS俺	����t�	L�P���Qȫ���U%V�g.�m��v��۳T�����,�9�'���%�9��@����Z�6��ec0�S�%���ƺ���D���(�Z���P{��֯fI�:���en��b!� 8�1�/p�+m	���]G(+�ȟC,/'�r�@� �R�?!L�*�?"*k�^Z���#��ѹ�|��o�{�ܙD\�*#��˱�R�fNeѹ�	X��}~WK��]v�u�.�7��z؍����;�뽒.�&Q��n�^��F���;�aS��^�)��?^Bԭ�fS&A�g-Cn���� &�o�c4k���c��v8[+!^Xؑ�^�C^���f��vpk���EE��b?m/��	�(���	5�W�0cyer�$�Ƣ(���LMߞ�)җU������Cr��bZ���P��?�5�b�m����kIܳ��:�JH�
�\ւӵ���|���A��.A�M?6d'~��?���1�ļ�OUmKi�H���Y4�p#DM_��Q)����)C��Zϐ�tB��pЕO	���KE���T�?~z�1
B�)�Xn_��Oh�۽a�W@���4�sGB��� �+)v���r�<���Ӡ�ƻ�ʣ�[9��2�@e�l�`�m���~�K
�{�~Q��$'�=���=��ǀ_AjI�0)�OI��V�,�^��i*�4Ӭ���/ʆA�rE!�F���֩6)ZLH� ��f�*���ɚ��{\�eN��](Q��3�� �lρ�@�n�uG���ΧAp�����	��0_U��:u��U�Sü�ǭ^��B��e��3W�2=
�¡��I����vEY�`�`���(u��v��ڤA�Z�/�7�]:h[7N[��>��E�ݽ����J�M<���%Af1���M�3N{EQ��i���r+� fl�h�a�Z\�w.ĚXV�\|��_��PZg��GQFo��Ӈ��4���<�d�ϋ�xO&� ��6�C�o4�g�����c�^�;uyl���~�۠�������_ɇkݻ��#-IjL�p\ξ��]=3�JUg��kP	��t�:�i���I�!�1r%�"�&���%Tq9� ��s�)�C��V�&Z $��DQ�7a�ֵ�bY�'�p/B�hظ��]T鏈��$�.�sʸ?�Z�<-�����ˤ�H��7���B�-�������� �]}?%细굯��V��[�YY��
X�&Mm��AH;�6pԢ�V}v�|&�Q�T^��4O�#�E��m�Fك:��S��ĥ-)�d��,��u���W�N��[��w�ϧ.U"�\!�<d��:���S�+&�Ҭ��? d�� lva� ��v%�tbr:���ӎ5)��A�o�+62���1��ڳ5#��Y������u�8���Q'`��`��FD^�[G�	2`�B|�R�x��9i���!�u����=v�X�\��a�Pj3l���r�7��G3pl�K��c�:N�A>6"�F����0qk~:b�^��m��69+%T����P�=r�A���j�B�&�x.�:����8��ci9���Z �!+�| L�G1Z���΀�찰� �Qv�\�����/�+��(�7��K��!��<1)�z��f4���y�^��I?ij�
]��Z��?��-�
3�0���I�_�7�X����ғ�p>1�������g��6��	(�'PU�s�q�d0���cSi=��a*�k��INx9*�J6��Ci
��ub>�;�M��(m�+�{�Q�%��C�ΛX��Xz�
}p ��Q	
��t�%���M9W�
$�;��8�E�o�7#��(����c��D�.�b{�n�,}�yZ� w\�X����T.�dQ(���Ք/��s5��� ~EgD0�V��c�d�f���'�1JS)X��G>	��J#�����%~�8,��fz����1�B~�¿}�Z���	a5��2�<ۤM7v����T/�?�h$C{��=W��C���=�s�f�}��`9�?yKÒ �u��|L�V�w�\1#Nt����M����TSlamC��0<�R��k!�Ƚ�p�6c1�\�I���D�+�lC6M4tS|���j|��-���>��'��9u���dVT��3��H��3�=��B2�Vz��G��3���ψ?����_�ߴ)>�*Yx�ĭ^�� ^�.͂
i�)r<$4�̐�[�'�=+it�!��&&�Oʝu���d���(�N�`��L�옓!T���qy1�M>�+���KR�oQ	Gc�F0�&R,x����'�L� Mr�7�)r�giJ�ȪD�Q�3��nZ�� .��=w�1�X7����Um܌ݼ�� Z��YuK�e�X��� .���m���n���b��;L��	빠vrȰ��	���'UL3T��xt�����XΚ�N�O�� �IsCBA E	̽:
 <���l�sbz,I��
ӒGiP�5��g�xƬk���g���,7�D���G������k������to�[`O8������,�Ke�&\�Oȱ���aس�l�w��U!ݕ��Ҏ�x��Z΄h	�o2�EѲH~mL�K��E�z~0�G����-fO(���p�hy��Dr��zՕA�p�������h�KE�,��u�׻P�E���)h�Ϲ�e�Qڹ�D�+�� ���ۃ�ـF�\h���j������9��]�3�H�u��# _Tp���[V�: ���χ�..���h�,_����(�Z�xz7}E��D����Gm��t9Z�y3��j/e!��[�aR�?�<�2�F�q�������YK{b�[:�B��~_�0�@��)_[�:*Q0V��`]}f[�2=?e��'p6+���v�U�����n��{�w0`aAߓ[z�/�x������N{�N�|�,�;Ɗf�˖[�ɠ���C�Jl�r���zj��c�F�����@��p�(W��H�\����On�I�37��}�eH���ujG�z#1��7e�X�,�&n@�H�B5+S"��j-Ay:P�Tt��\`��B@f8�N3�8�<�B�����D�u����.z\'��j.��M�C����1 ���S�)ӊ�Z/MaJ�����l(�
��� ��߾��	Yiy�����<&��&����M�83ve̉c��t�x&�!,��<s#dr��G��x8q�=�ePc�d�|���&/e�/�0�:h�G0����y�2_,'�t�� #1�򔨁G��+R/99�]]�ͻ�F�<�_���%%��{��ӂJ�I XA͓�G4O�cHS^�O6^��Ov���'�O���)�CQm��)�
R�e��׉ �����~f�'������E��1��r�v�9�:�%� ���θeV���c���걣{V�^�� �G�(vQ����#aa-���u�㈡�K4Cd�-?@� @s'׀�F�����|���q�u(CQ��I�V�;l�r�y�������Rq���e�F�,�6��5M˔���ک�;�ܕ��B�A�W~[*��A���ba�8ST�Uk�NP�H��k� ��GoW��e���@ʮcց뱟����G��@��'�.LK�aٛ�E%��<��#_9Y���)�U��1+OTqx�>6|'�R���w���[ɻ]��	�D�QZ-Oy���iG�kh/՝fn����i�f1U��~&��W�\��Q�
���as9bՋ����%qA������t�Y�Ueo����o!��T�{g�����"�A\�s˜𑢖�ei�;���ǵ�7�T��~�Ę������;�=Y#�@?�Ul;)?xL�zD�.r/t�`�D�\1��sW
1Զ8ۑk9B,��/O���Q��7�%���;���zڒ���sp�ܡ��c5��J^W.��&��(���='�qc����,��@/�GazZC�$t����nnX��x-B��&w���Һ�I �O��������A�S�N׏��%�I��s��jEM?����y��7�)�2���B��#�p��Ӌn\	�SE�5aV�I1���C���@�#�g8�T������7&HL���4|�e�<N�`mkE�9��mP��P4y D�P\�t�'t�Gp�)�N,� h���F�/s�Z�NK!�M�E�TCˡ/�k�H��6�
H&�*�ݺ%X�9��G픃`��ܓ�M6�1����s�l�ǿ��iM�����9�~o��Q� xUe� |L��En�_5�,;�v�6m48p_�|L�o� �]b.�4�^�N�G� =%ʹ���d"^�x��\�>�8��_po��£�z��N�e?J��o��e������J�,�� "�e܀�D�B��̦�퍀Np�����b��T;u�T�\(�=A�9\S���{T��1�q�U��Zm������W:��\9�6=�>��4�/M����MR�L�e����ܖaT��\��>��,:a��Q�Cq��5���;�r�E�e,Q&)�ʤ�pd�+7���2���h�*�Z�'�y#�`$�h�?�|/���D�
��;y0#$�b��z�t�[����##{�@�Y�c他��[�b�۷݅Q�f"!Y7Ud��{����`�'fS1>�DN}��n����/Q¦��kp�=��������a ��5Q���y�nX:/�Ozȷ~6�9���o��^�Շ�+p�
���� ����t�����������Ո�m6��J*3�(��pks�a������4���l7Ck�ٯ��}B��Ȧ<�Թm+���I�]�o�����9��kb� �y�_�����/��2`�րq��lG�a|�Ģ�@���_��
�S��l�����C����S˖T�g3]'������ƥ��bH��?��z��3!�
y��V��{0e<u��S���y�[
���[����C��̠�\�|w�--M?\F����_�/��΂���P��"ԍssb�������s�kT/<c�ى2F$���D9�1���5�S@�+:�����n�F����l[������C�?��B��25��~4L+� ���p�5�¨\�(��F��ۏ\��T7�`�[62C�M�;�y��8T�!R;���1�!�o�<�f�������+$�%����,�A`�8t��p���o4���>ڶǕO��P��~�[���y5IcV��D�3�[���9[��Y�)��ƍ�<�bU��o��8s��	\�oELk���IMpϪf�~*s��z_{��q�0X臠pi,�~�B�T����.�<���c�zb����Ey��hO_��+'^��و,�v�����{��^�9�z��D���癄��MCDBӜ�׾�qN��6�����[��䚆0��(ooC��$U�]��E�2�I��L��M���~������iNU�e��4�C2a�[�00246	���Ȅe�*+5�&�W1�P��t^��US�K|<(D�gw�BPN�R�����'�N5N[����A��S�%N��Ӽf� ,�O%C�d}`�1j/6���x9��T�@���ۈ/~~;���7�?(�2H�rcv O"�f�/�k��"�\�t�X��@��e��d�9�g���.������@���%��i\ww�-�EAMu��1	�8���xT)�/,!B�w2kh��C�h)�7�8]��w��%��|'L�3jp�l��A{AL%|����6������Cܳ��뱝jb��"��z4Z~GZc��^�_�9����O0~o�1������e6[Ÿ

^�ֲim�
��tA�އ<�Ѕ�[����ه-�T�����,��Bfg���_*p�7��{�hX<�ve�Q��R�`q��ͯ#�]G���C߭����<beW�)���O��]D��_���t�<�/�\]�禍�kg�w]E��3��VBZ'�-A���<&�'�k+ޟ���\��4�uqZK�ћn&��@��iY������u�l��dqH�_7��L��G.������-�M�U+I�{���|Uй;&�CS���U�o�6~�Գz���⺚n;e�X��� MQw���2���8p��|M��� �8�>I~��p���+ÝuY$Z$��K\����ͅo��u�Ո�Z��4�&y(��R��@'�4өJ���DXjd��A/a��������)�;���.�O�M�#�.���%Z���.}���"qRN"�ƈ>3�h�X&,�}wiM~�L�Q�n�j?Z)Bʽ��d�3��V�:\'�e؇���*]����� �s�ؾE7�ӳ׈��E�R��?��9*�9�H��{���l��F�>es����U�W�T0��>Ti?�"�G�k�Cig3��u.�~�sȐ��A�z��-�x����z��X%�y�CX�h���$'!ڧo���I-�I����Ϩ��:<OF�P�����=eu���X��U�Wq�K�����J�s��S�C0}4��Z*p"G�a��gD�Ƨ���.#�7����D�#�����'m_�Ze�+ޜI(�ʁ`7����.*��"դ�Fju�4uTX��}إ���1�q�}���LXG�*���������#��E�[SG�	�B�&�`nL�3�Ԗ�lV���%J��q���3a�^�g� �<�꽧�h�sm���tm���w�9jBĆ=�a�d���3Qf�����Ph����n�\��,������WvusS�� cb�lI�ધ���#��G��O��˼TВ����#�u�h�E0�L��g��� QV��H��z6�!�YCGv��آTu6�@�n*?y�i���f��z��;�A� Mn/��BɊ#7!�t��=�5�H�aٰ�Xx��M��Pv����J�޼�;%n!���;�i-�p]���ߞ_.�6U���Jޥ����S�W Op�Q�w�w���${��C5ۏ9S�"��O�������2��oT�\�nF^�%�3��@=k)8r�2�u0�1�g�m����t��B���;���J^�f��kH��0�U+�sD'=�W������p�gW"��0�C�ADN�&��Ex ��6/[���&�z\�����PQ8
�b*v�]Y���%Wz��-�ʦ�Kx����(��Ev=���7��D'N"�E}��o�g�����U`O0�UR"sƽ�¯�5��).5�2X�%���4�x���S�6 �l&n�l���q����8�d�S%�2�e��NR%Q� م��C�]�ʨ�������ѱÐ��K$ <{We�ؐi�wۅ�^���є0����Q�G�%�e�g�9Z�FcÝ��r��<H�UQ���{�~���h���[�f��UD�!y�2�u�ė�孅+:_�G�a�`UѠ����⠩����]�:�(��h�^c��H0F��̲��p�՜Ty�D�5��͇w�&O����E���$�'�25��[�=a-��n��x�k�]u�t�}��R�u�+���y@y�o�z4^L�)�N�"�.��B��0g ?�����zi#�R��C���>�YoLv;!u�2�b������:9��)������"�U�<��K+���0�Xc5�'�c�s��W��{)0-7�aqc�e�f�0���Ze�-������M�dٲ�8�#�Bծ�!���c|P��İ*���9J�z��[���6�q�
�-���;�"�W^0K�(n�ᤙ0P�St�D���n��h Uݽ��<8�#����"�2�6O�M_��NCc �SӁ���?Cr�_�	��ҷ�O8�P�u�h���&����]e�d��F���vL�%��l�2��H��ت��\C�b�N�9<������s��=l��C��o�	�q�W�@;RmQ��������
��\��W�$���6&���5q�O,J<�b7!��Q�:��_�rOS��"�$k M��l�:���q4�g�<���ÑLw��-tv������o�m �|.��P�m|���72Q RF��_�+f�����Q�kz��^)�ъw�z��05k�\j�=.9�r��ف�QT� ��.��"�)V=l�8�E�γ�N�H��luFK5#�6Z�O�;3[�"�
M!�� �>�U�г$egl-�
�b���	���{����տFa�쀸|�)�cuz�� %&+F�-4
��֐(�}L�Ç7`6E�7lK�[��-*`(�)���9s��?�/ΈQ`4���խ!�@�V4�����NL~z��j�a�}c%�U�!�5���Β	3 ��?�h�b[W���UB�%-�w$r��J�fT7Y����Z�C_ϩO��4e�]�b.����"�_5ttdwN����*7�Q�[/�Vk%��t��B�pW�v�u؂���n�ouAl�Ne�Ԣ*D�?��|�ֵ��d2]�z�&��X��f��X7GnhQi~����n����˧��jx�����"^N���9T'U������4��yI�����|ʟ����(��~�U�C��s��'���e��n��Zsx����xj��|9G��Ͱ�zwHz�v2�*g_����'�4&
�@�8k�St�i����D�*�'u��ED�����N%��������"<����Y���\Y��K/�����b�RA�16����cb�ifB;$
y��3���)��=�����y[)��?�����;�-~���K,б����Kۧ�N1y��[���}\�� =�TD"X)� :xQ����I�c��ZH�#l-�z�%(�����/�f���fC�E�bgU:��ĨܩL�t�8�u��~Z����猢�?��l<�h��Xy!fb�Y1�yb��L���m�TF�9ƃȫa����2iW����QT-�"tz���}�3K�>/K�oo��t�M9�
�ir`�rHV���h��d-rU���+�����IHT�4[�	V�����O��,w���::�5�<Ĭ��QRc�(i�I����.�e��d?/��;[W��L��a=M}93j�����y+��B mB�L��X���Ʒ�{�W������"�)��e�A#�-��U�]��w�)*O�g�QC���6�|��~��퉨�8IH�H�3���?Rc��*˿�"x��n���-�Qm	�R��X�us����i;=����v�a\B}$| D��9��έF;�+�����-�%$Z�a8�>�
~�~<�GL��;*�`�wl~���[�G�â*�tR� 9�	�Pk
z�>	�a�,i�B��6^�i���H#�\RT	p��O��1�Ƃ��1�Q�#�����o�nOX�<<�皅VŶ�`��}��^ɀ64u�$���$��Te��f4�C c���e�(�|���N�/�D�_ا�Z��
�ҽ����%_�CW�K�QFi�ԋ��n4Ȣ%�Wh�/����Jx�QM��u�N0E����ze�����tT?��J�}sR3fm�ŤeJUd��x��M|_��E��L�k��l4w.O8�qY�%�G(���ύ\�;3X�25�y��
��
���&YZ2y���<k�G�����&�(Kʝv���%÷k�(�Z����bFW�K�t��KGӋ�+N+y
2*����~h��f�0ľ����s
)�����;��D,����ͦ7��7�yQ�qs$SW�=Y>�U4��D��0"E)�����;�K���y�F�C_V.����ԏГb�S[U��d׍m�^�ЖX�lFi����ip
wE��W�ug�ZK �ќZG*�<m��}5�ؕ ��zŔ�*Z*�6m�ϴ-p�}�ά�
>�`���J���5VP�ٯdE��&p��l;��Ȟ:��»�=G�dI��)���B �t���4y��4Y�v=�a��"�6z^-�����d� c%�Z�+2;LA�a&�����$޸-��ѿ��˥�ݙ�|H���u�$�<H�:}BȩTkV%�m(����M�����	?��ґK����~�G{Ã�F��n-�7ny�b��.�&�=)���If���D����*m��K��֜��*���-�u�5b3"��$��	���0�XW�zU|��`��@'�����X���H)Ӑ�Oc�'�;������r��:�`��/ d#��ΛJ �C�2O�u�e��L0���BE}aq"�~1��Һ�����=�;��s�I h�%���W`���a�#��+֐C^CvXɫ����6W��Hּ��ȎJ��.��Ag����UU���F4��ͭ�waƹ�XYגby;hIux�mY���
�\]�䌕T���;ܷ�>;.�l������]�&�����"�b���Ej3�J�YY�t!GË�#�S9	���^��5Q��5o�ɱ��SG�l����㛍�I�H������$�\���}���h#N�6i���*�Y ��W�\�
.��T��G��u]��Ԁ�-:�9�]��y��P_���֯�7F
��g�[1�E�-�+gk�����g�,�^�rǖ��*�aC�
�xXxx��#(U3l:�H��	�͡Pf�:K���U,��p';؏�<����W�,����h�$��L�J�ӻ��D	�0�A�䜥�Ҿ���fe5W�J���˱^�=z̃��l���ɭ�������<��
;,��� �B��}�14^�\+Oan�"	���=&p藜܋`16_b;٬e�"�ݓ��-�U-��E�ސD��WSHF�2?nÒK��2H�J��wQ��Ύ��!6��*�L%7.�Zl�h�xsQl�\�A�X�<C*�+�$���3)�)��rk�
��v�
��+>�6����QP�I��{0XeR���LA$�"�D�&�9�$U��OA�^��(QK^zWDu���ʾtVu��d�4��*���9r�l뛵��*�.�~s͕��Y����=�����2W$���͂�{�]�̕�)��L���5��w"A���&�H�^�)���CHeGͪMLtfj����@y?�$)Ϋ��1�Э��51�>��M&�y?DL<��蔋��v߃�쿹��(A�f6��4�w/��J�_K"܅�A'>�� v\�����R�N�Z�]�H��4M���RX���h(gP�O�7hւ��v6�$����K�ml{}�K��kD!cm��
��E�I�%�:��^�l�#�m_&�Fa�v��~��}�䨔pt6�Jp�@u�'C�j���d;���e�����v67�#-?��:�%Ժ�6������1o��P��T�{�Е$$���hV�Y��	U-l�Ekr��;�lrN�a����!��8�-�t�(�µG�'0�L/����4ȕ.�-��2Ef��#W��~ 7c���<���:�F����0��Z34�c(>u�4��X��-^�F� ���(d!�i1�4��-wH.�<�Q�H�7q���1�h`̍���?��Z��y�E�������;��1�������"�O����3�����^���q�ϭ� W���Np�`�����V�"�9���c�_n���V?��l2������-�Fz �D��(�&��!�����3)/VV��u�C��\Wvo�<q	���Q)�cb���g%X"������Y�
�}ɔ�a���ծ0r	�E-k���jƠ�P�1_14�]���߮���5 ��>�ʟ�j���:����\(xm���u�0��S�wzvavS��&��]�S	߂A���7�3j`.���F���wY�9`����`�^#����Q�"i��|/w��>�^B��b$�U�ݑ��]��,�s/TO-���
u�g�w�Uй8�B���Ż���^�k���`󚖒�T#��3}Q�k�V�ƚ�ni-K�F����
Wo
h���󭘸'/��A�p:�B{t<x�m�O.�+�j�'�%�OU	�v^�uk�s$�w�չ���F"j�"����=C�7��n�IE	��D�KI���Q^����V]x[5��'eDߡ��Y�J6�x{�����7�>����#�^
��WJ*�u��	�WO,ʦ(�}��$)U56e��n�k��T�4�O���윱�R �8�*����t�P!KI�"]���9<�I�d>���'��p/��32��|�^c�D���2�B|
)�Gc�j�S�����i�ƞ]��}��&�)]��]�rG��&��O�22M+��S���ͱ����%��2�Z��H�gh���K�{t'���лwL�_%����G��aA�e �bt� 憪���:�$SM��v����i�F��sG� ��h�ӧ)GU_5b�c�?�؃+�ػ�JԵL�t�g�ؽj�L�+���-Ԛ|7T��I�뗇�4�_lXH��[}kȄ��`>ҵ�~Ӕ�me"�^}�΢N�"4Ӳ����eLz����2ӟEΐu;08�ï���~��z�G��C#�A�~���;�����O�#����3��xۋ�)c��5n�;��	�Mc�sP-��l=Y�������������X���|�a��Ș���T6b�� y��{��uܮ^�n$-+^�b5���K$������ژ ��t�\��H�L�a95	ТC��rh5����yMy���f��Yٙ_�u]��7f0�P�Ȩ���S�Ff�����o����D�t֑؍���I�e���*`o�D�'��AX��I�_����V�qD}k�)>4��ۣ�)t05�"�^	<��m��$)	�MF�*�&�u�A�?Om�VX�)v�<�F���*��U:����G�ݎż�[R�<�@pu����{�O�}T���h�՗��g�P#c�ϖ��Q�
@��0������2"1E�}�yN{U�P���#�3}1]��zƿ��Z�B�.�ߏ��,�Z�e�%,��n�#h.���@b��ܽ�zBb]$\"�:=|�~S�=��ae�S��/b�:�aH�v��asX��;D���)ɷ��(la�IhJ�V�}&_��Wʒ��.����ѣ{8�!�q�L�"lVu���<Иi�P;k]	�Uқpd�o��k�wqQ�a�G;���a��Ư�Y��p��Sh����32`��3 7~VR�����@ ��0��Gޢ�:�[��
y�q2J�emܒc�^��l��3ȚJ"��_J����tC'�w՞[7���K���T����g2��-0�"򣭌+�i(3�H�y�&t�W(��,r��g��\���Y_�x�{���j��FI����V����.��ֺl�gΝ��ѵv��0)"L�Tw���F'S�8�W�g˞��P��;�����������4�q�������Gu ��)Bp��æ���Ey{.�<=f�+ݕ9���4 ����_��ٚ��Mf�.����\�L�.l��ڌ�!zH{P��ځ��Pʃ��6�J=pTd�7s�g�A�E�������L���Ɗ������s��!���)��ν��؜��i����:X(�����ct�n�*�15\�#.=�b��m�0�05?l6rѡ����f�S�ѐ��Q�/�/����D�WC����C{t�����YQ��˙�1N�t"�	�j~7��!`hV��W:����s��\�{*,���;����)����)rvDÐB"��;����cմo���&�T�H�T��*���
|�6��Ի�
����e`ܵ�,���rO�Ӻ5��:)��a���c�\���R��r�b����#��{)�������9�9Oӝ? b���p�����6T�Q�hѵOm��p_e+\��_%7�)W��Փv+'�.)����&B�\�NB8�W1����+��y�>x9��D&�Й&��9e��􁮝�P&���+̆ފ��ێE�UGk���.���X�z�R�z��%��(�.��7��k>�cӵp,��%2�R������[4�!C�����U03��?���<d�l�tXy���S=(�Z�d�p�1CT�T����H}of�3�2��m=fu{�/).-o�J���yk���o�CH��v���$�<R�#�W~ˑL���#<t�
H����?h��"�=� �~~>#i�LX`Z�� �e�}΁I�ס��j�����uC�N���p�k����v�YS~-j����l�.���E#��z�Uر�n�a�I��HG.0|8���0H����dsà!���,	�Օ~�"����?f�|�ZA⥨�˔����v	g�B������Ox����jP�3�4���!���L/{2k���f���i�Ϫ�,����[��j\�G�ђAY��"�������FR�&̛y=��qm�ZY|h�w���w�U�t��y'7Yn:<�#�����Z��\�"c��m9L[��b�;lM��
�m-���e���n��p�LU뇤�΅�R����	�_N��ƿ��;��Û��Eh9�V@n]I�c�,��N�NV�s)%mA�W������=	�˫�i`�S�ߨl�`f�Z(���Ft��>[�ؽ��{���S�&�;�J��9���'�c��T��׋���K���s�y)����V�6KE=̖���D�W��F.R$�s^Za#t߭�M|��,�Ș��_p����{Rm�n��B������0LI$,P9�Yt~��ZKʷ�ٸ��g��ޔ�۩�-�
������A3���g;F�<t0Z6d@��n`1�oXWoS���,Y|���(?A��c���U��t=
��O���J+jKZxc����>3�?�Ze�s�5z�O�	6}Ei%ț��e�>:1yg ��gۈ��$O��A%B�d����TCX�U�7��Z�ځ�W�4�:�`�V��]�Yw%P�v;Gv�����p�I�ji����I�2d��l@�m���3&)�D}���>%��Nt�G��*�Ǿ 9��o:�T* [n�+h�����2'����:^rN8G��U�Đ��NO�sϚj�.�x���`���5���)*!��aZ\*�F��(��y)��4H>�_yr���L�C>f(���v��%)�ѹyG+��ovs�X劀�dC�@P���
��������tT����%��ϲ��>��ZǬ�1����i6��Ӷ�����"A��� 3�gX]<�7�a
�輸����$?��<�8Q>�}�31��%3��wR젶�&ex�	\�O��n([1�a��v�.��e�J���ٛT�ר�aR����;X#1�P	�T����T�ED��g�iA/���eq�y y�(��f�D'IuU:R��qy���9�lr�P����k��H��`:� d���$";��l� �x���"�B�ݸ536EP�qv��{m��gΩ��*��ޭ*ϐ5��*!#ƵM�K��@ԳVUk��3�~�Q�n�	 e�c6��#=�_g���e��߄r�0W�PT����ڮ=�6�b�g��� 3�5ɻW)�ea�j~%7Me� ���1 B'S�^�z�^q���&o�r��q�G�Z��mk����;d:�ok&�B[��.1�t���w��'[}�-�4��J+vj9F��I8�ܯu���R,��LC[n���?`=˻�\�5�:<o�k��R�Tz.sf#��~Q�dS�j-�.9W4���H��U��:�[	��Rc�d�Y'�5AzNB��n� �ҭşP�G&~q�:�qd���.{�t�+{��A,DU�?ֽ����o3�:"O�l���J��+�XY���-��me!:}��1�_�Ykosr=z���mf0DhN(T��Aŭ����y���#����KR�$$c;� �Xo��i�Ǘ!���ᛆ�mR�8���S�53_1:��wj灧��pI^�`��S4��3������G�v���|��_��ϊ��9A�ɑ�S�2���:G`�-�����r�
�.B���w�,:�sRA��#�/�z���P�2��+�8k6P�$_V���p�$-uǪ�J�[~:ſ�f< t?�x��G���yY�j��xi���z�8�T\1:>�\��e�Zӿ?F�L4���XPv������I��I� ]<���vΗrŸs��>��o���,��@NAW���
�z7kڲ\�*��_��dߒ����Xƨ�M�����ï=/���W�U����y��M�tN���ǖ���5ɇ�F����K�-l��d�0�h&�D�u`�:^��~�-d�!&o�����/ ��u���JBH��,����_y��=N.&{���X�� }x= ����6�Sn�@ۿ+7�j�e�8���,���Ϲl�?�0�f[~.+;�CVh޿^�uR�O��!�����k�����&B�����̍e4=^-�������D�)��
XX�k&��L�h����ʑtQ�}V�ә�HR����c�����@a���{Ln�2%�KӕV7D&�R��t-�x7D��߼*U7��M�n�`�	o��#��kA���܏��0�W���a'Q��;����'�ݞH��vdC������5�w���ʎ6��*~�j�샆���h�4h���-�Y��B���Ir��L}f���I���D�_�k� ��9�j1����t<b���5e^p�hh�L�>0_���#u&���k��{u����&�'�M�_�T����G�(�2�V�e<���=�ۛ����~��h��i;E)�� ��m�юPp���_\�j2��Gs�A-�����Z|�$	8A��'X����]R{���D��M�-�J&g@H���oX/��+���R>�0����nqzUb=��H����3��dZ�|��F�)�����I�T<��x���<HP������%���В̅f,X�=_��£�j�	\�,� Y��מ)�ܞ3�"Oŵ<���Hg� �&�?�eD���(���E�qK{�R�ԭu��]�9��n+x���C*��˻���Y�5S岳�@!C^E+bmѠ�J��l&�H:��Z��5�r��La���?.m��$]pS����� �њkϯx�1��� �?VFZO���;}Y�n�u���E�8���p-v��%�Kn!h5jmO�����⡧*b��&���#�����UT�"����e�:Mwx���L��DK�$�3�&$�c+ɱ�G$#`����n��фWE�N�@ݒ|'A��u'x1s;��8�FL�x�BR������{kCL vk��#���uЕA��30Wh�eü�I�@�Z	@:L�ԡ�гg�#�W��ߊ�n��7�\e��ȼ��j�;/7.#jp��%�!w��7T�Y"�b���CeI>�4S�����u�E$���iK�}����==e0����g��KV��������-�eA��k�NYR��1�Q�T�D��5�+�v��)ƒ���&���{���T9/bߥ�_w�Y��5X �}g+[X���޽��E�����TG��%�(:ɥ�	�DZe�ы����h]S)Wj!㶱P��/fqS��?z��%�sܠ/i�Z ɅH� �5����i�n�C��s:�ɛ�?
)�$Hn�-���ٻl��?}������Z4^����@�dY(��0��o�/�4 Ұb���W�~��$l��M&؃cӥ����#���~��6�۫:z��6�ZŸ�K��q./���b"�˒;6G�ņ��/Pa_�ЃZ	�p��"�>0���z���ģ`��-�~9�:��Q��<"�=幯i:���H_�q/(�AV۰
9e
��Y���K\�*g����1��|�Z�_lQ�	�l��TT1�%����*T��'��[��������z1/^sV �m����/K�=�+�� �ѧ�]^o~P��:��0,���Um`���v����4�<��(��s[6{��0h�Tn�7%۩&֍������YW O��YĞz$���f�,I�s%�|ۄs��澬O� }Ǎ�0�K��|+�D�0���ε!�xi�"�,���kR-}��ޮ_*�����rվ��z������������2�y��w��H;�/�b�|)�]�|�?�6#:��+I���{�$��%17��o&`�;'�"FA������S�uu�k�~�{����K�TMp�k N�x�M%m�b_����F6U�^�2��gYl�����|a�[���ے����tG��L}�WX�&��h{�T5��kR>�z�`:��}$�Yj(�f��Oq���3'w����1��%�n�h�����C
�X��?B@����{�4f� 9 ��}��G�!�$� Eh��q�|��ܯ�美��)����]
-3����y�s;V�4:�����kAlc!@KQ\Y��
�i�X�}���k��/�Ͳ%ɽ�>���W��NQ�.��]S�<�aHd i��PL5H%��>���`Y���;($9\x��o�X���f��`�j�� �m�E�x�f�퐌�|��i:�e�a��]��sN�rd�zrݺنG)�)�˩;�F�BOGڔ�O����2�ؾ\ߙO����`k�� �W���k���#�V�xb)9~X�D�`q�a�܅e&.W����k������(qiocg���ݧ��V-��1�3mz��7B�76�lҳ|� qt���ո�'q&���ȹ9�38ν$�1];��Z�V�n�SbЛ
�H�(��`��)�B6��t�F�K���\AЗ�RD����n��/B�!��0f�Z�?)6�=�eu�K7
,�n�v��w�cBgA*���\�4b��{,Hr��X��� 2�e���Q!V�+Y��OįH� �P�|s+t�݆G}�@�n4��u��պכ�W�~z�`�P��OS2H��)v�oӃC��˱r�+#��wc{������M�W͘"	�d��A��.f�V� �:|9D�0���F�5�O3߅>�}���U�m�Z����t�Im6��\2��=������9N�xY��o��W&+j{5c��u���7Z��;���xp�Q�~9��ɗ}�f40�Ƣ T�����TK���;��{���p��w@&�=`�ށfƪ�R������^3J��w���.�HObҌt���� �3��[e�/Ь�ht�/ 0���B��ε^,Tl�ҬG�4�'8}��bwL����oM�9;
hپ*��$Y�p-Q
�V��D�#�;�cR��o�Rі�r��@��H�3�|]9}2M[<E��ӕ����{�S��_6a��ww�[Z��E�$���>%��RA�]�����0�@t��
"���2�G�Dm�c�|���h�r�:{Lφ@��L:D�6�<��I1���%mP�Q<0�)��Nq�ή;<�&߸�z�q)���,��Q��\�Y��$�Kf��⯇ y_{�Ǆ�M�x��v��O���gI���F�6ồ[b�⥞<w{�+l�}Gf<�SQL�`6mNh_���j/�,n�pl�͝��	Qܔ�ۿ�����t�M����]�^N��,�_�����WKG�V����٢}�ޙQ����Irvy���N^��BnS�FT�kGt\^bm<1�Ab�n�B������0�gD�ӡ�|�3��֬���R��I�}>�}�D0���%b�w�+a3�G�!�D,|� �iA.�Y���~sMA����ݸ
:�t����7��R�_ȱ���_7�v�l ��'מ�d%b�A��������-�ۭ��N�Хr �Ȩ2�# (٭26�=�^��H�z�%3̖����Ze����ro;"�s��pS��D���A����?�m��q[�j_���T��r~L�K���G�G6�S}i�y]|�`�	m4g(5�*'$�v� #�������� W���x\�4�
g5���߭IP�5��Ub*�$���u�F#^��?�j�a?��֛�ORM&6�WgZ���Xcf��!�]�Ӑ0�`߰����v\�4�0������u�ۗ�Z,4u��{��n<�0K�eل|����E��O����	_9����?��O�kD�K�%�%���e�Eu4����L.���~�~�A�!��bi|*P8B�]ī�Q�O�0�_��L=������tȀY�bu(L^����P9dH�O���'3l ����;�X�/[/\��#%O5+nz%���I�c_?��>���MD�k#��U��0Q����-�~o
�4Ҳ��`Kn�Ǻc��."�Zmti(D7)$ı-�e���A���Ӷ�m����=:�}/�����l�3�ŭ�7_rUj��dE���*RƑ�������"m�g>��:��y����t,��>]̈́��dk~Ro�OW7J㫅��J�>�.�<��Թq� 9$��v#�T����v�����99X��$F�=��)�o�|�%������O�g���I,�r�Ϩ�.�)`m~���V<�i�]f~r�a ì|���l���e�e�m4*c;��4C�.'�3��:�۾V�nٷʉ���}�Kߠ7zq�@�"	�ֱ&P�e�ꯂ1|���8��a	�fù���1�b�B�]���A���!�H�L����|�cC�Nl>�axh\�2pl��NC�$��Et������[B1Q�:m$`�.f5�}֓g��b�ٞawoؤ=sw�x]aX��u�Ӟ5}v�ݾ�4 �u2A��uN�F�8�f8����������؜M��&�!�X3�w_E߲\6���=!�Bg�ε�����f��V�/���pے5����L�客�Vq�=�7v�^�����������o,[
ͱ���Q�ځ�Pz"��y��c��t�C:_������jW�YI?���VRd�D�kvF����o�SU��� i��6{�Q��]�3�j�_�4�4$3����"�H�x�mgbY����)�	&������x={�;��.،��2�6����N��Ȕa�g�>�x�m�����@f��8�&^��^r��a�1�Z։OH�& o�
M4[4�suȭ�sf��!�ДfvP�3B��!�"������}!���c��@���2��(#]4�����@���I��s�)0c��Q���
.k_�����S*Q�\������*jԚ�*y��<{-�lx?� Z'ٖ���a}����K~��z�"���A�0������(q���ҍ-�d�DI�/���D�{�|���r�t�f��Q2�;Y.X��&SA ��u��eU[?��t`!6�j��Ǟ�A8�Û��'�"������䃚u�o�d2h����O�����r[��J��<u/���yT"�s�JL�K	ұ�E�L� �

99��F�Z�˿��5�X����,�H��0HT�1+��$��3����s�C�3��q�#"��~+C=ua�(%%J"?�:�Þ.����X��ڨɴZ�N��^G��XWdj���V�[x�'�'R ������{˭%��U�_�$���q	 ����17�M�+�>3D���ؒw(�ϳ=WH���á�@��GQƸ>��b����W͜#{�1^�Ȝ~�f�8LJ�J�SRI��1��a��K�+	H?r�1
��پ�Tt}�/H��A�7X,��c�hQ��fsU4! UQ�AI!&�#%)(�V��h_�1ލ�z��:����������r��_�q�D�k ����x�t���%*�Se�����\~�[@���%?��o�5Q�/j�6�2b{QEG0^�N��|�Y�ͯ�:��"�P$ Nʦ��h��+}�
[dd�{��w�B�%�?�HYW�te§l��w�5E�N������F��H^
�81�,sŸ�HgS���U@rd�6�v�7�}7��0LV'�3U�q���2���	�)n����.t��86��U����)KP�X�c~P>~e�V6�3k�Z��O����h��tY���?��X0����XYj$���&������-Tw��m�������)΁]jV*��c"(�SԵ̀4׊�X�62A�d3�rj-Jq�/o�x�j��xsKc�1Cu�3���y�U{�h�o^��i��}vmco�+&�j�tC� �~+�4���_��r��T��j�(ez6߅�D֕�A*����#����/�w~g,���4i{��x���	aYx��ђ��8�_A6߅�q^6
������Q[�ͬC0:S��P�r��p��qz'H���Ci�J�Yf�"��;���n�o������� �AP�WSQ��	��_ݑ.g��?Uy�/���R�;MCZyD�����(�����#���
��<|��w^�UN#����
�m/��� �86�
�~�� �Z��2�]��2�%!��S�C�j���H�vA�+h@�mlrO>����8']M�w�ub��������kbvә��n5q���oTS��Djh\�79� �'����f��$��Ogѩ"��i$!N=p(W4w^݅��,5g
�*��s�-���t#ߔ�ܧ����yC���:���S����tS ���9�G{��(��KP`����8�T�p�=�-���xذ:��ò	UYng7�~�[�u�:����E�!j��>��z!��hJҽ�F�G���Y��b2~�"X���ϫ �j|�v�!~�{��U�*�_&�1�j�����hj��B���tq	bA s2�9E��y^蓹e/Zq��$�O|lU����S��]�k�.����h&8���"�l2��-�D�$��o5S.�6pxc����4Lg�}0��!�����>�Q+��)��8 �ZNu����au~qb�CND��R�Z�Eƪl/k���
#p8&f^r
����o�j�F�(�����kY
7T���R�s;��>����jT3&�U�4�?؃�@�ӭ��y�S^S�#�Eۥ� ���j��9������c�B2���@2!�>�sŃ���G,�d��R�V��*K�H�{���}�rrU����;HK���S5��'1��m���Ј�(��60�'�}�׵.������� 2�� D4��5���0%K�6L	4�O&J���צE5e�"�]R�}<�t|�.��m�s��'�ݯ��"��so�$�#�`�hЦ!�a�Ťda��6�C���雌#��H��0u6"a�����Q�@�\8�C�����9��g�RD��9U�>�K�Ybcp+�g[(�f-A����%���_���-��<x���r3��:�+K	�����f)Z�N(M�����{Ҿ�W��84��P�N�^��f�=u�Ñ@��g
mɀ-�{�p�A;�q��v�ݜOX?:\��B�mh":�1.���P�.�/�:��<g����G��ޔ5���������J2A��v�w��\�V6R����=�b��C��h�ק"��*$�� � ��{#R@�Pq�����ɯ����'0��S��ŀ�$ �clIR���V5�����gt��h�r��`�n�'u	�ӈg�:���O�ڬI�`�qwXw@��h�{*���uE�u<^��F��r�o#���E�7�|���)>H�ȿzZ2f���&�v�Pw��"��]�G`�5F���/�u\�(ȇO��"�1:�<���Q-�N��8�)�aߟ���RΘa(i&ރ "m�yALz+����'�Ҋ��2�W��<ڂ-��PE�D�a���_2a찃щcK��ا�񦣴E|������P���hR��H��KY�)c��`�(�m ����B�;!a�ѭz"NR�Q �3)ͤ]wDS���^.�R�.S1B�]^X0�^�(��v�!�H�g��|�`�ѻ�J�EWU���E-}_��+\�y c�
��މ��)<��^�M�D\��7��OT�Ɏ˸,�����A7/[>�G�' i��s�{i�)�LM�[	lGd?�0����1̸ve󿰩k&�j%��ɲ�h,�K��4e�������ќ�a?u���b��W�%�)J:�X!��qf�C��T�J�3�+V%�>�	������1n3VWb��	�@�j�m��$0����z��H�� 2=7L��ܥ�ʠ�L�J��ޢ��a�o��զ���B+֔H�9@/bN�"\��hF�<F��"�w���e�4f6!M�oh+f��⿲ϓ���@x	���c>s-9��ٴ������yrB{z�3Zu~��6��1o�E!aĪK�>y���e����P�2����n�.䖺%�1��W�()9ܡ�)���7�z��%���P��g�����L��뒄R<SN���cP�����	�r�`eL91�Z^�������8.����㚒 f6��N�F�K���
�s��	TV����P��B$�qܕ��6B�M{���H?���h��(-�2�~X�jհ�Y?��-�W�|AgNʏg�k���	�E�n)ݱ���b���[`x�8����ۻ䞹�۫A�?�+�;��+LsM��`w,}�f�M��;�[/�d�!�G��i�΂�`�ЬF�n�'L��&�W���y�7ݛ�ngF��F�_����GDu�«%�2:�T�雩���
V��y��(�~ucDza�3)/��2�p�yɝ˱�*]��E{[�SX��� ��a���q�H߅�x�LV&�r��Ɇ���s;��
_o�mg�w$��Jjp
�xQBS�������ǔ��Sl"X���jTC<�;�y0���Vh�7eo�}מ�}�=��Ŋ�!0b���3�^�db�Wv�^!����H��oho=ۼ&qcM�-Y�-�ƒ�Ѐ]wzE���JnZ:ƐG��G����; Y)���&�2����C:�9Iﱳ �
c���!��:n���0x�:�q
`��/���Y�i"�Ϟ��a�+��/�(|�,�hIǷ���w}�P({Q��Cb��ey���E���ӗ^\�t�D��>l�O&��I��������/�X�[�"�d��S��N�g�tҩ��=�MP��^�Y��ʖ@G�mM����e�ʠ�&�}և����]�T�zLp�qւy����K�A鋪�mŐ���ES������p��籠	���~]Z�㒛����T�|�s��0�+�>ү���Źo(��-zH�*�ť��(�+��1��tl�e�&��i�h�(�������N>�ƙ��4����5Q5_�b��� �T�����:$H��8g*X<�b��kR~��eҙ�G}�JA}㺠F����N���낪�GY
��Z����%s���:�p���N�S�;��X}œ��X�8�:�^ߝİH\��$He���TŜhN��IJ�n(��Ò�%t���o�r���O�2�K��.��95�6^�Ml���"J qF���H��Z���}�z(�I:���3Ú�vA�b��D�劉[�yٚ�1#<em�h�3ݺ��Z��
3{�������vK�?�X�_�F?n�/W!^?qQ0��x�J�o)�-^Ǯ�,v`)/q_u���]A{2�q��uaڃ��5�W�"Ke
�%�;��R� � $5�F�S-�I����?��+�L^�ou��Ӏq�1o�䥇o�� �s|���vF�{섰4�4Yô�0��?wP(p��6�]T�^�pG�F�pn(��U�me�g�쟭]ɿFg(���\��ʘ�u�Q�$�@�*U�Ŗ��հAqYᖉ) ŀd��|������(�������<�� b�N�kt�Pj=�ƻud��g	����t�/_?��<;5���`k�PѱN8�q��\!��*E�ӂ��S�S���#6N�~!�+��lFbtD�-�+ȊR�� �$���^\0cVL���-��	t0;���.����I��()\�*P��~�7�����������>�̗���g n�5�7U��r�D�������-�։}4�DHC��*����T�{~^��1������� �/���J�D6�PÇ����8���$H��<��t���
7������f�i�'�}��|(?��'M.� ���+����<���:��N%a�E����i1)�w��,}l�i���C���Ͷ����?����o�j�m��_f�����RAd������fTs�R��"Q+��(y�