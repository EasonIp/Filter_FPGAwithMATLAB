��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5dδ���KdXyݕ�2�j����B�}��AlU=w��m�C�}�S�[U ���c��6��u�������K���ֵZ$�<���?�ޒO 	��ȿk�Ƽ�o���n� �����4D�������;����l�{6d�0
�Z�^�^�2�;�D�
�UjR!�1�2>��Lb�`�D�l�W�?��9�J�ס�Y�u�kK$�ɓ�#�NA��Y�o�~8g�!'Q�Qd���1��+j�i��|Dσ:���x4����j���g��6��� n�벙s���c� v�f�GMcˎ�����0���6�R��$́r���E�^vq8g�O�jl\	��ч9ݢ���/�p-Zo;i�c�at��zb��M�պ@
�G{���CM��0Gm��w3���Q��ɛr�v�^7�<��cq��Z{ۙ��]l���gw��Eh��v|ۻ��&�xN�I��X�eъ�_�PB ��'%xRWh���e}��w��X�ə*J�Q7�j+#�1Q"���E/n3L�r�~��(>�,^�"O <r�b�?��cN2}�8��[�sA����+k2��\�8�YҐ	��~��@�D@�|��u	T�IU���|L��Ms���<��ˊ��U��F�5КkvП=5Ǩ���-�a���ow���I�@нr���\��.C��JxNV��IO�,�{�F�\��kR�[$t�c[��ܘ:^�� ߐ5��nV��m�H�p�m�:��y!o�k*y��P����P��U
���܂��BQ���,�O�/a������2B��1�f��oĜe7�拙���{� &���"�G1����E0Ja�>��񻺼�\�z�aA�=a��2Oq��VG��6�H���c�1��`^��uKr��Q�p�Fj>�ZJ.�~�:�4F�eV7�^�q��Md��E������,��wT�5l�}'�t��ȿ����+8�Y�ͩ�_Q�.b��	���Y�aG�>9Q��ǎw����(z�݅��o�{�a䵖��0��]�(X� ��������5�j@ �G�4�&.J(\�8�#!@��Mc���-����&�H-Ѫ�N�"MӦ���tqƊ�bP-V۷��x��÷oa�	����/����V��6t���p �-��;����П�}B�ؠ�s-� ���D�g4���ТϖhNc,�?"7m���<�+tj)�V>�5o��}Bl����0w*��ѹW�
'����1�Q�=3p���5�F�3Z��=ܐ`�j��|���U���&%�m���b*ɝ3Ŗv�V�
{Ӓ_G�Y�}i�۝5����}�W0�G0��>�7[����`�ƹԢ��̾�u�k�L 
��K�T�C˗Ċ��3��PJB���} y�i����c�݉��C�|}��C���$@�������X�M>}w����y0����绘��(�6	_t(|��*�a���
~;�^1;f�Ǧ���
h���{J�aq�|��Ԥ�Ġ���ò*��A$�3��t���SԞl�?��u=���E�?#nr�O�r`�x~�U�a�� ��I�}��U������� +���P�#�ǓȨ�Ƀ�A���y[��K��*������:X��v�_/N�㝏�o��C�Y��GZN@��=B7g#��D�Y1F���o�$�����o2>3�.fx�p�.��O)\�ʝ�r�Rt�X�]Y��U[p��.� o<$��V8�_G�VF�M��am."��s��Ўy�|�6;Ga���>[�]�fw+<[b�K<Q�W���>�ev�ɻl-�7h'G���'8�`(YB*�v>RX�y��0�mf��$����pg;Q6�V����-E���ޢx�6�X���t��@�(�9Ѵ)a.;n�_5��o�u�qA��z�,Ӂ��wɶ�\��R�r��Cl��;e�Z]�g5jP�e�[=�ע�#�:��a^�g����-�A$�Y�7!�X u�A�Y������^|̠�6�ȯƼ��kc.X-�����M�
k�\_[�-�_Z�vU%�-*Y"@cT�P���w�'�����J�sBE?
j{����Q�=o�ŲqtK֥�@8����߮Z�9�~�o��
���^�H��'�t���&��ﰩ]�)stÖ�ZVB��G����l�do-��FW|)@��Pۭ5���?K�y|�;`>'�Y�v�4)�:��0�&-�ڕ�a��9�-J�O}��"/�D�مD	i�pz�x!b�Q�QW4¯�Rua��cg������������m����'�()�pi��G�s��v�X�焞\
��+�\Xj�ܺ��c%�.e�������T�K��K�k(�c�*�~����Gu�.e5��9Ux�`�*�ʋ��β�/�$�m���n[A���򝫰�s@2��&OB%0AѱUU�HY�S7X���u��[=�b{_�dF��z���@�6�'�y�	/�kl���#c�.�P�X�r�'h��"��mRVЀ/)�gժ�a���6M�ρ )<;�yl"�H�Ŀa�ې����EVG��?�Xs��vc�4r�nE�ᚸ2��ڼk)���~����W���ʼIFCpC.�~d����#��-$�[Eb����tl�!X�>�������,��:Z�6-�������~]�H��̵�������a��-}E�~\v��fbpv���d�����ů�'
H�*8H�!<�蚓�ǈ2T�\��;O��p%@Et3�B�����R�^�R&���2;�Mٞ I���jt}���G���i��/]${�-4������r[�CX�L^�)�)�	�C�I��h�@+�Ҽ�s�꒷�q�"xEdX:��/��կ�`�v��V�B0 ",t%0WY¿F�R��1�8�qX̸��u�����v�ji�&����P²A+�V�<{���|[�ʉ>v� ��y�j�z͆1�6���/�|�0"p 6����I�M��V#�$t��҆2���X�F�`~:�iEl����Ƹ��8�����{�)�뙆�
v �-6��E����ī]S4R �A%Օ��0��F�-