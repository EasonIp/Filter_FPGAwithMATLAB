��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O �ٝ�l�������V��fE��v�-�Q��Rj&	ڭE�����<��1`5��o"�l�&��3J���m\�tu*&W�N[��H��j	�����[6ҊZq]ս"�!z���z��r5����nk�/�v����~��8r��,��:ƛ���M-$��e�~4=#�g�L�C�� \3˂��M�~���Wξ���G��Iǎ�S��IhU�_J]��;'M�J�ӕk�g��b��v��ҵ푣�~���/O�ׅ���08n2�B�
|Rh�ώX�T`;<�/y��m�=q;a�߸h�{���ð�t���f��
*tLb?�S
n�Uj�
�J ~���lAoT?�!d$��1�-;�59�C@YO*��x6S�����0��*�?��'d�>�fCŝ�ug��ENm�HKj���i�@�����&�F�kZ�8���E���b,>�#z��Ƭu?�_ͥ-�BH�k>�K
 ���AS���+�����>�E�c��?$�*rJ>&+a�#PS\�-����r�٭|�!��S����7�9���[|)���
�;>(i�>����Z;C��>��T���:1x��L;Utu�S׫E���.�ޒ12�Ꮠ���Z��|�*Wټ �iVr�+��<wzl����d:�:w�"����:Z
�Μ���IU���~�w�HJ��P����#�>����2��Ms��_�'����~J<!�
?V�9�o���bM��0��� �E��S��k�[�s�L�O��WX��-3B��O�
+ʮj��"O��P~���Q�_����~�����ؽ��̍ϲ�=��e��I�n1Rn�YDy|�/�\��v]A�>����M���z�v�s+�a/G��TB�w4xnРCҪd�����iV�sB�郡�1Z��������0~��,K��|(�{�| B��\
)����b`�j>j�O�
��6����|z5&~萤�h�����Gq�/�!�`�'仁"0�q3�X L ��+ ��_�-I�<��ܯ����F.G��C<NdĨoÝ��F*�T����PE��<r�5��^��E�Jd?@	I���/HRd�X� 7��z�t���M����d�
Ƴ�%���[v2�5�>��8�h�db�l�=����n�+��)tr�.��� �[��4C��Q#�jD����|9��1R�"��&�b3r��4i3Vc�WP����w���*�z���1�!�o���!�#�w5E$�۾�1��י�*ng������AF���L;e8_sq;jsx0U�����+�#�q �p�y�bS�M_���"���Y�������[�nU�����K�5��@e���N4`i]9�9 ���0i�S��aL��&�]w��޴�.��_K:T�Kk����4��2�AА�t6#�<'qIg���к�JM{K����!z�{pĨ�0A��걞��)XY6؍^Y��ZG�����9�sX��E i�PU�s.�1��D`F�zy��=����o������۬��hox�cV��3��+=�6��(R�{��ݱ�V�� 
=��?>x��#y�kSGS�ɜ��_�E5>����"����S�~0��Q�c6��?e��=����o~�Z��U�k�T��]�c�<��'�o#���7�Wq��������!|���8G��T�����TĦ�19v��8���3��f���+i�}��a�t���d�/�F>��al� <lhƒ?�Kw�a���b�W�f֡O�K[w�^V�,-��{r��j�3���u#A�c��
��`������.V��bP�q���#������	�4΋@�+�U��C��Jx��� "픳��S�&�X�ڽi�-���i��/��*�6i�z&2��2��)�����rul�(�f?:i�-�<D8���w��/�����zf&�h����8��<�ʶ� �R���o.Z�ϱ��X�9����xzQQ���w�޻#���:9F/Ѱ-f`��{�|8h]�y��!��P_���+GǍL���M����r:��E�G�N�������{\!���=�RD��8|�����rf�z���xW���QZh����O&?dS�.���&O�q�:���,`d�1�����O���A��!#��;Y�<����,ڦ-�?��VI�h^���B��>�*�:HAöD� �n�y��5��^�.�p;ۚ����7�'v�'Y���	ᕪjx�b*�`[�MŽ3z7ǫ�x!ʬr���K���֕��Ȗr��7`�b%�k¤3Dy�����;���3�YpM$�ނ~�GD�%����l�ҍ�nkH;vL��[ �X)���$��;Ҟߋt\�*�P�{*��!�NiCOnFT��#�t�=��u�؉��=z����7���
�g.I0S�f0xS'S#��Y<M��O�O�4:�F�6��f,�Ϧ�%��=ٹ�ʵ�b��>	�P'" ��H�[9=� (�n�rs�ȑ̤qf ��C�h��Y��Gg�0>zZ��b��`b��a�8���?A�u��F]��ZNwv<(��쐯
���fk�g73w.���J�V�An����5��7dp��)�;и`��dZ��]��Cp��6��Xa>}�B!$��	��.����_���PJ:y�l%���Ԗ 3�:ЅU;9�����)M��t!
� �鳚�ٛ޳Z0�ɀ���T{�u#�q�}���,��#m"��(`�����R��Y��pH��S���a{���9�,V
}+��ǁ=}���A�ؓ���ĩs�Xi�-�VL�!k�ּçE�&[/J_4��f�a 3xd�c����+r6��'o=����yc�H5�dT�	�����,+��:�R�T��ɫ�����^?T��>G���]��\�]����Ak
�؅������Xؕ\���2]�ǆ�ݟU�H��t8AV�Qu�
U�V��c�����P�S�@˚�p�槨R�����~q�s=�+2� 
��(�E����D�G�&�-�ԩ�b�����č��+yw��Q���pn�ϧ`W�`ŧ+�|*���\b���
�Yw�x�#�o��-��|�P�g�<���+Qh�Z#Sq���uh�ֈ腒@�&��y���r�a�/z�/��vH�	�̐�ϻ�?M��4S�O�󇊯儲��8����'n�V��8p5W��F����%��3I����񪫰���d��+'�Y���3@-OH�Ƙ��Lk���њR��-�S���b��� �e���6��|���F781n�u#�S�tW.ւ
�&0�����@�M*��Ǣ]"�싾��CWA�9�8V�oQ��{l!'�2l>�<o�ُ�Q�PЂx$�ur�$�8�م �N��4������>r3��e��Ɏ�/�`A����_�p��8��A�j]����Q�UB0��_J�r̭%����C�~:Փ���h�HG0�]��4��7�*N�X}��|w���k�֔�B`a6���=��[��W�e����9W�ҏ���bWt��9�^�RMf�/q[h6��UZ�%��"RQ��>�4&*���Ĭ�w�c�F���L��TAmm�ʷ q��\�E<#X��~�v=� M�w�<k2��<-�P[[����ϴ0��vt���X����J�3_�u�N`�iM7b;|��o�e�*�Ԇ�s�ǯ�7>����H�B�^�aX�6vc�`E�<Z���~�[�����-�g��J�C�LĪ��g�@Mh%��&$�B���
�������&���W�Q�0Ӄ߳|��"cc~��Jl��G
����9��gZ��ù�jJ�Ƶ^����$m?~��?�1�C[]�)�M�e�A��u�U�����o5��` ��OĲ�}�T���FZ<�!��̸�"8��*UT1n��+p�ew�z3�ly�A�]C�Iv:4+cCKDM�9�F���y�}WL]W,���h,���pU��\�S�
^��0��D����}CZ���;�J!�D\ ���{�ԻE�"7���ȣhif{����ʐ<ÿ��C��վG�?$�V���q�*�/�$���RO�ʴ�H��8�rG��٣oB��q	og���WE���R�u�>��`�H��`�ub�Aj-s%8�GG㼡�TB����E��?r��.�(���q+�V
֫�ۇ!���GD�0Y�a�L��cpt~�Ϟ�Ε��im�a/�b�P��5Sv������e���H�\A�w���Df���5�%FI�{YO:iq�����XSFO�%�H�ي/���i��;��x�Y������U����uig#��vU�(�?����Y5�&��Va/��Wq���u<EG?[��v��"D�8�5�+�(�U���US��1�y�]��!
,�m?R�Ȇ���ȽŔ��!�[d�#
4�E�� LL�u�m�Bm29e����T����B�!��	�N@���f0&^��g�!�܍����8���FìQ&��2W��&��@޿�_�����k_�-���k׃K2�+��I���v`SB���H'g (E�B��J �-���z?��1 �qf���/ҋ���S�ً��5P�����Mn�Xv[�V�j(���".EY�Ւ��r�t7����9m�l�'
��#b-�:��5׌�����+!��VE!x�&��Ewqg�Ɣ�m�9��Xyc�y�ސZ����ݼ�%`rq�g�_�_� ��B��9OO���I=�8����X�`�:v���*��O,'��z��݅>\�:/�5*�ǁ�bQ.ƞ�\���Tz�#0{�zf�fkW�5G٪�t�i5ϑ
�W̅,�6>�0s��[m��>��.Ɍ���hi����OJ������G�Ѽb	�iR:��/|�1#�N		�Q1e�g�ǧ��<�N��(�I��+AP����%�W[��:g8W(��T�"��訴v����>���͵|q�oC��.�9�"��`��g�o�+q!I}cJ41<C�������.gT؛�,�u�B���k��2���Y��Q`������5�FΧ����L��Ȱh���L0B��o�Ҧ�D�G�R��faL6殒4aG=C�c��<ǩ�!r��f!�ZQzI9��D��B��i)��GTN�e����ѱ�N���3��t�d�4d#ҏz=�,�pJ-���H	89A�h�BSasɟ����ӆ�1�{�]noI�γ3�;���U��%V��\l�ˀ�'��0���V�)¿u��TId�j81:s�0��ȕ��#$��3��.~���?�x~�@+�Seo����X��j���"TxhPSפW��+�d���1
}��O��-|%�k�	�Qe	���#�[�~)l��S'�����d����D�w���j�ZmhՇ�K���'��{w+�GҺt��ʏ�!HUgN_��}�q�c�j4P��Y;��]�^��4è�"��O���ԥ�B!�#ב�r�7�ev&0K`lK���0F�P�2C�D ��?C�L�@�	���
e2�c�ٰ��d6F�.(�ݗ�"Ju�tb�9+����l�)жf;��V��ݯ�t�s�!��4�{x�%�&�,��3�E�Y���X�
�u�fT����ޓ��Buψ�^ ���d[0�C�4�$�;���dz���/��kW����T𢤏��
mҲ�UQ��6�i���#f>�����F"��g`�lC8w�6ו^C-c MY���W�U��]�\�f���u�nX�t/����1�l�jG��
^3M�u�A�APFD��%eHU.8P�C�	���]HS ��p�i ѓS��ƄӅ?�PR5E��kI�v)��;��>�>1�)	���� Y�n���@4�.J<f�#���&�غ�q?��B��/��T���oL�TN��q��uQ���q�Hl�i���=����}��whS;����H��O{��YE"ؾ����m>��Z�"�$_l�R|5FO�Y~(5�Kp�� ԩ�H��;U�q<��c�}ы]����/�P�����ŕ	�V$ud�d��$�����/V2qnxC�ˠk'#��7����ޅ��� ��� ��{����ogEXۻ�����aw�<P�T�w�Q������%�b����|*�@��n�f��k��I,�A�]�@�R$x�X��a�O��:�@2e���K�����t�z �A׿%հY���V1��j���(cd��2p� ���g�2V&�.c$XP��������n���q���[��c^F*���w	1,z�]����6�z�Y�J]��wrds�r�[w�K�pj"�z��1Cvqf��W�DW�q�>��ޏ.�H������~��.�bj`.MU�b2���	�"�|F����!-Q�%�"�L�,Q��..�V+f��h~l��u�X#ylz�H��MA�nX��U�`~���
��\�y�Ǜ�Vs�������wA�}GyYˑt䧊V��nyū�"b�����l�,~aqp�P6ʫ��-�u�%Ī��Đ��c��CʊG��v���	�Tm�2d��{�u!��=�Xu�����n��lR���򜋜��%�㵟-n��Q$�u�E(S��^Q���}%j���ɦNmw�eֈj���_��T~+n��M��32�<<�Ś���o�YEQ@5>���ވ�[�:|쯻��<���+4��Q�	�hu��ZT��k�d�T�}�{���:~+Ԩ�@�tp��*��y�6�<1�]}����7ݐ�����α~G�t[*́��NVsi��m�5F�~t���9�);��)�R��+�a�A/*)��UB�2B�n�Z��I~�J𦈤8L�>�Q���8I}��_��`kp�����=L�3Ʃ�J����/�;�|:���(]y�a���j�� Ƞ�v��afDP�h�� [���'��׿�\sH>T��a����z����玑]~F$�ű��q�]~[Ob����ΰ��n*�iSO�����`��ِ�DZ$ʑ(�G��R`VϘ&qʼy�ͪ���'$-�5�}�?��Z0�W����g���M�Frƹ�RCW�lf��j܃CS�c���������g[���� �B���N�����G�Bx��8� �Y����4���J� ��	��n{WEQ0+�3�t>�
-�B�H�s`I��(o��0����Z�n.������h|�^��/�f�^q�b3����Qݹ���ǓO=�5R+|�5i�:��$X�*z