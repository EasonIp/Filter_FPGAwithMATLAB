��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ���L�����I&V~u~[rR�C�XT���o����۟�V/]�@�!ӁUټ��)����؊������I�Xa-�w�H}�T0�me��|_��������M��)��H�BK���G֓�r`6��Lg�6�ދ��׌�ŵ�G�0�2�!�J��c]Mw(�C�����Af=�Эh�c��I+ݎ���O�� ��^1��0s���=9�߸K�V}9��^��*!�S�����p�QtVx]�����S`�)|e�_R ���bd���_63Y��UgN��l��"l�����I�Gɏ0�4��<vT�5���m�༇�µ�U��H��z�4�n]����-R������ބ��I>��L�� 4):E���V!����Q##^W`(�
�P�CI[q���Y�ӕ��Cp�5뿳�p�3� �agD oa��EčgF:K�=/��R��MV�ٳ P�"�:����Zk�Y �{��W��ϗ��ݟ)m�F0�XFk5 ����V�ӹ���:>�H�A_!��K�� pxH���КϿ''���H���%��?H�} VL�Wj��	[��WUt��6(2�"��M�2��d�)��*>\o�䝮6g̍�u&���;AV�{joНgl�z�-{@��oߕ�����W�S���i�f��5+��l�u�Q�vdy�-u��D�d�~�W��QX,_�_�IZ��E�]���v,Ik�5R̅<	�{�B�v�ū݄8��Nf�x�L��_��amY�A�A"���g�.��0U�8W�Y5sgVu�e��s,�	Ә�׹�+�YŅԘ�D��9+	�!�jߟ<��$Z90TOK���0쨃}'Z�b�Jfg�D�fj
���En��n�A����ߡ�S.~�vZp��c���xw��v'�ҚM�Wj0��~>�^D���^���>58�"������`�~���N���P܊o#�����?���uc��D�x���ekJk�8���ʊ[��ز��@����D�{t�3+�?�h�7;c7����#�����)@[�6����c�q)�$�_JF�~��E����6�a���
��y���ڲ��h�7g�v_����jp!�x7�M�l�I������ů�*�����pSX�/���қ_�dnb\�u͋���9�_��9�jD���g�)���쯋PU<F��5���B����$e}���r�Qf_��`�Q�[��eX'�/l���:��)�!Q�[v�	�^�f�	�>sp	�:�~������`=���n����2$u⭂���Y%�}�A�V�Ic4�x�+�%�x��'�}�S^�ǰ�4Br���`�{z�3a�}Ӿ5َ��H]J�H�wKaEN�
G<���ܞ�#�h��ɛ˥Ht��#�]N%���#�z�lc��N�H��v4�7g����6��z:?j9��-#�*s���eO�'8�I�WO�SCE�u3�lV�ѱ[�>Y1�/��j�o�)�Y72��Xo?-N�>�&п��-3]vӐh;���`�������z����h�%��X�v���~��r_W���u��}�[�A�JVk�,z�DMy�K�n�&W�h�\������5ޝC���x�߆�|�TS�p�	[���I��B��W{�^8��*��,^T�[刍�	�>Z\�Zl7��CU͋�5��|qt�*��`�d zx���9���C�*EmG+o�8u>;^�cE:w�lr�9w�<Ppq�A<j���G�'e�L%xt��s�����D��ܕ���'ȿ��C�b^�8��{*�m� L����4��0��My('iӊ&d̉��ȉZ8w�`�����!���<O,|��)3{��:~U�0��Mj�{�颀����%�3�/�?=S'��7��-:^h��
��V(9�p=m.� ��`U0�1�]�>Km�f�r��߻87�UR�o����`�u�=�b���0k����Ox�b��R��T���4ӥU���	�;��Dv�w�3��E7��[�x��ݖ������c5�+�3�(O1��at���z�z�s�cI���?4�}ƽ��T��`U.6�=�P�q��N�,^{܉l��ޘ85�S��/&mw��G�>��H�۰��:��B<�F��8К��e��Ntl��P(�������)r�^ꉽ%f q�dq���3S�� ��bEg|��p�8�a���)� ~�d䢞q.����.�v�Ǔp8��}
Z8���q��)�)��*J�V�S啽tW\{��@=�fQ�,Ȫ8Oe�%ɮ[�i�~�~�-pr�����Z�"�<���Vk��跀L�!�<�[�w��n���2<k��*����<r?�_PR�� *�|~;�K�[����\p����\�?�0�6~0"Q���Tج�����N�\�.pA�*��_j��=4=�<W�yv�afCx�+���Z�h�w�e�'�f�\��"W1"1�$�l�]X�@pɰ��J6b���km��"�J�ϒp�? ���'O6�t���t�a[�(����P�Lu�R�nt���TL��UR���}~��b�#߻��P	Q M������]��}��L�T5��[�]�� �Y�ud�6G騜=��UT��ۺ<<����|p���jSkf��%�L�{�,���!�J���-/-	�&�ݤ����h�@}�7��r����C���,Å�IpZB)� �ջ�5i���w�����P��N��	=�˞N�%=u�d\�(�s3��F7�>+��h!�3�	H�io��(D>1�S�-�
�t'�d|)������F�G��ϝ��B,�
�%�qV���l��t��c��ʁ	��	M�G�q�V�� r-dQ?VL��+^N6��Z�e�s$(�vwt�!�_ i<�;��l��Tjծ�9˅��-������Pp֐�?�酵���/�����I�UT+e��G���E,�����K�}�ĪI�G 1�
�����k�D��]�Z��/��~ٻ7�MV�Ib���d��e-����X��ꝭ�ҽj��@�B��q��������D���W��!��%�g��v4aݘHȑlm�����j�~�*����m)�ν�)d��^D�B�P����S�%P?�ެ�bq�s*��Ã��>ݥ���Aʧ��I���i �fi`-}w��R�о/��toL)O"7�6)�.�}߽�?���U��(Lw�(��2�*�Wܿ	�(P=rI?߫�;YwE(��C���M�Q�RB�l]'�;�Uwz�$j��s:>&���r��M����1��Y���g�'�(W�-iz���k�h����e1ˣb�29#��=_�Q2�grp��D�&����:�[y:�ֿ�L��~	�~~^ݢ����X