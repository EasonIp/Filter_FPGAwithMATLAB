��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5o�h?\bv������Zr]�M�wM��a!��6���R�}���h���ƺ{K5I�*�q�p~"^g�3��j���;�ul��:m>s_`�i��wi��2������hL��ۭu�+U�u�.R��_�o���%�t�|�H-�*��I��x���yiI��`�iJk��B���e����O6��k��;�q_�׆�Y+�M���´}��E7!��J�Ż���p��_U띕Pݻ@�݅'"`&�1�`t�z��yE�W�z�Ͱ�NBi�YJ���VM���T�y�f�rf̟	�-M{�>!:D�N�9��!ċ��A(�j8����n[	��W�u#kNn�.0��$�Gݿ?&i�h����0�g�kq1�;���;���D�,]*Z���3�>YɬK��w�c�hx�]�B�d��ۈ�b���Y�C�.�e[�芬%!-�~�Xa7��ؤ=��7X���q���z�(��Q�P
�!_m
��"y�%��z���^�PS��N�T;������o�C$��No�qP75a�yHp.=su]�B^��9�u�oP���Y�VƎg�嬧���^ʑW+�C�BW�52K�?$#j�PXƝ�LGG�c�B�V�s��l�$J����*���1����h� J'HUg�|��P�������M�{@.YT�Jb�#�Bѓ�refU!�7��A!P-�O�Yx,5�u���N�Cي$#���v�հ��.A|:��Ec�-an����!������^�,3�"��ӳMp�T�֜K�� �#��/~�� �gvWRl�L�c��l�\Y�Z�'��R�"�>�<^���?�/3���c�_�]�EP#YDc����5@'�/��r-L�������^e��pH��G ���3vO�)��Mx�ܞT�z̀�#`�Ye}�8���c%�{����0]��������0v]D�ܕ�j=��<���yA�'Kb��bNך;�km��g�~�E�������<�7(#'m��:�2q��a�I�C�
�tx�i��mN��9]'ˍ��h-_^��pL���xn�vd4�7����k���ff���d�,�g�������J�b�R�:���R�ѐ�=~�L��r�Q����f�-d��|?�GCXJ��j�v=���J���ў)41���:��ؠf�
V>�v*%��Y�c/Hb���+��
,��4~P/�8��+M�2�0-f�}�+,(z��b&z��}Gث�Y���m�O�n�����g��.����?�ʌn�(�:z�~EdWf��@� �կ�� �T�'����sL���.L�C[+9\��3ɰ���+��N��1��Q75R
(�"xp���/��LAkC�rxG��î��xK�3ڏ������{�gj����߈I�$���Т=��0CVIF(z��(kk�i(����]t2 w?F����&Q1 Śn�1D���@Kڜz���"|.s�؜Љ='�wA!X2��54p�(E��CO~��8�`�����4��/���rO3.9��G3�����b}:�e�g��A�%�Gk4z����J���H͒焅�W���r䜏'�q��ֹ����w��io8�Dy�n�����!$��Ɓ/���/�u�x���oH��'	81�]6��x���~�S$�;�ԅm�%#�4S�s�&9�!��6�!���u�g�pz��ݿ��7�D��7��2�<*?���v�K]��V�O
V֚����
թ,�_|	�䄨nH����K>������:i �L�uv���b�k�1�R�.�.��|Q8�x�ƈ��=�v����]��N�y܍Ft�A]p$���N��h���5�5��u��b� ��nj��(@���	 0-o]���	�6�.��ޤ�$<��q�j�n�=�n~8,E:�.Vv����H���E��}`N�G>|"f�E5�A�$0�@��E �c�.�̉�凴���(�Йa:f�;������J#�� �ٓ��L�7R"4(Mp��fNDO��&�A�a��Ԕ;�d��.��̕�#m��_��>�n����:��/���JP3dj���W�L�eF�-�L�v��Q���<&{��F�"/�Z��`��gy��B��"�՞:��(��i�ܢ��Q���匕"Ϫ��w��<�vS\��y��>�,Q{�1��Xv{qDK��/�m~���˵"u�BR0�ƣ�}� eCmF��DG�$B��G�ə(>3S�ٯ�h���`�Ce�������a�Fuv��j�LTN`wkI�^�ѳH:�j��(���8cj���h���	 ࣰ22��ůo�E�ƋK�雅X�P�����5�AD�'�o��Z��Oe�tM�IߌR�0�C�n�����.A�����
����3�h�N����%��I�w|L0���:����ꁀ����0��TIj`�O&�uG̀�~\�������6ڎ͓R�APQ��/�aY=�OX���~����n-?�� �Yw��u\�T�?oX� ���^(��;��w�d�	�o�43��}��}�%��x��A��b-�}����5k��a0LIhA��?�5��r>���q��c@��c����� EzO@\��� �jV�ʼRH�+�Dd��3Qᵭe�<������*+����mʋ���L�F\�@���=�� #IH��#ޡ�%9�$��s�T�d��'�w��"�Z�_��{���!h?w�\����ۦ��B�Fa�p=H�ܢ�le$I)��	bZ���@�T,�zݩ�A ud(������i�X��*������x���z��x�W�'�D�7���,	�z틗mɶ��tVN34}��,�|�a��>$h�a''h���"X*��<�`�=��
���R�'.�6��c�� ��n���f��
�O���ks��i��M�e�)v��|B�$aqߐjo'���������( ���h��.G�Y�F��/v1�<�Ć�=�ߊ��f��wLb �b�r���ҞT�A�+���]�J���jnX
��}(�KP���F*_�߄w <�T��X����*��+�!55�'��U���?�C=�Z&g��xYZ����2�x�X�C�ʍ���:�K�X�$��X�&�A�u�u!��I*T˅uG)`"��D��|K�F�\;A��m�tx����+ol%o�LV��k�7w�uOsdլ��J����3l��%���Bb���DF:ۉ�r��JgW� ���ȭ���f}�ڡ�$��-	h��p?��Ex���������S�)9;8 ��'M��f�EP����B��tܬC g�C\�c���V�}X>3$M�TmA�ˁ!^�y74ݤQ�E��A �q[�>�zW�~�1�
 �BU�>�^3d�wгA���9m�61��YE�h<?;��qb�/�C�����5�U��!t[�//�kiP�S�&+1l}���Q�8]'���t�k��n�Y�j7)x�V*�h���o5�M����	Pp���q�D�u���R̪F)Lҝ}P\����t1�u�<��lj�:F�����d�9�uq�UM!�����@*)ɟu�wYb&�Q�����3�c� ���m����$���bÊ^y]�@�T	��V��a���I9ή�7�HW�)W���JI�]��~hs���}��9����w=)~���pg��C�b�<(}�����B�x�d��u���BJ�G;%�o��R|ߝ��MÕD$�1�ˊӹ���끥��2�o_�6�o?�>g��Q�D8�,Q��l�����6��Nia���v<f���8���:j��H�b�9�x��F$۰��g�a<7�:��P��X����q�.j��;A䋶1	<E"�5z�{���*ՖX� 2�L�-��Ľ��3!�[,-Cm���W}��̊z����� !��Q�kFL�t&Ev�q^X�z�X�X������O֊�R�2�����3��Q�F�������;d��-q.���vjaf��[�Dvd��X{*�=��+�4��@Kr	A��2��9�a�Z�d���ġ�C#�.Ю{��O�ymN�X4ȞHA���`��,o�����_A�E�P7{�=]��W�Vai9�j �v}�ZÌ � �[A�nb\m2���_(�@_���>T�!� �N
�%�&�D?l���!7��@Fz��y���#}v�P
G:�����߀�uyh�2]I���a��
��FU���5��E���>6P){�ۍ�S;�;(%0�&Z�$r�U	�Av�H(
H�Ǧ���9�X�2"���T=���͠�ԏ�
n�fC.��B�B����Y��WՓ�Z�O3M\�8���8�;_���<0����-o\?ܬL���6�	"�� +�4�#�RkF7�j-�1����8Y4���r�s�z����V�7�~�ģ�}�Jf����o���+V;)}���!��cd�����3g�:�(�ҲD�؆�\�0İ�e��