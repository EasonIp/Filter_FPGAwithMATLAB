��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+@e9wR�܄]�-N���w�Tf	��%�9��#�Ac#�3��@���q��#��e3(s4e���^oV� ��bF$)���LĻ�R���a��V��:�V�)������7�K� |��'�y�ѹ�i�^��ы��L=��6���ja�9�vf�X�p2���fq'Wp4cSyt)�}V;����i/&fȻޢ�(�İ�>Ľ�d��!�襾{r`���s/$p�����d}���&5ԉ�׋E,����r�{�h�e�n������AH& ��d��D��i��~�$��� (h>�8��;F�R$Fo[C�^��1ug��÷�ek����a��:�����l���Kk���F�.�C���}Π�q����p�m�������';X/2s��m���;�/4K~�d�X������'~���a���ҥUF��BK!��\���f��.� �w���k�\{�uӏ�p�E"i#c�<lnh�1F|�-�8��]Ka8�ɒ1��_p�4������z��K�����	'/�j���;y?�� r
�`�4ǑU�у�� �}F�|4��i�G%^Ɂ�.yO��� ty	�|�=���ʬ"9�
l`�PKC���3Ðv���ϊ?��=����J16��~�����Wْ���f�e�2.�/'�R��|�ʖ"j5U1���+ ����
��T=W��o7�rV�����|��ZC=�pz�΀+GHT��5uQ�J�=SW���x��G��x E����f����]���A��y��K�������d��k�v*���z_��}׋��2�id�:QEʶe/d���O�E�`6�,�?G!��h��h��X�ak0�k8�0�M4�X��{:�	;��������'�D
Mʰb�E��A;Z�"�@s�\~�X��_X)�{�l�-%V� 7�
���"
��tײ_�7�@wf������I���r�(W��d�>! 飔�;H,'S}a����ahMRsN�W�S�!�s<k��!P��w��i�������es5@�%�LU��sB;n�N��`��-�6H���탖\	������S-�B;��k;h��S�	%	w����"..�څhBW��o�_��ᩪ�� ��y���#o5j9O��l�ƹQ|�hM�J��l�'^�XW�_�@��nc�;��4�{JĪ�-=�f��ó$��z|��ޑ�"}U	ؔ'�Cjv��hx��s|0����ր�l�}q\��,����� >���<yq�B�34}�WU+�8��G9�t�6i�s߻��y7_࢓�y�W[�"k�Iޛ�&���\�]��<�ͦ��'��So�y���($2V�̧a�6@������1<���5������^�hFn$��9e��um����v�6I�V���Ǉ��J1�Y�q���5���W�%�����;��Aϙ]��.�,�21 A{���B���2�y�3�m0�%��Q��nX��Wh��˵�[����ȇn�T]�'�k\4�w@im[l�s ���:U������Ա�%i����T������l��u�V�X��!�����Z��J��uW�HV�Z(w�����4d0�6��ﵤ�*�R.�Myo�տ,1��J�)���N�q���e~7~<9(�n�I���f��Z&(�/��74�
��Ƒ�L�ҝH������X�vNl����E���3��jQ�͠t��'Z���H��[)*���'�h$#�wr��k��P�A ���F��,�ϐ��7��R�����O@������lu�e�2�F��Ɂ�y>w�Ƈ)>����n��Rc>���>��qjn��{"���p�\A��:��E%�8�}]WݦJ��eD�;��g������f�B*Z������x�w�VWq�.M���|%�����#1TڽK��������C�����p���	+�Bhn���hfs�j�KJ����b���jZ�9M���������
#��,�<��g���濶�v�<|��Ѯ�3�V�fپ�ۣ8}o��D��R�{�Mq�<��ZX�������Q����N�x�I�`Z��FX9�(G��Q�(FD�'�c ��Gay��<��cQ*��q2c�G�P/��AL&N|���n��fw��\"%������&p�&9RWjN�{j��R��g��	��`�\�Q�0��P٭`��i>>u���2�v����D�@�[�����O�&�|�,���$��)�8`�˴�cץ9of���P�1z�M�3���1~,T���\Ўh��B�����I��`���bKN�y�a=�%hI~��C;���!˾LB�/�\â�=^�*9�EE�Xw|���]�/QͫG�G�T�ƴ1؉��B��TN���c�0\�C�o%���8�Z�:J��[[��uh .�y�u���0$�88����=��!uEZ�ΠB�����j&,�Ni���!=�FՅ����e�H���B��*?��=��EK��Y��u����LG�@Y�x��Jcw�H�LX�ܬ�W.�-aN1�1�H��Oi�=k��%-sI��U�<�F^�8�O���zmAO�К�i�&���q�Z	��i�҈3�Th���gad~���P\���72�қ��HH\����`��}O=ӯ2�l����n����oݲ���)A)�̹�[�*Yc���>Ņ}!�%~'��᰷�岌���w��?sN���;o	شeI���/|�()��qs�����-$��<��k��9�+��6i