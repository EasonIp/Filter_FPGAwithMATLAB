��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$�ʿ����Yo�1Ҕ����ٗ?R��
Hj.[ptU��%Ȗ�L������Q]���IU��ՐSv�e9������4�?��qօ�w�,�&�{�!|�(���D];j`~���Q�E�p!�⠜v��r;�.e��.-�y&}}� ����N2#SHl�\:.��e�(��TN�Q����n6pZRr��Q�U�M3¬,��������l��8\��B�3c�2 ��Aޡ���<��9mO���n����� ���J��?��w��������2�N	�8�*	��f��Qy�O��~ۃ,��p9����?�PС�q�5�a��V_+��e��Gb�ҭ�n�Vօ6z0w8�!���e�	�)غ8�����\��y�5OJ�+R9	o�_�3�N)�{����b|�2\W���;�L�H�y�dT�R���u�����R%\�րq�
v��\�A�wZK�t�*���z3���]��Y���6�J��q:̖'j������b�,^\��}���v:U�as8���2��f�����o�4�N��j�\�#K����6�
��<���d'�,�T
!�����F���o
n!�)$�P&
�0Cw4�Ƭ��S&�m�~��*�b� ��(�'	'�W�Ά��Y_�2*�jG�4�RT����l޴r ��N#r��=����J^̟�z�-�O�����@�S�»���Ai������]�e�ᢧ�/��#��U����*c����:�Dbt]�u=�}���a\k�"�ko���<w��^Q$��9\xu��l�k13�ҩљ=آX*�����S�pfL��=_UB}����yc@�=$�FI�7��D��4+�*�"&����yT�K�*7k��pO�"P������/��Ch��S~�E"���U��D��/�O�\�Ĩ�uu����դ� �c�G�o��i�$�f�JS����������y�f�I��<;O�wp��$&��g&�%�Đ��%���&W��r@*X�mA��Y��Sg���S��\�U@{�u/�Q	�7�i��?,<��w lzJM�x2�d�=1�5A�扏��xS�������"/�'(���T�q?t2�����@F�H�..�Hy��H�?j���BBF�Q���H�2�RXy��u2���5�K�hCax�5 ��R�w�xl�`]_"\3�iN6���VB+�<RB�O��ac�P��jic�����U�������>׍��+���#m0~W�l�,/+��?����w�>�.�]"�r"�	!����њZt��������Ы���K~?:����,:���ĊK�6d5D*�E�8X�Sy%��!VZ��s����ӓ��q�j��E`��Ȋ��Sq%��o�����J��U���^�P%���V4��E��7���n`D��^|�H���V��#!&����V!����|9�a���9P=�FdQ���$m�|Jg!�D��=��ע��g
?�����4�	���	������Y�$����Yd0�_$�^A��6�~���r$#��ݯ�`%$m�:c�˜`(h.� r�ӏ(0G7U�pN�|C&�E�NWO0
ϴ�Gmށ�kW0<X��� '48m� 1��Z�Xi�"�=d��+dN��Ob��+��@NF[��D�z�&c��:8�x�l.w�,��@��v��p�j��4S@��e޵�@�z7�فl*���WkU~�;L�X��}F��ei�L�Ǯ��l��S����7�֚���񿿣���CMwE�k"�}v��	19f�r����l29-����jS�L��p1O��8ĭ�Dߘp	�M�%�C>��B�]�.4W�����N��F8#��
|��g�;I�D�}$�s�.ˊ�@��NSىĉyӐ>�j�IK�3z'��l�WN�Uv�-wh+�ǌX�i���G�fx
���y,n��j�i�m��/�%'[��q{��E���ƽ@'�vUo�0}���6�ɛ[��xx�T��o��Ep�Ud��m���)���@�\B@���HȻ�����c�)�?+�����i�#i��3���R��~����������?`}�47S�Ֆ��24��t��y�j)m�`�&�� �:�K�l+�D*�6o*_؂�A`�P� �. :�
r*˲��l���F��B`�0k��am�Ԍ���7�x\���ۋLM��3O����G��餘�w�q�����g�y�A6ؤ}�p<g��B���v�J,y��#�(�����zD�9��{��ґ.�4����2mn�ǧf�#�^k{I��S�~�9N�fggCX�}WU;cɈ�ɔ��p�v�{	·.$Du��FcEC�bS]w��6nǫ�o\�d����}��}5�oZ�wH�铫����8ǯ�Y��l���֎���7����m۪��j�L��`�~l�?�<�߾��8DO]�ޡP/>��jh������L������4*�IE�c��צ����23�IF���h�=�d������7�9��T���@:�q�8�{�#b�y�W��_�%�/��o(-@�������LM�a��=,��-I_X@T ��Y)i���5�X�e�o�N���Q	#K���Ԝ��m���Ɵ�%��A�Uof�6M�'����[+��$v�>�a�F�B@�M������}ޏ-��O��?M��-A�I�HM���׭��qR"r����Mk4��a��p^�ǎ3c��ݥ-�s�'e%o*���n

ja��Mn*�6甏$DC�k����I�`���g��3+kڦ:�F�/�>?�?�&��/=o���,��:|S*�o%��`��o��r\A����ҳ�����`����M��B[3��}�WK���m�nS}�_��E.�IO3�02��?���&_��b��Y�a�
��q<��n�$a�h98��3q�S-���q�㕽�Į��L۫�z���yM����g�q�B�.w��^B�5L��<�}�a��߇=��S�*́�����!!?��FG9�#[:�[�FS�*�V$?��u)M�bw�o ~)��*�x��N�#ii����%���w��L��4
�Ů��8z�	)u�~H�T��2C��K�-k ��?/R�SG�+)��KK���a+�4�Q�ю�{�1er�p�0����L�Ao� �O"�W�A� 6�|�KX1�G��'�G��DJ'<̧��������9e��.W�]^0bIzW^�ē���� $��c�vtH8����l_���l��I�p�����U�?�[����"Ƽ_���hY���ៃ���&P��S����39����BB���nG.·P�f�����ﱾ��K���Z*y���<�8+ �i������S�����1������G�ŊC_���8H*����p�4�ub�
1ߝ�H�[��e 3�����i��l,��=ʞP)p�R,��T��
�$Q�6Ǧ�p�;�w�v�j�&��T�X���v���8�n�}^�ɆM���N����eJ��5�qtUʌ`FO�]�q�RTW�Ci-������p��v_�ܕ�(�K��%�*&���{jW�a���U؊����(�*���wt�g����t
��'�����x�.�	|�-��jXe�#�����ai99�b�L����tq�!�ɼJ�?Ҟ��5:������Ö����������6'���5t�K\Q[,� ��^U���jg&QX���)KDN�3�^¹��&���xő�+VζV��V���y��Άk
{=GQ#��9��l�P0c�2F9���<Z%�4�m��陊$�2�Q�i���#�=�gly��q�s��±������8��1�E*Π@i:�R���.�ЎЭ�B=@�;'�__xJ�pc���$��77N7���jfvw2�v�M�'h�F���8�����;���.��.��}�{\�Y 䶝t�B6}���i{<� ��ɴ��q��5d,	�Y��s8�F�6�7a�&g��d�Zƨ�oTк�!�"~�h�����g@�o��g������>~ߜ�hof��_�	�ւ<{i��dQ������%YM�u��+M��} �'�ɡi��Ȯ@�")�0|Y��V�WF��*n��9Rr �4!bjf�$�����VJ3��+g0-bR����Z.�l�	f��ሒ!K)�T�hp�/�p���ܡ�R�$���s`p}��>��Y9m���G��	�k�2�S4ګ���ޔe��0����}w�A ��}��pл�f�"D�גL��pm�S�X��/��.M� �,���oڗ�Y�M�z�vk6B��C49���:W?����4>.g�#~})j�t��Ě�%���tu�W��:�����a���?�)@#l�R�P�.�-�i����0�-���n��P��X���l221�;P�[���2J=[M;;�y�S1���b�:�nȤ��K�W���%���q� �GNcgb�S��5�/�u����ʌvoɺN��k�1�!�h伂 v�D�_>���{�Sz�(�쥆�����V%��1���d�!���R��q�u������(���A��c�����_���=\�D��@�Wl�KA�!|#�6��̻�([ F�^6CP9�ar'�:fb*ţא&վq^����V�~���
j�Fv��s9R��?v6T6�U��j�o���s��>5[�������q{�Z��cbX��'��縏p���ꋙ�E��1���I#n�$�]��7��{���XM�[�i�l�<��Ц�{��t[��\������̂�W����y0>(��T(B�]����pڹB;2�-�Y\�����U�XvK�
��|��)B�;J�t�����Q��^�Li059���j�#ۉ�f���-7o �{~~ү>굄1��v�:)���M��e�݃���" �7!��r�����m�P���}u,�\؁�z,�K���v�<���;��ɧ(�{��fyq��1<^����d�{A�a?�l�My�0Q�'/�߰4��*e��/%�2zq:��َ����	�E*6� U,�}j�h\��(7�A��R�������h��a�C�G��o͏�gX"�"�,�S�v��|H��3��5���$4k��v{5�_z����0 ��Y�FO;���	K�!����#6a�/�l����������z���\yzp��6��)i�����֢R�<J2�X�*�,X9���1�("��P����~�w�ߧǠ�2�_��q�;��������S�0���3�=H*��X��c���ҕv4�.��;�&f�+�	Lθ+P�/d�`"�W.���W��c������vôH_�&o�����l|y�w�X���+:��P�D�k�5s�6�k�4?�OD��ލR����8t�3?-�3�[�4:-�p�v��M#V\��\ZzD�{+�ŵ�}O+V%���!E���R����S���=�7e�QC,�6������	� XC�/��zϔw96�>lnen�������y�/�[%�S5���2�8pg��bö�O�8S��(Z9�>������[���N��;��XZ��(���I��r�6�5
�!���K4{�&BpmeA+yE�!��/zV��V:�%�>�>�|�H���)�\�(.�*��?���`�ԱL��=x����R@s�L���jst8~����SzV��ݎ�!�d�`6�C�§�s�/Am"��(���"ӲP��x��q����莰ZHðیA�^2�x]���%5�>�JA�љ�M1_�.S�U���.�T@+@�5�h��7�Yr�C�Yы���XB�|Z�+�c�`��pB�(��k��j��b�����͸���|0���ꗢ�v����c�:F�iE{<ɓ;Q��y��XЋUSiݔ�x�dM1��ޜ!Y��e�x��a�� �R��y*����x^+�\@,hE�'��t9��x)U.7T�!�+���Ƨp��v����;b,��n cK���m��n�O<<���ƌN��a�	�_�b�6���zg��AO5�nލ3L�/���oԍ��g��`df��݌���'k$�z��������D O�v�&�ᶌ�	b@�b.]���m����a-�.Q΢�_���Nv�	5I�6�ؼ�͂���U�6癰��m�>#:{��1�-fqP�t�9ga'�z��_D"kmH�Gd?v�Q %*�Pa�@�,Dӻ��Q��.��Um{G?x�nޢA��(�b=��_�I���	�Cq����f�kO���b-c����`�����eI
D�1��t�b�/ߴxL]Z*p��io��p��w�X�j>M�3>#��|�pi��������E�o���7�]O�|x^���ق��N3�2�����n'��p�yw��+[C�I�)�e�<b� ���>$~:Ǐ	yԧ�mn��8�3EZ����i�,���u�-Џ��@u��Ç�6b
��:A���:Q�<�֢��۶~_����K�O���%�y?P��:xM�����
��ı>��W{}�C�Ο��o���~�.דk+iK�>�@(�H��|Pnh*����VL���H�B�2�}�0t)�����x�4��L��@i�!�P������E܃��,�-��>���W�)i'`���eh��q��
���:id���0U���U��J]Ɔ��C���E&���+��DW��xR3u�y��c�3/.�w�t��9>�������}�#/����gr�zy)�6�]K�7�� 0)�4�	;. �J��U�Ę����c:�e��#b�h��1d�]	��9|����[��5I=_�³\�d����a/���+)��Ju}�TG��ZcN}n��ئ�Y.K"8	�ϵ�*�����3eޛ&�F�N�>�!*	7��X�R�!K��߻���v?C��DN�/�߽ۆ�E�Iz�����2�q=Ҡ�<�[����2v_8��V��g�t3��"8u}#�-�w6&[4뉽�F�h�k.@!ނ�{�;	�^(�[:\��Q�1��`/�G����f�&�y���1]�%@� �^>a�lO:��_��I~~O�_VNN}ͬ��22&x�7u��tٞMw�b���r�b2�-f3�i��	�]㖻LN��Hvn�h���e��!f$l*3�mH�
f8��G�Ϸ���q��g�{�-fɼ̚��)���j�#����@��ܩ�B�	�7��5s��h�Ļ��*n�Dx	kܮ��,U6�R����l"⨚�ҫ�l��kD��N=/�����lT��Y� FO�td��uyg�� �g��F�R�Bŕ4�E-#�XL��-W��m�L�%���.���t��c�%�-�*�J&	e�2����'�R6���a#RP�>��9���b
��e�b[�d��J�O7�ښ���#�EG��ˀF�L3�t5e��%GD����@�Ic�k��1�1�$+���*&g�2L����B��;�(�c�އ��P��9C���O*wR�P�!Ȃt��l9��0A�'}�oZɈ�ٕx�$K`���y�a�.�/�  �
7����C���-g�W��bt�������Gx���xڻW�8�U����7E8>HE�©�ypP��y��I�w���Zd�/6�tܝ`�������:��L��hfe)Q~��y�7�̕h	��Tk	�gϥ&�#)����7\$��Qt�A��E1��i�WIAM�*Q�;��LP��)���y��~U#�F�m��� (�ቖ����1�)��Q׫�ЯTy)U9>A+%<+>?�Ÿ��Tڼ�y�Z`OuR�]�@���7�����kI�nO�D䂷���+�6��!v}9,s8�ao��qCk"� ��ϴ�L�޲ܿ0�$QD���D)2c��q��X�ad^���$��b]w0�{��w݋�zD/𮪸���E��)z�@isA1*E	r����;��t�E���xi���S"f���Z-	m�ƪ�1?�hr�4.Y_A�����>���R\��"�\��l���O�b%�?��z,��ho�CKfxg�	Ś@��}3J��ԁ/|��0"s��ˋ��d��0��z�E`m{Y�6zQ�{�7�o^�_��	���t�����n%Z.q�	�%���;5w���f�1�����E5��{K�E�A�ݎ�fx�`���御.[$�n��'1�1�|e��i d����G��bwt��`�#w8��.)U�>��gyJ����?�_~�m�����z�}�����WN��6���Q�@"�ۑ���7�04�V�����m���ȝ}�6�Z&�܌���M
a銬2w��R�JI-Γ��R<x���<�{|� ���tY��m8�ȁ��,Xe<{߇�D�N�u����N��������Gs>�Y�6�RN�1g�4)Z���l�ڸ�}����`շ�
��>S+A�w�|)����Hu(�%+��*�"z�dj�������=�Ln�.�H�����+�gJޜ����E�zt4�}WX�|�$^}�8M�uG;)y�H$Z4'V�8�1�o����5H���Ε��ɵ#�ά�������-�"tB�`�(��k<��T�k�HJD�=^t����#��E����Et���tz]Y�N͗c�D��j��L�0#A"@��҃��7o�D��M��O�[v_������(����K��:�~�,�=��{�J��?�2��}��q��S�f��vZZ����=r�-�9+P"�@r�'���Y��W�{������L�c���]TX�eM|��.�� s�; �0�a2K�����8��N�$�� �Yl��<��p=Y�lG��F�:B��[9�������W�I��A���P����QYx�%Wj.o�(pn�DUȉ.����qK�Wȯ\���?li��Tg�\xj�*y3X���9��#;������N?��nu�����)��j�X��x����1b��c�:)��YɚP��A��'A��G���.Ք,�|��Ů��˧�x��4>�ZQr*�"�:� ?:q�rOS�{?�����ܬ$�_S͞��c�o�R���aFWfǦ�I��)��;�o�1{m�(�.`����&�nU�xSIb�@0v�f=�Ȁ�`Ǧa���ɱ5�(�$�)������<�Y��!<C2��WҌ\|�5�>�bv#��1����n�)P5�r��#5�ۨ��3���_G܅S���[?0�N��t��.�N�m�X��=zvŁ�X�@�&��~������m"��1���+4��M�H��ѻ������b�ϐG����q�Yz��CU�GE&�-$��Y�'_��0������鞛�N���V`;�Hpe��I�o���p��Ǘ܌%��NNo�nj^ f�;�;�58��%ly"�>�����	���6�HH����y΀���xQ]�SrS
ML��X��1MK.=�R	�`VHkVx9ܺ�gsI�b]<��pt͆�o���\���Oz-��$Rk_��
T*�
���H�kn�mڄ;��I%.~|sE��W��ˊ�У�ȕk�K ����4���y�r�cI#oM����L��``~�"�(�Q�Ҏ�~GR�� ��^�M�(���\ �m(4�뢱/��f:�30�ӟ��C���߄H��Yn9>my�д�FR`�P�ø����닓
��Z��ȟ����I��¤�4�""�Z|hU�!�t�̂|Z���p�ֹ؇�#� 76G½G�l|�Knf��7`"��'���-���Y�DWt�/cj܂�X˨�bF�[n+�E�4L$*���6F|��ta�bغ���r�eS���e1tX7�3��Yt��[�UQ�%g�&5"�'�:v'Hf����/��Ez
��
�,��5��ћ�<��`�m�f��*�$`q�[ Q�������[*N󾧲Z��q����P��f�g���hE�T\�{C�(*��K���P��[D�jS�'W��+�	�:�~�(���B
��9�L#�[\d�����=��I��J����g���;��O�ÑN��b,[��}{�
��[K�t%/���H s�Y�gA���q�n��	Y�]��R�G1e�� ��C�����;໕�~��|=�@��mDw�G'��>�W����ƪ�ƫw$ir ��-P�e��_���:��_	w<��8%��2P����n��k�@-6!X`�%�-��?	�p�� X6�:g]�=���i]�]I�4v0�^:cX���J�9^�a��,M_���U����
�K��L �*�T��eN�7�<���sp�*�ȸ����y�-~V�xWC��{��3Z��)�������0$?��4<�I4x8�6K[�yED=���G�U�Ӱ7�c|#.L ɱW�z��+�o�\1G)鹘GY�	^X��ZK��z;:-���[�?��?gӶ:4v&�v,h;���̌� o���Y[�'^l}�*�����V�n%Q5f?{:��Z9�;S٩M��`ME���iJFt���N���[P���Wl��c���Q8gL�,��݆�JDW�_ƞb�.6t4�<+�{���Dźdm��b��e��>/�Ν�w��8mx�@E��{��N�L��1���������"�;�9�[R(&%M�ٌ�L��������ǖy^��%PA c:z��ӋL�L����1Y�	^rimm�j-�G4�M�
%Fs����]ǔ�}:�gK��β�	�~:�8�����u	j�0B�`LP�L_յ/ 33�Ĩ^��>�ow��1���U��d�[ɓ[qi�ߜ�1�r�E�V�`�A����|X#!W�_�$~������?��,���8�����q��*%�=�t��N�ҡ;�K���r4��%�����c�}ךbz=d��/�bD88�W��V�s���c��0�CWZ��5t����!��ф��+�R��-�����Ү�H�����8�v/�;�S�� ��P�U���c���BD���T�.C���
.�5�UU��1��%�$M��>
oH/�1�Q�Ұ�T�ĉ����>{�ͻȋ�� G�I���t��V-˸�7��N��S�Q�F�Uݿc/�%�.��g�#����e��+B�|h�~�ᐛBp7��u�hK�x�W5�ZQ1M"(v���/�VyS�-&����d6���>�V�u_�B-� �GK�h�f��YX�"}�rd�. ;_��0��J,�<�أ�h2��ğ䊗����y�T�w���*m�6��t�X��)u"	�/4Z��^P@]���#��)�Ж���vb�iu�FD��ߺ����:�U�G�o}�|�����(�:^��7��F h0��t����iӫ[�1�%�?�@d�[��M��1`޺�ɒ����Ϗ������K�/�]TV�n']���
�����bs���ù�R�	�)i�¯H�kKa&�$����ey���/���I��Q�1P��R��vה��������$t_F�/�!`dr�h��,�9�=Q����nd���x��c�AJ�|�
���b��"�4�X�^�40!����}^J����=��H���-��O1"H5��&��N��mO`7s]�r�E�fŭ�)ݶ�L��)�.��lK+�
{:��ȹ+k�^����L�K<}U�A ����$a���bV�zbBea9c�-�yA±q//�Et�,�sF�fS���2��{�ag��F!��'��y �6��kȦ�%©��u���y��*?�VRNCŽx�A����ײs�ߖ�-;����ێ���>�N�F����cp�� |:B�3��#�PO�A��||. X��_�x<d���������?Vn�)g�@�Ʌ����XN��z�Ǉy���"z{��8�r��ck��CfkA�g���k>��t.��dD&�~�ы�'ӛ��B�f�T%�����P���Z��q��t�FI�+g�w�V��~ʘ��x�M;����ȏ�羰� q(``Pv��&(:�H��,�p��Q7j�O�/��%�(����˲=ARd�Yl��uo��������BH��������F�"}�^v�Z��t�-������	m��(#���L������=N��fjX|i��@����Kq���HԌ��W�w�ěOg��D�V�׼�(�V�	�X��0��ap�'�4�~�MA�o���W��W5 ���ݸX��m���&���;��P�q9��c�S^�~{�R77��@C ���xc�HN�!n'_F�9���M̲.�"��0�65Q�&���y��_w/����%���)�8E�vX��I�ӎͳ/0�f�(N�R�*^������q����&����"�ܮv��$��]\6)��{�rp&���wo�2B��Y�)���5�����ʮ2 M�w�P}W�@��C��:�2�4&��#�����������(��3E�u.c{37��!0����!
ٵ��~6JM�Br�^{�ƍr�����w�!.f}O����GY3�߼*r�'��k����t���9�A9�S�%;[���O&�V��:�XKe+��C�s������G�e ��P���� �V��?�S�h��L�.�e� �����q@�A�S VGk[�.3���;#?4vj
A��:�5�q���"��ȫP9��%��M5�&�o�s��ɰ���Ќ3G�@&�S��Z�C��ɭ����|9@>v`�&�j=�r23fZ��1�5�~�_R�r�H.��\X-1d��������»���$�՘5�Ϋ.+y��]���Nio�X,m��Tە���k�/��@�zܛ���h���b����bv��h?�?{Iْ�Q<����L׹�c|#E^;u6�f�F�L9h��Kf�������Ӟ�S����4w��e���"�1L^(�qcCe���
r�S�_�P��3�3�ww�\j`��>�PD	��i.�Y���۩�D_Y�'M �?�x[�Q &�|4�����.O����9-v��:)��(4��[�;� ����b1®@+UB��	�!��傕8��,�]8okT}%{0���Z�|��ee}Zt9��8Hs�2�K����[gn���Qy�y�z~�T-�$u�����\���7t���/5}y�I���S3]��ņ״Xn��8fНU�+EHbr���4ڷ����8�I�<����	+tֺ� ����!�;9���
�9jzM��i c�UE�>��u���z&��˜	�x��M��/֭7x:�:7���_x��~zW��`Dr$��)�D�+���$�_��:��h}�z�z�vL��8����T@l�$ו���\b��φ��;r�f1�3��v�/��T��3�����ѥ)���!���:��+ͯrl���Ţ-�]?�>&�n�`�:E�����@�J�?�^�
��x�V�IwO����p�?D��D  ���ᝄO����Q�٤��b�{��r�-q	w�:2.���"���Qn�V�7v���Sa�e��ꌒ���㟃�����&˕��.�x!u(�E=�l�{$	�&� � �P�qVs��g�y��]�Cj~R�z]����#�X���I@՟���Ǚڥ	��)~z��/��z��kvE.�'I�dT4c$@NT��ڄ5�# �8򐿦�|���K+�kI/�l��� d�8����`��ے����&f7��D���"R���!��hm�@����6^�� �6�Q��|.�&M럒~�\�EP�k:�͔��R?A����*��i�~�$�朧�5%�v+<ۺ�R^�D]�����PA��V��"�;�$�f��)ac�\s���g�����$�6���`�J���)ӯ ���Gc��P.ni$���N������	�N�^/���-����n�REul�����m�[|��!�!�OKwj�䠊#xQ�ʸͿ)����k��㓰�,&��F��
�E{E#H=��ZG|Pޞ5o��(�txa������	{��bm����NGn:$���̼������&ֵ�ϖ�xW�V�O���_ou7���pZ��y0RZUtD�K�:b�^��Eی�:OL`g�(+hNN�l@�C�a��74늢�VQ��N��uG�ϓ�:�b\bνԔ�Aε�ì`�-ܓ
��I����Yos��4N-J6�N �.�T5I��
 ^���	�I�A�Y���j�س����i����B�P�=���N1�ܕ<�lڊ|��鞖RO3�!D�M������V��I'h�wLe��MW�dfG`����L&������(7a��z�U��fQ�lN;g�N��Gk/�\�
�r��>���iݿ\O�^����h��Q����Bۨ_�X��_@&�7�?֟Xⳍ��f�E ;�W�xX�b��?�����X����uS���Y��|�p�@�b�8�p��_�i��F�+ۄP<Y�(~9�������>�f�G=~�}������"��d_���̦f��(ɷ�:�d8G�Îܸ��D��/A߆J�4-�m��Yq��px34_���
=I���<�j��3����7S��G�NV��]��� ]U��k��ڌ� h5��آ�xm�c�SyNMnXjQ�� �Wy|��ۼ$�]8(*�����3q�}W�WK��<w��twr>�'�z��3�x��=G�s�E�%S,��w����ؚ��iQ����l"i� Jy����K�h��;�)��i��
<�H5A��Ts��N>�v��Xس�u�u�2ˍI��{r�"3(�4�,�ޔL{��`������5�d���e�k��%�\8�d���w�"z�`H<i3��EWd<�N���P���z��S���8��ς������\��P�^"��j���z�+��NЬ����_g�V�I�PC��(���hr:�I�x��5�8ߢ�����Y;����[W��%���^��˫�U�H�sx-r�J�)&����D��K��|�V��-ޝ��"�L�3�є�"��=��P�f�@^��NOs��de̕�q�I6�R���� �8��2_�1~]F?�m�tY�hm���T7��p�%�G���x�ub��'�|`�Le�`c�`s�U�``2tI�ړ [iY�`&{���La�!�������ɩ+O�Ӟ�6��i�V�ȷc<Ѿ��"U�<��4T����4�)�,�_�lC��)�=|�e�N|-���r��M�h����R����_�R1<�5Tr�����Úw��Q�#E�a	����TɑN�9�z�E��	�E�X+���{-��4b�����	���5�/��H��9R'��<���&(Fy"���W.ԕ���#�`�@��@�{����X��Ɣu��a7��h�&�o�
��1_,�&��I�dY��� ��5V
}K����z��j3��[K�=\���Sz <6=e�ۃ�_Da�(��#��ny���sx&Sl�9���)��o�vR�q��,�����Bg$[���;^Y�l�ɇΚO�[Wi�w�i��e��w���ک�V���%;tAɇ�.�-
��'�)y_*�9��BsL�4��n�~�s6��+�=L��\�G=�9�kD�nO�[J�gҶ�����{� � �
�$)�a�רY�[5��<s�8�:TZ{�N-f+_� ��~���:	���[�T|H���O7��d�ZTn�v����dc�P�QT57߼�9�K��W���|���}��@����qt����Ҭ0k&��І��W��W�WG ���BR����'�_z�{A���/$�Mp�(�r�V�щ;Ӯ�e	�E���/����y]�@'@�/�� 2W�q+U�T�Bb[�=@8��@#���.�����V:9g���w|�&�&n.�z#\�`��囅`y��2q�Ȉ_oBP��Y�'����h�y��6T'�Q���d��O>2f�y ��$^>�s�8���L��U�E�=�uF^�9Ӓ�5�Lp�Z%���׍9��NO�T��,�>�qr0�.Ġ������c�m�ːa�+{~f��~$����  \0h}_[!--TCؾ�@��Vҽ���?�6��M���#��W�.g���u4S���Ze�
�0ϲ�+��Z��W���$�'�H��.k[��d�������<��9��`��'�^F�OW����m�p_X�'�K�|@���U9�>�Enb�=QFw҂��>.�?��ڡ"��MXشR0���]��C,�1��w*�MwA������<o�{�#Q�t��J#ҍ��_�g��'dGBz�Q
���q��%���]���)�c���,tB�\K�V����As�!@�q�� u��ØzM��V��!����i� ����R�����_�)�NH����^�v(���8x8�0B��4���� E���ٻ���j�<́k�Εp�(�>a�I�p��|����q�뷀�.k,&��� ��
�G���{"����_��h�o��s��$�\��(���v.=!Dp?9u���	�/�Y~��OY���L&?�N3S�5�wѯ�Gb���FYJ#�����X:���\�j6�hH�$d�url�h��'7e�V����	�lp�T#]�@�}����_��Ql�<c5_�Y	A�}��;;F��,��f@L"�^Y�u��\�1F�H�f��_q'9�OK�w���ɟy�zD7rO!J`"lA�/N-�8sYQ�q`���S��I�]�y֨09�������N��:qVV�xUxL�ӑ��x�T�dv�u`�/Kv���y�]7gM��)~����g��0sݭ�FC��2��V�^�4�ն<����g.vu�U��P7�4�R��,�jQ�8){mr�w�����!�R��M��2��qsNdE{��G�_��ҷ6\>"y�sh����$�|�D�H��nBy�Z���^3�k`�[�.�&[����qe�e]��\�_j�I�q��W5�%�`kК���_C�a;O���",,�#�>Z�D[!G����.��4�n�����ّ�T�Ps�-vC^䪃�i�ӑs+ve��p0�.}BZ��[\+(�C�x\ͭخ�Y��Fa\��ܙ�YN��{�Cv��� U��Z/Q��7l-����S��$?��P;q��f�;����8CnT4�y�(�,���^���Ն�#�5��SD�ܲ�-�]�R6�Υ:g�51]�FUG��ɡB���W��k��Ta��%8Xb*�6�I2�!^�O���G�Z�\!����\q`<	���m�ct�+�O��[�_�k���2�e^a�����J~�,�ֺ`}�1�D"��y$�!u�D���t�ek,���L�zX!{�R/�]8jG��V4�C���,B+z��ɯ��Ĭ�����\�G��˥�},r����Y��v�ݚ���Y3>v�Y}Yp'�e|�/p�ۻ�GA�J\�]�8I�_AWN�p��&�E�yC�@q%�5
q'���Q��ӥ J��؏�LW�gh��6ޜ�j�G�f�
^�ɹM���J)����A�4J����N ,��j�l4��7.�!�0�4Y�1��w̱��΋�n~K�P�އ��@'?�9�M<��
����K��ܟ����?;�ZL�ųP(��m�+�B{"��nnp��F�@	E*�����/ ��� �_0�.c��j{�[����ʽ�����ٜ�ȼd�7n g��ױ|I��b���pZ��mMJQ�٭��P�~��~�as�_=��CP�rW$3k\�+{2ZJ`P���s��ozl�|9�uf��U�h�s��Y�C;����x#�ͫ���\��guX�i��_��4A褪_�W�����:�C'-~J/pWv�����\��*+5~��b����m�n{��cm�N�'���nz8"�������v���F��,���S;1�t7n'
�^�BC)�
UU��|����z�jQ��y���V��p��V�w�\X��qA~�'X�39�Aڲ���G����[��Χ��ġ�4����5}Oǖ|�T�U��v]vu��)�<k��-�;f��s�h
P�h-���;����*�%<G�^�/f,����K~4ٙ��r���Ӆ�����,^R��s���������>�BR���?Qd` ��@KG
2���QV��)�H�XZ[�g�<���~Ң ��z�:����;Y�,*�}\��6�z�YF�t;g����T\�|z؉�����%9k^"����Y.,�
�s���"�Y��$�ׄ8���=���Pscww78��K��pnz�d2c�=�J-f��+�%��b�M�)�!�^0l8u��?}��-�(A���K
95�o�㕐����Dwߞ��͇&�(ϸE�$����zJ��"��$[����Ϯ"���*m���ֺp ��ȢH�e;�r ��::��rH�93d�sZ�~����)�� B�:�]#�"y��:r�`���	1�d|�L�@���Y��ln>ԗ`C]�d�k��mn"���u���j�L�����W���&n�˃�<*����
e�;n�Np-�{ֹ�l�Ӎ�z�����t:��YqF��-#������r����@�#�D��7��E��{�6.���]>1�5ɣ��^�kγ�?s����&�D=d�|�RB�F�D�Ó�&Uz�<'�G���S\5���y����d��H)�Ս��v��X���X�!��z[����}�<*�!��?�װ�t��<m�{~Z�h�hK��X�-tW[zQ�H������)i
H�K��s;΢g���n��a�����M!�'��Z�Tj(�w1
��n�zf�dȢ��g�NXj����T�?W�LtĞ�J���s��W�Q�`2�@��E�+�Wt��s�6&��&BThᠥ*���A��x��J�i#F5�Q���;��)���X�䑮�c�|�#�@4zY� k�\� ����qCF�[w�Q�n�{`�j�`Z�k~������%�W��Mz��kV��l��}�*� J1�)\�M�~�}$�r;G�/5��YGNs�!����g�
f�>�:����K�'��0��^2�vx1O��}��ꤙT��t�[��������J����K�e��77�e1TF/5���*>�P:�Ơf��W7�O�1FI�Q�q�$��$�M�P�)s��1��i�[�6;���~�Ш�}j������6@�(�H-�@6D�Qy����0���}�8��0v�9�Ρ[�FX���xH�����D�<�f��%��S���|K�� �p�Sc(^�}��\��?���=*��P�5f vde�0r�qK��l����n�y���0x������E�� &�T�CB����5���Q��H���n�A^��%�G�����p�n=�W��{���V���*Q�p�	�	�SՍ��AZIK�������H�\�lI1]���)�Q�W��"���r�D�D_����M��N��	�8����4�y�n�vb�#��� �����u/��R:�0�Z6����.s�d�4љf���A�3|��~�7��{��Y��5��,[,:��F�9�3Wu ��vA��;���{�lc@e��x���F:wRfr�DU�X�H霟y]�c�ôM/ciA�,]���7n4].q(Գf~��C�	�%��-#e%L"ȅA2f'���E��e.����3in��n��W_���	c�JƼX�c�d'}رF\O� Λ�,�+{�{j$�L���� �G �odc�v��*5E�1��3��e�L���w�n$�{ �RΓS(��~����ٰZ�ƦUˋ�P��Ès�X��3�ev��x	�Z�'s9�����l�²��8.�k���즻ݚۜ�Hj1���|�[?s-[�߃:{�ńD2���]v&��t��<�VCO7�+L�e�*��?��#[��?�ZZ#�G��0L̺w���.�p����$q��jd���C,�k�5����s�5*�b['g]��F�ۤ���J�S�nM�yXB~�`��B���N��fQ]h��V�F�����`���;#��xw�!u�yO�mK02<q��VM���h���R�N�	����ϑ1�Α}��6F�9.�M�U�����7�Qb��<���E�����R���3<����2���w`��:b2�PZu����7��Υ�"�M�9���}o�9�e�g��9�������j��9��+��4|o9�Ѫ\��T�#�qi0C�Z1�P\k���3\!��H��)�o}�5 ׈���J��)���eyT�k�������F�x*����/^����������޳�"���<�D���E���䑵o.Uu0A��
����T��Κ�BC�g�|�$�狙����,]�uB8p��z7������~��C#���&5�o�6W�g��\��8�> *�U__��,b3j�O]�&�V�b[� ` [�#�����0�%��NS�;�DFEp�%�ي��XU�v�+N��j�*��b���o��[):��g��]��E�'�3Gܚ`��97��z�����<~�oh���ȧ��|�v����D�&{@ve6>`�}������r��P\������!qw�vO��۽�>D��
p/�SX���tx�.h�M�!|N[�m�7���J*z��2��O³_�s��[�� ����#���)qrR��}��N/ ��¡�H�i@'�M-wb�!>�����Cc��������޲�		96c�%S���g���['�-)���[����d����rk����PV�	I�N�)��e�fe��5�<Fڠ=׭�0`��G�;BN[T�[U}i����{��/w���F6�M$ �)�����>��Xg�w��C��k�ߩG-��͏�A���Q>��Sk`RֶHoX��t��^��5
�:Wv�C�c�nRX*���o�3R&�t��L��Ef!U�TU݄�,�Ԉ�0]-/}�)�K�Q�qɷ��7�D�o��x;}���IPT�;��D(0L"}.���pT@�d��*(��X��bV�[�A�a�؀](K?TxW�(s��X�����âҧ:w��]���rD�zE4�K�F��4B	���	#:9��7�A�g�����|���@�-��rNS�
�S��/Ĵ��^�����N�eYQ&L�����׷�����r&J0��
�s(�D�8�4(����ƅ�䙌)B-��ih�KÈ�	��͆�En�ƜBژ��	k5q�Pd�i����'��Ms�z� �fX�@R?���Y�������fGň�����_1U'��$Kl
��A�@R�+���%���Z��t���.,B����[�!�E��!�R?���h��؞�t���O����~;�}�C46"�w��>�Q���#9�4�_ۨߢc�A.q��h�A�Wg�	�6�@��+��(S�q#(#���>Fw�&8�ir�KA�$���Q�cf$b,�	$�(���6ѱ������	d0㫓?�������3<���x\�Og��@<����{إ�������ku!�#&X%�A�'��M`��������,�U�ġ�`&
E%���C���
�ur�5Ɔ̼���\�K]�F�����Ch0�g��{y��v%����w����$���6̋fQģg3_tiבA�1M��K������Z�z�P�ę�$�?k����\���������o��Oa�g��(*/p�k����(�	��'�G�ainxV���o<��eu�*E;�́	����7�ɪp1�LG���\�����`���͔�igݸ�A+����·8��������?��:��V#6-LhO�5��*b<ær��r�3 ��"A��ש!�5����S)�m%��ޖd���*�mԬ�n\�J�b�;)z%��gm�VǍT]���`�7�[A��#U�4������ՠ��E�[��/) л�\ ��R���y��Mfݗ�]��6�7��6z�����l��(�la��A�)��O_�&��� �s�}u?r�-�~`U��c�(�)�O�����e%c���5�]�O�F(_^nQ�C��/n�b����n^���Ct��&��u9���'��iӪϣP#�*\��!n���0�)�0_׶��?}�*k�/�]'�Z!�w��r��XF`���B���ܜV�T]�+n�Ja'�:�{�3],���G���*��N�AO�401=*Xw�f�n�Z��*U��zsĈۿ�խ�F��/1H)7i�M���gU��8��̥Rp-EN��7Ǐ���(b�F6~���j:V�Z�̹��wөТ�q�[��J�$B�� YZ�Rm.��I��ս��*��l3�^i]<.���#�,s�Ky���ҝ�Y�k�e�i:�{���Q~I�By>=���7T:��P_E#�m��)~�n��a\X�=8p���������-ڳ|�,Nظ���@������~M#�V<�ү1EBDl�&���	!S����h3&L0��9)�d\�F�1n.�lMjI#��YZ�}Lm���ӛ�ag>m�|��;�� ��f���4��HRE�� H�nLذ�xI��l.��Jh��'*�q$���F�	+leՐ0`��$�r|!��/.l[�D��=x�ë�ڭ�L'îc�ba8�CR��)kX�T�	��wY�V�[(q/u�f����:t��~�N��ҕ2rj���E�0��.h�9��������Y������W
�7#ԥQ8q��H����e��r���2hc�n�7C5Z5=��J���ʇ�8������3fEX���֬=�-M�\��$�5�[��r�	�?]�8j�u�+E��eTX�^���/�5%�(X,����> 2�N{~���W�w�����QZ���?�QN�����49�/��?��19��4D%f����.V�T�q�X3�����ʦ��Z����g���A�O��(���hۭ\�e�#�	�*�����ǦZs��g �� %�_zg��%eF�18��u�������p�m�Z�Xֵo�&Jܘ���̸<\6�^�V����_+�>��&r!T���0kd�Լ��J��a-��,�����"��2O0U�޸56�/?�e)�������R�T��6+l�.g�f�{�D�Օ`b�,Y�`��"���>�A"�Xu�&<1�����|ٛ�C���F�~��C��\ߊ{b�duAhI��a�&���V�Ӄt�mXX��C�)O)j��#�Z���s�I��O��m{k$�J���6�#p��^o��ڭs֜�!�Q#�ϥF�\�����g���wҊ7�+x��oڽbQZ/y� P�U��|������o�$`SҦ�bd[,�B���hRty�_�zަ��t�J�td�M)VeO�V�`ce�%)Eϧُ8h_&�N��w��oj��~�����1������f�?F�޿��}1I�.2�)ݡ���%U+�s��#/�c@#l�R�1A"Mk��hG~@m��m$M�S8�4�Le��6~�/_��@�R�w�h���Ѩߊ�0<v}<���L	�f�>����nKS���[�U��c���]qd�f�X��J(���%~����f�� ��B�]�}a+ C��R~5,�>Ӈ�r8N~C��
�;�c�����.]�?����~
��?�YQ��z��́g>"�C��Gc��>�ޠkp��DV��#����D�p�-�/���ςx� 1�H�$VW��uՈsC���ѳ?GT�y8�����OX<��V��&�t�z�B��H4|��RJ�(vp)t`�,�Bys�����J����6��OZsy͕������ѡQ�qՓg	�'��B���Rf_��Ƴ0���p�j5ai��I����z���D�( �sS@���P�1ʹn�3�m�-��۳��!8l��:~�vn�h����g��G2YW����;�i�n�#TH]l�=\�v��bt�)�_��ݪ������*��);���M�z.7u6��~�Ȍ=���C�p�ߺ��R�YI?�K����"(��D�nm�!�8R���^�j�UJ�x'�5~�v�L��	�f��N��K�eSI�)dͤ���p����@1o\��{��k���	ח��,�ŗ�#ga��V ��gp�i�F�] ����-��c�k�*$~3�ϡ���C���9*�����s���g�*��e͞�\Fr����r�vp���7Pq__�X�f Ƹ	f��A�?R�ۍm� ������ �m���H����~��[-��}�a�ц�e�~j����ک�z�/؀��ŇU��� K�M���ŕ���O�$\���[�(k��n�"΍�}p����5D{����'M6�Wi8�cqb����jW����j3�@�[(����<&#9P�#� ��6t]g~�'L�ئ+�h{�6A��,�\h�,�2��T;�
s�ؒ�ē�}4Bk�"�kD�۩5wX��;i�]�� ~RۛqxJp�7y���$W�����O'���Ta�ؾ�`ws�h���ۃ�(s�W���k޷*� ��P�z�x���{�ԥ��&7�M�A�U˛pe���>ˏ/�yM�s��D�$'�6�AfJ�k�ufL��d���F�ݺ��]k�=>K��a�O9]�)�u�]�Y�Y@;��s��)�=�0��z3P��*Б�|�f!�IN�]S��B���Cf�;�	��LF�f?��M�u��4+x;�6��"6#e�����2�ޚ�b�<��|{���������/�4A���6ʡ�sN�Z��D��Ǿ'�Ci�[��r��-�6n^��z���ۮ��#Y���s)�K�C
�)<g����wzJ���*g���e�)*��ueMP��o���ܛYYC�'!�tH٥���T`M��gD��n�x���/�]��W�In��zw5]����'B&��P&��=�r.$���J<�,�<�K��h�n����	$"�M0���H_���Jc~N[���>����Ğ��@���#{�xy+?��#�t��B�	���,�Ld��T5��h�#
��֓`�L���Â�&L5�(-��e ��}'G�����`7����Al^u�ś�J^����?���>��Va?g�s����/���yx�XԷ(�D�n����qMn>����P�r��S|�?a�Ԯ�� =�xƥ�33���`6=�H�^�IP��o�\ oXQ�;�P��A�S�u��B*A�?p��E-�0�����A�q*!d�+*�#��UZ���T�a5v��L�ߋ���;�}��+
h�#�}R�&5�v8|��'�(������-pv���ܨd�\W5�v�l�9t\��m�E�:(��ăɓ�NZIG탨V� ��83�tv?���W�%�!?��h��mT��H������j��5��k��P�N�RI���mT0�
ܲ�W2xѱ獿�Zx�i�&$��x�*�%���Nצ$��0�1B����?d�`ƘhV%+��� c!2K꜈��8��M\!�ٔ��4��1/�N�RG��D?J�o�SQ�発o�p$��G`-{�r�ԝ+K��rz/������B�Q	�j�]3_��	�i����ݒ-��n������t��YNDe��x�d>l �U5>D�4"RC\������/���r��g�>OƑ~���`����Ќe^�U*ē���)�G�<Vg~Q�)�N�gh5�`pw������E%��ť����r_��@�.G�c#c9n��yp-������
��͸�3^
jng��:�֙8%��K�&����$ڌ8�;���酔�t�^ie/u�[������f�H/������K� ���«�y�Q0��a���J�����u��N}d`,-"���z<�lK��ĥ�ɗH�A�)��u���S��`{�W`�
�!�Hgݸ ߢ!�c`�O����Cb����y��xC^����@���J�Y~�H���p|��,�W���[ ���}v�+ζ�
�>�\��}�G��U�Ϸk�J b��C��\ds�p���)�
��A<���B���a��D)A�<^>��A��`��a��� ���������s�Pa�x�IJ��_.VJ�d�7�3�E�}�ӫ��M�D���Vk_���@8��h��/^��`:������2h-�_m��--�
_�͚	��:1 ��]q���m���P�9��Iƺ��`��2��Ͻ+��l�~�V��<�����"A��1_�
�ŀJN���c������D���Y�%�2*�#�P��&i1��c�v�QD,��*�fI3�6~b����?�29�.�A��X�M�N5:8�|F�@6q�⋷�6]씘�
�[�`*�]��;Y��
�<��o�����q+�$�Կ�3.��S2l���ί���� (��FD���)���B�S}�?������q�K7$�6�~⦶��n��,����ԫ{b9eP-�V��C���6$��x�>PU4��&Z�Hm�fm��  �	�K��w	��:h����k�TG�	�%dd<r��p.
�\bUq���=j�d�� ���l2�wא���i��TA�>i���f`�"BN���gW) �L�O�vd��%�نҥ��}�qc�j���(�
�#ʷ/N���^���H[v���x<7�%���a��T��bJ��6��y���g=��m��-]-v��j[UHu뭫�1$7>��1�,���]-��eJF
fV�|[��:{.��.����s{�ŋKPV4 �[�7����ĨQ9=�ܬ��U�t��`�s:(�PJ���~�vVB��֚4�ۇn
k����z������ίK9N��	V�tAv/�=�~��""�:U����d�ߒ ^�8[��`��?	�>~���,���%��ϟI�/��w OuYgdw+̃���e���ޑ�F���:�;�7��C^(W!��Gs�A↺���n5$���ʚ�!��9ק�H�Q@a�e.#�~��OЙ�O�����������W�.%�j���&��9o�K`�	��q/3�H���%~7�)��d�"���R��h{_����E4<.���k\ξ�b�cx�<��
A�<��?�<�S8~����΍�JQ�9jtL���?v�&�G-|r���h�gts �>�
�ʳ��_r�cmhzB2$���U~0h�W�{9,�����=�v�߄�����s���og�W�(!r?��.�Ei��A[�iy�����{H56����I�k|+�Ҽ��o�(��X�10�!�-VK۳��-�T+�]3������Ì�Gak�|1��k�v�|[�bڰ�s!��<rA��rY~Qк�����rM�֒~������D	D�`�e��h���@!�������h���C���x�^�Jz��hk-����˭?q�*U6��	������@(�\��L���69��X�Ly��MS����PS��q���(J�7�_�h������цTU��F�<�)�3����__�:��m�5��-:����p�������fDb㦫�8q��H2�!
G���1�c����EX��lq�\)�*ۉ�?�ø�UIU�Jv"�vA����P�2�N?������t��2#��X�們�r7Qʦ���'�XwH�Fk�=��=ʼ_�R��7�~7<�C��ɇ�jn�].�zE���2�Ao
�[r�cL׌���T��wr�Ƶ� �R�ҽ��n�=��œ�Z��]p�����4rkV���/�C�g����f:��O�%@aO��u�D,�˦^,�m����[ y�vQ��b6P�h�S�'T���3�>�	�%vz���ߚ1��C�,�3+�ݨ��0a���ɷ��c�1��0u�Ӷ$v�Y��P��W\X;�j��V	'["�tY��bד&_��d��қ'���ZB>α��!_u'H���š�ՐڄS�B���^�5T�2���0|����H�/P��B���U�p��n���B:9r�����2�����s)j5f�L>��	2�9��v�8o&��9}մ���w���}Q����}rꘓ�ژ]SX�P��b��=�ل������d�����7pȩ�b{Q�c�=P�0
����A�&r��i���UH��M.q�ީ�7��Ɉ��!I����=%��f2��s)NTg�EӸ_'*B:�}��� ���,׾�{��Yd���f�ߓ�7��C!F�}���FG��E�x��@m"��;�7�5J���S>J�R�� �Bg�K�SW&O�-����I>3&�t�=���RL�,AF����;����P�)
1뿣!>�M[!Ր[� ��Z|k��=����f蹥���ǖ�#�i#E.z5T�S7���9֘��#Ub��^s�Kq-it��&tp���A<����1N�>5"[�u��2L��gQP3���k�P�)�g�H.��������y��R��eAұ�*����j��ʮ�9�ֽ~y��FFr��ˌ�y�&�7�>+�4����c�Pӌ*�����pQ=�@+$}p�����)�%<�k��iT��cD~>Q���p_s��\��9$���>;�+�1����/�h�P�3g7�?���YX�9@�s����T�Ѧ��D:{���/_��G
��o�-/ū���h*L�{�x8�Nd�%jz���8gb""����a�2V��U��iQ�?�c�خjG���?6��ؚGu�B�`��� q�1��x��F慦��^p�`�� p=��Ɓ�Zc���z(qA�/Y����R��(��*i�h��3�V����?���l<��2:~�iK�`#~��g�%�JX�B�ܐ4���h|��\4m�;�i���٤]`]cp�=B�X+��Ls��m:�:tn$5 ��x�P��C�6��I��>��}�9���j�P�!o���z���;���$�9�v�j�:�2$�G�k�%q�O�ᑨ��LI_��<N��kD��9lX�Gn�E[�n��5n�G-]���F����L@vBn���U���֕B��@o�}]o�$.�H��_Ѓ'��_r��hx�ma*�Y����[�L|Gpkm�=�3�{K�Ε�u���!-��uu�^��E�~3���]�*�U�@k3-���˕�}%�����aUf�$L$Xݷ���G!Q�RrW�K�qp�ѝb�0i�r"J���@��Q^��JZE�0Q�M�Q;�^���1R�����IKh��$g�i�R���\U�ą��8��u�O�%,L�&C���U��uQ�#��-Z�|۳�nh86h�4Pa>#����.���|�t^3Ȥ��n)F�v�1��-|�o9��Br,�M[���A���3����
�ޗ���	���J�Aj�K)�=Z>��X�P�����"[K��U6�6F�ړي��N!,��u1���S2b`p�!��u�#�Zu�hʜvqe��vZi���w9��h�30�<m���B%J��M����~c��CI�Ƒ#xw�	P�_�x�o�g���R�H�gp�x�h�s'��:��3{����9čk�P��DYZ>ty�5��P���姝��)�S����s/�W*�m���5s�~N�fм���43�c ӡ�4l{�MX����&�y����uÔ�Y%�i��\��
�F����g,�'�/M8!nq������掙�#��ʪ�nBK�lpV�#xރ��ȭ���'/*�7�"���6�Ros�Y)J��}|�D�c��=��;*?���W]�Yr��[�ݪ�H��t�a#���	� ->���K�W�p�~l��%ؐ��Ɓu9KL���X���lA��%�h���dԕ� g�G�����N��lG	"{�8%��Tp��z/ZͰfP�ք�/,��\!�[E�1`�hKg!��3p�I����P�|?���1�Uq>�N4��sI�u��_ �܋Τ�j�0�!�ъ��G4�����sc(���m�Q���$�W-� &U��1Ҳ��M��l�I!����E�����R��0��opg�Тf�3�QP*(fxrT#;6����]�@(<|7�W�-+���<U�~��RX��@�WsMLv9&�s�|]LY�$�e{�{Nf�R����b�ڥuf�c����~>����Lp�Iy���"�l�«� OK���y�\�dpUf� u!�iL�M�u��-xJF�o�����֥PBh� ���{|�WL�Y[w1^������]�/�#�|/����=an�h��G��ŝ��ge�e������+���ů[����L5���;b��	��,<7�'�*J{_v��5���aZYr`�nЈ_�E#����^��ra��}�#(���2�B���=K�9k��Л?"�o�N�@��@��;���Ms��=��	ѥ�Oq��<�U���0�y��V	
$e�?x�c���ξÊc�b&a���Z�A-QZuN7��q�A��L�H�2=X�V�V�G7Mh�D9[��J�-�v8���@�\q��s�p*	.���{U����*��Z��V b�=h�'o�,�"\y�F,� 0�[R.Wn��7nc�lH��W���Z�Q֋-�Mg#\���o�C�J���7�h���nI��	�aP������t�&I7�"����>�]D㐰�a�V��Ր�w@�Q�)��
� ����
��K�����M��Uj�g|�⑊�T�c��g�r� +g�L=dP�|�AX&өo��goG�!P
��o�7��w*�-�)7��ǐ/0I%jD�m`����Z!��|^�#����A���I^�Ԁ{�<QmM������gT3פy�� ��������*�$7�۟�o��b��Z�SyHz�E��T�0�p&��✈\��H�vm��e((z��H��_�\���+��Nm5�dw��3,��+D�$��(�/�CPva\�w�=��m0���Z�����t�`)Nm�aN7<��Ŏ�l沚n�!���x+����v��o �_�E�6��"1������4��4J���No<���v�<ES	¡v���(��-&�`�W���Sg��=����}5�_�'��7�&�4��T<\��Ȇ;	铊g�E؂����L��\�9# ��F�b���/�)��J.�%�&���ͪ:�_�r�L� +D���1%��	�����7����t�T�lX�,hD���L�a��t�.vX=5�(]�+�crY:�_O��:qS�2@ڨӊU��W+��	eg���}�Tꉚ�g��.h���o|�����Y)H�p�BN�C�.�۫�9���'�8�}E7f�e�pxZ��j���B� )t�!���e���x�V��	���Z��hB�&��2��".U����<p�i�J�7~Xf���A]�.N��Ki��d`R��� ��.���@&�qD趨�����r�����TH��+s� Ï�4(lV��yS5���1���X��t%�ʝ��Ю�By3�͇������A�/x!�ަK�s�	j�!����E;%T�r��v�"���MހukZ��af��M�]Ƞ�k������&�>ul��e�m��R�W��~�b��� �|dg<ɕ�*�&lŔ�{���0$t%T㫩Y�Qq�/����w�Mt��
��9�N�뾷,r�Q��k�P �T�ODD����ݦ�Y�^���5�Mdc�?]�g�G��F��1�L���I����p/ �X��q ��a�N�l���ʔӃ�k��8f��_
և�0��n!>��%66�J��'��P����(��}�J<5�y'�F�/b�<�R�?Q���V�
Z6�����3]D6�kQ�D8ď����W��x3���V��m�ёŎ��t�?�BfS�a6��0f� ����7��}EQ�����=�AJ��JJ��r<К̎:�����M�ϖ#�(��d{�Gux�gf��7H�b�7
�� ̙�u���(��f�)�qƤ��]���(3�	cf6\>���g�Ǡ����A�k��i�tЅ<�GJr��6�����$��k��!��s`Y�IV��?&���W��h�/�d	e����h�!�<�m^�(�$��i�S�$�^��b]��AD�Lb�R}}�5��%%�m4澰6-r�[�DO�<�K��q��6���S���є��]T����U���:��*z��GJ}�`���X8~�`�$�>;I :�ƞ�:R�r���9(e��Q�tư{��_����z���l<S0�g��V�j���(�7�dMV�/������LF4o9��E� K��}"4?�S�e�F�T���b[�d�.I����r�;��{$�P��Q:S�S�<[������]������;y]v�Q��G�ۏn2�P��-�hS��? ��?���s=j�\
[Y2v�і�#`�-�c�o|���G�`�$�r��\ҠB�4@�1���j?�A�f�ޞ����;I�����vSX�l��ʪ���������!9���z���nJ�9�z�8 �8laU��:0�TL�s"��	lc���#�6A@v�!Y��x΃q����a|Fp�v�c=���	���]�������:��֫����e60��_�B�S���f\l�i��%�]��H�q��0љ.`<����l���q(����ŵ$��l_<�'�o�������L�B��"���V
?��{�b,=��oɩ�7�� ��'����X7C	���U�O��\�D+�;5��b��ƅĤ�&a߳ǅv�߼
�f&W.o��8�<��#��bR�z�,/ֻEo�O�:�*~sc��[��*=���3��lM������~-QL�V�OJ��.��xl�l��B>�� �Y}�R��.�cǯ��z�:԰B	�$�� ��`4*O4���a"=9 ���O�G�L����Ì-2Yޖ6�%��d=��XK@h1�~�*��{�,O�o����i���G�����<j��+�$\���A�> ���q�}X�:�xF�_/��>����>[Ռ����wǿ��q��z3��pG���-�bVJB0\��vx͍ʲ-�Ve.�SW4�)f�w��}�oأ�[Tykrt[��{�U���R-�8$:��F��w�d���r��ZT��h�A��t�ֹ y�1�˂��g�4���8~<�[G�Xʌj�Kc����C�b9��^e	u�iN�a8�$�Y%b�T"e�6I���B`�+��I�P͛����?�ؚe�4����U
�W'�]xI5іS�
��k�'ƈc��r¥�@��Qe�W<��%��%;(˼?������5��2;��[jl&��k���]:��I��\dn1�=��09^�W���_Q/f�;ɧ�y�E�5��fPPƷ,Uv�|zZ
�	WG��m�f�	�e�݂�bf��ڣ;�7�r[l�]#�8D-�H���CK��<�`�#�|��}�9�S�M7��<F�d��@�6�)+ ��9'*�{[%}� �|��}��7��`ݐ�6	ٛ���s�������������GD�9��!A�����,�Y�c�w��ςw�̪��G}I�n���|0�>0��8�AɅ>q�fQ=�I��[]�0�He�"�)t��C�:3*8>�����k���L���c��դ�6G�]��-��(�g��M\י"'�&^Oů�HV�n��=eu�=�WY��/,A�5����.��""m����дK��A���m!޳������OT�C���P0(q��O|��Z�@3�A
]yz��zU�<y��a_gkX�����2�/ �U�����?�r-�'���� 5��µ~�m���݉���l�F�J3��x����,A�<dK<���Ɣ�o,-69��A��4�E1�G�I�&)��x>!�3�En0��a��c#����"*K�~)}P��R�5 U�-��C���'<Ɗ�YB��P�`ڋ�������U��pD0ye#+	6��l�F�t��'�2綰!6	8|�_A�c B����h�j�`;�P����A[zz��<��O��S�!�S�5��v���.�V�ζ^	`;�@��o�Ӂ+yM"?�~��H��,'>B|
yx5??1��̘}�()��u='
'T��l&�~�mռ.E��{d��7��U�V7�!m���5ʜQ�1䍨Άr�(	tt���W�Q���R$����Cz��#$k^�Ǟu�lC�_��F��A�^�=�� tvC�j�"�Zs���2hk[�q��HF]�~N3/P�����;�_�a5�� ۓ)�r�FxT�,��{qf[����h}���,�KYgqK$x:���CA����ڛXu"y-������HS�t�i���8�N�b�L	 )C�0�K�mX��@�[x��b�*�Y��L���S����j^-�gr�U��Н�i�t����O��<�-aO�T�RaW���+�"��gD���0�[i�����lvOL���$�&��y��T6�5b�[`莗SgSY\A{+��1���֎�n�˚�E��rUY�d"0�������Zv��il^��0qG׆�����ܕD��X�C���D�n|�&�Ӕ찣p�u�Cڡ�ӳ�{���҅�Hĥ�eu����<m[>��:+X�#!����@ob��%_<g�����8jG��KÎ�+qh[�ޘy���[/�ӱ׋��ʜ����a`	v�87����5����'횲�I��]lt��}揦c�N�^2.��q���P"d
�_#[������g�֊���2_-T��ĕX�ԋ&�sHA��A&l �������s
�B�V Pi���&S���6ؐk(�L�	���M>�p�BtN�9�źjJ�\����}�͔.��D�Y�iN-	=R�h��]e�|b�M����輂qb-��,����i�Ho:x�j���ˆS�
ֹz��f�j�t7��n4�p4��̼3I��f�>l�m�����a�Ia���|����#X6A����d��2�7�uB���9�w�K|�f5�:�=0N0�]
���2wc2|Ph>h��X~������<uG�0f
:\IUP��b���-��`8�T�y����|~��^ȉ��P�p��0�? �[g��rE�<��ෆ��1�k"4�u�[_�g���T6� ��#sh_r>��\����߼ʘ��
���ZYG��ue����Ց�j�a�b�ݮ���������5�lo��"N��P��o�������	c˰��.�܋�95�h��k؀�G�T>M��~꒵�>x����ʹQ�ܽN+��Wg ,dL/!����;&�5t��NN�y�u��#�>�,�k�w�j��۶�1� A���>�?����6} B}��cp���v��l�o3m&�!��X@�Ǒ�5p�ԣ:2"�ֹ�&O�g�R!�������ryߕ�-��bEc��B����:z	���/��p�	����P�s�P�����:�2�Cܨ�b�k�fI?�^�ۢ�Nm���@�0x!O&)ޜ^z.�H�#j?ݨ���_���h�+\��l�*��nd��ێ#̖����_/i�D�kC+��2E�}���*�<���]n�,V~0N:���- 3���|PROAY%��%���b<���{�B����"�)ڑ�A��ۃ�edzC-�ݣ�24%0�6vnM��IK�/��
ɋ`@�$�v\���Sg��#C. cW��S��7t��.����:u5�5��l���ZRV��G��q�ʫ-%8YNv��U�rj��sl=No_��R�d=Km��G�-[:4� �8����=�Z�'�LnC��(�Z�DB�V[+��s��K��c��Nzajm <J�{Ò�Q*�T�e5{��x�(3�qC:����T�����R��Օ�Y�g���>Q�ޚ#F�%JVR�<�f�:Ia_������;~`����+�n<o����-8�W&�/Ÿm��(����^O;��w� 	LDR�󡳪t�/�(p���}YږR?�}]�2�
X��J������\�u�c�4dZ�%���nbE��G�/��d}���2�;z��hH:5�<r.��[�� WH�����1j��~x�H=�h���&���������Z��|�����On
�� d�L#������/��\���1\��AF�pR �oh^l�����B�Y`g�gL �it�I��^�����ѳ���C��o����'S��V-�D���G<'c8�.��x	z��'�ޟnR�(��ۇOmr{F�51"��d� �|�>�S�;����U���	\����1k]�k��=.�\���\�Pk�K�5�ނ��wT��W��S��tݮ�h3�mHCm��;F�%_b(H)�ɩ>?!Gc���C����f��I�������5P��-����D�<��̈��4z:�⭘��Bo��g3�Wk.^ ;��#cQ�mU�=-RM �Ǥ���V�,�"�r�3���n3G��0�0f����N�e�+��%���8�|�oK��~d
ʾ*�����ϣԬ�Z�j�4�NhQ�e�o��7�1��cOU!�Umz ��>�`zN�,���0UO.���Q�r�_x2�$و�+=cz��߯�6���֍ �2�dX7����~�0I��t�9��x&�z���Մ+�u{J(Uo"kѾ$�9�������#�u����������b�I����{+0�O��l5C���Q[}�TɣXo#����i"�TF�0���B�HB���łN|�o�j!ʩ�f�D���u�Ɍ�y���Ł�)��1��m�p��J��Lc8�7da|L��TE;���-�3!�1!��uٙ�3���ll���Nb�M�荓tkwmؐJ� CÅ�h� _k��-��`���L���mPbQ�7s$槣;�=Td�i�|-P݂R����;>���s2v	���h ������/T!N�Z��/��0��R�M�N�vpp(�M_we.�<��M���/���E�
������@�2��dY�9�{"G�ENho�pCƎ�G�Bp��j��9��-,��F�h���h
[[�x�{��(_~�^�X h*��0� �}�s0K#$��? �ʩ�ç%6k?����f���dd�䆏u�nӬ�`������q�ؕ{SwsU�f�d̀�H*�fMa����32��P�*�iĀ�z�	{�����C���Ģ��35�e||�Yp�js�1�W�R�Qo�E��s;����"]�6"NэS?�}��@�6�6�z��@�L��S���z뫹L\,���$����n{�A�+ҙA�5tZ��3j�~�+Z>U�0����i�7�Ug����.�nf�	���W�h�v&����|�}"��.}.[����N��&���+�:H�)��Tʆd��&��W�{�;��o�<x��x�-3|2���֜#M�߼&�oF�9��8}\�����Y��tŊH�F�\߈U���=�tz�m~���Ô%0�8�V��q�|ZUpho'R���I����,�R�9��-׃��=� �|={�?M̻�6����DjP��3����$uJ�kl�	�%�ֶ���W^����qX̑O�l����?�I��q��,BS�������\�d����<-�<۳�l��v�����A����a℣m��N!H7��5z I�c���Kj�d�3J�>qh!�'2�H '� $As��%k^S%�����6�jG<EMA�e��B{����՘�m~ñ��IRB}p��ȓ:h��`V�h��~|��R��N5a�V-�����O�#�)���͍Zcܲ�4~ҮQ�A��M�ȼ�3k��>@�^�
�~�x@��襐����Q�KQ#{�K�'E����3ۃ��J*�R�H����bU�Jؼ�ְ����g�_�&�:MP��)T|;�&U�A���e�{x�3^�0߾T�"m&�"����٠�'o*�HB��On�`g��O�:i�(^-����kr�d������͒Iއ��;-�.��S9NA*�
(ɋEջ�9���!@/�A�T���r����oW�6$�X�%x_�E�H՚�`� �����X�����eeo*o�F�&��ʊ��8�;�3Y���2P;WW�h`�OIYDչۗM�I�����MN�B+ny�(����uȵ8�<(��Q\�)"�}R���g�{��d7�Ln�궗vb�p��ϖ:I��.4-��A���}`׬����z�9��&��M?�u���M��.�.����]�{v����*�;�L�4�����Yr^jne��V"H�q�Y��\_��!ڏ `iPq&I�W1oX�EF�>��aF���j���4\j����t��tW��>��^j��JO&�@t���ܯ�7����\j�ÖѺƿ������B�B �הOt/y�e(d�1e�
���՜�0�D#�Z@[�;Igx0l��D�� �0��|���`��\MJ�Z�:T	D�#�-�h�}pZ�~-�B�	��d��(S���>b�V�/������	���a>���MhNк.�,�M��u��[F�į[�	��7Ѽ�#ظ��[�igt�p=�:�m��� ��3�9"N������Wv�G������G��k�����~�l�O���!��oG�ij5���>r*�-�+�N@��%t�8f(y3_	���)4�5�{�b��R�jT��t����!�`�ʀӦͨD.��w�swj�nso�.X�A@�Yl�
�n�~R�1�Q7��kfH�"�o�����+g��7]�5��������-���z!�4�Ph3���q�l�0Q�z��;/8f��P��4\J= �.�Uc�o�<D����L|w�(�>&ip]j��J��N��4vӳ%x�$�+��F%���ފC��e��Z�Z�ur�c�˰�CJ����wA"2�1�������r^�i���\�vӁZ�al��B~۴����q��/�����1��|�B��W��#�*�J��f�������,���1�	Pdg�߻�c��9V���ĵ�ց;� ̟	�ĵ;��0�nV�t
Ĕ=��j��+�� <t
��=���h�Wyz,<��3&����m�|�z����/�s7"{Ǒ������,���5��d��������#(��`��'Y��4|�y��y[;ce�J��4�x
BrC�
X�oN��+֧vefa�Y�(!U��n�R���^�~\N��%�.-g���
O8j�Y���hk��y�5���5��6c�
��������P �P�Ɇ�#:v�uN�l�@6�����ͫ�Υ�{���?%� ܛ�m�F�:�_��kđڲ�c��8v��(|��}�֬��@�&�-D_=�z�!@`i� \���_����K5\���c�f��Q֚���0�r_\�<e�5��󔱵��"a�m��$�?!9۝Z$ X���b-���ˊ��7(]]�4XG�;�$�h7�y2�
�&��� ޜ��!CH���.2l��&c�|��L�GfIKd�#�P�	p��Tl�IJ�5F��OI�6Ύ�6��.nC^Ag�@�ո����M��"��v2p��4G��BD��Њ�QnA椭ɦn�>�<s �(�gd�	�x���Eם��������PE�T�f��pd.�Q
��4I�W`˞(]�&6ݞB���u����+�Ý�MbkcN�+!L�淪���!�sxTW��B�6'\T�
�\�s��#�-w(e~6�,{9��@���sbD�E;��f��M�R&vj�ЙsB��ת�O��l�Ɇ��J�fQc�2FKb�g��5@�n��j�.�hYґ�����������/�J�8cNg�<H?噒�+l������]��w�A�f��,�;,���=:���m�l}�af�p��v:%���fpd)3"��K��%�;W
R$"�v��S�d�kle�0��N��x3^"
J�'Ꜿ#�߰� �J����T�3�����ں'2���S[_��Ə����뒣�����ކ�bO�X��A� �?���p���w�U�BCb�����Ps�L���"C�
 ��K���^�0)��I���Q�F���q�U�	0�g���ӡT*�s�EO�!׎��	���2��4�*Vun�vALRA�xgef�.	�6��ye�2���-�Ƀ�ҌU}�'S[���'ų�}�o痫�b�C���Z��R��6�G��q{~ɰ����唻��U�Q|�d�/mF�d͠��'�0�>u�?'h0�:�Gn�Y���M��Ð���,����SMa����k7�jE9?����~�&����<��;���)���	^N	1ā*�6)��K�i����CGFr�-�cUԿ�<��A�E,(�6c���4c[�_�X��I�"ҢT�&�@s>����J��W|1�:��]T���h�ˉׯ �d��BBv�n�ȅ'�:�%���OO�87�?�]�q�������T��v���5 Ҿ��4
�i}��Y1����T�6-,�����!%�MD�Y��h��G���I��%*�	לrm$�cʻR���ޓ4�n��{������ht�>�;�j�� �)�3l�
J�A�Y1s�:�+��m;�wMdR7�w稏��Zp�4Ez۲5X��
��.�d���0GY�-�