��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|̪��q[�d�v�?�X$���C�O���s�#��\献l��ȸHm!�R�����<gʊ�O�W�}#�4I�����:�u�5���`���1)���V���͜]w���B��<�+S֮AN�G��J�8O�ER�����ɾ��gt�����z�O;��v39�3�f��L�f�d��\�Yy�"b���������ӿQ��s�3���&��m8��)��U�?�����܌|��n�`��>��3�9z���*@̫��C��)��Q����'�q����@8��ؚy��9<����vk�Q'�t���m�4 � ��r@^��Oc�*4��>t⏘�n̅�2�y�	��4���*ARĊ	�m��������p�Q/�2����L���\�����q�����u��ְ����&9��~����ޫ��t��Ɔ��C
�5uy> ��u9�����=u�J��%L,�3�"T�[͉� t����R��z�N��������¾�b
y�n����~����q��TpX�߾$y�炂��������'0TLiZU���O�Ԥ��G,٦g����.��`�Ѭ�1�]T�Ⱦ��%klQ��5�9�8�/��e�����1�*r���B#ր�Kx�`��m����
�0�٧��<6Ā�v�������Q����1�l.�^�����~@*� ;���ԅj��p�v㍑Y�G�]���g�>^��]�#��Kޕ(�M�n�z�������CZ�u,��	P��|�����
���]���d��bcl��S��r߿��/vi���w�)ش|ı?�n�?_[	�����i�\��Ѣ�`^�'�]
⬀G�5aW�_-��/Tem�f�M�y�;��DPv�o�s�u�>�23����U��?�v�]�CI�6=�����~ɞm��-U��!^(��i}��lM�cj��t����uX��BKkr-ss��S�9��{eD��U-�_�ܢU��~	v�i�I�X6+�����ִn�91S�������Y����7�����)\�<c~v��i\�t�����(��h]�<�,t�B�,�����~�T�l�?�<���1�Ȗ�J�#��Me%,��q��R�`N�^��<�t۩_M��.Ѱ��Mхl��0�����eo'��,t㤳1&Z�P���*�D0��`7:�h�p�7z����u�H�ۡ,nHg�{O'���Cw���h\���O5JG�Y�����%h��h;X.e���N��$��֑.�3�*Զش����"Z�8��Iʊ#���n HhV���L$��|�A���܊�\�T���?�q��óܧ�tb�����B����dk�X�Mvy�ь�:JY��*����� t���cPag�-h�ֆ�񺺫��^�;,.l!	Y���s��7J�`p��|�٦⿣�ł��T_�'���x��h���^�> Jg6	D��ie��\�������g��ݔ >%Z�F�t�c�/nr��p�f_Qӌֵ�� ���t�E�ky�<&���[�bDJ5h9]�@�.�U��	�F���� �\�M�4�nB�f�����h������N�%��豢a���B����"��P���!S#���N�e�^��A���UR�R�y��J|��U8��`��s[������I�̕�tln.wǤәj؆o��3/Z�$}�%Ӗ�(�DIW=.}�f��:=�gHU:�C�g�d6QTTR:̤a��Q�,؞��vg�uϑɫ��!��tg+,�����pXa���n�a�p�+�h~L�@��y6�j,�P���wL�1;ǘ��e6���1l9���zV�W���y�M�O8����aզՊ�^~��UB�]ǉ��'&K#���:+�<�j�{yZ��l�=��>���ï����T�o�H�R{�j�Ws�X���.��3I�b���sbD�R��㙉ի�@e�잗��V��#���"��S�y��w��$�<3��n��,E�x�\�ƚ
���5�W)	�d`�[�� P:���$��6V��fee_�T��xT}n��K`4b��((q�H�F�ʹ����7���?De����,]5���.��q:��*P���hҶO�(�Ζ?W\ኣ��0���LهD�Sv�4�����z���Y=ʈ�Md+\~Z^�j�^86�霜��</�����mPD1"�w`َ�9?e=d�ILR�ϰ\\��J�05��+�V&.%X���<���Jԁ|_��L�%�GBv�;�D�M���t��.�~gܺ%�,�D� �V%_��w3YMҘ�kx�6�wd��Gz���i��aA��}�LҠWv]!{�>L�Q��z��5_9TG&��wdB���R�r�{L7�k@��G?����jG�$�L�
��^[�\�lfe;6���S�z����*�Wu�1�h�R.]��Ow�Ei�.�2�͞ ޱ��t�k�n��O�쬭x���La� �r�[f"���G2�J�(�rV�f�SF�ˎud"|)3B4�8E�W��A�tKT����	�k\�R>��%K�r�������*6��
����%���o��,���j۰W�K�/�aۆ(���	�����'��Gr��O�;�9Mqq�=r�Q�	��J���,I�2�ў��7Nq�VC��^c񊦼��J�y�q����2 Q��2+��˭�3��V���� N��2�r
N�������G�k��k
�'|#Q�8�����oY��#찫N�KUԭ p��@@<+6�>򡵫���S3�P�V{�6ِ�/)�L��t[5I҄c��GƂR�FD�~&�/R�[�XG_Ix�RY��%���m�����خ��'{;U�������m�U�7�	VP������@����t)�0�pQ��.�{dyrD�Q!�*i"]�.a��h�R��8�9�J�����)��O�&ٕ��՝cN��
�dk�^���@�%�d7Nv�V�1�obt�����<aX.qP��w����'��[H3!R���g�R�-���s&�dW�g��N:rJG�e:H,m����٭�p�b+9wʙM�d�|?GS�"%�Y�ǭ���r��46#wf�-�*!1S�lU��@���}��"�6����<���	G����.g�����1 �ݏ�
��h���:]#�L���>T"#�z	\�,VDڄ��S/�r����^�O1��9&h>Z�ap�q�:俇�`��򽉉yT�����P�l�:��ǲ�����z�n���3�r�c�C"uN��<�Q��D~���}��f�]��\z0&k��@�EF����W���ȯN��o{�.c����u["D�3��D��]8ι�� ��� '{|&|p[��	���D�sL���K���Z�h[f� #���+w}AP"�g��Iܮ���@�,�!b�Ux��/���Ml8��%F�O�cm��{=~���=-��1K�ש/�����f�)E��U>���2�Ů���|:M7�Ϧ� ��k�D6n>�����jp'&�>�*'\ʄ�(�����9uD:���%�����u�>U�	hmM�� �������x�;�'�#��̚�f��t��FО���H͂���&KB��?+ĉHX۹�\�s6L��-��9�������h*�0�)��{� t9z|��3���~����[L�����/YzS"�.۴�z��T8�x��J�'9N��h�i�2�$u%���~��scu[B�zR#�(��d�ĥ��+A*�b�IvLd����6���!��E���_��㞼	?�RÜ����T��&ҌYZ�]x�ʪI_�v��x��>���g�R�X#����=��e� 
o\���-�����<Zp}�l��]zu�gt9Jn�k������yy����Mq�"�C˸�J��u�?����ڈ���j��:�A3 ��ݮCU�_�����y��z���'՛Ql1����ݭE���}�NndS�uV���X�S~�3���Ms�
*3�����|OVZ�Ko�����!���=Y�Ӌ�� �,�qch{�5r��F�HTdz-S���lJ����C�f�|A%h�z����:�
�� �r��Z�E7���B��ɳ�h�����"&�Au�(m�~�.E��E� 3�p�_���:`\�/l�H��0Fߍn�?ܖ�����K�y���1�i��Tl_�PCA9,��6�\I7/�E���T�R�Pq�~�{��-�k�����qB��	���-�\����+�����㒷1f��x6Ľ?+ �H>3�$�_��� �vi�N��\��݌��3hvV����V=cw<8h��Zw	���\O���ᄪ�e��=����6���O����7L�xV�ə��0
�)ߦ�*Î�i����@�@�t%��Uc	��{�U����=��Dho3/�����/�js�:���h̓z"����E�m��hS�5��N�	
������J�B�T(z�b�s��zt@#��GqЏ'D)����b���#�0עf�(i9k���uU�9W~É佇�ު$�\Wk��0d`���Le��)�}<�츩9`�-D>Yhn��Y��׽K`��eg驇-BP��+kl%���0����0��&d��觀pL��%�~t��;������+�[��m	�)X'��̮����4�Ăc��:��<�$-����u)dD�B2�뤔�}?���	y���w�+5ҟE�R�vS�E�����$�/5л�1وS��ђ���l��q-��Q򅰶٨v�H�RI镀��U�Q�@6��臆g��.�LD��{��\'�%��~����\����@�M
^��o3�c�����u�e�ST�_%�=>������[a�$h�!o�H�魑N\�x���b�L��)�VP���T@�`�|�@*��*-;OȊ�7�J�S�|��7ey�f�K�l6_or�`����-Q[I�_ˉ�9t��sD��޽�TX�L��r���/���{���B1����գx���F`�J�4	��#�\��k��m9ڱ�6�9���Z��.����A7��D
öq��U����'~_Af^ex�%�r�F0���	uI��_��m���e�Ax\�Y�n
[Cy\�ŭ�L�� 2�"4#����Wa���7� ���b��NP�P�:I8�v/�U'0��hn�G���B���&��
�#�.���x�E���p�%~�,�*.�6�:�����8��b�PE�ef��	L቗�ס�����(v��֨�9����˕�4e���<�?�e[5c����7zd>�eޙ]�$�������Br�%�H�����