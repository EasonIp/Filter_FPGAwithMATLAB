��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�&���ڴzk^�2�\����糿|!��g���!aXZ���s����?�.����
��NT.��}	?���-�$�a�G��m���E�E71hx^���x׏D���!���N�� ����H5*_X{����e�hCD�C�1�B�@g��3��;Z����z�Txr�LVr-_xL|��$
�7`U{�sn�uO#8W��%jt��*)-�-�^Q��S��x1�|������RU��N��q��nB����x  ��
4�N���]��7{Rͮ�|��[�&42����|���>�"`�;ӽ�U��;{�G��s�������.8ܜX�Е��dɯ�����ʃ�K����/���
kgb�W�wV��&��V9��n��2�YVڒR\c:s�-�hB���n��^R�Tf����˔I�ʷ⏔}S��V7�ߝ���c+v�olk�d�C1N�{e��w'��TE=�VэП&��n2.>I*��Amaۼe+�n�������?\]#���k?�w~��Lz�<H�*}Fb&f�sz��Gy�L��2�y߽>+��j̕/���M��57	�E��-�Fb*���Å �Q�ݬ�ս��Ҧ�֟�~����G~����Fh�0N�A$p _��^�������٪n*��{77�z�-��2�w��С�Z�Fw|"v8#T2YsJ�����֌2�6��I��\Jt���ʪ���;�C�;�1Y13	��)MB8BF���i!�Z�ԞN�� }1���9�SD�$$}���o��r�Ǻ*�U��p9��^�V�������P����n��0-���������@�o�ؘu�ڷ@�6$�O���Ə�aY)�1��۰�����?��ސ��u<��G	��|Z��F]N�J��O�X�<�c�� wn�8h�u���LՎ��RHK�R�ݓ�0u�,�i�8���cH�l���t1M�F��s�]'����N�(}�$i6�J�w�Vr�5�\VxK�\� ����^����
7�t�[��*ש���|'A��0����Ͽ᳕��;�� Uښ(/���X�V�tA.�	���X�1y���2�JOR����Ovhft;�ya�^����TK腹��@�|�t��!�7S��D~�$�f�{�B�V岔u�	'H�j�AD�b��rm|��k@fC�k��������O���LP���8����J�U��s3��`%�D�6[�������������up���wp�M �-V��7�Dry�ަU�2�t�s^�' $�.ZM`?	t�Ր��&�� ;�G=�8O�#�M���.���LT�m����d���Ue���A�r�?�����SzYc���[i>C9C��Y�$��.�5�����` 럭�9���u�)���� 2��Fà��R����m?��������JkM<���g��Fm��O���3y�&.1��@bTE�4����)���i��.z�cS�]+�R�b�(�r�Y��Ab|op��U��$G?"N��A�٩�"��T�
(b��\n�~�K�I6��V1v&$��U±��P���n�X�4��� �`73%�._f�B�Uw_vM�#��{��1S� �	T���2�Da�^�t@m �;!��z�&,��p[F�MU��C�<�G"��M@�H��o-I1{T��٬�����IY�S�t�1��}�d�fG �������W.���q�D{��Y��,���{�����Ul��a�ДsD�P��oxf�X� ����
�v��`g4����OlZ|��+�dH�b
XK�Վ*���_9B�ƴ_�~��u�t\71A��D#�6�]�ڟ;���֮1n˨3>�z��a��gϛ|i�Y}xkO�&���I���P(��6��}�xV��V��LS��"��ˎ���hH'�x�3��I���b% ���J (�Ӟbx|2��H��6	>P���}Lo�u��|�I�y6�]����eJV�h�I����+�,?x�#��lQk����w��cuQ��]��\�bv�8$5Grc�|��
��@"$O7w�J� �Q(/\P�2�ىہ+Bgp7O9����x�SZ��%i���l���ܐ�(��$�]��i�>P� ���O�S̮({��X8��fOP��$���wqE9��E��h�fYiA�ޢ��A<sq�^. �G��]���p�7�5����5��:�oCs��x�f��@T�hC��2C�s6Rl�+�O[]Ka��6�;�����)��Uu�-�ܠb����3?��N�@x��a~�_�nfEI�(2=L�
�OIB����HTeq��ƚ�l�����_�r�s�a�d���0�n�R������|�V�ϱAc�汢L�D�7� )B����'�N��>������/���:#":0�Ӝ���S��"�!���TK�W��,�q�m#�ej�;/͒f�.���kj�����1�Zc��?U��!#J�cuc��6����2h�-!bA��1ޘ!v��ݩ��q4�+s�!j���p>b�����Wj���w( �W���q½��|�|��3����/�ʃ��0x�ˬ������'�"s�/ǱJ��:M�4F���v�}�p�Ɣ��.�>��٩�y�X�"�9�� M���`˛��2�.\�+a<�;ȹ�˝�8�nZP��:%9�=󱞙i�O�G9��Ǜ��=V�����bM��I[hk��(N��8x�*���y�Ȕ�I�A�e;���9E7'���������bse����N�ɘ���T��Z�hWO�� f�X�0��lxIJu��W5rW"��~>[�w�?�u!�.�����f�mꕃ�j?�ΗH�A\���g	s�ߴ5$4��M5
r�Xۣ���ٽ�]���*"w_Xz��õ�Dr-����:߽�8j�fC/�����)20�A����J��L.�e�e V�����Q1G�dMl̏ *K�d{�0��X�g$#���x�ʺ�C��Z@�@��ށ���>:S�>`R�7v1�7�T3^}�wr�6}���=�%f��3W�B�f9@
qCV�*���鱙e�0���Q/A���_A�@�P�򠿖3�i����)(�a�k�4��y*Q.hO.��v����Q/ֶ����/ZOz�y&�=�ho�.�~/��FW>P'�Wg'����X�Km��H$G���eJt��|�]�2��.�ɬ�JK�?4�=_��-}�VC�M�e�8��M�@�2�ѤR��ŷpc�1�G} ���;�n@�=�|K�ӛ@�o�{r��j�:���r�^�b`�'�i�12�)za$��X�]&��m���W����{��5�Y��A�O��q%���k|�q�r��Ɵ�܄��ܡ%�Ω5 ��I�h�Ŧܽ�e8� ����P+A�:J!u�����{K��	��Zh�pO��W<���"q��v��O4w3H:�y1�ڜb�V�������j~�����Q j=h(�>� ^���'?� �e���D��c�R�J�ʅ ��pW�}]��c �;�k���yQKK��|���#K�}����@<�-H�����wA�A`x;)�h�����K�*�]_�j��A���vXD-�2P�\��U/x?$�7*�`~I�!���O����A�&��5"�T_�+���ћX�<�<G�h��R�H�΂�"���!�P����.f��;K����A��w�U�u�Go��=�܍>M���8��$32��ĩ�P��C��-#�5˨�I�-�1D2�;S[����Bq@i\*��k�ߴ$],?9���Qh����2��G���$R��jǲ�S�6�P��O&f<|�Q"0,�G���������)YoK����{��Pٕ�Hq\va�-	��Y�>�v��|�l�$�|��yڞf�a���R������Ca��+��+�l�.ߊ6%��ץ�'��Q�Kvf-̪��y*�>� T1�i�3Q�pm��߶��\r)3N6ע�$�����ְ ��d���k�L�$��*8���`����A�q���r�����|��(�4��i�1c2{����0�1cr�(�f��r�u7��|f |.��E2J	��ȴԹ�Aa�k��r��(��q�T����:�o`y9 ��4j�O�R�.�{�St�H���W0R�Y�9���P��h�j�a�\��d���3{�8��E-2��".������	I�
{�	qa���90}���~G"�J��.�Ra��H����ׄ�܈p��G8���	f�K����X��P��m^��)-���I�]�+U��Dn���G��ɑ�Z
�����g�R��Б�g��'F�T#�Q,3���k���$��	��@	C�|
@t�A�G�K�aM���:�����l����>��J$Z9�b�:�|j�+)v���b��M�^aИ�al�B-*�F��֒:�T(�/��:������߱��xDa���ژ���Ř�4"��F��<#HS�)�-I.��Y�v��B�_iv������EX%�6��c����/�k;R{y�:����L�3�9�����{����|��,���,'��=	>d���T����h�a��<����S�|ՠ7�}_a��qH/�VX!u�/��"�98aH�?��\���䙖N���v�r�y�$�rgLUf�W�ws���I(�9k,O�/2&	Iݳ���� vw�M����Qn�j-���L�׈<��ꮣ�[p���i-����(R��.��5�PÅ.�,I�R"bn�BV�yG�!���%���$"?�&��}�57כ2��[P߬P�ؿA�q��+��ܺ~�qT$Nv�.RISw!"[����S�JHֵ�#<����c!�)R�K��%n��Zz[�W�"!'��]ĉN��m�3� �����
�ӆ�:�;p3\{)��[絔U�{n��h��O���;`q%�>I]o�eԁ��?�1�Qc_l�F�O� ���i�RO�'�1+Ba
�i��6�K�w �(lᯅX26�i��@�u�Af���M�U<_`%u �o�Ql�T
B����
�4�IʃqX}&�nk��2'�&:*����_M��Gr\��ۙ���� ?�
��70_�>�:{j6���q��
�X�x�l�ɥH�����:���Z��Z� ����ӯ.���v��V�J/�.�",�~͈�K�2�do�W���xR��CY�0�e�뚐^����+gG�)�Nv]=�\��_6A�u��#���&~Z3���-
�4���p�6�i��:��C�:���LpY��K�%���Ao�~��0�v)����#������K����j�n��Js�3��L�����j�S	R��Aޫ�D%:'�GZI��$�h,���
���]Q&�.��~�F�r��ub��fO"��|墎���m�.��{�O`��}mvՕ�x�k���D7+^��2��^S�8��!�~���m����<�۶T���ߘN�z*2�����_���������b�$��в�@6��K��Vg���ջp:G*��C���N��!��(gEW�E��nlPw��d��dҴ�4�6�n�$Y�����7�@6��1&KA
 ]�9�n��d��$����o�i'�_#����y�{�f[|�P��`q��[��u2�FF�*~��� (�'�Y�����g)h�� �|��R������fGŐ�H���x#kg�@Z�ʥ�0�z�'�ē�S��_�M��ȯ+PxU/�	h�Aܜ�o��Ć
O35�4Q4Z���,W?*l�?\8����=ʸ���y7n�g9�-:oD�����<}r�S���������P��*X��C��R�:�A^!7��|�t��`����2M������S��dQ��׀oL�Nq��",�����W���H.ٺ����Z*Y�a���D{���?����0`)��m�X$�SK	����<���"t�ΰ\Kw�����4|�����w�t���c_�W���mq��_ޏ�-F���+]k	W�Y��?���Q��Wj��A���O1X��簹������2��@4<F`��qj�7d%�B�г��wK=tnX�����
�t�F5�S�{0��q�]r*�U��?(i�S��~�s姹������*����[�o	�*��n�apQv5�� ����Ϟ�!�W;�1 TW��ڴk�kB�A�A��5�������V�f�S���A����*N�;��Y��-#��T����\	���]�ڣ�\�	|�h_]{�;��Z}I�Nt������蔄zs�*_�%�(�)㊋��%B�~�e�˅��ziX