��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��I�ɖ�P�	��[�&�T�u�L �����wR�K����Ҽ��<�X�L.���[��"uq�`fm��\���t�u��Пwn��(�7R���o�M�q?���������p�6��s'��%!��ğd��B�yN��}��C�� ]�v]�'Ϡ��E��|6����r�R<��@�1�TZڊ���C��Y*��MNQ�j?�w}5\���F�Y5�Z�Ư�fR�VE��Z��{�Xr��^ȵ��v-3@6抵��b�7�&Ϸ�>�����o�<����![�F����d
%Z1'�c=�^��p1������6N�J���P��fK�Z���|gR���f�(���o0}+��b������'  ���B��@#K����+����5�|�2"��5�)�F�4T�O�U��?��*��tV�d��	3 �m������*����N��.�SOs�>@ם�R�B5�t�)����O�B^��Q^ֶͯ���P�%E�C�O=ё?�P\K�G��]�?:Jd\���r�;@?�lOզ���Ɛ�=�8�o��%��{�<�lւqYM,��K�(��9���� � ag��/��Rp�*	�T�-X�"�uZ��hw>y�?�&����@Y�)�D
c��)/�;���"�7��F@�`��!��.�9.���"'�R�jl�8�f���M�$Ԥ�n��J�6nը�wG�!0�0^w���6}�k���.e��&Mu��R��*&�{�0khތ�e�܀P����,<(ø��Hq�Rb!Uϯ�Oy���Wt��fۮrMNq�L�P��a(��)�A󛦻��:����6ZY���f�yētg��|��	:���Y�����A�g��d�5��Չ���:�V�¥֢�[UV����w=�4��[��@[��\[MH{@ew�/ ���[>QY��V���j����~E9d�[��:򊝅"rY"���ǅ�*�������rC�E����`�����&�=���K>���!���^�`TZ�g��(͆\Ƿʬ�ƬXzEB���P�ة�5S�Q`K�e_V�*D�a+-�Z*�V�}�� �[3W	�.׳�(�sBܕ���1��u��D_�/��JE�M4��0�ods
�фf��C�Q�Xl�~��-ҕgkI+��� ���zM�X�]�>�)�l0�ܷi�NŞjS�U�#qe���KV6g�ڰ���|����ԑH(J�M�ʪ��V���n�@�(a��L��ʧ�����������[�x�k���X�nMA!��E����i�xP�5��ܙ`�&KR���U�H�ʩ�=�*a�ʤ8�~N{�47��,�����ѐL��i����U����+��6�f]޻�= ��LҲ=���y3,3��'UL�HMx�el���%�pB�<��,�YV�	��6�<pD�w�ݢz*�聇�h��9}SvA�d�C��i!۫%�w9[��[%��_>���^��/AL����c�Q�����pH��L|*��FV��dc�ƏY|�%�v�$�~)��q���[N��W҇�X\
���J��H����F)�ǐ�IL��D
��
?6��:�q辝@�f�F 4h u8�� ��Y`ƾW*&����Ӥ�J�6t��@�IyH�l�L��$�֛3ŕu��b�:�!v�Hf��߇~��9��B�jf��4NL-�}�}5��_�b���������΅�P�^�:%�M*n����,d�o6���9�Z���۱�0�U���`E°��c�m˼{y���ö���NЍ���*k�X����ܯ���/w{cw�|s2S�k��×w��֊�K0�aG�q�7�w�Nt������c�|�D&{X��Ω5�oY���_�mY]��Vm�	�@������~�}�SXL��(p��?�S
�1F�D�g1t���8�ĺ`4���������K���-�k�����
ZO�,�ׇnH���TH-��z�o^�`dMѴdI7����7�z�!,yl;�pCF	�k�J�Hs�=�r���)�;�Dk{�+c-���ޞRm��C��1��)��|W{:7�x�d�"h�h�J{}����B��M�-���YI3yX�k�f����B2���6t�������
�`�7�I�"z�9����#���/=z�$�ϭ3 >�G�~�]�}���}��0�UE�-�e��͌�^���^�0���Ћ�a~���fEc�W��,���K�a��9`Dh��|�Auk7ֳ�{�0ۇ�a������Px�μ��A���&�%!�8v5~U⻪�������Gv���#��P��M=/��px��RT2.�w�8�9)p�C��d3���\5����>�hK~O~?��\'�=4e������gl�/Ҍ�����-��!����ɧ(��jU<O�!�}4Q�8As �'��7�g	g`.��_4�e5Ǜ�K��e���\	I�����D�/i�V��4K���BtUh:����m��vXȶ�x��)r��s��v�pG�S�eԉңm�wF�;P������Nf ���j�G�v�\%
����F_5��/��������Gރ��3���n�}�Yw=��J���3r �1T�KK�j�,��u�ٿ�?$h�U�O���+�q�3d��u��h��ߡ��UVD7u�ɷ``H
\�VaN���Ĝ�h��3n�Mk�Y_��ݧ ����7r�5��c��^����̐�\�!���tQ���ɹO?D�{8%3�X��%�0T[�C�)��������lf�R��5k��WF�����I���Z���x����`И�(k}�ĪQ�����{���~�ڪ��Mu/6�F����$�]@����M˘�t@ēX�Lr{�!�w��˯(F�U���Y�Gt0m�D&S�c�].i}o�s8O��{����wM2�#&��3G��ϛZ�tEs�vn��A( � �� i�]u�Xه7�9�/��0%t�/g���iܖb��S�U���d�s��zd�4��al����!	��3��%�*��ճ)�t�Դ[)N0%�H����W��t����̖�g9V���¼��˧V$�s�^sY�Nݹ��1�wm�}���eʜ�óu�*�~���f"ӢG��L��?w���<��o9���^c�E���u���S���r�l	z;�b���%:�d��QSr�{r�+_܊v����=�:�3���K�-��e���ń�V%�˥j���4K�Bp-�0�#�����$��w�Q?u�։r�N��OD����mc�=
�L����?��:D�L���ldhy��8��m�T�#�|X ~ă�����র���f=ǉ"vϵ�$��"f��!�d�!	8CG8ф��^�M�?�����>�9���a?�'ά�r\��ӭ^�5�Ŵ6L���AQM{ҦV����� ���OL'�e���A��{�[a��$%^�A�y\���F��*%�C�N�4�o�r(���pķ^`��L�/"��#�A�Q2���ƣ�y�~kVn`h�@{ X�ыeQ}�$�^&͔,7�.�S�s܋nk<`�j����%d����l��ʥ���<����Y>���5u�֑�"^C�g��Y�ή���Ӷj0�7GS���EQ6P�w�8_-��N͝��F�:��QL7�@�t~�����}����)Z
O����ܩ�H�&LS��iF}5�R���E �e����)וA�E�!��k�<���:���^�T^@p�j�{Eb�%{��#�]g+�0��