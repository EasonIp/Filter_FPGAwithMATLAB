��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$�ʡ��s`����_x%��J��f��Uz�"�a��������4�4�)S,�G͛�H������vw��o
�x���ڋ"�Js� �F�!��C��*W��QB�bWZ%�	���sQ�x� �+W�=@"6kqUv	� ,��/%�U�o\)�b�b:P�Uc�j�S�k���_/}�����)9B� "�o Cݓ��w%�W��Z��3���N:1~�h"}y �뷧������S��b�ɘ2��C.��z�S���ѧ")�~��:�W�6QYl��Q���ܖ�$�W�j����������t�L~wfF�e�@�F1�q���\Y�-��܋�b�h���d�2��$�^P]�zR:����ñ��*'*�����h
L���2���]�M�;r0�_�-�fQ5�G�PK�+}箹|�䀺&�j�V�pUK�E<jf���R��83�(��g�	vp�P�pE����opȮ�q�X ��b��U�v�\���4�3�t�`,�R�.@������^��t��+��S�ND�aDO[[)�J��0~���N+���b.U-|ao���ݶb-��h�{� �� 흔v�״���@a�����4eՇ���/��h��W]
�m���.5�"@��:o}�#��|�	���T_.E�@Ʌ�"���8v�[¥��S޵�9O<�^��	����H���)��R�:ҵ;�c��{[���$:u�l�3J��)v�~��2J�K�p�J�)+�-�s^eikƘ��Ո�,��+nk��$Pqs�XүR\�D��'�H��Np�EU� 	�'���c�9?�)B�
�JؐшCG�
��M^���Nm!mg�ˌ��?]3��<��x$���謜�2	\NO������
?�i�TV������i����V�$�� {��&hI5��
Jk����o������Ny�`���	�9�.�a8��L�4�vנ�P
%�.��[��Z1F��^�?!,�sW�fk��&%f6�Bkn�o
O��cG�Z����X:#���+^7C ��|ګ��lz��n����b�p��ފ�Զ *1����Z_d8�<��f����^�0Z������:ϴ�����nr�U�l6�)�ԟ� ���w�y����U��$�o�!��ZL$�E$�5������7]���Ԇ�{�e#��i���*�]���ǥ�M߁a��M��1j���$MPH�6Mz�N��� ���l�����1냉O�+��JK�����F�H��� �^��:�$��V�O�o�5}!���\��#�����y�a��3I�3�ޝX�;cKۅyt�a@Ѡ�z\� ��t%�q��C��e<��Tݻx*��s�4����;�3+�e0F�D>+�<e�^=��q��\K��|��Џ��d�G�?�#� R�Z1�HM��f���Pָ�3���xh�h�[x�v��D�o\
/��v�^��ih/�@���.P��xd�"7 �j�Q]~�\�^gO���u�ƻn���G:�\�;V��ǌ�7Y4�����Bg��:H��%\C�E��<�j���Z�P��DΦnZ�x�4`�M$b��J���4�OѺ��R�t��G�y^���5�@���N���WK2/NR�&��2�Z٭���氟�>����+���R���04DB�j��Nu�(�g�\�y��W��.�Q�l*�B����=��E���PlDEQ��
D�89�|��Pi���{ޮ�����G��O��)�G�oH ?4�x����":F�#Q����%����C��
�Β8ҷ������M'=ݨ�3�~�7ǒ�7z��1�#����}9/�g�.w�3�NXpH)������vY��5İ>aԥ�s=_2JC���Ǣo	3]c���0؝��:v#��Q�1���2Ҧ�k��KA�Rk��`�a�-�΀Yl�b�^�Z�R��^��"��6��s_���,�ɘ��I~c�{�F$�oA�sȵ#$gr� \H/�����xB��E9��b���tǓp��T�h��2��(�ʳ�[��,\�{�$g%Â߃�"�w����&�yk��}�8���@��"���/d?�vk��G�0���޽����&�S<;�g�s4ޥ+gvVg�J���o����CP�iՉV�J�^2�Ul�Kn�O��2</����Q�������07�L�*��J
�y���֊Ԅ�T�}zq3W���f���f5p@k)�qɟ5Jq�wxaX�� �n�;������Q˥��χ��S���H6z9}c�!�2E�4�t��j�_�Y�;4������cB���
P�iz��E�b��$�6%XFD��<�x����	�D4SsR��g���#2���|(&��@E��&�X�"�� ��H��z;�7uD	���o�lo&l�rA���I�f�
��^!Y���7���	��:��P8b�B���]ݓA�������D�͋PCC�/�[Q<4���Z�>�Ġ��;d�ar5J�U��hV>�������Cᾼ��zw ������"�R�q�6f����>�E����	������+%>�1�`���ЁY0�cv��0,���3�!�K����8�/@ ��@���P5�e�sO��fYLv�����8���"�R���>�W�����ټ}R�������
��D��טD6l؏�x;u��~Ξ$)�ֻ�q��*��vz�y=3j�{�5��wa��/�տC�G5��'�uʉ�6��9�� CHs�!�E6�<�k�_)�B�hB��n��+��Oi��eJbw�b#��!�7i� `95�X� }Ig��u90�3�{T�r&B�p���|�_5�h{�2sE;A��*����O/g'l�����"27�#�}I��	n_�*ԃ�-{�r6�D���Xb!�H��G	�ZAP+�t$Tf�����bi�4��A[�<�T~�!ҲH�/� ¼��\�ܐH�4(���k.wT=D�-o�X��R�q����זt@y~��ծ�o㥀�~}�{�%�����?*.�4�qK靊��z�\�����������3�k&u倡�>&��(W�D�I�&��V0���I��`6Ʃ�LS}?2�ĵ�ь��MAnw�V��H���=�2g1��h�Nq��q�O���R!i��K?����������W<L�Gb���R �e��h<8��+�3�5}��֖��'��#;�}�݈�!�O�*ۙ� KDF�f��$@y���5��̆�`��,p�f�6����P\��C����ۣ�,�ֹ�o6���άK}�K�s��>E%��{�����%�v=��� ��gr��h��.f��g~��*�y�}�.��%�I��J��(���[\]�����T���]yk~�O�%UG��U�"`�^A���2"\��p��f6|ݝΖ��5�г��[{ 3q�'���Hn�)�	Y �9Ȯ�^�V�NЖ�6�0���@�
xE1X,�Θ*U�T���8�ST.�6y���2�6�54Ј��Y;�ԫ�����=4����&�li�v0���F�����<�uwZ;�AAT��X��Z���B�O�Q�pGڭ�j7(d�M5oZzc���biC;��l�g�i�b����Ϡ�c���5|M�D��~�Nݑ����Z���>���5B�#�8���j�2�RΚx��Q>�<�O�y��h����~Ϝ����;x��{���C\�cH�<`VJ 7XR���{�����S���:_�EF�>�ߗy~o�����E�6cS�	@�Q��ñD��{�o�f_1�u��-�OL)[R|{�rkv�R�nd�~�쿮��*,Bl�:��+:#>�m���%���)�F��FQ7��i�(�0ͱ��:�`[\4��!`!��x���U���;cv���W���V+���z��**_�����T3�6r��>��D�v�8,�qu���ﱻ����	Љs~��9O�ȵ�BR�nʭێ]�O��'�֨a�V_��;�X��'5H�88U�5�E2���
`Lr�F ��~~8U���/��E^��
UL,D���<w����%lQ��J���Y3��l��*��+����vk J�ͧܨ/ü^uW[П�:�8A^r*��P݉c�������i~�����w�"ֽ\��Y���V�iʤ�D�潥lw(Γ.W=�������3���(@���!�""*�T��1��m7. ���r+J�����Ɠ~B�3�\�0�P��?���5�Ҹ�Ɋ��^﫳>>�$.�ݖHҺ@�S�Y�cOA"�H�\��@�j���L�?>���j�*�Xث:WE+��,
e�>'>HE
��o�(;�;ŗS:�ۻ�f��yW�(߬ێ�5��Ϗ����f���@u�T_N�}����8>!H@(��w*��?}���8��k%��[<��}��[�^4z�]�mF\x��OjX������%#d���\n��������فE/�w����Gv���L�C��63�*�F�y��|/����sufNįr`Q1F���U>��T�����$�fo7�)����!��V��M����2�W��%i��Aނ���
u��L���?mc�=��OL�?��I>ȳ��O$Q��C6��h��@O�M�R�.���R,=�^!c�Y���*��^��d�>�D��V����q�4�V�t�Y�o��m ��l��ǿOw����m
4Y��}I�/��u֐C9�?�?��t���p\c��`}�RWV��Fi;ِp�FY����+@'���ҋ��1f�9 �UѠ<۠��Q嵤�\���ݱZA����2qC�dCg.�l>�(�ۛ�pw唞��|��&�j���G,���ӽ�L:�<Đ��?� �[��m/=@�?��k~j,��  �Pv��~�! D��pj��ee��֓�ʠр?v^>Uָ��`��=�_ݚ#����O�8 �诣�K�c��)�����9����]H�lf_t܀�0��\mP��=#. �B��_�T��`�~�L? p���Ґ!�pFa���F&s�p<�&�iIb�_a��{F_
�i�iG�x�8�+n��%�a�F�)�k�OT���I�=]����h��|q��|D�CBM^�ú���i���}��6|�*m��G
�w"����1���	~"�[L���6�zWCb��p%���l���k:�S�����V̰����~H؁�f��{�hjn�7��=ԪcN�Ѓ�M[��:�8�k����0$���Y��Ml��C^��13�FCg�&{�
���m�#Ͼ�y�J*�15��EU�㭔^7�3G��z}�W��ɹyp���D�6�i�������d@�CB:N��%h��G��S�8���1sے���s�>�]�c܁���z����Oٌ����]�����A��q��å� G^�S�9F �;I����l�&Q^C�W� �4�b�\��V�{S9�^�J�O0m�P��Y�����6����X��e��ѭt�(so/,�E��<�iT�)�/K�!�e�aƓ��HU����t��y}����$��P��eD���w����r���E�hP��]����!V���պ�}�ig� �QY-xG���'�k�D�~ZQ1��ϸ�0�$��u�P�	`B������n�aZ��� �{�	)~{k���a�S�U�}a��=����L��1��ץ���^��͹�$z�Sc�&ޣDc��u��8��ˎ$��	�[�|���7@ӰD`��O�u|{7H@� ��L��$�V�#�zfO�?�o�U����I{�\�4-��	kh���RF�?�ߪ}��i@�1��J��@P�o����9w�
G X"�)������|��2�ӫj5h��ad��h�h.�����Q�?�n�Gz���?�p?�pbZO��M�/R��m�;�kt�5�TZ��yEds�̻�םiҬ[��p�`r�u�¨E@���bd�S��zc�G�v�9��dc���`$��d3?�kTN��Y�����:�Y�YO`š