��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�uwC�5�b ��ϴ�	+�
Ct� "�J~���z����<
�����'k�z��ߵ,d�.��Z�Ӝ��2�x$ҟdL��h��ʔf��#
����;�;m�ȋ��[F��E� &'{=u�3jg�b�)��LA�u/5{<	����oiܒC���&�'aV7������~^��ލI�e͍��;W���������R��DI7t��9��1�(�XS��+3�l�ɤ��{T[���L�l�vH��7�*���}I;nF���T��7v���4�9X��DﾚY��y���g��_�@�w�vY���0q��:�c���p�*'n��h��,�jC�3����2��3���v�.b��-��x.'z�mڶ�T*",+����H��;t|D%�c�?��2��^�&���R1R#+�� r�-�->�EYw������9�93��t���v#qf�//�&���@�"�֏hpAa
�����!4ޛř�z�|�rXU'Bd{��	n=7�Z�3#�*��X6�7�3��N���T4�� $Ai�91���I�,D ! CN������WA���@�NVX�W|���>�&M�:m�K��y��4�dz_�qY�c6 ����m�E����M~/rhٝx���k[���=�^XP3H��7��D���d\�-��?wg��&S_8�ee�l��؎n��B�y/���K���!�D-���R]9�� ���"e}8��5g삄��_�]z�$�����`����;�T�@�Rh�j^��ʍL����"V���`A���rP14^�sgˢ�U3�M�@���I�2�-�rp!�.!���g��Ǉ��H�*�}�(���R�&�b4����$�ػ�ɓ5���yΙ�����y�]��r��J=!h��pX�&2JxI�s�YB(��wo��f�a ���o~�t/U���Rⅽ�bE�L�t-^��!����2�x��ٽ5� ��
�F��7_���n2��O�vE���˺�XQ`�����?��l�JJ�n��cLh=��T��b�y�7csaɳ=7*�� -�K�Dy�M���� t]�ȅx�i��yI5�ޏ�
�4���#�<	�'�0�INf|�ʲ�¾���ķ�N�m� �?�V�!m��f5�=:ف���j�� De�̦�r�6)4`��̀�ӑ:�W1\c/��@T�"+; f��m٤-���6��(���0��d|]���~?Io�\��H�C�o٦�q�
��'�C��nn��j2\����� 4�WLL�T#r<:�m�_��b�?vL=>_�K���)�������]������2���@��2��2WB���^4�xk�p�W��/~M�۠y��KNŠ\��G2�}J����Q���$eF�y�s��*��3>�J�ltF`���xI~���<ʯCtg���2��,3�ӿ�l�p��_$��䍎������&�k2�^B���J���}�.P5�b��ɍ�c�>y��{�od�~F9j7��A`�KA��X
H_c.� �W���3�.'ݧ�|8*8"��,���j�k�i��Q�"v�z�q��O��Rm�6��M3���+c%'�&�{{(�)���7�|!��1msT�9��~���[| !V3����S�|*�y�o{9�,�E%ˣ枬"��׎��ĭ�.���<�~O8�����[��	���h5AC<^p�E?+ ��҆"�{�o���Q�����U�>E�{A&��`M�*��'Nn`e�;�y@�"R!B�kF�%
��~�7 n����M��8��N���sGjz|�����cs���Q�a#�E�H�������is�@�란���Or��� zd�9���xh����"Z_����G�Tp�$B�]�.{�}���%�=����/l�E��������+��e��vp��R�k3$�kE�$By�aH.�?�dn{����`���.x�sR�8B�5*ͬxE��pM�_��~t۵����}�>��z�M����3��6E�?m��Qo��Q��Cg��R�CGh�k��kr���/�5�]���b�b�m������$	�
�N��чύ�)�@X,�K�-�>�X�H��#j�8g��c��G�CDM)FP\W/��8.����O�gk<8��ꪒ�jYq�Kǆ�Z�a��#�ʁko���1��rD�O�{����i��@��<]�RVx�#;l]L���&̴���M	S��tU=�]���ȵM�P�Fc�d�,l������&>Ӣ��[����F����9
#6�1l�6�|�_Y�Yl)�����q�5p��|`�i�9�W��0w��-�Pm5����b"�m�x�c��k�	�O�������*6�S���A�`��aT��[�6�4~�eE�,��Ӽ:�zI+�[���D5v�ۼ�K_P�[�$P�5�r��qan�A��H"���C�}����@_x�C��ڂ³���!7	]S�T��n��TP��y�n���ms��|�y�rI��S��U��� ��b�o����Np6TG������ Β�_{�u�3ťO����aF=D,�E��G����-!6����w:��@��%�E��^��E5slD��PV00W~"�K��\��b��t�;��c4p@���d�]:1qA���cb7�U��a����#?(��f��G�[鑟I��K7sy�]��duw�~�S�E�i�U�WX|������q���"o��%Vv�
�s �W�+�� +m�m{J�h�&sj��r�D'�V�-20�q���9_�+�C�\}�#�z�-�`�qP�������5"!@��C������lݹ�g����V���)�v 5�{�[�����)Q����D����4?���GK8,k�n��K�6��5����T[E�-�F��/B���+���_�tX����\[c�Iɝ���h��xŔ����r7ou@��oX�?♁��8i�;�Nb���D.��f}7�A{���c�ށ˲����]��)��
S(cۦ��^MH.N[A��'���B�&'��ͅJd�u��b] ��.:�O��T�R����Q����u�VZ��,,�*ls=P��B��qn�=���ld����?Wܜ?�#����ɿ�K��U��/��1�&v�`�gmI�BH�/�7j�����У��1@�:6Ȭ��"�-������Q��Hk!�d��j��
�{����h�MKD��Y��T7��^�cϾ+�b���rn@-e��]���+K�A$$x@������2n���7��y�w�S����D�L�_��50�E3W�Y�,E��I�s�]E�`m0ld2S!Q�l�ёQ�D�֙����,�.\����a�I��!�>>*��_�9��ǥ!� �����`�[D��zu:۠X���<�m�.Z��  @�1��*1T��6��#[�D�poP�OYl�RҲ������Ը�I~9#Y	��a�6�೶�œ�����a�j���,l�N�5��9xY��+M`?'����Ԟ��û
&;%���ߑ�o����F J��L7�V)S#�&�dp��=)�h�F��(��F};�̽G(:��{���0w����M�
��=�0�1+9�}�N��tl1��ܑ��0p�a(�g{�OF2fb��a�=�'7���Ё5�צ��gA3b`L�4T7�_��i�!ѓ���rf�X�?��W�2z(�`p�����o��k76}�	��]�1��X�T%}r��^h�K=�\�M�W�.lE��,Z=�((>���3��a}�M������	�s���3̙�-���S��+B�R����^ �#�	��L�Z(�����Te����ww�,���B7�c�B9z�	6��J(��O�þ�o�^ �6�Ҕz�~�şR����Jʯ����K����˨���e��AGKAhhP0���?R�Y��rڶ��g�Dm;(��r���-��4�[Q�{W�"�9����E�T
P���P�9A��8���l�'��(�$ћ~�+��������+@̼���?]5��`Y�8��x�br���5���M51��)'�hcx\m!�	�5�B�jDi"#�=C�{��}�o];H�I���~�Ve�@�Rz�����U�_��L98ͫ���ܦڙ�I����mLB_��vՎ����گ��8-�����B�+dl�۬���[��J�Jek- �u8ػA���t�Z������:�xDC&�n�.�K�J��Ws��I���"Z����m���51���zgaC�7�:��av�J+����H6ǆR�@4�(���d��у��MS��|B}�sp-FZ�C6��]m&5��I[r�&�!�� �ޟ�M#4��b77<FG��D�N%p<�����9�me�A�����j��`����V͞2�i�~����ʾ��;H��pU����sx��w�p�N'B;�r[=��A�7[ق^��ڦ��<�DY��V� "X�Wo^z���E w�EP�-�mj��x�m�A
@����/�w���o�R�^x�}( �����*�P��7.E%���"&6�Ɣ���o�-��/��u���Ѳ���	�<�%s��@x��G�n�+-+�|���3Y�~&�"\��r?$�v7��2����x��i>CNG�Ƅ{n�-;�95L�?��>�i!SH�NN��o�@QE�
�;	t�����a������=Ʌ�Uh �d���ԤP�b@g���Ȑ���B����F�ۇҷB�����?�_�UmcۛM��W~�wcQ`�C`��wCli�����ˈW�&8\w- �02���Sb�oT�!��Ц3��a,|:4q�lc+uO߷F�U�&�\,8�BY@M��AR*���'✽~5Y��/�?s��Z�&H�ތ��#t�y%ԋ�.ٽ�u��
�Ua	YL���8H-�ǈ��+�NP0MSo� [z�$����rdҔ����K������8�cXgEf�g�d��-��}D�CԐ����n�#pP=� Q������"�x��4t����j����pIx���D]��]$����(fD��
�������`}P�n��8ݷ�M�"����r5��?�s8g���],�z����s�����y�ﳗ�C�:0�Ik���v���+G"t�a�!�!Yv~�6��O6���X*�V#��������E���h ��]��2�iBVV_�+�� �/�*������5�h�$v/�xm,������_^$���|҂ǜ����y8un����Ij�#�l����~+6Y~�n�@p!�+���N���\�N�,��	�K�)��S����$oо�x��w=�^�������F�������+T�У���7��`-���i��n�| hF`��� X3�D4%����f~+WF�$�x>�~���WDa#.���C?:�5�qV���#��B�yjI�W����b(G�Th�%Uu���5�]܄��J������9uc ӰTG�;���
m��Um��LxM�P��Q#Pt2myg���O��c�$w�/�U�^�`�{-�C���~��=-%�U']�j�K�<ꉊ�+f�Vr"�`[c����z:\�z�<c���� ��K�`�	�_����@O`����|�K��$�D�`�H���Ҷm3�P>��i�$r���
��&�u5zKt_�˸C��IM3�0�;�����)$�t��p�����b��н�߫��.�s��C����s��d�5Ƣ;���-G=�>��z�x'��M� (J���{KP�) V�`��K�����33R�j]Ӈ�Do��y�hI��Ű�U4��C�N��w"t�?Q��I�$*�5��>��5�l�:�S;��]:lQ<���b�o��:�c>��6��JzZ:�����:Jqk�� }�~t�J��?��Lȼ R��g����SN\ٶ������N���S������8Â���:�^(e�eZk�AsdI�9�N^Uv|�tJ/�ϱ��c%�Ȱe��J���o(�3���Q]~�{	�;em�u��M�K3y�S<?�޺�L�mG\�'��B�Q^�4�ι�_2��s��g��Ǭ�@뙹�zD��C��gs�n�a�h�P��{��Y�[{�f ����w�u�L���wp�Um[9B�ԥ��oc%���\ha�е��Y���]ވ��q�/�M-V��2K���H6�'���s�S�ۺ����EX�A=�xX؊rkˉۉ�|-�e�{�?I��&���ke�A�3�4u��W�W�xa1��=��e��j��YXn�Nx�/�����ѷ9�*f���q _�rOG8� ��w��\�NġS:#Iu�G9]~��Q	�H��LR�'��9�;/o�imrw�Z�����ZB�(<����;�(@��JIS��G��W
62,l���z�3�4��y�T�f�8�a�ɧz�h+ŕ T���M!�[f��w+��Tʢ���#j^Y`xUƋ�G���������~��-�QID%eׇ4����.q��������낺/*P�?n\���KP;	]�A�Q��!��(*��#�)�z���3s�AZ��c��;�^�R
~nH7/u�BP�O1NߔXӓ}$�6������htY v?5T��uE����v���<%ƒ�q�����2�ٚ��\sIf��뻟�4�rBn�S)V~���o���o�3��c눆	T[�^sچ�>�B��s�A�����	r�t��*� ��ӊ�5�Vr�>/zҏ	�*QkƝ\n5�?��O�"���d'��EY֨��Ǚ3��/!V!�����>�3h�sp����A�8�ӏPj\1ת�
ʈ�1z�S���s����6\��/^!���_Q^/
���Vj��'ׄ��:��i���Q�d���q�ެLJ��� &x����,z�z%��[1+��9rIy9-����BSy�d�UWoD�EO�ʱ�j�CR2��V�Ǉ�
e�p�b�\�Jf9��$7ȏ�ku����eI��#�og�6�O��#�Tմ9��	
hQ�Sȟ��gtn��=���ܴ����ǰH޾W�!��>5�
�H9y��h�3+���+"�w��l�Z��uG�4�HN��Qz��8Gd��sI+��	�9���r���xh+�ui��� �"���Q>u<g�.�m��,��T�̇ \�����=DT(��H��ɠ�"k/g2МݲB�Q���kMt��P��Y��<�EZl,��骞�X�`�.��� �cd�B����+��@'�q�7N�i�ڃ��_ ��ͭEG_�Ur�Qz�Gܤ�fUI�I_�c���)��"��5��H��0�#~��t)n��%%2p������	OA��!l�38=%�cm���1��|��O����,B���9:{�C�5g_m���v׌�`Uo9���{�2�e�|�)���ic��if��o��l�q'<J`9�X��!j�3Z�����2�<"r���9k_�~;+��x�c3Tvl�"��Ty���@%c�=�_�R��A����Ĳr ��-�޴}����;-����R3�hE/j
Gj:Lj����k�:e�y��#�'ygFuWJO���T-Fývh��ͅ� !���c5�Y�[���S��s�a��;z�zS�Z��Ea�����"���ӓ�䫗j�QFc��y��	 ���W��&^xm�+�o��}w|��`��n���A&�6nr�@����
��$������A��8F5M5�4�_����P%T�!m�5�^��8��4fȂ(������v�
�E9������K��5�г�p?x�t`ݾ��R�KVb7�+�j?��;\��	]��ǒ�H�X� x��XFNI<����3L���ò溪��0��CS��.7���"�～�n�U�B�ꯍe�U���C -!��-W��t"m1�/r���]s��Bܰf6�_��gF���K#�W��?x����3]Bƕ��۬�a�����6�JP? ��/h��B<����i�\w[�!Qܷ�4{`g2y M�#�pC̢p��b]�3ar�� |>�c0�:�/��~3hv���k1��.�c��W&���Ёqb`�p���K�ȹx$��|cg[�
�a���ֳZ	�ďl��E�� �4� �#0/��J3<�ϽQ����g��4yԥNC�db���	�0,���A�E ����N���Q��94�χ���+\QGbPY9O���-D^#	;�?1f:���KW"��aIS���WZC2;S2�
���~Q�4�'g�m;��k�\O���^�gl�9̮8`��0��b��Ԉ�;�}x8қ	��"��R�Pq��MQ����5�&������-+�Da���l�}��z��P*�QEE'8�G�RB͜�Wd}/fk\�8YY�_Z�H6�h�}�)U�"��o����t,gx8 ,�F,�"g��U6o wR����EH�
ן��f�@٬9�wcllw�1��_�m����~W�wZ@zrq�ٽ��Q�&(r�W���Ya�b���C}�xSi�E�*
�@�H�:a1��2(�\{����=�I�-9q�:������=e�Z"�l�g��#�C_n��ζ/�����%�洺�/{���%�IU�D�0��j�.Ope}�F-�.�K���hB�o��o��X���G?$áj3���R;��~{Y
���Gk_xq�@���Ԕ�߃ݦ� ���:�A>$�L"g�˗�Ĩ�pdl�>1�G�X�}e���U~~�q��Cq�\��K�"+@�Y)�>q���Z�i^�����s����F� DG��"&4��V��;�
�Ŋ���NQO�'����:��%�m�Y��ĵlō�<�~�Bn�]�1�[��_������?�?�Z��v������gP��`B8�ѫ,(T6�ߺ"4��0'3^�hj
9S6����(���?�dʥ4��G�j�m�c�p�����5:]W�ygg�K�kґ��f�6��C�QoiBh� ��&������!ޢ�n�Z��䂬��z�-����|��Cƭ�s�Jg�PR�MK)+"�`��62a��g 	���X�s�t��o�%q�t� ��-a]�����/�,���̻�2��Լml��4Sg.��z��.���߼G��W�b��õ�;��h�6��9��SE���;čEȡ1z`*�Gv=[`*#�X������Oٴ(������X���i��떨2�4�F�>X�۩Ü��(ZA|#�4�"�Hagp��p��e�ў=����l�K@�|W#�"���P,=U���N�8\�q\��_1�yݏcW3%7g]�U7��o�V��kO��f���xD��P�H�][��K2�M���=��R,F(�^��b�T�,�ꆏ��|Y��4w@��_�'흁t�:S|Iy��T O��Q�g��7���9�0ƌ����U��*�UU��s��x��K��O�S�<2�\\j}�p�>�kCoXz�'�,�R��C��i������W��!t0���(J�ߏ�V
hjs5��#�_���!�7��A����9��>�9�T@N�!��B�t��`�^5�5��A�	��{%���`�>����@f�4p�@����Ou��C�\��j�����v3Ȧ���P�� !����$�X5�y� �~Y�=��z���~1�;f�
���q�#�q��\<,�e���V�g�!����t�(b�o�G�qw�ϱ��Z��#����$M "c4�nrCIH�Ln�0��{k+��za��7��(��:yy��$l�V�ݞ*�W��V��"�ӧg1�
)�tQ��]��O%�*lk���@�`¸�r5c���WC�^���mW����×'�oϏ�_Y㪃$��0�r�p}IL&���}|b�C��W~�%��~����iR�f5�_�`Ӝ����D��?��&��,��cz�N#^T`h�$u�'_�San� *�w�˝s�n v9;-~�=�>��iK`ָ���\�~�G�vP�_L/\I)Ͳ/��d��Hz�������oF3n�鬊GlI1rV�@f�J:4��!7�+��,u|��%u�5a����|I�BvNqМ�]�(ҹ���^�쁤]�c"�$��5�b�vg�)�(�1�)�+~:���4WT;���0磌<��`��s�i�2`+��~,������j2W$�ϮcgL�ئ�I��j=�`.���q�$>�4�㩥��Pv�*�zރ���$��`�mq��"�?V�Ңʺ��h6-x�>��������U�F����k��R?�L���� ���YƇa��`@;���E+�����=�m���� �I�84n���mn�8�yb�0;z �
GTK�]b�9&�H�]����;�$,��Yt�U�9��TO����l�������@���H�G�nb#�c��c������#J(�b�!�b�Z��"��P_��[� Y�^p��C`0	�@��~3b���r���m���Ɣp�[�X,_�C��a��E�ZB���]�7�7�{��IHRo�pj�1�{`%g�
'%��<�S��Z��ڲ�5*_Q�q���&5��­�N��?d��7"�|��Ss�O�������Dl�Koa�����h�K-n.�a��H�9l��_�Ϥ����z�L�P �{�.����x�F�wuL(G4̫��H����b�GH#3J�
�*5T��Nv!9�=�WVI���b���ቦ��N�+V7bjܯ�?C���-��}/M�\�hD�����6߻��\|��
��O�,~LXvP��
��������68ڍi�����~J4���tĬ@��"/��1	5,�D�&��6�:�.����Q����]�ӓ<��Qn��%��x��2os���b�� fp�{m|�ӫ�Z���Mq3��������E!Ӑ%lMM�2���v�na��s��s�j*���Y?K�*���oz�2'�U�-�kC��{T���O�wm{BL���b�1�r��!�},�%�z�����#����lKԆ�:w.1�ģ��=�$P5>܃[|4���JzC��<�7�`Hb���k\���%�S�_a��X��W��d�h����l1�l�B���Y��QJIo\W�Q�g��C���a�r�&BkN=�7� az�+�]�91�=W�(N���s�B�j�0��t˨��t%o�dut�^�����Y���|��F*�
;���M<⺛�h'�;=s�',TIG������8�2��:މ�[qS�G�JB��N$i2ݱ�沐�j[Z't�a���}\ח�K<�~%z(L�ΌOL5�@a�tҗ���&,��-�����n�����9>�ct%p����W�O�z�Fd��VU#���`6�/.J��
7���Z^V�<��T
��(~�8d"4���K=�ˎZ��̭�J�e.鬨W7%g��D]��e�lm����t�Y���u=��Y�-~�|vD����ە+ޤU$��]�f,<�g$M&���;�
e:��=m3d+Ҥ�LӾ[�����{�Jk7�����dR2�7$|���@uU�(c��c���������Ji�G�{�j�%�L�؃}�'�礖�b��"_�leE>�e��(�����)�R��&�m9�f9�[��8��O������m��/�f����uR��#����\�Z�|�1%�˻.�>~̠�M�N�M��f���_�_#]�T���x�U�}��=��*��di���؛�^�����b�55�v��E�Q��-j���rq�3#�V� ^� �WAX�_���1(�f��yCV���faK����F��>ۋGm�c>G�=��j��g@+����F�to��#����a7blV�a%�})Ҕ6�ϡ�vT��S��d��> �P����vN�϶�`čX|G'��v��,.��~z�s�R�]{�#]�� s�,\r
b�x��B����+ �%&$�5dV��"A��UD�����E��֙�h\-:�5'��B�!1_)$�_�����r���J����購5if�L��P/� }PDc�s/�8z���«�T✥�q���jq�x��w�Vkd̓)�_��_�qB˿01d��O���~���B�����F�yP��\������_�@�*!h��P��B��p���,���/ߨɰy|(����r�zx��n�,���3e�WT"�k�z��~� �$�x/�� a|�%Y�䗴���.�U�s�ӡ���Id>�Q�����W�k�e(�������.P.%\�j�=��
ej�7.hq�05v�V�T�y�%�����7���h�ͱ2!"9��a�l�qs��|��PC�+Au$,�����&�/Y�@kq��y�� ��#�0�����8W�A"m/X��g(�w���� 	QH^�?�qN�������T�#�7�I�H+��@�gw;��F�t�N9֖��3����<f'.�Q�y��98,��?G��N>��V^�z�/{��_��	v��s�s8�Mz)m�i&�3��9�6!�~m�3@�� �=�
Y���]^iC+"7�ʬ��/,[������ V1����3��64e�ȯ �+��:U�YSw#1� ��~���a�|ܖ�,��}:�~�g�����WQ��9�ڬe��h~+5$���JL/� ��I�p�x��}����1Ҍ�p"��8d6~W�oS���u[�Rv�!��k�Jo��8��@��6��3yO|.xr=rSJ�k��-��:HK��G�����_�\|X��c&��T�}���@/
]K��KAXlGj�l���E@��v3����<�{�`δ�ulT�gA��I�C}���ㆥ�b��v�p0�D^əb�"e�oN�q�WJ�尚������r���Mpt������S4h��k(!��&��Ȟu������۷�]�Cp��������,4���2I�����l�[��ʾe���0��Ư	�M]Y�����e�ɺ�g�5w�\�����8'> Uc���䶤'I�^B*�oܓ����S��6�B7�ze��W��BA�8�v��I��S��s�
"����r�q�q���'�/Iܳy�-���o�
��ar�J�Cg�:>��\�l�P��B΁�b�4���E�O\�0���eEp�¢&!O�3V���p&�'i"�
G����B`��	?;&'��9O������#VEO�����*��3��R��TL�|ź �(�㍐�Xvś��=%�z�
f��ЎM6�i����\%PV�&'P�+�qz$��.�&L�Z���e�K�pQ�9�X_V拦�W�)�`���5���o�!�%�-t��=���	З�׽ l����g����-�X�˸8����׊��<
|����A�~�!�A�9��A�0�������r.Ʌ�������Q����@���^*�{B�\)�)2���/��z��	p����*��������eX����X̜�w�e�v ���~�*��K~:б�mu���oJ��,�gp+-0����<�'�H$+�Ǥ�L��Bd1��)ۢ���J6���\�f�Vd1Nȶ��� ��SZJ�&����wv������&tz�%���󩦫�<�z�	��ݎ�!�G%�%8Ti�Yq�TgDV0
I�%SqH�? �7Z4V��r6L�[Y�r�NZ@�6#�{9��[�SL%`j�F5��N�o߸�"�(��'�5ne�+������8�/�~~��m�G]�#���	�#��88�?�N�n��?Eq`VT�<�B�|���bz5�	_<#�9���5�"���@:���\*�Q�ܝy9��n��{8�s��cV�t٧E��\O~��Y��q�9y��-�گ���a��� CJ�@�md���f��A�⋣ĳבR��;�J�F�,w!A@��>ܑ�8��:D�a's���#��3�m��Ǧ3���ܳYR�����ڎ&��yC�u4Jq%'$������:<��䲑o��w��ӗ��c�E���Aʒ\�-Y��ų���s��Q�0څ4}����������l~�� ���*Ʉ��;������Y�^ҳ"�ī��~��vy���10'�[}����׵������c[���՝ҏALFÛ�?��3~>�B�b�I�ea��ԿA@�6�rt.�SVo� �-?)�,��V��DN��>,2�X3 �q��"���b���q!�MŪ�ke�m��D�ǂ�)w��u��Z٦�:�Jv�~Z���D��IAw8�<�F��f�1_�C�c+PBp�v�1y[`N�_l;ٜ�e'���^�����]ƥs����K ���u<��Ü��h��;�')�6����k�=�#�T�	<��n4.�#�8F���r0�4C��p0�KK醊���[� �G�T�-a��]��♝+i�%_�O���@ٯ�X>܆m�ᗅ  �?��_�A��e�^V�m��d�����7�;w�b��ʑF������@��/���ڜ��LqF$�Lr�Lsxőq�����;��=�:����h֟5�[o�46->�v�Ő"��|�{X%�ƌ�4������|~�LC׼Nc��U~�@u���>$�LCh3F� �+H7��-s
�+H��x��ٱzk���Q��@1���=I�����G~���Y��;��O�%f�V@�)Ȕ~@W�B?ȵ��H����f���A��r+j�&u��2G�I'=�2�i�ۜ�,��כ��!!���R�`.h��B��l�ssa�����,Y��B�Z�y"+��C��a���zkFJ$�A�5W���o�"��0F�`�B��kp[m����h2��j���~�P��/�x��(�,��S�����AV	N��*zlZOA�p(\Rt"��,
�Hb�s$�x������a�@(mqY�|�q�tB�ow�e��X�W��1���r���5=�4��]�_��MF�I����޵�1����J"M<Td�e�E�T������6����9VX�G�uW�֛��r9.�p��)�������D0=,�ޜ��@����*�XN�3���͏�Um��	I�@c]2Ul��<���F7xx\ǔ�9��l�r �-�����䏚�h�GAU��H.�"��Z��+��T�f W�+���em���p��i���:�%�?��Pk*U?2����.�Sw1�h#�"��d��y��B@���Z�M�ھ��LNd���Wܧ�.Ɋ-I��F���-O����3���T��\����@�����_��~����b�q��)r�����0Na�C�GL6���y����Y�>͈�i��M�g]�}�)�g
�F��� ��y��P1��'؝��{Ж��&�,�g}g����߲���Ҭ H����>�gvSktV��S-i��cR�ݗ?A�e�3B��_�W�g�'�%y��Ɖ{o�]ʷ�W309��s���zr�%(�8��Ж�C�u�u.�3�'�8#�_;EBw�o�b��l�&ͦx�YX��pk0��G2��zشjjweJ�1�dQ=��M�<J2�3^��!���������P�ѓqB6���^�h�`���8��鮠���q��/�	����O9�@/yng�U?pt�U����!�\fd�[R�S0��5c��/b��IY�����e/H�&hd�q4U��!��6R��z���q�e}��UH7L�t�H�r�=��;n4{Jbz3�%�ؽEa���x>��8B������������Wp��r��H�b@|��~Y�60�?X�a�6�ˣ�/��4�r�t� G�m�ƄR�H���`�R�ڂ�T^���)�eN�bi��n�L�� ��(	DGCz��K� �S=peb�uBt�����,�[ńě�
�*+���4p�� �$�S���B�L}t#��g^���������0��YZ�8f�����H?Eo@R�h�S|�@Gv$�DYj��� ���b��^�jvpȓ*w�;�ʨ$h�����l���9�;��&]�gs~�3��1(Is��?y}�k�."���Հ+暘��B�[�Q�?�'�\�ۚP�����Apr�fn�ڂ��#�3��D^�iGQ��
w&�{�2�:���_cI��+���뢴~�I���� �{!b{��$Z��T-�Ǔ3� ��2����<�����=��S�*����M� ��Y2Kd�N@Y���~��|2|u���˰7�Pj���G�%f�~��UZ3�
�`�6 ��ζO�#)xЬ�_�զz下8���9�aC�G�+EKw�<�Nw���`�z���qrR�?%*�b��Y�û5�������X%����2���C/��+�T�ud��1U�_���y0������L�zϏS�1��a�SߑuN�s�[�>�W�X5���_�hS������R�ߎ��ݰ>Y�_Tk��Y
�S	�FI�j����׃�P@:�zx��C��,�n�|���bӥ�F�INK���F�釄fC��H��?^�&�Q�xR�Ȑ�n���(�'IX��QP<�E�d�D�v9W�h���E)(,J	#�P��]��u�T;��B;�m�s�v��@�m�`5\��M8�7���_������X��Pe�%��4�7�{�{�3����W4�/ �y��y��zm�n`��1�䐐U'�jf���#�!zpU�m��9�5�wl�V�8ӗ1̕]�>����G)}�����&GQ�0�Cd+4��`Gw�ӻ#��B}�� n���I�Ƣ}rF���&�</t^�b�mO"���n�z�䎣K�*?��D�!OD�Wzְ�ҁH �ܱV�|#@X���D�s�!$Tp3��/�D��W�h�_���s�p�j�:�C���̶Nd�[�/��R����iA3 Z��V����M�xf�7$��il��Bh�'�g�ޡ[\����I0�T�-��o��c�}�;�  �P�1^�����$�r���{Sv�^������=�����2�XF��l��Y����O7H�]��� �~H���D���u-�2�+�7�E]����{y���]��Y�PCN��e2�bIϭ��U�kv<[�]�N�ST���qkO�m���0ŧ�3^A�,8׺Dg�g�Q���dV��`�x�$Xvb7��lpC��鈧_�ϟv
���D��b���I9ί���>�C)���k�N$�;��3 {�v��e�n�F���X�U�t
	���H*Z�o~d$��qW97m���;Y)?��03(��}�H?�ܒO%�l���j}R�m�N�����`�ծ9�����'$mx�ҙ�ED�ZiL�2�[Ԙ�K��׷���@).nt���[R|ĥ�V�YGp���'��+U����$ےp�*����	�{~}9�X�a�$��)}�Q�#"��N�� Ϳse����V���a��R�&N���Rw���X֬:B�Ŧ+��mb�m&�
{=� 5�t��+��ļ�GnC�6f���ب�ĺ��n�5��rcsL����
�㗡��xf=])%�QQ�$��U�q9gw.DǼ�aQ	{��$.�N��۰r%������0��6��ky��'�U��m�G+]����@��?���?]�"p`Gy����8��S�H����ה+۱���$Y,ʕ��Ɠ�oXkQ��p(���6TO��E� �}uJN����o=I�2;p��ڶ��/x���朣i�0�~��$B�9�(R F�CN��jͥ�`o����@̢�F��;k⛕蚇`����g`��4%��3����v*\�&G�r&�_G�Y._�ɟUm:����Bc�5�iD:���g=�0)�Q��s�����b��ï���i`������vr�om��v��y���^�'�-n�����ق'K�i�yk�6^�OXf�H+4{���UK�A��*x�H\_H6?�_�j�K�=��r<~S����[n� )��n���nx�#����ء~][�g��(��_0~��grA]`%j�=��<[¯��D�	��	�Q��5۫?��ŧ�=1[	�^PsN�@:�v�!�x��} �����d'9;�QF�9��e�@���f~)�q�����(��î���ŝH�Q�
�]��, ��|HQ�Sj+�_���@2d�[;�}0Y���ZꎴeZl`��Mb���m#���1A��΃��k��m2T]B�W �$I�o�[��N)4Q�KM�߰��%�ܹ��-
,/S݇�Sc>�Ш���D*h}]��D)O4xV�^h�қZL=�y�A�fHL���?�
V�M����3�Zy��W S���9y�EmkG�q˸ޯ+���p�������'�y��N2��u�j;���"��^P��5�9�'�d�#P6G��^�����l_������n�l�	X6<��9�Ls�El��x�_W�����P�3G����v�o�����u�%@-&ML�,n�B����'3ѧ0U�l�&$TW���Ȗ\q���w��@�e�U���J��sG��;��!&�@Ǻ!W�4��l�,Q�����H�=�g*ݨ�{	^ĸ��Ʊ}`ܪ+wB�8;�)YG+U>����en�����/����.��9�F"�3"�0�"ù�&�k�-QM���"���*��Ž�^T%g!��'�Zճ^�.��C{\���-[9�RhK���sX!U��륈��X�|�x��Y]_���	�CfsCـۖ(��.��ˊ[����~��>�8Ĵ�C�Q���J��aO�̼�ߓ5��!l�M��H�.%!s�67�Ǽ`�7k�� ��~n�bX^׍��1S�����4]f=0b�zt��?F�UY�yeaʈ�2�\CtF��E�l$stT`0�3x�P�a��HJ�Bh8tq�Ȗf3���(/\����%�҅�����e�؝^c�s��]ܦvG&A���j�ƾj��f����K{�FV�pJ)������ڬ�S��n�kTT�)�I^��2Y�riE��1
���/�ǀ���c�V����0Ъ��jY�f�)e{�`Z_}�)�^H}��iG�B�k"LE�Κ:�_*�����]�9W�i�b��b�Ah��	�x�р�KUV�JN�ću��e'����b�x����ȬY��Wn{F�h�a� �۞�0��b���h�������2\�C�����0��&U{�n�m<R�������:��O�3���웹�)�W����С2���^Z�.%�7�fDE�OЄ����zRc0���b��E[�SA�ǶJ~�eOp�Mq-�k�U�Z��<���u������I�vaK�+��] }-��qV��0���=&ޫ/uBE��(�E C�!f%�S ��13�m��h� �J����W	\�7���|��'8J��@0����"W
�����ظ�3��b�T{�x�<����ɍ����U
 �����	 VP�4t|@5�]Di	��}NH���R�3�s�`X$n
��}�@�XF�E�̘v���(3� ���+̐��P_Jh�/�#��^�
��N�L�l ���xo�#�����<?#`�4�\�#��MA՜�K�=�/=�6se]D~��~��Iu��껯c�}��(J�����I:�6�ƣ�q�w��Q[g�&�s�l������:)�������8�������#{)$s�6���~t�(g/��ֲ=</����?ap�}닯l�y�H�P$?Vq��o�7�Q�Uor|ӥ�$& �c]0`{�w�iz^r�2a��t�$���M#ΚV4�Yԅ�E�*V>,�������f'��8��,��ڜ2Q61�3j�I���o-�����C \m$��o~��0�Z�Ochb�0L	����|e��tMO�g>�s��ϟ^Q���E��1YT���C<S�wD�Գd��b}��	���?
�P7�}����%?|t�]d�e�:Cr���-��j���3���;���z�7������ɿ���=��_����y��z8ZEn�>o����h%�˵�_���|DSR�vy���W���۾R�f����R�I����F�%U�3!������ٱR"*����7#�<��r���N�e�*�8ە�GZ��9��D��qy���zxݷ���r��1q���4P>tC�\ ��f�<[�vSA�3T%z�5o�M�C����[#�s_�|d�$@ykx���x���>��]"N"�2�[5�T�0�nh�^��#�m�Ǵ��!'�'SwFd	�t�t��Scr���1�.��3֪����W@�a�k�?P��^T�CuΘ-U�G��������K=sv�,��$|i���ھ���D��_yJ[���h���)#�E��Y7���88n�Ty!HIE{֘v59�NL��@��H��3M-У:W�]�#o��AS�kN#��H�a}������lEZ{~�vm����w�R�=�kc):�Û�֛W;�٭6����}T��2��������g��Ƚ*�����������mef�٫i�]eُ���63]���4w��W����:w=�~��AU�	�k�Zk�)jjc��x��].�{z��Ƿ�	*"XC@t���}\���FNA�:��/7/U|N]�+=l+7hy�^��� � r�9�i�~%,
�Ւ&�̟0K �R�| ��gi݊�gpʏH����(��W�$���;��Q�rR3�s���z���I���&�l��M�����=�]��̼�U�X��@5g�R����t��#đf�m`��@�pv��_Η�\�6X`��O�/�m5���[6�.L8��*� �1��+��6Fb���7	��i���#�M����i��F�4��#cE�[����?1 _̷�q�c�O~>�����d'nE�'�j(uN��]����9�}��>NZ��V��y����M�3��bg�l�5hC�����#2�t�wZ�B�y��]�/Ʀߨ[7��JdI�2������|\$S��ƩH�܏��^�՘NG Q<9����
���X�`�xk�-�C3�<�V�'�M�A
�
� yjK����O°(��}��#�\�T�a˒R�c C{hsʧ�ޥޑms��M�6�g�?I ���/'$�!�R�6��N>�0�+�)<۹�1��9��4�-אǬ�\��b4�?��7!.�ߪ�L��������Y��hZ��� PԨ��ʵ�:ા�kB�<]���l�G�e�r��NV�P��҅&/wE��ZxŢ��5�e�AYH��>�3pY���M�h^���'T /��y��ˇ�Q���B9�������u���_�)�o��\�7m����4�`��tۜ��.��<N�9S�������ܷ�Ա&���0�ڒLt��)w&�H�o�����̛tp��5��H���xϠ��76z�>a���2u��}0���Y,��`4}��nΧ7?Sv�t�h�aÑ&�m��'lB\5�A�ǡ����Y�鶅x��)8-���]��G��7��Q?
a�T�計\�g3}�-4�M�U�X�6ŕ3��{A��9n�.TE� fY6�^���U+��I�Y'ͦ�B�;�nHG2��b�%�{����5�dq&(�Q�k��uƷ��.�#���@�䨬����	2��>���(1}K��5�1u�#l�oC�ﴒ s�Z�P
�z���|Ԫi�󭮺�o,�M�� ����l��I���'g��E�ץ{�<��[�I-����K:/3���-�'F�4��va�������}r��?���j7��Q�`}�S��h���R�st��D2cӻ~�-�V��-4ޛ���Ͱ�ǟ8i�״����	�%�{竍��X�9����u���"��H,\J"��gkC��jZ{�@h��&0�v�Y��?>�g������P��K��:0��f vey@�GxG��~m��e���t�֯n�^�Ld�/bP�Q�$"ҙe%����.��)6�'T$St�S���i��;Pi	׸�tO�_��V�e��H-Ÿ��h�h�D��c�H��d�5��(�J���Q�ٹ�aj�aB��Jn�l�e!ߺ?���������
��^rZ?/�KWv��RA�Cg������{��ı�64-�#-��殁�)�!�W���X�*���Mm� ��0,d'��p��{9��W#���V���ta���𕒃&�8e��G�+�7x]X�����r�)h	��+�s�"�X3G�QzP�j����5d�?��D���Z�1����Ł�>,w�pc�~�����e�%�H��=f��Sɮ�͎�_��N����	�D3��䎝_�}�J����v{��H�/���v�LXp���Q|����q#�$�����n�+H �u���z��dJ��i�E�*f'�@LT]ȯ�� �|�>#}���g�!U��a*=��VO|.n6Q-�!�p"tW@MB�<|�t(3��wk"H&F����Qk��zY�������� ������Դ�3�Qm�&�,�ˬF� 3��R ��M��4P�b�@�J�j�P��~M��QY�=�nww����y��H��=�˙����=��t�����j�T�db�o8�Ⱥ$m��kl{lA�p8;f����G��n�ML���F�.TC͓�B�����蟙��V�D��B�E.��O)z5�Q掁��L���ѕf�!��Ʀ��ydn�;Y_���\� *��9�C,$	�,�C_����V�������6bؿ�ZC,J�US�VB	�"����ǽZ���i�$�6ib(���g�l�ҵ~���>�1>G~��͕�̄"�N� �D��C���j(�G҅+���5q��qP F�bч�Ѡ
mB�k�]�W.���Nbq#���L��>��G�뷭��*2d����A�E!o������C)�ee_)Q���ox�z` v�K���t���k'i��Ǣ���ё���!@����qS�wޱJhPxj�W��W1��u�X�I�(�8t�����KG,/w�5�Ye���B�k\ᆪEb}d�K7mc���B��C�I���ف�B�ι�z����G	��x�����T`�m�6^���uC�+��L!:6sF�;[���
���t�Zp�JJ�p�ϛ$%�5�5[ ��v/��mD��]c.�'Z��B��,�����C����6��Ji�e,�rR�pXK�V��^"��wy,_��a
�ۻ�Y����껧Wل�>����-MȘ�gӋ�b�����/���0ƭ�0�b���}��qQ��!� ���e~��޶G!��.�5�Ps�`@� E/���t'��G��	r'c���N2�g�۶�d�����r,?��N9_:����'u~��|y��;��E�#�k���iS�O�C/R��#���Z�E��B��^�8�1q�`�T!��R��@2R��C�lG��
˟M�2�Is� h�VD�E�nĚ,��s7X󱓼9@�w�����	�o���
�R���Z�^�����N���~���P]����n>��uF٥= �kv��I�v=D����&9#��2n�*���#�'�/т�4�3w����Z���V��ю����T�Z|��N{�P����e�,>��;��$��S��|�D	K������!���'qY|`ja40��J�	��7(%�����M􄗩�����߇_j{�e�'�.�a�����e^u���l�Ǒap�/��Ba��v^����WO�
ιX�G!Cu�i�W����F��}�G�O�����(�����@x?l���zJ���>8W�׬����݉5�f��U>����r��8��=��xO=X.0�]�l2[�{Ͳ�3
��.�r	�w�HT�{�wf���T����<��h Pw�~y��L�]�I�1����z�i�r��/J�h�#�#ǯ�y(��яp)B7�m���{w��z'P�t;HXm���r^�N��͎���0��cJdl}n �eR�>*�ᕏ�3������/�����US!$kþ��%�d<IGh�6Y,��}����X ���ĥ�%⦔�OZ��윙%ez���US+Ώ���`L��@?�Nñbmպ?���.y����x���Ų�������v�J\	�I��@e��3s0.���H�$Ks�*ǲ���6�M{�EC�2�zW/!t���v�tuG�Sy�"���5>����>��z�b-;<r��)oU�[�'>!�Z�=����RǑ.Bub�z�b����H�)�Oy��ۿ]kI�t'�PQU� +��d���'����j�V�M	y/蟹m�v�7�h8�'�[�-�r�1ϣ�-voK�����;\�&ql�F��}^�F�z(�мp#�����{��ZDy����65�`�;g�L�!���-a�����j�ZL>�}�+0}U� l
@
�+�m���\�u&���/�`>G�Hi����z��.L?�;+�����._��ai��/����}�ɋ�AT��ߏ3�*7�^��7v�h7��]��<�����M.Q7�.��Y�xfz�Rhߢ�$R;�QF&'A15I�%�Nh��:�����&H5�0����.�-��|K$={��z�WH�JtM ��_�!PB�J�uj9/|���5-RCqCUZg��B,���-��aS�8D�'�
�Zp����<�C����ݡ�����O��V�n�b3���_���%@*�l�Yx{��T.Z�~��{%Gz�� ޢz|�*\CJ��#�X�ܽ��a�gi�
���Ҿ*�5�0`W����]�c������K�R�Ԛ(�A��e�8��2jC*o{�a
��r6�e��UXЈ],�����l�_��/6��L"��E�R�N�-Pq7�Lͩ�����_¼b�<=�x��jf�]�w'P��(4�otg�� ��xf���RUmIbm��#� ���M��k�g���W�ߢ���i�Q�lU[~E��H���v:kE���f��Izm�nǮQ�l	��
f���G�vB�g��c%%G4��)?�@e�	�D���� z�;�����_$�?PG��@�́,�A�W��`[��iӜ�V ��=
/�lλ�:���e>"�N7���r]�� ��`��������ѡ�h'u01N͚c����6�3�D+�K+QT�Y듷_}�Ģ=_?AFR~hOREFE����p�B�6Q����0������_��D;6�f��Р����}Z��&ΈL�^��(kzQ�^��K�#���~�A� <��%��P�˿NY9|Ō^����ѭ3��ѲH:m{j� `�銄$fG�ÞW�D?���R��Jo�b����(uᨑh=�H�3�*C:X�؏1�����XdD�g��)wk׭��ͯޚ���.pG��=�vX���yNC������6�Wb6�m�Ɍ�5#�R�q%W��;��E�}��~a�G��Ǯ�5j��+G�U��k6

�W��e�ܔq�z�"��H�c��7�ڮ�������A��:"?&�o��~�tzV������q�7E�$�ަ�T�M��Ҿ��V�>�%�X��:[�~�'6T�p�>�E|����J�����-l��ݚ{�!�}n+�tzF��0mAtt.c�]���=��9��˱u�Ċ�0�5�ӑ�v�X*��b��M���
�	���?T�˅����W�-���7N��I�p<m=ez�Q��%��1I4\�|����<�9���>��C�х��cȢ`}5��k���9��A<[��]"��=+Ek�9Z�fܴZ˂�L�IY��jW��b��N�ȑ�wPh������jE
�((��<��[�4{�M�c��"h(S���� j����ǌg�٦ �O;*I�h7"&$pT٥V��#_����qY��l_YC��1{(�� vaA��o��^�`��+�<�>�m�GFn z�rS�.����E��Y�\�u�c��vv�9�f��"�~���l1�t�L�F��?+4�@��veVa�`��0?�d�\�Po�:fB���M�8{�Jp�2�O�Æ��2��Q����1tP�/�Ah$�2�[�
 ��=<<�ӹ�ôa��:�'��N�\��I�{�s�3�+@�N��Oz/罴�2*
P��P7-�"*wd����l��"�=D'�ۮ�+Ux�:t��� �����f�y��F��.'���$��-H�^���FeAo�i_mq@��E���!)`/e<7��*\/(`�ހ"�xk#k��:�7l^�S���cf�0�jV���Cx�t�.���������:�R�w��ʯ�##?L���I���eѴn������Ce����R3IΊ}NI��9��� �%��dW��o!5�e�1��t�DVS�K����n��9g��ܩ�{h���A�K� �f��$mW_Q��I��Z���߈,�3@,�	��P-&�5X\i�X�Tm8��/�k�����d��K����O����:�m��:?uOK2f��	8"�o`����Y�ܾa>{b�	 �YF�i˓��� }R1-מ�S'7��?��W�r&Ъ�O������?����F+�Tf3#[�q1H@�g�'nx@"��R(z�E�l�\?^gm�LQ;aQa��'Z���|�v7�.�U91K�ɒ]C?�i��ng<�Dw����������6��u�e�����烎9�ܮ'�j�nF�ќ����%��Q<Q��²o��T�ogV:���#��}�G�����)���di���#K"]�Y:��A�6���&�KI�Ģ�\|n��*�^��K/��-�6m[p?�t�4�t_�$V��)(�\ e�DX���2���H��g����Jc��6�tҤ�!yoc�+�֓�՜ xU��"�>��@MQkH8�H�ӣ>��*�G�6!@5���*-�-Жí9F�<��XO�bDl���F�3�eK_xV/\ayBx������Yb�?��N][���aƖ,P��N�m�'�)�M��P=�8�4�~� 5�5������|+��Clί.��]M�U#�1ع���P(�� >�/�� G�y���-��\���r���$-]��?F���35e�C�B����:
�FVU[ԸY�ܴ� ������ɦ�	�$w�*u��w&�9���Xu>����O�[�����.h�/n��$��'hX.a�:�D	k�jjC9�� p�DC8�����ZU�Pjhv�-��}`=�R�g������v�[oc(�x��R�g�5g���U��6e>\r8C
���N�|Z7��{\�>4D#�c5���yf�Ez�!�m�	gZ�x��c���a�N��y��t�&�z�
_+P��R�h���g�=�u7���[�O��܃#a��4?�C]�ڶm05ѠP��z�ڑ�J
X�Z �Q�_���"�=-�^�M���{�}��+�(&������s�1q@l��� �g7����y#u�Ą��Ű���{�4��uJQx�%$�V�yHo����'��co1{yUz���!r�Ǝ�e�m�vDOTJ˫�V�C5�a�6�b^.�� V������Ƴ�7$�ĳh����?UKj-����M��Drs�y�<H�ʶ�~.�Gq���i�s�K4�Uϲ��~Wn���XvB��nԶoNxV��G{C�n7�����X�����S��i�$t�E���;����B>&)7��v3_=��
p����?m����:K��߂�.��w��.Q)k>��G��O�<VPi�w��n�ˀ�n[�$|;(S�u���Vo�B6���k�ԽJ)�r����v�q`<B�����k���E��dM��i�1�~��r���ԪL1��^1M�x���d��г�����;B+�0 c|y���ąM�o0���H¾�Y��q�?��MW,2�:ej����)��>q�3}��i�)\�2K�j34�&���5�=�9-�-W=����k7"{1b2I�F��ko3��J�i`�H� ��MĪrf�Y0�ow�I��vY��SmSd��E�|�eEX�$M~�ت���yJ�T��\�H�ڨ�;���?��L��&P.�#u\�����ں��m���3kJ��w�S��ލ'�!|p��dJl�5�wW�A
#�~��� )c�W�8	+��;�R$i�S&�e^�<Z Nu������E�����W`Z��V���E����?��e��9~l�e��Đ���w�%[��K?��e)T\̇I|)��`p�gޞTBЭ���619bM �B K�.����H8����^����^a�VS˛�Y(�É�8�6�noUz���허!~��3���Qh��aU�ӓ����|(�qa����Ow_̮��������eq�Z�f�Ky��0�����l���_�)n%�j��
o�(fT7o���鸆ׅ-���	Vs�w�{t!g5?1<)�� ��c�ޅ��{�!����Wg�y�5ݨ�C�cތ��e5�Am�`S� ;�Kc�*�Ê�@��Ѧp� ��\�򎀀~�E���S9���- �%��3&��χ/5t�t9�ͤ'mdˤO+�K^]"��p�݂�g���+��)ǁ��X�q��9�m�k���x�p��j�]�;t�(��Ҁ]�]D�%Q���$ �+���E�&��������{����4���/v�$nf�2��u�����a�����W����V������m��5Ĺ�!�K����o	�������F��h�@�JgCC�Ю���� ��$�i�����dAOFr=�I5ŮE�~�fZC����Ά��q���P�o�z6T�M\��s�r���\k±�̺�B�S����;�(h�-����w`V��>���w�*M@����\�
�X�����ѯ0����CE�P �#p9B&�>R�����)[��4�WvU��6#&�{k�|��|��d5�d,�YV�����b�{���q_d�׼�Rt��Z=3��ͼ��b�����Vp{�t�g����I�ѩa�)ꗛ'��bN#FQ>W[�bkM��q�A|K�[��]Ţ��s���5���_9~�|��OG��o�7UV�̉�- �!3�����I�q��Giޜ�
��vwc���f����j�h©�)I���y9�42����T>�mP�f7���+iϴ$�˕�b��q?���d�EGW�k���v���$?��d<V_�8S�j�&��R��LP&�y�����Gp<y�Nщ:��xx�Qu��w�#b��{�庅j���%��}�� M�	�tv�F}�	�ʥńܮ����h��r'�j#WT�Ys1���.���
��R�I�̓�����Ru�u�?���r�����E�۾a"\Ɍ�~1�խ`G���WGÃ��z(�G��2;�4�	pf���:c��_��z����K���:�ﬓ������ �OZ s�Y5���Oj@��Zl~�6�4R���r~��Q��O<%���SfS�<�|;F�m^p买��q�k'�慪�X�^�/���:���.��
sq���o���[��6��˘��>5�A��c"��ڏ��f���Ea�u�a���"y���\��c�%�
�O�Lfa���Tf��5�Q�V>�/�q̓�j��p��e�̉[?�& ���@^Y`���z����ϡ��7� �r(c^�����h���� �Vv��5�#�1�A�Ύ:/F���"KΜ-2Nü�8���)3*�����-�Q������8s,A���0N�P��~s��L�o�)j�)4����"���j[8b�!��ܵzչ6�S�,%'��E#簔�)���)�"i��c�=s����B��y�+O�JD[dġ71�&Lz��Ǽ�)�X�4f��*�.���������E6ߒQ��c�>������# ���k��(M&�{ �fV��6� ���jm �KS�)��*\]��ܠ�������6�F�[:��)m�%KP�������PŶ�l"9���G�����$-Ʒ��qdz��s<5�]!����6��ꪯ�"%�j-T�5�~����x`�S���K��k��23�;��pї��p�E�ɸj���-�S_�c�����mJ�P��:�=G�`2E��X��n��$��+�炑{FFl;̉ö�F�_�g��b��ns\�֌'� ��LtoK��UI�n������w�,�@�_���X`MS(��>��؎m��8��G�d�ӣ�\�l�&j��{D}�t��/ņ����  �u�R�n�9�΄:lP��Oz+� �������׺�x_��`t��=&̶�	�X6�8���Gl��xͿ�������K�!*��#9���a�������@=4�	�e����[��M��K'�7��17�e	��ru��P�C�O�.��e�V�^�測j �t�����.��	K��yEE���N�_��Ɲ�����s	����VC��h����uD^�4���=H*~��"��
T��XYቡG�V�D��j� �H>�?mG؜��Ů������Kn���*���M'��>Ѿ��W4_���3��os2�<"���d܈:;*Uͣk���[l�PX^?]J��o��4��� l�u8��$�K�y�/��Inṗ�p<���3�+�<��x�������ш�a�,<Q�P�����{q��g�O�>��	��[�i�-�I�Ǣ�5�)Sx�)r/&�#��}#؊��@�2Y���m��!F�D�0�����ѵ$C�A炭	|�0I^\55�J������;���e����c]�,���I=hf�c=Ws���ၘ	���CĒ���h��*jѳ���ϭ��o��ĝ}D��*@`���=΃t�ja�=�S������%JR#IϡZ�Л^�<�P%��ʅ@>���w�������
.N����c���F���w�>��F?�7���d]�3�;�q��0�ȱx�S�>�3g��ZN����Z%%m��6We3s2S%&+P�٠��]�I�h\��I�_�eó�i�|�u�B&�� �8����%��9m}��ްQ+!��ߜP���-�dS�S�<1JS�9�l[��Kg,��BEn�akuu�\��\p��5�<�M��.�HJ7P'��"9j�y;W��J��-b͋��!W�U�l�e����w�{8��)�B�-V����%E���ڙ��t����[��3�Y��T[����8
47Vk�~��"�}��AB���Ti�!v�!�qf�e+[6��W��W���Ny`�-�Ƶ�Yq������R,���ך.ɖ�A���U��
�enwE}c�\���;.�9�����V�5���#�x"�eG�{��9y��(�,*�����$7��귌yצD�/��x~8)v���;mt���P�Ev!�@=����;�3�4�K��)���7�s��|����O��nk��چjȓٻ���x�@��l
�H�0��C��9����[+2�٘Iiy���1e�Le�3�q��]�Z�K�Q��z-鄿�
�߾�y u����:���YR�P��[F�>MH!�4�@%?W�f�I O�Zv��#���@o�R.���o^���x��ϜuS@h�*@��Ě�=�/JRYQ�d�M�ʐ�,�QVnfUߔ`=����N�1h�����H;Ǡ'����]`��4���n�ɮ\M�6�ȫ�	h`��f^��E*�~��>,E��Xʶ��[�*굢���T�8+��P��E�ad�t��r�����Y�z�n��X���9>�-�j�
nr�����D��� %���+�� "���~�4eMX���`6���g����ܑ��C�s	���m;9ji�6����~�h���{����D74�;����ڄ���ڀi�"�O綛M�{
�P~
�Cj& e��M+�W��L���a�F3n�#���0�|�[D0����:7D�Ϻ��z�F�4�W������j�נK6Oho�?DIv���q� �u[�Ĳ��^E�YgRͰ'�r�G^�)��*ο�4���3�n��ba�0��A�Y!#W�K#��g�#<OV��>����c�hl���P�Xj�f�5�;�j�\gգ��O9�#�:�����q��I%ocK�(�Pj�RagK�{oP��_ �}�Ҋ���*ݱ�L�DI.PA���%��v�~/�(]%?�N�K1�&����#��x���"VF̡{�Xw#b��EЮ5�������!�]�}1���Y�/L�$U�� �cH���70�I�v��S)�^g�\Y�*���W��0��f-�y7�m9pyKa�$�����Mu-I�!��f	a	�����H�:h��pa� ��S�%�x�$�4@|yO�mt�Z���qF�p����4�M"�뎙8�'�Trv<���#�&%`����/>�S*&H��cn(僇�����ksc�>�KR$��{ix��l@i���P�e �� 8�m�� ���7ρ&�k�T��\�����58�b�b��p)S��A��Ӹ��k�<-������5s"Q��F�Q��a��w�E�3�qcb3����lpg���S�x�I�/�d�D�"�]6n�"��n��s�7W:�Ɍ��������(�.i
��r?�^�$��Y^�ﶈ=��1��{'r�ct9)��nn?]��3�T�B�s��W	g꼫~k���[c��.�T��U,B��%Z	\vz3��fc>(���3Yּ�hs�������锷�O�k�-�)r�D!�$�U�	���1H���/E�.Ic����q�#��N����G��ٰ}d��U�BH�����_o�})��U?��P����y�k����@��Nsi��u�:�0wh�/Hx�8�A��8��>�Kk��)���(� ˷�}b`��B��8�T�ls�,��_��;d�*���X��=M��m�P2f�6u�KGs��P��2C�������t. Q ?,&龤���W�(zN�X��_j�Μ9�1���Xw��h3C�3�\��zi�/Mjx\!�?��e��Ou�
���V�(\b3z��O2x�o���]8f
�����{:�i�e�B�i7�]z����- ]�ylD~w����Zљ-�'��t�𱂱�^�8���_`H�3�*��8	�@�����.!�6XL��Ƽ��T�Q�R��,+�/c��0�k��O�4�3�:L�.��6�,�IDC����ܩ�"�>�q��ћWn��@,W��^���Xn6rp��7,��|�n��$�^�1ğ���Ϣe�\�%��hF����H���ݸ�9=�uY1�`��e���}Rl�8�~�#oA��s�F)��9��2Ν��t]ʭ����2�@6��I��1�;g��G�
��]p3��x}�uB��ɰ򤈊G>Y��X�t�/�S��T�X��S��H"���Њ�V�vSk)C�56JmU�d>9<�IY��
)��vS�jnB�l)��s
���xDXMR�X^�I��*)��Y����(���[��KH
�ֱ���#�hh�MM!;�/5q�yZQ�F��u� B�������Fna�-�6&R7��A�qw�A�4��VeP̢���)�=y����H������:gscL�� ��7$s�]��+�<�0����c�%�Df�,�L���0>@�}Ab��>-��t&N��5m��������-��dg�jvs&9�����s�)<WG�(DI�gl��ݺ@�$~J����ۃ�͎�h*p=�hX���͘�oYxk� 7@�'W�!;�d��b�Y1�
��	ղE��y���56��^��Xt�i���\6a�����)��^��J�x�3� �0��+�}kkN�B�i'��=2*a[X�� ��[,�AC/@&�M9Vh�x���xj�h+���2dX7آP�F��9�� ��wk]VS�O�D;��6M�Q�8	|w��P�2������tvjѸ�`�	9�C$t>�-Z�ElKH��p����㯓�:��K2��]:!����FI��6��)r�C)N������7�:˔R�@ծf4���>�&��s�f[�^U �H��L�b��������*i�PL	�eGq0�BT����'���Z}.�W���r������P7U���G��=H5Ak]ǁ�)89��9~:Q]�3�/y����
<���!�[$+���3�y��RZ��-�t��m0]e��nvI۔�q��.`d<�{$�W�}��������=U�����َ�	Z��~�<�vj�q~��%��ۡ+�UC����`�{�����F�_F�f��CÚ���KZ�)�>/�TB��٦ nDG�T�FI��ʰ�U����E[ӬL�hǊnu׉]YT �n{w���̏�+�W����\��vkܜU�5�o&

dM�r^n'|���_`�i��VW"���j�܂�4�W���>`�X|����KD�3�
����I�r�u,� �:�U�1[�tu �g���n[���[K���J"��j�d�bvL����
�;��;���YAL-G@���;���a"���r�g����ڜ�(��VdY��} �GU���5��6g���¥�W_@�R�D4�������W~^gN��b5/����9�1 �.� 0qS�!z������-�!���=��Æw+ž�@}�o��O6�����W�9����>3���5TU�߲<	��W�z5C�2XLVPJ���2��5&H9OZ�2�=��^%P?��~� X���LK�b_��PW 7f}�f�Ii]�έJ��O���#�|�������(??�"-6~��&��|!/
/nv�g��;:�n\2�i��1��z)lhL0Kl^���� ��>&e���rw��n�T�=>>t���d�#�>�j��w��|��t��Uȩ�+���e�u��Q�,�jK��Sʳ;CI����j V����z�9�͹�d~��r<Ic��Mg�����I�:vˋ-�}ƭԹ(�2H%e/偪��+��¶D�B�dt�;��H���$ګ8����H�X;�m�X����Q�U�	-�ӆjh�N�޳�5ưL��b���P�,�a7�^A �O��8�j������6��o=lFo�ޅ����;�#V��(�T��ٙ((����\̡��c�iɊ5���G�jɂu�y�跼�iQ= ��cCw	�z)���5M�$�s��=���Llv����,fSr�ub�D�ߛޣ&]9�m`At��I��U�~�a����WQ���z!0�n�,USa�8Կ�P(_�q�����ؼ� ;_�*<�K��Hm1s���(8���%`x���^zߧ�
qls�F�a%.�..3�J0����6�9��تE�̳�j�V#k$(�H� ���Գ�ͧ]�����Ǽz��T�9�
9]1 �|���{|#!H��P��D�@���l�,�/k�]���R�kt@b"����J����6+�b�K��[��c��}\&���>�}�<Pv��~�H�{��y*]�o��!cv�0��p%�B`���ͼmrO	-��\�
�C	{up|�����EҖ�J��3о�Pn2����P�����]���g�_S|1���+�ɶs�ʗ8�t,�(J͆{{#2��7�.��9�/����l�����A+�<9�7���m�SXb�3ܐCn��I��	�z��l�~�,�~(��G��'����ue�l򦐒G�P���_�������͂4S��}EE���s�Ib^��(�D�ZwU�;�T��]�~���L��^�T�O�*2&yb��:�ǲ����~���院�O���6�V��l�G��hPrɹ����Z?�:(U1�d�"�=4�����˯���!�*��'@�[�V�?��Ʋ-�j��L}��I*+����$.<'��Pճ��9ۂ_*����B�ϟ��!��iז��p'|�����g�67:�AS��TfF��Ih���E)�w������̍��Qj~��j��-�|HH͙��Ay��I�H��`���Lb1跻6Ff�߳jYtv^݄����h�fb�V,1�{9x��?�Ć�jZ�pJS�zw?w��md��A��4�=�+��B�Fl%�4�+��Wݙ�H;S���fӷa#�	e:Z����)9�*�i+O���ԛr�F�&�jq!��|�����9� >}�U$���OD�#AV��JD.v�)���:�/d�c}�#��L$�x-���ɀ�?�R,J�uw?~gt�g�[�����#X�������DLB}�ZK2�X��t��oD7���6 �B�b�O/���Ḇ��NW����7��q�R��%K��K����b��|��O���#���@�t�Q?C�w�j�H�n�c�W����RvcT5ﺬN+Oٙݨ�xS�_����cN�_��ԋU-vzS��7�f(�s�`�RsN��Z��s�Cr�SL|�\ý�8�}�E%$�C��@̹�ꆶ�ʃ�?����a:u��ߤ}�J��}�@W��)2SZ4M�A�`��Zv���MD	�o/�{�֟i9LJ逶�)�ŋm��q������1����Hn�br+�]�Y�V��M(ۡ�q�L
V�2�:��`w�B.�o��&�,���U��rk���n�B��X�M�zv0���z�	_�oj�~�*玒��R5�Q�&W`��ڞ .�t
H�|�k	��B �ǟ�l���Qq>#k�$*��ptH��t7�MbK�v�rH�,c	�󺩂И]���j�X�e�Od�[`
�m�j,_8ɠ�N��U�7;�C.��Ze:�&d�$q+�t!�U��섰�(�WE��v�w�j�n�GxlGS-�ʞ@��Nt�T���b���ɍ}S|��o���"�QM �XeB�ɃY�ś����=�m�^T1��n[1�w�6��pG������i��׎��js��֚)�3�a���]�O��xd�u�88K9x���xR���3��*S��%���~�o�U�30��8�� 6,��r���U��$�\'�Ȟ����CE��]�*~�mٰ�2�PZ�Dx4���w�^y�cN�Hz3y�a���Z��3��k8z�"�4���H�6aN�n�u��z�ޠg��{`H�ޛϮ������p���I�5�ߺ@r����>�0$XT���uv-�aVI����t�\?t_焆��P%}_��a-XX:$&f�
�G�
�q�e)^�f��v,��p�ۥ)�
��ޜ~Eӂ�x�ZdV4@:�;�&423 �0f����@��9}�����'v.k���l�P�T��c�����ڃ�ȁ�B�,�:�\3��^�P�J�C����KK
h#� f�KܟJ� �����-['КQmCp�8�t�-�2;���e��(p.��S��� ,����DM/%Ž�U@\⩌7K����w*X�g7���t���f3�A𦀾eo�E�2��Z �� �t��V)��5���c]�Ӵ���D�Z,Dx�K����	����,�[p�\[�L`	���n�}X��$���s�&�^0��*B�,
��09(�������kB���q��93��U�u˷��a�^7�v�[��7����?�1{_.jf� ��s��� վY��`�r��i*�Ф5����3Qz2������WaN��m��A�z��Ƈ�!�P"L������V�e��X�µ���
W �`�u��2�|[j���C�hl���敷}/[�<��	���l���Yr|q����gz̖���U�f��0+�Y(t���~n��(�	�.��v0
��]��ໆ�:o�Ĳ���mJ�L����B��l JF��̪�K��&��mE�^'�l�/hk�m���t^���xm%.�3N�0���|ƕhZ��r�9PPٛ�[Qj�x��1�@���ߐ���%#��Ѽ9��/��'�\�M(��N2�,F2���r�wW6i�Ů�
�_K�y��%n�ع}�Y��N�'���;��b�c�C/?��;?�n9Ȅ~6ȵf�1a�4/_��������Z��ܤ�����_w�<p"��v����Kv�'l#���#�ԁ�Kt� �ES�"�[)T]�*�TI'�[_�S��"���[���Ds-�ֲ��i1&�D|=}O��B�}b���	�%kY[��R������h��}R	r��ۛnh	7(32н�������rI	M�n;�ن���@_C�Ú"�_NMZs{�it^g_-�귶<����1o�>l2v<ʤ�{�f�b۴������s0��'X	��-H�\K������`�o�k�R�~�D�K"Z����6��YX�\��k�
^��)� ��HקId���T�Y�K+)�*K���T�� ���)o�Ə�0'��NIKH
brJ��@�}2���=��h�*&ʽ��KsO)���XR4q���6�u���Q��d���W�4�r�¡�9T����p`|'˸�Fz��v�m62�&�|��.<х糵oE8fu��̎��墻�}&5�[$y�H�v8T�!�}���@�,��!Kl){؈�B��^jM}��1�A�樋����u|q���2f�mt��Cؚ6��ۦܛ�y�	����z5�	Jofq�~�e�k�'�5��\I˗�g�v�"�0��s������Ƅ��\m����l���P;=>g��4~k�9p�� � �(�P;��W��
Yp"8�Z�j��i�D��^�}�]�&	�	%D�N�C!�Dҝ	݈��ׂ�g��B��b�4I�����K��OE	��x1��[���D��!�4B 4!��c�H������;v���vW��ɆT������	�Y#��Pߨ�J��\y�-ZOX�|����Hk�T��r�,�E����5�V�) ����AY����#�v�b:��MW$f�=FV��ót������x�&"��t�.�m���7A������Z��`!R�� 9I��qH�[6m�Е!�'� 	Gl���߻z��M	p�U�;��jP�%�4�Fad�Sm����{��@ �Jo �
}���9E����u�$T��Q�̸/�;��8	�2��o.�꫾g���%��m$�G`��>s�e
�����\;�,a�r�-W�jò�F�h���$�0�t��9w �~si0w	8���o)���T����Z�$�O�-�w�.o]�h���Y��߮�A�=�ǐ�xB!1u ����ƼݑE�+�Hu$�h�y^S;�����=@CRM���m����]0s�y�XL"-r��W��q��ꣷaѻ�s	�o�
�OTzĸ�e{t��E/��j����t�^/������I�AXgY!�;����k���D�6��N mk�T�[���t�s~+0Ë�S���g�T�,r�x��
��]c�5ul[�:���ԩ