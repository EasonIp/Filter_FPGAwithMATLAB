��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� f
���O�Q��Y.#�d'���J�"����4���d�"�Ŝ9͜����
�~�a�rN�����o]y����1���nJ�]s 3L!��,���zَaw�{,���{�b�[;ҙ�u�\��������.7���}����H��ΰ�&���ے9��y��y����͍2��ё(��7q|U9��1���i��$>�[�G���^#fU����S�"_a[7B��7~ez�#�5��-������>[{Љ�v��G]��Ew4��5`�|x}��4�y�z�f�|#�դ�e��5p���1��L��d=�㺔��y���h����V���Q���t�̿�rբ��6�j�mcP�iT
���c�j��5�j�KL��tlV��d��x�Z��"ks�kCK�|�i(�;�����6��12�XTeP��[��'�0u ����r/X�<��/�]Gȥ���%N��]84����Uwp)
���un(c�Åf��J��f`9Fqv]���+�<�w �N��fѧ�h ˞�C;4��#�i��T6n�Q�T�����ڸ}�rS3�*�x�٨�j���y�~E�s�~+s�G��'��%`+�w+.}��(Jľ�$SL�2-�M�M�W5~���/%��t%���0;��3��G�rq�Ħ@];
!}ˬ � C_3ZjT5�ъ���29L��>ԡ��I�#iDn=*oB'R�؍����v��< 2<���oc�M Yx�R5��ܡ�����2=ړU��oLW9oq��4S�um줂f�X+��t)�a��� R��M�Ć8��,=���LIQ�n�Ҟ�ݔ޼C��`���.��!�i*F�8����P�X�v�7I�i]��q���=)6��n�I�p���")&�73O��(	�������Ovg��n�C]�g��2
�K�Ι��ͨ81��E�||�,���Dpk�J*)��9Kȉ)(���f|�(��f,���/� ��V�R��	�fp�Yk���J��������j��j+f��i�x��J�1�ɆʮL����Ы�x���lQ�+/^�+��/�I1�Á̈U�Zw��F�]�
+�8#(.?�(hc�ZC���T*)�y�����l�p иr�W�.g�����l�q/��%Z,�	���r���}�<#�Ϟ�E���,�884�ǟ8��J2z\�z~��C��MŨ�3_2�㺃V��8�ϕ`�%���k"���k�z�?��']^��>��A��#
7��9��t̶8$�����0p�.����2'n��I�ǁ�r�`�쿴4:KlQ9����ƒ�[(���`�C�#�@�Lw�%{xOR��>Uj�
��|��`p��e/�����Y��$b�����tljXx�	�ε�}�Q�3?&Im<!8&m9�_m�����>C��hn�<��k��8^�̻��U7���4��:�!%�'�o���j��'�!/b����/u�ƴ��x:E�nr��!,�����[�صե*�`��7���z���@�͗��.��`.y4j�ǐ�x��҈�V�� ���g�ѡC���}m7�6��i'J0���D,*Z3�!��R�%� ��~����W��
|R01 #3�)��,ŭޠL�
�sp��������L�%4Xc+�����'ǂ�2o�uM�%���R�� r5��*�N��i
I��Tk ,lNA�6Ȅ�Ăp%���>���E�D���B���tp/�EM�����&���8�TH��s(�T�����k�;��>����!��z:���n�Q����P��(�=9�\�~}fE#jخ�-h@"E�_u�㐸�~��[}����q����L%��(����x}���Ͷ�-� �*ĵ���J��-͂ġ$�)qah��E,bji�`ܯ��핼��<1�
`��3(�����sS�=�B��
��6�Z�n���źC�]]u�/C^�nlӚ�+#�����uA"�����8�1�x����%����I��_?��dk����#��Ot9D�����@�l+qG��:��&l{B;�A��$ߧ�mx����\sN��M�j��|t-�7�:�x~���딹<�B7n;>����z}D4e�t6,-X ;v�u�AAA	�J�V���+��+n �@t"���k�f����QU��l����ے��W���x�ɦ4��\'<�x ���[M����Pt$,�N>Q���j5p����J-�A��핍qS����av�	ˇ9|ڰ��BfYG�	�ŮE�f��Hղv�<�Q(XW�^����)f��-�,�����>��R������HS��u��7>	��4NV6����ʽqcp�������M`ި���,�?�f 6�-޿l��N���� {���]������[��*B�;�{�v������c�wf�uLRO� ��⋓{���m�Q�b��@�$u-��m{@S�>�-*��J>A�K"-/5�\7h�k��E#��1і�%6���6�?��qӞH�]i�E^�MA�X���{���ҡ,_�h%%9�*�1-�B��1�ѸW�H���
��d ���;d����ܺ8�O��_/7�궇;��=�S>¨�KN�Qhj�yB_o�w��x�H�Җ0���R\���_�����7��e����Z�^rL+,�6�9���
���_8�Z������%$�$3��U��/�H�/�˽7�XJ?��I043��2wR(6D�Zt���%��bjNY���B;�����)�#~��=�j�6dZ�����ԥD��
yT������z��f"�,�g㞌�}o	I�82�Qj�N��iY��ӎ;R��7��	�k�{�l7I���x2���h���dq՚y@���7`���Y�:n����J5�m�6��F,3�
��W�ֿ�9�7�6�|�k�f�4�7��1�B������b�;�D�5K)�R��?���H�q����ݴ{��q���}�K��?[�l����k�ѵݎ�zX�m�U��	�O�j&��gDd�Z.Үy��0�H�o�3r�]?�y�li��¹�83���twbO6�0O� ��F��)�Q`%���o��(��TP _5��1�-���o���x����)�li�����o)�++�m���