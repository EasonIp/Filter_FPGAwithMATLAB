��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�J��"4�=�7(�T�JѺ�ő��,\��s���ӣ�F�؏���PlI���'Ժ�0L]��-/��1P���n~'�\�eƟ�����I1eDC��:-H0�-�����hNl�i��V}�p�#!��!�@甮��[p��
6��ɣ﬷=5�X�L����2��ξ��*�=��A,b�d�^��ZDL�|��ʼ`�Iz���?�pc=~��Ii���������(aA[��5ݬ�y�#Ǿ^���Զ�m��gŻl�ؾ'Mb�B	�,���3��(h��^����!��7X�H	���z-��4sv`�j���X.,��bwmfn�e%x���?��X�T6ҹ�������z�\b�2�-�)��z�q��GU���*R������`?,�s%X��N�<A�O����^	@�T��8'�\ob|�Vg�Rm���x���ؘ��hy�� [aǫ�_#���~6����A�[J;��ˢ?�vOw!��5�y�ڏ�=�����O�	39n�Jl�󨗒���1E� �j���q,co�,�j���|V6�#�!*y�^��5TR�L�;T4����
�\�}�|�����+�he�C�{�N����_�[�������,j� �08r�zp(=�{�ϊ�>��u<���%�Z�K|�8`�iś@)�y�(1t2�e�I5������(���������1��/�����Z����b���d�~@P1�xB���oo��a��U��n�u� ��|ݦ1�P���X��j�׵ +��AT��{k��u�	 ��\F{.��'��Zޮ��Ixd)s}_�0qY��4B�7�˹�&�I!Oxi/�^��������;���1O��|�]<yų�&K�U�a�����uD�g��\�*�B��P(��S�r�)'��7ȹ�+a4b�PnK������H��{S*x**��_$w�]B�M��{A��w�;=7p����IJ�_ꄰ�ӆ�L��Dk6q���[�O=$�	�­|��cW�=W[_��q�I�1C�S� �{�qT06�M�Z��iP���3,����0�׈]#X�"T��g�s�ɠ��Q��ǌ�����ޥ\;n�i@a�ʾ�}����K�x�G����=�s�j�M�)]�Gq�A�;�j�'%��x�-�����dzW�*�8+�7u�g�Ƶ��P��^y�Y��\Z��Bî3ã~�v݅/�z'i�o���c�-z�ʫ��������*���E��pĸc��x�2��C^9|�#r�BXw�y���D�W�<|Go	I6�iIG��P���G��O�XeN�ǙC�sÅ��Yb �3��ЊԥҒ��I;��V��S�&�߸�6�>SƴЭ�A�����M7�+/�	;� PV�}�: (�P�4	"}nh#ޜ��?�H�o*.��V��:on�q�����?���(����}?��:����\Q�>H�_3l�v;�Gtټ������<! Qk$�9��M->~{)\����U��C"����O�N��Y:nG�*�oy����<XϏ8b�9���]@^��}��R<�f��A�Ң�d�z6�N�J�d�����:�Z?:� �3�k=����}"S8���: ���DƑN� ��;��5V2!;���@�DJ����}�^�X�r qULp�H�#�r*H�=�lK�Q	�ݤ�y�ؿ�A����"���r��n޼󸂇�[�l��̆���g�]ԼcR(*ɚ�Z��Ã@�^�
���V�[��-tu�?l���ט�"��e5���� �W|\H�>��1���t�%�[/w��fO�'���A�&����5�*��N��E�n�{����}F��I�D��>ގ�#�S�]��q��� �L�YL)�X�0�sÜK'���$��~H߇�~��ud�y{b�����ɞƦ<��ɀ��Н��C�������C�q-�l3��6D�v�,%���\B�V��?Z/P<]��`�(K��B��ڭ���X);����g���R<7Vk���љ��l٘���@p�5�vƪ�U�1!a$����֔������j��������na�&]�e0dt���wؓ� ��1?V+�l�����39�s�=3?ɹ[%����".e>�\� ���֋���3՛A)9lp"|�����b�a"�%�(G�c�0K�k4��j�K,���R�@
��%0��ңA�a N�V�bqPZf�|�qC=�Z3kp}w
�	gZ��x�P�ƶ-L�v�I�i��݁F9�u���t<�bnP��0\���Tn�!magG�m�r�Y�-��V�k->`Y�X���{��$Q�
��}�$U㝆�ܕ(��� ��S�<[竝�USܡ�G�|�!:\���Cus���.�Pm+m�5��v4v�Vq98��м�HP���u���FĠ��94h�?C)x5/x�	��ۈ?@����B,\+W��|I�+�R�tm������׸HM;���\��ʳ.p��1H\���LP\�)�Zi��>��=�$�>�����*�z��s�s�t�a�*�Rf�Jkr���p�(M�\^�	~�Jy,n!}�~93#��2W�(�{�J3�Ǐ�ȳa���}��K<SL��̤M�ZgT6p��ڂ�*�Δ0to�򽝻��E*���?��.���� �g�&M�f����Vi5I�w���yϧ��UZO��Q����d��pfE`�J�&$��`�pR�i|d�DZ�O��Y7hIɲ�V�>�Ɛc𐏦��a�ؼh���Q��N��vF�A�V��6D��~H�?���l�3G���B)���J�2+I��X�'��������"S&]Q��)�I�$�T�}���3� ������o���������� x<�ݟ�y��ƑM~_������Q�8�$^�%�P5h"{r͌$��P���wˏd�&����m����dUH��I�� Re��9�����`=	�R�74훫������\q�*��C~�?�W5�qys}P���k���V�=��j�x!|�sb!�E�U!����9�|�