��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$��c�\x.-�M��h�T��ȡ��0�s��	��>��,-�M[����ZAy~C('_�v@Վ�E�AݛOf1���WS��A��6+�e�-���0�S���	_~й�/G��?;�Z��G�-��v}'�(�o�������"��.T���$��.��(X� ����-%���o�@k�<ת4�$��4]6�n��A��NI�0���i���>
�� �OE�W4P^����R!;f�70+_O��ĺ�b��A 0���p����^�3�Ú��L5u�Fx�����_�43�a�<��BEIݢJ�R�����8R��?��
MҰ�ö�fO���O�)�#Nf|�In:6�ps�.�y�BQ|���/$�
W(�U�݊0��x
ZӐ���Д�oB/�OQГ�`"ş����ցOk��G�۱bj����֥�Pv`#�By����6Ed�+{�(�!̜-�]�6�v��2�]�뺠~þ9�m���|��E�)�r� �6���� �MYd��Q=�qs�L�FL�a�_�"��OT�mz�f�}����</�㭍�H�`��v马���<��_�\]�S�K)9͎�?�*AKW���������oD1PY�@��� �qX΂,M��{�}��("O8Q��O�{96!`2� �	׫1����ܚ�f�T��M�T����:v�ΤK�P�l���:�t�dH��#�:ߖ]��GAʊ:�Q���5=�^��>����ӺL��%��c�|}̈���zi�G �C6K|)���r��z�.]����X���~�Z����:��cg�7mc�Z�y�8m��~�\s��ݷp�'�Tha����:�L�6��E�6'����::��u���b6.15��A��J�H�-,4��W:lh�f��	c�b$�eRr��&�� |$���F�9"`��i�<��#�wp �L_��xAc��FcU���4�vG�Үe�����L��|��V��7���ne%��bg���9ay0S\v'�NY��5g���2Ǣ����G���P� �4ꗥ�yÃO���;�,7�E�
���@T�ӈ��?td7�B��Y����O(Xϳ�=<���`�C�B��֚��ۍ]�x��'['8J�w�,-�!�<�(�e����DMF\pF8�r0�|H#k)�&�Kx3�(Y�|?`A�2�)���9�LN5���
	���lEn؛�1%ryp��>��Lx@W������B�g�F������0(��_�3Vg�c>��0`L�F�u�AyL$������%ٰ�w��b��C�R�@8�OٍP�N�ɽ�e_5��ԝl@P��bê�I��w'���C�;�;
�(���c���4�S�p:�J���׈lźw{�L(��3�b�P*BB.���']g~&�3<?�-����	�лw��O=�tg�Ѵ������xӖ7m $�f"٘�pC
'q2�+��������47�'�#\���-�twh����$B�,`��E�u��Q��7.ĶYuH;w(�}�i3�7Eן̷���OQ��1ܯB��b�Џ�W*��Y�l}M�n`WG�����֯,�q��(+DN&�0����cM�x>��>@/2��g0�����	��%��/u1�m��wD�����Fq�����b�,�9A. ��r�"6�0���Л#2��e����R9\jK�Je�D�7�
�QZ�{�c���ޛ� ����l��N����&���^[�_�Le�G��g#�v	K��ay� !l��+A ���8��\)�؅UZZ혟�4;�0��Yeglֳ��-W�G�Hk�1��mG��4���غ*����_r�zMI���C6�&��mͤ���f�$�/� ̝eS���⠢Z���9U�z�^�H2��:�I��˻�/��)���󸷛�E��Ǌ�&c�ˮ���u��ni-�YI�7i�D�������V�|�x M~�F�����(������>�߽$���<u�U��Wh�1w�@)t]6nZpj�;䢋�p��;�K�[�U��4=�j�"��(륟�.��g@��"�j&_��k7�xk�gcgiڣx�o�U�q�C�j��k���8#�%�(���S̐���p��!����`1H-�m^�a�K@kIw��,�QDx�||��c�<$�o�[��(�Z��͝��d9%@ ~\��������/L�K+�c� ����ͮ8%�_"�PD�ccGQ�0/�y�#{�(��+z%�GA���e�x��������N._�c3��|zl�I�v��������W=~Z�0R�R�̆��e�Ϳ�2���������p�kxHAǫ���|P�}����������C
�tjW�2w}o#��r��c<i��!E4uo@��e>ow��'a�������C�l��^^V��#��Ҟ/��)�Hn����'Yf�p���Eju�Ӌ�e*��s�-��M�Kh}�:�G)�N�=�������)Ⱦa�9��/)�5���6�'�Z�&f*�K�  �e[�����"�j� -�k�ь|FOggh|vTF\t4���JW��s+�Bw�
=$75�čـd%\�݌4 c�Tu൫�<�i�J��?e� .@�����1O���cNd������� *!�I����?��jG�88	�e�]$�����n�ǁ�3���zM>��+:�F�+m5vR����::+�ǒ�C5`-�'�C���d�b���3TH�����6<.�����m�w"/����C�rh��0ƞP^�G���N�Z�:V��v�r�oy�h�ӌ5���U��g��a\6[^PV���,�l�ȱϼx*#���Q��	�՗��{x����W�� ��LWXiׇm�y�`u��q�u��go��b�uU)���X磴����t`&lj��=��&P�c�������§>;1��(�o�4@p�@������.�q́/?Bp��6C��o��|1)ʘ�҂���`.��\_z`���G�ք�w`1>�慾��|y�|�mF����:=��������r�{q���s{�E̪��ӼOZX�"K�`;j�h'A.7��r	��.�<a¾;�"#�:�+Ď��]���W��C8}���f��$�.t�%p�S�UWF��M����T�H0&�J��*x�|�\��:� �����-u�	,,`���d�e<(�"g$W{�\���CE�m���dˉ4z8�m˚�0ى˿ε
�p�ɻ�)���u��M��׃��jN����M/�#U����!L���
~���'-�w5e{���y~�7ٙ��P��7�qwr�N���p@6�:Өﻃ���crA�H�}�8콚�9�in�r/QR�z{�� +�/S�it[�n�����Q���U4씳��(#���b#(�-L�e�m����wlTʣ럔F؄�)Y"�po��!2�R�G ~�q�5QS�o��i�	���2UXZ�*�����	��纆�퀕:sa���Ļ��2�qx9r>��0����O�{�7��xefRͣO>
n
7:�j���\�%�i�X�tJ��cf+�2�Z=��*\1��^��2*��-���2���h-���tŅ:_d��t8LÓ�����~�D^�����|���	��e��z���|��ᨩ��P�L�2�i�w�?�/R`[V���19�u�K��^��%z�gi輠҈�{U��n�]߭�<tr�:k�&�0�����#��ˌ�T�f�{|t^ �����Y"���_��7�=�|�"��cU{�om�<�Ɠ�B�D�)c�K� ;pYL���y��ΉD6O���n$�4����X�N�M��\�Q��8�+�����a�w"naV��7��&8Ѣ���N��&��K��9_����w1Ht)d�6�/� �xL��D	�A{�m�ԯ�Rz���P'��5�xf	J��e�p���SC���k��d��
=wPi��fn@�:��.(�y������{���$m�Bp->G�اQ$�>T���H���@8P@���B�d���_�+�M�:�L!��tzit�C�	�3J�LV��N:�jjl�zv`�飸RG�6�w(����'u�;�"S��+�m�Lu��8�ۅM:��Z���_�{�ܦ�yޔ_������=A��e�R��$�M�q N��ٛ�l!�q&�]z��q�*4Ϙb�=uB��]/\X���xa`���]����k���*�ÆuB{�o�'X��i�?:�h�������ګ��9�r��s����r7���w���*���\��@M�N����@G캔�����lAv��Ad�%^Y���f�w�OV�T�凬K�l<��m�;6���aF�	��r^���9�PҀ+��dS�Ǘ�7�ts"^1�b��9�S������f�)J�m��?��غ@J��M�s�G%~��
w��ˑ�i���2��k��مҫ�Ė'��b�m��
3���s)Y�EK�q�4�_����:�
(~6>�)U�X�uT:�����{���C��G�L�TK��ŕ��/���t�>�D�X̱1���Uq���^�+Y�]�}�-�k�5��Zys.�W2r��x���uEC.�f8ɿ��x�1N��{�+lr^�]}� Q��^#�ٚr�G�U` �t����J1[�L&�nh�1��͋z��('ˑY��W�'�R���IE�W�1��D�