��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$��1h��w(9#�z��Rѹ��q�-O�?�ƴ��Y�B���D������b? |L�G��+���x�q�����"�L�:*��K|��&�@����~���ȄQ����Ö[�дW>�����@
�v��Ai�f"ʋ�9�G���s˖ۊ�w3
� |40���1-u��p��F�$4�f�{%���U�Y5�緌	A�5����HH��@Y�wОM�4@�M�	�D'���~:��^@X�=�L~l����տq��K��	ԃhr�G�X����t��9��F̵)^s)!�0���a�z��c< 
�=%�ug�s���j�疻?�+u�2��Bo�vӖ��8�Y�����s�ь]]����)�u$̮}gbI�,�W�V��_5e���}��7qS����I"#P�c�l�	j�WEZ�Le�vo�x=�U����n�vy�O�jf(�Y��"Aoۧ�Xr��öqσ�q?eB��
�T[�mc1���Cr�ͷ]-��fk��l�o��>�q�[�k�n��%o�>�;t�Ù���Diǵb2�	����a�:z���~�\c�>�3YB��1�A}�pK�57��9�!��n�E-%�2% 9�E?c'�p"}�H��S��_�9ᨘc B���7A�������/���e�3�OI�v%�)�በ�g>�V��M��8Øg���r�ȩK���6�r��iw��\�ܩ�EM�7��m0�2�8������(w#�I�rg8�	���T17�F$�b���*E0L��d�եe�T��c�m�#��O�N�a�=�J��,y�1�}B��~��0U2[���v!�yy���	��`]Z���Vr���G�oA��hsNb�ss��gJۋSG�k"����ֽ���F3~f�B��/~y0��-|���޶X0#"6r�%����B�j�����z��rթhb�����#���DW�AzO�-`�tw	��7ګZ�o\:{�1 o�Q�*2��@���첯�ԫ��d-�y�/���QP%bu�&7(3����ֲ��9�i/&����r�W�^�:�������0D?�I=�Col�-�Vڙ*k��$��EF�\�Dl�����ma�2̋���!C��a��@�8�w*��}G\�j�4��2�I��PP����?ؕ���������
kZ�!��;Q��Ue�~�Z��2�;���	7va
���⨏IO�w��M�gU�x$��_�^��be��*X�V�:K�E1�yٕ�1^���%�=m��Q�8Ro�e�p9��YdH��O~n��{HI�6/�'U2�����p�e�df�n�>!��5:��Bm��m�'*�О�������7�I�P���P�!*['�Ơ����J�׉t����E�g���������
n�Y�+!E3q�g�%��0�q$�������ۂ��T1�-=��U��n���>�5�DDR�	�ɜQ��>-�>��ʙIN��F(.�J��g%�O�'����@�TRw_g52C��@��7y�D� 
O7J�ˏC���T][x�yo�hj��s��4�j	�r.�ܳo	db��� Q��u�n�a�0h#�C��`1|�j��/�	�B��/$�Ki��{8�	�� �.~M�D���邙�`& ���@8&U�کkq�}-�y��E�d����ܿ����Ԛ�M��lT�<���i��M�%�]��1mi��IK~�hfr���92ʗ�� <sQ���V���t^b�k�~��m�4T�y���0�#ӵ�<g(u�S,$ Ysҭ��fv�ѕ>ni�p��*���t4���Z����Pt�h�>κ�ӓŭ��&�����{A � ��):����]��Q�_�5�!�q9�KP�ڧ>'�
��ݑO1���(6����@r�נNX�@w^ګ�/�`��D4�?�}xV��9�/u
���V/ؠ�7���.��s�����ش��H��.���@�WaV���\Ѫ1�h	<%�f�;�w����F��`}'Ӏ%�ҩ��=Y@M��<�H!�W5�_R�P������:����p���Q��rո�y
o+��t=���Mg4-�e �Ԗ�c,l�����Rws�&���l�_�X��
�hɶ�h{���l���E�O�n�c)��&#��"2��x���Tm��t)�d� GTgm��8�K<#�:s1�8[�3���0��g��S�xA2��з��A���:��\��X�T`n�'ʜ�zO/��uv�6"��\��Q�6��O�y����d� =��+ �&I���`y]S�D��lV���s)-����jɈ��TN�Fn����+���ђ6���%��z~�)Q)'�� �T�Mk摆kܐ��+f&�њZ��\{͘�w=�K�s�X������J����BT�_�+��-����u��W��p���\�=-��T���P��U���B:� �1�S�> s��
+���ӈU T����m9���èЦ�ԯ��b�Ὺ'(�<#6+=j�̉_��ܗJ�����A�ȫQ�P�����%7�R�r�-�z` �����B����pv���!\f��@ԝT �����+�u �H+	܏�m/���L�J1Z.�.��H�B9NY����D�\�t��a�����tj��P�����3K����>.̓c[&�jE�>���q]��G��@5A�$M[G*[G׭��Y�Q(t�=�޹�8�<��	�ءh�ud�]|���E�49ި�
a���O5Rny���3����(��+�s�>���M�˖D�>9�/����p��?9���l��a�4؀8�#D�;�q������M�?DL�_�����vD! .ZW�� }E�T��ht����j���h��5��F�M?7��m�^w�����BO�0@���8F�%p���/�8"�5���9-@eAWUN
ug��j)ry<Mp���UJ|B���Z"`ӻW�n�d��"�pў�S��y�U^e�����B���밙�=s�O����d��6��i��K���\���0�F���TE;[eP٬��?���v���h�(�`�,���]�<3Y�ra�0��!��̈́�x7���̝��a�H]�����v�%��J'��EY�E��-��x]�oyk�;~>($�B��/՚^�T�E �з�`�����-i�M�o�l�����`s���A�;�-n-�>\>�����[U�/��(� a������K��:C��^����Կ]T��t�@r�RK��"� ��hȮ_�m�}U��,R��k�����!Qr{e��<`���o����nl���Y�H�����$��)D�m� �m+C�� [�aӛ �\����kaWi��fy�]�����ox������,f��Ç� �TpD����A����Dv�I�Qԏ�q^�����k?�wC&���7'��w��=+r�4���=��(�i�&���zi�Xtd�"��7�-7�".SW�W��^�j�՟�Z*TV�����D!\�PBjN>3r��EA�kVP�-D�_���<�꺑�N~%:�bh����5�M���9�[=�Б(g�762�L�D!;̇��`���-3��8ԆP�����	cU�P!�م���m�Al��v��$��I�y��2�����`�K����c��X����Q���0�E]�����.��A�����{}���	�TKOX.��R}�\�՚�mX�T!_ń	�඼���Z��B��J.�E=g.Tħ�<������M��"��Y�:q�|:��<&��B���E\��4�^�R���Z�XЫ�S��F��������g���3v�|3̧Usj�O��[��*o_{�$��d?��)1�D^7��x7�l��>իp]W���e@��6�H�[~�	�����rj���Ǻ��r
���G�{j�۪r��W���Q���]I;k�k�Z}R����&!�h0�x��*����b5���)-�Я�a����ҩ˭׹�.�wr����N*��(�iW����G�W�P�7,�_:���=�#�S�(E�c���m��s�|{]l����@�19�q�@EU��\��.��"t��(M�;s����C��s@�~����a8�ȬR�%��,Y�cq.�k �d_�&j��(�t�\������;�A���f��:6W[;ߑdi6L��ÉS����&��F��Z����0u2�5���S� U@_Mt�b�?��>�p$��܌/r�҉��}���Qy�.�Ҳ:��w8gW�Hx���Su%�,��x/�����.��ǕzcdP�8�	vbI�!H����'��꼃8>��HZ��)�cn����I����a�-�H�y[�����t��'L��	�CN
�<�e|�F�a_֊�%�}��[R��]��y����a#.��	:�ɭ�"q���	uJvn 	���$�L�@4	!F%KZ)aA?����W�|��^��;ϑa���`k�{σW�̼2�bPڗU�u�5��,�lSO�L�t�6��p(m-W��^-'31q�)l�[�a,�ս��X�p(��r'���)����i��p�����_�'�4�3�c�%����:�H���H��`D� A�o�T�������3¸EY�O놛h��ɳ����@�^��B��.�;26���4`����蝁;�s����L�3U�Ȓi=�ȁ-1և����xa�GK�v'����i����b�XQ�SW]^�Y�f��T����=�N�q�DB`h-��;j�v���/�*?�t��3�əOU(]n;v��Lm���V�@��b1*_�{�u7�®);������J��:m�K�.���G';cj�����Z����0+��6%�[�w�b��������=��{�	SG�Ƙi�Tl�C� �r�<<�ᴩj����bm޳�{0Kێ��6��p��6S�Nq�ca���lu#H�A��Q�W�����er��:F�qs�T�D��&����M����nMu��.�B��X���ot�V�!�\0�ڄ.Ȳ�!X"o/�=��|��S?�lf��	���(QR41^K�z����y?�Z��m��X��c��LH����5�Z-Cf׊��@!�s�E��c�k
�@ۊ;�p���h�;�߷CV��*_)��ò�)� �	l�l��#$'�;�^����R�q�Jk\�� _��S%"^��/Y����"&��+1ۃV��r�k����l���I�?a\�y��|(�c(�ŷ}���͐��xQ�O��Z�� �!�hpa(��Ļ~/�JC\�_f��w�n�|���q}CU��+�zU�udjYA��
�t��a3	�R���6���H��\�ZX|�z0�F0����>��ᮦ���ȉ*|��u��K��W������T� XӍ*6;����]��xY�Y!�~�AFM�#�9A���m�UĠF{��_���3�Y`w g���(�=Ce�z�fk`o/j�.�����Fm� ����G��1�\ �*�	{����)��A/�*02��,�I|��,]]�@R�����=��H.0Ӓ�L�������s��͹<�߲�b��>x2�	�R���-gp.���樳�*����Ʉ�����Q)C��v��.Si�OE~�x��0�m\�������$k��K����ӈH`�/H=���p�Փ%��|��!̅-�TYJfy+o��q���ࡦ֋�2|�F�p�9u����?Թ$�����<�C�($�9����C�S�l���Y�.=7���(��5E�ȗ�d��Gi�_�33�*����wAu-E�7O����L�O���b���H��H�ɥ�����)z�eJN�����:�:Uǝ��2�W�}t���p~͛�~}����M����/E�|�Iwl)������:�H�I��6
�mg��8N���fY�7і��9�d&2��?���&s6�=k��jB'xeI�u�������<ld�����)�.Q��֜��Jp���Y�w��T�Y>�Qr�j*��x��MPmz��J�Y���3��(��<ܹ�Z����@"�zw'#V�ab,}����^A�ڮ�qʅ�*����^�"��P��o�q5$��]��-���C�S�y}�8g�%������ߝ�Æ�t�H��'�P��#w�]��D1�m1Ug��ߛ�X�AЃ"��Dj6�
e6�⥿��_�}CE@̹�5�ԩyTm3��J���Y�X��W�Lk�m0�$E���b$r���[��%�����ci�T�㔎cqS�}v%��?��y�������r� ����b���C����,���1���G��樦	BI�=����E�'6f��<f�,+�������lTD��e@�\������+������> _"�/�:�����@��l��(��.$s@�D���t��T�d�l���)/�t���#��N�R�$wXC_����b�ZL����uǕ��ގUэ���2� ɀ2��fM�H�o�TI��
X�_p�X���l1�6�{�)�,��Ȕ�fk�Q��,�O'p�<�v��!����	r���S
�kK\t˛��oOj;	Vt�u�
Y׸�ġ5Xp��=S�t��H!�׵季+�5�%�4��Is��61���0�	�b�}mZm�0����ۿD�S�<Yp9�ЯR)Id��oz<|h-u��ɂ1�4����r��{ �!҇�9�8'A�@д��>����Ad����k��ޥ�Z*_�b�ZY(�Z�������6Ɏ���iQ^��_%����_p��e	�>��7H������F)Ϙ���a &K=�$��O<B
����h�m�.Hу��@|�
���&��m�@ rn�!�����q�{c����?��0d�ߞ��s�$X�K>�r8���Ė��@������[�Q `���E��J`�)�u�Y�ٜ�_?�O���P|sxG��t�ҙcch�/Y��R��Z����\�F�usғ5,��k�bZY]�C��0?e$����#�4#ge��+��-���܈XYc��4�(�p�[�fb�
�h��丮�Q��#'�V2U��/'+A(_'�̏��e��r9vK�yܜ)���9�~����d�&�e���azj�S����v�&f{f7����n�ժ��MX�����k�x�C6�U��{����x�n���=xU�������S72	�U�;��q\����m�z|U��#'�4���T�Q��$ǘ�/Omc 1����u$V��"�p�wV��`%)Ox�����0�+/ۢQ.���y�r���_ޟ�{N��"�Z��N��&�!B禯ۨ��}x(b��(���M^^�f)��$�>4�KVj߿/"�,&F�uo����u7��w�n	��(ߛv��D�=?���䤍v��i	$*�ak���j��	�a����װ.M
��kZ+"[�x�Jd;/�Q7Pc��}�1!�zׁ؇�k/d3�
�$=M�9����a'º:v!p��ޫ�X<E�x|��fE� Z����� 1�(8OP�6��R:��QϏ�l�.w�w�8O�)��Q��s+H��_3��}�#�<�Y�5����5�૬�/�sf��8/	Q�d2fuQ��S�ra�T�n
�$��#-��B�F�[ǫ����xO{z�Kb",?+1�/ˤ��BH��n��pu��(v�#��DNQ�(�� �h�09��֍Rg"���pѻ�K�u7D-?D�F�֫~\�e�0�jI�GHџ�.kƉ�q�>T ^�D��U��ԭPS۔�[w�q�2�B��(�]���j�j~p��q�o���� ���Zh~��Xι�_X����%n�������iX*[�q ��x^�\x�&�K��@�"�=����G��z��`w�c	8$�m����c��荝vB}��m3�e��$�"�GC-b�㧣�5�������#��Lހ�\w�zNqA��^5�$>a��u�h����?�)���e$Ty��cpCg׉�b^��]����������$�S�	��{� �q^�ٯA��+Ր��1� A�y�����HJ
��]V��>5~�	���d+PdɇVl��.CspE�����r�s�73xD�B�
�b�ᔹc%ą�T�ؼvD{����w���'�t�:9��]4�c޳q'�s:�?4��	R���������4��؁9��:��-.�r�y��� h7��R{�� Su��&@��o9�j���sZvME�5���iRvE±�-B?m���C"'������q��8=U@j�EK ����푦J��c���3��T�e�+��W�Av@wV%�?�:���j*y��v@�eg��y!c�`�&0��d@h&�z���3�C�f��Pt����,�b�Y��S�o�CX��\(�|q^�1����\ۙ+]�($�ML����|;���A m�3�T�k%@�� -��@t������I(Oʹ5�3S�_X����R��HeLFW��xI�cq�g����*6R��H�u[#f�>	1	!Ot��'�l �MMw�_���+ֱؐ�O���G2WВ�Vi����#��ld���$�tQSť*Dh�P�t�ѫJ�[�R���ao5
�� ��+��KF۞���{h��������a��.���A��N{E6��eK%� T�O��,O[�����]�T�=��'�%J`�(H:�Π�
)x�vz�Ⱥ�Ʀ[�jt�N�r���76�4�!����K�;hM���H��p6#0��k夊��?��{��6�jt�����N+��#�f'/Zc���g�а���u��Y&3+��"������-��oy`�raG�� LT�����.G�e�7���@�_ +Q�WtMQ1u��Xz<�fõ��&M�cR��^l&7���&��sH�yl�E�J��j@��}��Ҝ�J$�������7��n61o����y�����pf�%��4���oQ��J<�����w��Ph~f��z���S~Y����R͓��uY�l�L�K����d�m�m.us�@?�2��Eg�C�]�J��7���C0<p^ͤS�d��<	L��b])+G��"��M�F���M[6vAG����FS��d�%�zs�*��,fZ@���c��F�� �9����Ӛ#?ˤfW�m�E\˗źH���G$h#FU�Z��ٹe~�7����ʾ@Sw�+k�`~���_qN/Æ|��n��&�Z�r�&�
�&������1%p�F��Dv��7�@��8}2_oҫi>@�+�kp'�i�����=� �ZN��H���@�u<�>�G�l��o�֝�&�\��0� uYz�TkÅ��£�d$��"j�"�4�ͦ@g���$���q���V�R�1
�	� ;{�ɗ�Y�?��i�%S�͠��<l'Q�z��k�5E�;���y�-#�3���!�ii��j����W��S��i��2�P��ҥ�$րet�	;;� ~-$����JF��r'�T[��?��� �ʶ.�
�Yf��T����d�#^=dHN��Y��@��6\��Do�.����gH�H�0�Sfjk�Ӻ^�ϖƼ_T-b��+��Y����iZ�9� �S
??JH�(�D�&V��� ļ��8��Vcc�Q�9�"dTO����ڀ�ĕ|���~z@��'���H�R��4'��a�9ˊ_1�u�:Y�CR�c���k�V�ǳ��:�]�OjRY��\��¿�B��A�V��g\$�r\��18o%�w˘�G,�]!.�^�HZ:]x$�g��?��w�sU*X�X�(��d`K�T�+�e�Y�2���#����"�6XѬ�d���M�gK �,5Oo���9�*ဃp���$�Y��@�[��\���0���7D�r��m�]~C8���ø�/��{t������+Hf�7�������o��p���-��]���jP�������w�%��H��#ebY��,Vǿ�_iٛ��� f׋��>��0fK{���lH�m���R�z1�� %S���=+�����ŋ�k�hp`N��`�3�̓:���$��ۦ�li��C�a��"�p2fGN�9m��8ʵ!=^@to����^`Y�Y��ޔ�����km����,�����I�i�'�I�|l��>Ҧ�ڨ������.(nSe����	9�g��[>�W������{	��&m,}��<��Y�����d)C��&�X{��4�`���Q�n���))̻����gճм�MM}w���N1+0bv9BKМO�K�Ji�7*Կ��{����NM#������%5+=��P�h�i/@��M�3��(#�e��B^ �%�55�Y��hŀx�\�M���AD�E����\��{���Y�֞5��aQ�Dϻ�颠��/Ц��+K����+˛k���Hw��Iz�+�A��>حr�,݌1U3���x����GW��N��� �D)մ��oM߫��Fu�!����,^"4�nÎ8��֤ѫ��Oý�{�B��;�D��rBy����dA&7�.�QG�;����Q��h
�_�h�Ub5T����B�E̐�O�T�E�,�X��[Sn�P<����ჴ��~@��i�z(�ho�b��{�Gk�
3��#�Z��{�Q��2y�2��ȺW��V���xO`f0S��\��&�9�v~#����UcL���=�-~����*�Pn���;�/�8�[z�_/�#o0U��@�,}o?=�śM��2}��~_~��U=쎱zO|�Չ?�+ s�����=��v��"t��,T�t0�Vt��+�;W  b����X6�9f���+���a��x4����J��K�E��Տ�j�	�9��I�\��w_\[o#[����&�gZET�*���øm��<�|tg~� �p�7�#f�Oآ�*�/�'�U��%�&�A�Xゥ��d�t���k#�����ވ�:p�t>���T��b�؊�ev_f�\�z����ny_!v	���δ��\�{{��t̺ޮ9�e:��?�=��RY�jG��P��LfKGw��|�ӊE'dxm�V��3�qkea_E>]9YV��f"dݒ��C��tA�yj=4U���r�|D��`֫�ja=�gXg"��w�s�������2�BȊT�J��1]��~K)N�B�&��C@"�`�H�@�f������ͺp<8�y�J�����2��SF��������l�E��|�.�sBph��y\A�w8�VFL��6T�e$�mCMS�B�H�c�`��4\�$`���J5T��1�H�l���U+`_���D~l�GE���Z�o}
ʆ݌ZL0���J�Kٞ������Mٵ���u�$��ȉ��`��'ȇQ�殤D0����Y��쿦
,.��Ge�Y�f� �o2óg�X� �-��R��(��?���x��w>v�$��B�{>��~���ᙛ}��om%H%�w��F�{����6٦$r�^~I|+!y��r���{AsB���K%�v���ʎm�Q�$+�*��l3�1�By4r
^q�a�K��S6�zt���".	41�-�y�Uz��٩���}�8�+���F{�h�	���x��"j�^T�t�K�F���>Tj�eQ��hY퀲�
�ɞ�)�c��� �k����������T���D���:����]` 5	a����n��.-F�Y�V�����f��r�%e�.��Gc��+�]ڕ ��e�Xě-9�X��S�.�֯��%0��9�%]4��hChB䉦KԈ�2!�ꎎ��ʮ�j�U��aʁ��2�]�LI�QwG=@�v�ſhw������
�mk@� ��˭\mA�O�-�h����ǝ�Ra�Z��
<u\%B�a\���6%3�V�haN���`Uy^�h�Q�$�@W���9�Ѿ��DucR����:5{Gŝ��SW�K��
Dө�s憗hT����3��T��ʜ�!�µ�b�>�z5
lK���ux�_�.�Zٿ�h�y�f�Jj��#&;gK�4p�)��3j �틵V��6�#���,ډN!���r�vK!�J��H���ڜ��|�nYp'�4`5�n8�N0T���M`['�̋��soW����r�m�3F O�uu�[V�	�b����X⠃��/>�(��|�YA��ٰ&�y}i��ڇIʀ�����Ѽ���.��M�S.3[)���5	{ή�D %������2�I�/�m�=	�e�7;�'�)_L�_������K�0���{�Y������?�~�a��g��a\V{6�������]t��[�4�
����w��}��:2���keTF���sT*��;τ��9�����b�K:�,�Q��U��G�`u��w&,$#�kT�����b�0����ahn�N֤U�z����we�!ĉ>�03�w~w�ʕYȏ1��;����L-4��B��c)#���$~f+���ZN<zԻ�t�%h7�@^oiK���ˈS��!7�M�b�	� �^���wһ-!G^b��e�Oy�}y6��䓔�n5�.`d�DJ�h\Ԁ<�\5f�MH�(�� �	�WN=��'Q\��.�%
�2W/Y%ow�Y�	��CAo��j;�@'EB�����q������EZ��������y����M���gt�wI/�K�bI��a�&UItyf㕪j�ڧ�X7���4�>��D���;$�^�H�f��ʒ�H�0��7R��a�$@�C���D�0.p�ٿwY�;�I��E:����#eD5n[c��~8)�+0}�.��:ע\P_F��<�A���:wmK�[���
�y�ZLJ�U<�n*�f��Yj�k��eOC���^aޟڊ�3!:��;��+T�u���:)�����`�j��fx��<6]ВgZkm�͝���y�m��aMxѝ���x�&r��������5�ب��L?n xO&������[����9����������D%�)d~p�KH��[0������~���r:�=�.�L�>N���`��+���p=�A����*��;�DYH�k�%�;���\<ne�'?��$_g-s����� ����s��1L�����s@.�F���h�Ʋ���Y4BI�#�/��'*��<�Y��q��+��:��`��,:�o�#��kl�ԤVbi!�/�D0�v�;�t+�/�U�<����pa L|9��<�1�/ngL_�Ix�Yu�/ o�����Tw�~~�O���˧)1,	�)�e�-��)�WP�3�m-� ?�Ģ�H�������ѹ��q�V�oҌ8�*� @G���ݥ)����aY�]X�<YQ(y8#Z���܇����H'����;��U�#z�JR/:��T[	,(���x�*�>���U� �6���S��ꉶ7���A��k{{���"[
LlN�!!� �&�V7~UX��X6�m�(\9����/q� �O���H���DC:-�Rܥ�-l�6f���Wn�(���:%�
��?Kc\�d��V@*��!Y ��K�{Vج��~0���.[f��
s<4�y���v 6ԫ����(���sԼ�.�7����ϋTzó�Xb������ҡ��:q+��
Z�i=��ªǾ����tB �E���(��X-tWBǚt����Z�{i�\~A��`;c�9��MZwė�ȍ�����M���w����#.ܙㅀ'��{3<�|��ۼ������ ��_)A?؉!_�3di��r�G�j��}S�QFn|�'[u��|��>��YkO�'nƁn9K�����
��u�m
~�	SKx�66sY*�X�^k	t�$���Ҥ�Q~�m��V`���Q9Vt�J��h�lJx�)5���?�����'��e�r8ʹ�.-��v�a���);o�c��$�N+EHߠ��~��[C��9Ž�j+=pLs͡�&,K���c�Ԝ�#���jb����R<mYoiY��I1hW��}�ܛ�I��$Y�(#�{�U���$�h���$��z߈���V'�a��83Eq�pI۔�ζ� �ޭ�s�n}�~��g���On��U�	�T&u0<>�$�&h�Y��К�Q|�6#�u��T|ͩv(G�k�����t���;-�*��+	ª1��Zx����z`g�lF���nR����SQ��WԾ�#'g��,����-j�v��;)��a��	eA�!��"p1�nV[���<N����#e/���r鍲���ǯ��_j���_}[u|3�/������59F.�Um�=	 Ic�	�I,\��Γ�ط���6q�OO6���x��Ȑ ��J��!1_���0���χ��Z�u�wJV��a�D�Zm����	�W0��m����F��~
��Hy�W������Kes��w.l��bȋ�YZ�3�M�ذ�*	{��fw��3/%w����"�Z?�Wq:?G�w� <x��B9�~Ai�Ǩ�v�°[��8�䯳ϸ.�ɮ���iI߁����q�Їz��I�?} �Y�#-# Z!����M�n�Ԩg�漢Ar�Q��M�cY ����5�Y69�Ag<T�""�5�d�C0�70"�^�i��x��ۇzC
aV�Pþ�,@gw�W�=X���9�s�1_vA{��@.�2��f�l ���57�\��I�h7�fю����u�XZ�6S&�w~IyM�07I���@\�-H��e4�w�'���8�CQ
�Jӄ� �b���%TO_��Q�`�T�lI krz�YP����|���?�e,
��X����*<��ϭ{�U�<X�z�y�g��M�u���$��F9�	�*�4��ԗ�8%Gcٓ��}�h��kBF;�z��f��_F�I�SH�-�I�d�Nt]���ip8K&m��k������(;��p[������˧�rȁ`
��H�{�u�bYZy��
)�a�]�C��s�М�{�Tj�R�(��e�c3n���ό�4�W$)o/�>Ә~~ �ʡ�Mp19��9ր8�d3n�-c��j�a����?V9�s����[�$��	^�� �5�7d��8Qo�i��3#0�Ҏ�:�A-:��T ���VŚjD��Թ?��z^Ա"JK%���<|��7+�l�I�`}LTd�9�hX+=L,�mp< �h�ʟF�x��L���䡴 ˖�R���� >�Q�P��>����@>�Q�)53Z͊��b@|:� �*�����z�%$`��vNIi�N���q6�S�m�N3r�h�{"W.[�;�-?��J}�$ ��kU-ig�B��&��}��FO\�LA�(g�.��2>H�zQ�wM�#r�L+������o�k}mM&��Q� ������{Qpۯ"ϒ�S��mQ�P���B|,����ֳ�����0��E���6B��l�	�����ݟR��߱QM�k��J�ۭP63�g5��o��o!�(7v
|����! Ȋ2�hܺ_*�y��yk��l�������S���%L��A�7|��VF��<�v
u�B���pc�IwL�+a��m!��E��2/v h�4Nb�/�0��s��<a�������yi/�q<y���������>���'-�[���o�"��ӛPG��&k�݆���D웃WPO����5*Wy�����0	��c�aA��EP���ŕ�e=i����S��4^�^�`�c*���H�@�+���XS��V%����n)&D���_;�5f�s��OO��fþK�e�I���������� 1���8(�f�l��ँ��%,UT"�^��A�I#"��@9{qY��$��@�(�]�t4����[ρ,'�źjJ�Kt�J���.�Η�ox�'ﯥK���w���= �ì�-�;�n%�� ��}�d����g	�l��q��-&ߩ�"�>����7��b���Ck͋�H�4ɘm�ѣZI�(e�9=axB}��ߥVy*��Q��.�R��Lg�,��Hi�w^ܳ!�_'�$��Ȱ�5^g��&뼁w7+�`�K��w�Zoq�����6
%}�~���۷��Ls�b%���LԬ6���cq?\ڊ�N5@3���_s�Ư�_F[0-�������6%�4��5H�	�>�u���p2K��۳vTd�0"����X@G�sOD*�+�����(���Z�~eU���Bܞ}�E��\ݝZ�_p+?KėE���F*�\3����Ø�P�O��ǂ�cV��g$%��JI�ү�@�f�v��3Ԯ���b��˿7XI��ּ�e+ar�.A��d�]�k��O�P��}Hi�pZ!�Sͷ���B����p�{����6�D}��g��-��=�w�)|0�6?�lG��L�cP�b�.�/�@Bj��ƫi- j��ĥ�{̵xf�?-�ŪX�q��g��.f9�d}��x+'s"'%���[�����6��2�-���%��2���@L3�|r$s���uS����+���gȁV�1*T�{��[UL��P8}}{[?+x�	Sk�WQ����߄�[Z�}��_�;�\>&�e�r�R8���Ѐ����S&����� -�f�`5F{cP�iW8;���� �eK�ѓ4�㤒�$�m*�h�a �(��ԛV ք�Vn�su|a�������}*A3�g�M��,)������g��]�zK���X碯&���)3L��q_/{B�O����h.�T�-���6ͱf���H�1K�!++lV���y���єKJ���Xâ����\�����$���Z؝^AH�-a�ZH�ʶ��]��[��ߧ��IF����~�"+>��&i�:ÿB�U�!�EN'���ƶ̛��%1�,�?���x�ӻ3�;3�� 16ֽ�h!]�c���!��R�r�r}��3�W�H횩�W�&k���a"LQKJ9�xg����N���j��/���Z�K�@�l`���R��EZ..*>��I�Ǯ,v��'D�_��%�ā%�Ckؤ(V/��:�V4d&<(��"@m�3�ۙE�^^Λ,)%%�N�^��j�B��wdB��u�"�J�u��!q���g�_pY�=�Pt	���z��8��C@�5['�dz�iA2��5�Q�q0Q%u���Y'j�݈����8��s�:���c�<lh!��dA�|���F�o�)�`�����0����h��,d�6�;r�  )G�#$Q�+NYK'��v���Y��_�"czi��w
� K�dg�GI
n1(t��Ø���+8DbS
N�W���u���9�Э�S�W"E�Г�@+��(z�4��O�4���	�jk�G�.&�Z�+�TG�v
.|��a�8?�uB�	D{~|��ȃ+��Tz0����*$����e�ȳ�Ί�w��|p&H^	�/��y�U���v9CGgZ�T��^�x��=3�2���c7Kc��U	ݦo���0�䑅:�ȯ��
T�߉(l��te�(HƊ{=����l�-�K(��y�C�k4<<h�H���v�i��\������q�y�%H�� ׳�3��V��C�$�&b0���΄+��?�o�X����I�� �Bΰ��3���ꨥ'UW�\@��9[�����4Y��q��>�(�K7vG�!����/�g��2 �wMoi�i(n��*�M�M]�|����Blaˑ3i.-6-�Ϭ�tb�]�!�_S||�^���B�ک��>�c�����u�USV����Nv�'�.13�a-Yc}u=i2�|�L�i�]M������9����CU{9�A�
o�����RM��|����V���w�0ᥙ )#_�Lַ>�����c��3H���/;|���T�i�����x?����G���Y5���x7�6&�����@�J��.��~~c~�M���ws�O��y��&:�B�}P� N�˻>���ȣ_W�f�*�'�/�'~��������)�������;͒J����c�DR�O�go;?������S��-�������+}�������p�r*�T?�^�g�#7ߐwx`e�2���(�=u�Bw���Q����k�&g�#�sDQ�pn{��z9&d������c�q2SADzN�C�|���A���QKj����휘�iV��|��L�����-m+�"L&M����JȤ[iqNm_�Z��߹^t��"�H\|i-8��}� OhXz��F��KN�/X	�kHT�h6���EZ͎�A��]��PF�2Za!+C�)H�Æ`z�=���Φ�=A��v�+	��V��:A	�'dh>S�~v��:4M�in��=y�����AjC��HYQ��Nx~'����F��<X�NQ^9R�w�<<��_���b+����@P�+��ekt-[������w�f4�𭊢�z�ק��┧{�C�J�7{���Y�X{���2�&�@Z���u)��6���!7^��i�z��I��>h�ሃ2����VD�3�X�J
]�U���L�����%����%�c���|����A���˷�M7m�g�a��;��<C��F�r��M�ŋܳ��E�9�&r����!2NREA��'p� L$�J(-�� ��74;�0@��/�ys�0���T�5n��ޠ[�	8�J}��`��x|g�1��QKs|V��&2HT?X����cn��Ҕ
X�O�U	��9�د�[-r!m!�s��E��!VN,�0ː��Kμ�e��N�#��JD�M��ĳ@DN)���:
Gp6�te�<�6m`�!���'p�8t��?h+�D�u�B�Jde���8�v�B���!F1Qʁ���Ze�v$8�J1��y�����wy����q�9��OL�WCT&-GB2��QwV��w8����z���vg�cn<��n���Q��xC����j��p������!��9�
j� � �_�8o�����fpr�ɖ�3�gV��s��˻��5��nmZ��ht��n���
)+=+�v��r{�~�p�|�%��'������4v�v��^x����G�׼Σ�$�!0�Q'hmՏS7����a'�Y��d�����&���@��Yx�����A����{���L:�ݹ��s_�2C�&��J�����fgSCp����W�S4�l���݆T�&���p2܎G�C�f�"�� rx=_��'U�a6U��/�:cnKLz.9/�^�F�ﻗ"����(%Q�(���&{@�5����P�(��k��=����:�����;}Pz�HRZ�T#v�4,����P
�q��e)�ٺ����ו�%�r�T(�w!v~�iŔ�Ԙ>�ˇY���/�\��=B�ĿD|I�|��1ء��b��r}�E�b5k-�g�������L��B�� q.ߴ/�F��MI>0�SȨ1P�CD���	��ȣ�s�xj�"w��%_�|b��G�*��c�]Ҁ�@`Հ�;^ds7s�]c����I˼={��鸪d����լ��nI���;���ߴ�	Z�uz�&��U��O�Î��jN����h�����ΦQ�e��N=�z�-'�Yhӵ�}U���g��y'&��_>Qd���c�I�c����ւ���q���[M���6�����a:Dc���i�8��L< @����x����M���Å�Mv��X�g�B�䉋6��.���Qc��?��ɀ�JgÐ@�N�@_�q)S9�v�T�b-��o�ޮ�_2@��j�Vd"�|���s�Uت�O.�1 A*�F��~.�i�|�N��4�$ݶ:�I��9�B]. �	�7z��Ѱ�w��23m�l{x@��U�<��Ԅ�I�d��vRȵ�d}�6�֥�o��6�NȄK�?5��)p�����g�Ac�C7"��-�hl�Us�"!��Ü	�e�2�Nrޑ�udA�M�D$��zCj(�"?�A�6}b1� �`����e��Ү|�>����j�;H�|nOS(���MÍ HO�aI`G�铠� h
[������ɏ;����.%��%�֯�@��=�5��Yt��a\v��ɛ�	�Y��E��#�|ڂ�S��S�ѝ�M�Uc3����x0��]��QRXI�n��藢�+�#�Ԉ�p��^�]ʂ�/�x��c>�K�B*#��M��c��G���\��O����!�؋2}d�W�Y;��v���s+
3�m�:%��Z����if
���X�x� nx�z°T����3\!U��������Yf^���f� ��Ԑ44�6���迶��a1K5ht(ݟC�� �� P��]�W�����q0�`�!��elo������)�H�^GAQ��	 �r�D:4��� ��°"�ƖVoe����g��^8��(.��@��&Җߜ��M39=��8�����kD�?��M��7v,�}q;x��+�qtsX�lj�y[���[��8p����K������jK#���pA��dQ�A���t
�y���}<�"�w]ܤٟ����Z�&�j-��վ,,�,���0� ��=%2y��ո����94C��>.�Hm���>C����v�G��%�擈��l ��hxa��"�t������~Ϛ�f��"���� qn7ǶS���
9��IFq�ED��l��^�Y8������?d�L�#�ڹ����4�r����<�)���Z��^}����oA�~�V{���O�%��^�hg�)Q�$N�����9:4CB�F�9߰bѭA�O"����TP�E���%�ǒ=0�-_5��y�Y�j�;YV���pOr)�v_�gt��ތ�̴�
Aҗ��[7A�o�\*L��� A��*����,W�tê���(S�f*��)btN�Fh���{�c��IQ�w��z|�)�߯9!(ӫ�͙E��8J;�po�<��c��`"����s��B������ �J�n���{�Z��-$�^�#������������K���e�V"~��c���o�V/�+��g���8��1�1�;������Lת�_~k�x�ۖc��n����P�w�z�h���O�E�l(.��<�����,
)�H_�Ղ�`C�ڲ�a�m���k�J�"�GV��1�ȇb�%E_��Vp^.7#V��$�X�3<��6���)�d<_xp�
x��@>�Vy�w�B��/�Y�L��`�]8�:h���	�+��o�
�������"=�*��g��Kq�"!��w `f&�:�;fSw�y'�x�e4~�7
�߱�Jx�rK�ةf��T���8�O�����;A�oԀU�����/&�zl�����*�刔�QZ������ǹ�gS���"�-qx'��!��J��zlUs���e��z���
��a��:6���I��W��)#��E�c��O��2�:���O����ƴ�*tT�4�t٘�{���@$��G�/6ɘ���+\��m�g!R�VN�ި1�ih�E�(�fL%e�� O��|�)>��R��>����	�)��|H�{o��-�2��PpC�>�t�1[� o�|�Q=_7����&*;��GR��?�*c�@����p�s����;�^}�ʐ�
��*h
�CA��1��v{̝�G�~���b���hCTȝ�9,�mo�ξ$�m�~��IE�2��2S6Ty�Os��Y��� ���6��׋IZޯ�\�M�������v���G�8qK&�O��]?iw�8Y��!�]�����ۊ�h%l���?��2��L�n����,����).�'��X�&�Y��n��|���W��x`|@X��:�p��>HV�ڳm*���x?T[���<����]m��jc9��U��d�Ah;X�x�m[�P��3�Tj�H��=��%�+�eiECx �`"F�+�e����[�ь�>?��O��V�]I�㟘{�)�HH��ab�6�c2��"�{!� �I��S�J�Ї�5l��$T�T�\�@0�/�(�zt)����	?�d@���-zIj"{�0|�J����wr���C�U���/�u�69ΰ����wIT�P�l���J�����+9t�i�����ϕ+ش'�:ś���Y^�➯�ȴ:��B������B,����!�|/58*OJ����B�C@����9~rڀ�o�9������N����E��		nyyؗ��}.;��ڹ����V���y�������2QV&\U��\�<ք�m�u�q���U�CUDlD��O�kȴ��74BGgR�J�� sFT�Y|2LV=Tf�6&��(�oRP������kƘC�t����%>������W�B�G��c��v�&~�7��N+�5)��=�h�!�F�qv�,�]�'ܡ���+�����Cy�Y�T_%��3�g~.�mq|���_g��(��'�5�m^B���u��kb�-^�7�rqiv�
���g)��G~w��A�Z��w{�mr��'�5n�����6W�#���Cv7�Q��
�zϣ]�ŏFH�pF$MYG�͗t�O%�����rg�6h�P���=I��I��^���{Ӓ)�c[ �&x8�������?y��oD:T5o=B�Z����X!����ʊ?���EoA����/��b�4��Whj�y	�Ѓ�C�W#8���N/0��6VNOWF�W1ړ#�ޣ�~	�m�+f�-~Yj �:�V����24߹�զAH�V������
o��AZ�ڗw��<����/�̕���?!(�j;���wU��>���#JR�t]�oY<ϠSM����Ѹ8��Z�p�y�*�l�Ҩ���4/���#��a�H�ru�X��mu|�e��_����K�_"�J	3	��Sx�)¡�m"��[��#O�9�b
`wC�n,��p�e#��Ya�nw���d,�k�l�[d�ْ�-��U�?@�����Zt�p�)]qQ��*���7(9{h�:���X���x&V�?�I"�{�X�~be�})�()�\+s�4�fD;U)�p�==s�j����6��"-� �~����?�{�,'�0R���Z`HYZ�u><�R�����͸��`V��R��uR�*qD��oщ�B��Ta8�R���9"̪q�؝�b���S�����+�k.�� �2�[r�&2�;�[f@������;���ƾ/�a���o�H�W.;��z#�e��"�ȕVA��v�J.E5�L��,N~�G��)���..�/�����t��IT:=��}�0$���iN�b�8.m?�o:�<���<qk��bt�E*s�d ��q~K#�Vi-�#��@MjNT�|+0'}��$��q��u���'��dtR�0]�fi��J%4��O�;�w���X����dg�&e^�
�<���f��THj��VH�@v���6��V��Ȳ��}��Y<�Ru�f
=|��̥����n+,҇A�հu3��l����x��9���Xڊw�H���/x�[����\v�o�t��,�-�e�E��udf���o1U��j�Fgƍ\w���8��ź�ɇ�3�o�+��f�1|+N0KVG/�TμR��֊��ylTu���ѽ�^IK��h��PP���ݞ"6e!�ma��77�p�$F�89�(~F>Q�e�?��/IpҶ޾���&�R�U��r��51���l��G)���!yٱ;����
c�[e��`�{���-�4<y.����|��F��
�)3^�Ǘ����$>�q(���#q�@�)M�nO���Ax�5 {���p%w��{)�;Y;P�b9�`P���V���R�a���L�����(��lf��W���UDn6���uj@���F��j��_�|�m��6��m�����C��ʌ]�邁l��ƜM��r��|3�F��'�_<l�{�z:�B��SJ�%�
Z^D�a��n](U,U�$��l>L��J*jY�5��0��,!�WB��bxTa�1�	K�r�dά�^x�輤�(S; �@xC	�+�-��ڐ)� ѝ��*����̞��U�������[J��Ϭ���R"�8����&�U�]9m}=\_w�5l�C��݇ڲ��îl����j"��3��Jc/W�/��C��y��$�I���6���0v�ײ�|�-��Y�ңM4��� d��[d	�:
��J0Z����$j�r�<޵��~����ACXS�B��5�v6Y~:,��R*�T��(��ʕ\/�KH�!��X]c��^��!��|L齠*.��m�H^��">�Z��kp�Ƣ��i���/W��8�g�Ov�#wc��	[�/�k߆G|��F�ZQICG�`YCi�/3����s�������	�ZB
�����i�F��]w�\��l/�ޏ�lgž����HZ���xd�z��"G~�N�4G��?=?���5|G��:T�0�D �0��f!�� �_�3���U�Sz��p���;Ju~�'}���lL��m�坶� �g���Sΐ�B���-�bu�uI�Uh�wV���@bD�B�J4�e���'S��mqwJ�5=��t��/~-pt�T��i���a�U����gǁ������<��Q��co#�j�K r�|���&���y�:�t���ǮQDa��`�5DY���]�V+ti0�g��ĨQR�.�h]py�D�/2 -{��(�#��H�|��N Ԓ����p5��#�=���;�}�v׻i'�DQ!��:U��_��Q�[Sp�`܁��j�3����w�}��ʂ���Z(O�؏d��f�ޞ�{��X9�����5���*��X��_JSK`H����	���=�,O#�6��=����~ 3�_;R��Z��_3�7�(`!+�x����$�ߖU���w��ּV��&,l�K�y��k�>��x��K's/>Q�'v��(I��77\[F�:������r�>co��r_Q^Bd-��g����<�7๣�}��c����f��'{�)�����@̍�)��3M^{EB��oF�z��@� 5&r[����'K�.\+*�y�֠JU[��� 7q������Z�W�_�RR�Hamj��0n�Ci�	���O3�������b�Ɨx���7�X(�W�ì<�[AH��l�K0�N�^���0A<C�v@��M�6��uz��Zm"6�pY(R���N�����l��ſYP�����P����a{۴~� օ �&��������=ۋ%$�]��˃��"�ͦ��4Qi@�夣�B}e�����cB�����f��\��S�N�H�a�YV�b���%������vz���'!j�S>⃙&^�)s����p��W	�Ә�5��ک"f4O1��	
L7��ӈA�ܭ �W�UW�4P�y�0ed۰W�
���%V7z�r,>�',gN�\��qC��3���9	�{�.�p�Sٚn�;l�U��ʳb��� ���t/�l��0�1Uջ�_Fa��Cq���h���"	��i;K��ec��P ��Bi48|g�o�j���� ����x4�綌��Q����.Q�����|�S�Zw�-�#�
>���lU7�葷*��P+WqC��[�?��+G�B	`Y�Q����'-��ǃu@a��{LQ�H����`�7�:��AW10]�0�]���;�\۫'���#�Lr�^�@q��Y)�	�lYu����8%�>Vz�rQ�n�-3�6��5g�m�O�I�	<D�l{�S����ܵ�_A�9j~��u�!�ۿ����m��ѱִ;=���h0	�Q扴?�1/����vd-�>u���
X �x���xŀ$�2Ο��Qz3��k�]����\m��"k���=�Ҫ�r���!�	��-+��9<������� ��6 ���¼l�ѣ�v�Я����Q��'����B�{��.3џ ������5��5��[4�$n���Ҟ���.� r@�5�yx���+yR�����i15��6���+3�ꤐ�@Y�S�!boN�4RĲ���G���t.�Q,�㕴^�0�b'cZ�Mj9?}��L�Jue�q�b| �al2�3�������h���΋?��v

L@�����̔��{h�9�̓�q�´��T9��7A!Dnge��m`�I�Lg�#5͌�}A�H݃Dn�G ���0�zNk!�q�-�7��]n���ߎ�Yg=���D��sU�Y�?cM���KK��J,ox ���G^A]�$��lQ�	�8nZ�ve+��\r'5���,ul�d��q��~��������܋�V2����u�s������Sy_g�v��ڙ�3�*��:r��%��8i8����0pb�f~o�Sas5�ln�Ŕ�ف{�%u2���}�a4�?n�D8BH�l$Hɫ�����G\�aͷ�M��lLp��_D���C�AU�$�7���s%��;A�p��Ie卵�3�r�5��h�g6a���:_u7[FU��	�@�̹	�eS(������ր���z}�9 ���.���<#ö��2I2;&|��MU"�.�0�Riu������ XZ��t��(����_��iN8�	�����Oظ�Zڪ��,��?�[���}� �T�5�-����"Hu+!y�2�(%h�\az"��}O� 9��~���M�U1;�=���� �9�IGӴ��$�XKV;���-�ѣ����r2�$�7z���ײ�Z����7wp���s������a]|P�q[7�1�^��R���^տȆ.���E���O/�9U���&��4t�3kJ���S,z��$	&�C�kF�u�QS�"c\�?�A�H��
er}�enu�e��J��"~� ��|�=��A���b:G�Ì%��&}�^������`=������w�=��F�dAaNf�D�Rڨ�KΚ��u�A(��;��_4����y�cx����Ľ6��F�b��qӶ�4;�6�������"�K}�5��Mu���L�.�OH<Z�
�x�o���yG{�$i%@4�_��?J�����v*��E�ީ�ʀ	Ĥo����lɘo�s�����s><��9vVW�E4
uX��Be�v�g�}�E���&���q�:����0
���&OV�傩���Hǩ.�y�Ż���ѹI
K�Y`~㨍�]���L����ɋ�jv��r.���zc�6�~�op�,;����A���M��
�>�>��?����l`*: n{j�&uf�R0�M��*>V0����	� �r7�NRDO`m3�w˝*\�����v�7���Q91Q��.��>tMq������d'�Q���
�vAh�2A������_�d
0Р�~�0{�͵$".�r2Nw<��E���	�r(R2������h��������H������Tq��5)�@u���
A<Fbd/\K1׋ %�DS��c>Mʲ�
�;{:P��+�j��?9+�E���v�6�C�y�
�gf�픇U��k>G��'T�e�ga��oV��"mW�T��V7�b�Q4އ�7�]�	A�-~�d(��{���<I�,,pZu~��,���U����-�Ȩ�9�w�qH
|��f�|+s\��!�o~<�dvc�̲�E�ǲ;����`�T�o���r44D�WOr��)��9γu4ӆ����ܧ�$pi�	X�r����T��<��R1w�a.0C�{�1Z��:iV�X;�E5!����&�%Y�����*�'�w���90�bl(�WB-M�>f�Wܑ��+�1d�S�5�H��~�Dkx��"�p�Gt�`�p���U�<�j���^��x��Tz,R/;=n��Kq׫�A:ԯ����Б�]����P�eYN7eiF�ZX�_u�m����i�~�\_�!#R8C;�Rtp��	��8�ѵ�:W͑{�E�PS����s���n"b@)���#A��*
�+�C����<���m�=�0��a�g%��GJ�S��ֺ��U�λcٴ5H�. h��N�s��.���^(���aS0�"����g���,hi�@�
߇c'◉��g�� �
���]s�s�feGnņ�|a� Ϯ�$��ㅴ2���N��+Z�u��8�Fa����v����R�)i,�]뼀��2	Y�c,:���{����n��JA����:�\��Ȃ�����ġ)�w��o��.7��"�Z�в�)~�y�ӫiM�Rx}��uM�Ц�x�v3<�a鯞+˒�>��	�b÷ņ7?gY]�A�' w�Ie2C�?8%�5�� �fZ�gH/����ϯ�bp`w�i]�a3E�����8�A'Xw��LD�� ǼJS��d�Y8�W�zg�Y�bѧV�>z�� ���L?|0�C��TǲI�tS�+V��+�K��P^�oK4L��<h�����- 02%��{c �_�̷53k����d2�3����g?!i�A3�W��w&�����<������L���0ܵ�顼�?��h!4���ŝ 9䪃@;u{�7O�_8��&=r���B�/Po[H�����s�J�I|B����$���O�Ը����L��$J]$B=@�mGW �@ )6ل�ibԟ����1ԛ�_N03<������IW����6~]�$�n7@ ��5�DȪf�e�ɩ�D����~"&���d��ęy�l\Es��y�MF�|�|ᘶ�lXXO�ۻ�e�wO��~?�����ڌi�9������;	S[��x��2�u����K ��!��a�%BÚJ�B=5;"C,�a9�g(��[h:p���[�٫�8H_ �H�����b�����e�����U3w�g� 
_o-��	�����i|	�&�����������D�p�]�t��6��O��l�+�U��
��<!E���C��+�0�Z�Qd��Ӆ�x��-��`4lҒ�<��s>by�����gY�A
�*����s�8����S�G94x�����-�ڇ�����BƤ��-�K��G��mW�lk(��!H�fh��2-A���ӗӀ���@��)mL���l�(	�M'e�I�l�i��;w9�xO�B���G�"��!w��_���T��}�}���I�I��+Je�i��{w����48����`�F��y���EI�Fg���{Y��h��#���r֐������}.���g��u�����k��&Q9$��{�/��6<$��]sͿ)0�zS����S���Sqq��T�Rȟ�H���YO1t�� &Z"9�^�4���e9�	|���k��1HQL�}��7��ۡ���iv+	z'�;c�k���U5�[C+���樂�5j��r���h�>&����`O�K�������u�@<�k(�����J����O�7*:ڥ�c�4�f�8�5y�x(���*��R]$�D�����6I�J��^�" ���4
�Hўc�#
��p���d��kW}�|p:��&j�"$!(�U%�*�Z���LT3��s(��Y����jY)И�@��|����b���{E�RTZ<6F������2�Z���1�o�Y���%�IJ��"��O���dr�9��m���6s�Z�.��$1��$��3^���y�f���ˢ�)��:-��h�A�8��)K�bՁ%e���}\���+B�.˖8~����I�� 2� g� �W)���Cݫ&������P�޳9}�S���V��M�{���t��,���ǰQ�M�~��� �[*ܓJ�!���G��xfB̈́*�#�Xخ��;��cw�poBq)^&Յ��vz\��,scջ��f#1Vt��!%3�,�%��~�~ז��yͱ^��׫p�mT�Ŷ�I" kʆ��@���Z�!4�8Hn����g}��d���xH�r�Z?�z���y/_�Y�ɵ2x��	�Y����(����iz�kO�[7����B�GMTY��[YZ�[換,�$L�7�%��j���c���1}|�< ����s�H����=����M�	m�d�F�H?4��6�tT?p��_8�)7?��2Γ�8��벖+U�Jc�k��h(��2g�,�{8ޭ��M�������97�����H�qw�����!xBo� ��e'0�m!�Fz�Qrxޡ�)Η.h��DRs�Cru��rr�9��Q�WA�m��)�N��_!08h�I=�΂��jA��(y�Df��O�|o��w<-V�hŮ���lu��	��D/����KL���k�O��a��9@>ɖ����������q������ J��i]�oc�G&��N���Fv���\nt8MW-�x�K4vR[	�Pw �cA��8s���oS�����a�
	!��V��s�;�X��Ӿ�o�B�x��}��=U.{mp���V��bB����X�5�ݑ:c���yb�~_�*ߜN�+,�W}H5�?���Z���{"�;{�0	���I&Fe�\^�Ą
�cԪ�4܉?E��ҁU��Jo;Nt���C���E��u.�0�93c�RYJ]	U2x ]��H��j`f �"�ISCsH_|�<��vE���DN���H!��'��i=�鱽���,c1�l{�1�nL+�/�yh��;&�s�M�5���4�����-�ĤZ$*L0a�������5���U\�nX�@6U^��Hn�^����EW0�-�'-��n`;[.:Q�Fɋ's�A�7oA���3���_��R�1q��{��ǩ�nL�y�{o��%G�ć_4k�v�uϜu.�<a	&=���A[����ο���I�D�Dh>�qU� 
܇�؁മ�?���2g(VR7
���i�%��L82����Ved+�d�?N�E����I�mU3B7b��4��N�/(nZ[[���6�G��^+Έ{}����A�<��;��w�!���b�,��&�VX��zR���H���A�]�c�ۛVx+;iC�,���H������P��	J�&81�3-5a��i��U
���J�D	wīx�@��s�O3�n�km9�a�r¶K$�MQ.ݛ�כ&B�V��"�!�(�u,�m`UKf�:�\���u1�;������.�PN~H:���9[��h�l�x�8+-�����B���>����.>K��)D�*�1�ל��C���`0��F/q���ZK{��� 8	�{߂�2!��ʠ�A�O�E |0eI��'�΍�fe��A=��D�D�L�� -s�K6�O�)T�-֪�"JK>[��DZ޻���M�H6��En�
ljֈRӇ-|] �)��J����xׯG*t��a]�S���;��*`EK��� Bt�y��JG(�/hY_�y�'pm��!�x����^{M"����yt�������1&)�:_�f����3!����`ȁ(�@v����>��d%'�냳�tJ��y/�uͦ�@��&���)%�� ?Q���5��Z�l��}U�4�ǈ�q~�V<�,a7�o6 E�MɁDNH����v��Q�K���H���G�����W6��
v�,��.WtG�%�@��*&����4`��8����Q���l�%�۰�T���t~-�g�=S��7��:@� ��!F]���K�A�T��_^����t�v[��s��@	d��#/a_�N����HVj�5�3�Kd�z]� {5��Q�������0W�����I�{	�lM=�
���+jQa�N]���E:<+s��7�@_�����鬴	��c-'�`�I���v�F{ ��_�N�C]�!�oE�����)K�[	���!�� Nߓ8bT�/l����\J��.~W��.�L`���	�X+�K��=�Qz1��C���[;��p�Y�W�7��"e]enR�V���$��_4��h������hK���t^I�P�fiY�b�4qC��X�z0T����c����V'�����=C������:�ⶶ�%Ҹ�A���˼U��V�L���K2�e�>A�@c�MP�:����r��x��[��O7�a��q�^��2��أUBn�	�|�_;�;�)�<����t�/��bh�wz�/�&��JUYa*9��Ҝ��j��?����F��c��kV˵g����ĳeM���|���׼g�	޼&ʐ��s�U����X��5Ԁ�5\b3-���$�q�P������
�F���']�0�<љG��i�ֳ���*�lv�^���QuMm�� �#�G���I�'���t�q4R�F�.Bd]�����yr������ڝ���A'�*H�}��l�)�F4r����qǙH.r�|>B=�#Ӣ�q�w�~擥-��H8no����<���S�!˅=�3���3��� �x�lz��7�*��L��U(��V7u�R��q(������Yq���qheأ�e�����g|��_��� (DXA1�U��V)��.o �N[XU�f���&���*R��#H�~��"�"�P\��7�-U� t�T��=����Q�w�H�'Lp؛#�������};�D	��:��X3Ef(\&�E�YD�}��t�l	��h��a���s�K���.�+����v�J췎b�ҿ���YO���{D��sU��&�i�s���E���Nl�,PE:O�^��ǋJO��\���#(��jf�)��������@���,�r�v*�OӚR툏�b��XS�0F+3HʫG	8�����f'��@�J�|�JL��Qс�~� �R�lK���a���)wDA
��=j��&�E�ք���$�s��=b�n�j��2jd(:ճ�G����[<���:cJ��wE����������U�Yv�2�v�
��C�h+?_G�*�K~ئ�yK7�����%A�m��񲳩�Q��f���n���2�]W@��ی��8Jp�1Zt���LYG�.r�*��Я���my���Wq)�7E����E�& 딒��}�O	��C�m�8a��仺����V!���I��)F�Ode� 1>K>����(V�����i���fp1D6�Q{��e~Z��ͫf��X.�o��������#�|��RO
`��a�7�.��ܒ�3ohh����|�(��<�͊ln��Sm�������~� D龵F).��W+SHjD}��ߛ�A���[�� �f�Q���jZ�6#7�[�x�$�ut1m�ش�ɦ-"�R�Q�V�"C��_R,6
Q�!���x�B;�#o�t0�_�W���\��t`jh���f�����lԭ'�p?1�VD�9���������¸��1��ͽ,Q���C������T?�,��VJF�b��!a����}BO����Y47�ߏe1c(�D�X���V����J_�79ڐp��	�?��-o�T
�7�g�����n���Mݕ�#Dml%�CQ����Vë)��
��DG e�s��� ���T9l.uj�e�ƐR��-	ھ� �^������}���$��f��H#Ѣ��\w+�P��͠��ǆ��_���^C&��z�Q��6�@%t �qm�-Ed����=B�G�L��(Fw�@���Z������qb��p�g<�g�����vD)�P6J �ᢟ�C؀tKj�+��;1���� �ji��)X�{8�,�?�⹬m�����3���I�	W?sJ 9����\���e�y]}��`����ݻ�=�>p4� =�P�r�#�:�pHz�2�o�4 �:b�caDЇ<�4#�ɄU�=�.�������ᔸm\������ϐ^�y��,^�S�ȷX�w��<���>'qv<s����>�p�Jd*���h9!���|�>P�ڭ���$|R\ez�8�/ ZK0E�5.qaϵ_��ʩ����"��~sI�����2¿Jħ�|!��ֺJ���j���n}��0��]�-�����}BE!�W���Q���i\@Uƿ���$BFZ<:�1:��c�/��������5�{����5P�1��2SGJ��N�D��v�<��� ���rF�K~����9�����k��˭B�43ՋxE �#������"$%�W����w� �.)�ϗ��pv��
���\[@u���)&�i�����{�l���H������Ӄ�S&X��6�F���ށ5����8�%�Cy� �#k�w�ջ��0C7i!�{��yk�yb�7m��"؍1ώA���4㕙�p�k�Δ��+S��5|���ʠG�}�g@1�>�5.5��ٲ_;4";��>�-ަ�V-�LЬv`���S��(�ts���E�xO#1��K\:BY��Yl�Z>`��D��%��dg��ׂ�$�hM)���)��\:����Z?lfc!�Ћcs4Ԁש�[I���eN��Pw�C�8v�
�!]�kC��\#/m{�{ZǊ�	�)����:��ԫ�������
���	���dӳ^7q㫸��ޣ�C���+Ǽ�H9ogQ?I�c��q�+��6S��.�c�'��d\�.X�ׯ-rPr�dcM=}=���;��s�G�Ҍ rh�)�m;ISS�]�Q~MJf����bv�Y�� ȱ���~�]�|m:�>',��>�����4-��E���]���.�Ha�F�i�²�%�fn�S���&��\!5�׺K$^v,s�3 �"M����dU��h�qċ릞�ˀ��H �bD���f����ၜ�c ����H�?V���g�NV�,��0�����D{b[�M4̽���p��i:}wwK����H=���X�<��@�-�y���dD\�9�,�pE(ل9�	hy���au���I��<�O�����v��@� p��h���;�u�D�p����$�gSE�+�*�1�Sz#WVR��֌�l#oi�,�C<u2ֆ_�(�(�i�8	��Mr�+�uq�C �Z�������1�K��Qp��zK�/hө"�x����qoݟ��~p�Bl�՚�,oF��拔#*5�/A��Aݱ��g���V�x��wĳŒ�̓}�Tz��VK0�_`���@��g�p�+W��B1W|�;��p\�G=���0��f��Ѫ%���n��iؠy��5'$gn!L�sE_�an�zTW���e	��ؠ��o�%��-�Y����H�V׆�	<�������_�l3N%3����K�E�W���
Ȃ� !`y�>�q坧2��vuz#6�#^�#��C��5�6�D�A�7l�� �R�|���5�X���i-��
j�M䫸���N�k�	N's��kk�KM�P'~���������ʋ�_^�'��м`)��;U���UI���(�D�TA`��W���N���7�&�ޗeq���A��V^e��)�T���e�Vy�ID➏�vD��׃�Z0�b%bY�
����>��V�-g� �i�j��N�}�JV/$��h�
�m���0���~)y�"�k�wQ���ERR@X�<^�vڀ����LN�4I�ع�8�(iRP�א8��M/͓9�d����������=a��j\�l�e�W$�{X^8/,7�JP7��;����^o�"뷝|n��=��y]v. +o��s��8\&!�Y��!��B�s/T �uw��ӫ(����+��u\iy,O��G ���� kG���Y-�Y��` ���ae�r��h�SBuw8O����F$+-���&�JtT�z|��Q���6�'G����M���BI*u�8������'�L�-L>�_g�}�U����.-B8$>}`'�R���	=�Z�b<
B ���
-��>p����!�Vm�2���j/���r�5aσ
k��Ίp��R�TY󏝚�B���I
��5��� O��wT��l�Y���4�9C_�]9�T���;|�����2p"�B���o���i�Y,N�k�r~���\��/�w"o��܅y�L}��[��2\���b���cב���MkU:I3N����g���E�����a,������lm��ì�hsH�v�e�ě&�fɔo1Q"���8�e��¿�j�D��['H��Ɩ]�0�%����K�/2��T~i��D�E���g
�)�f��i��˙6�E+�����r��6 %5�(l�q~�+mH3q������?�R�W�~���.ţ��p/ l�_�%ر���/:��&?�\-����S@��vg��]�����F�/���� ����ȑ�����=�����q�SЍ�t=J��6t
,l{�>�6��:@��eە)��1��`�-ݎuo�o��"P�������գF�[����l��t��+l�>��h�`,�C��4���{w'��:�M��}UnDwT�e�T!t4��� R�1�b��+S� F���=6����ڠ�~k����6�����y+�<��<y���O�UI:�3g�(W:D\K]D6W�	�#��ֱ�{�ʡo���(2���������mp���.?�b?�_o�#V� ��.M&W���T1�)R(��zH|i+�"#&/��n:Y?���S��Y^LL��JL�	)+�� �(g��p��!�`3���ș��PJ8������9<�wi_tb���ͤ>S]�u,CY�j��O&3J�	���=6��r<!83:ཡ[Y��'5`��� ���yj9!p��6p"TL��5C���E���Ъ��9��`Û{��Ƿ`A�J�k��!�t����Z�jńs��B�z�J�#d٤����P�k��K�U�ܞ����+��������|�\�H 0`<�yD��i�qM3e'�yR�ʔ�������{��E����V�����&~�ok`F7c/V�������&��~�vS��C�aưm�Յ��i��D�E}�������q�ď��TV����ցw�ƪRc���9c+�xN�}�V@FT��j&�Ϡ!��p����*"�w���X�V�^l�Gqy�F����;�[P���Q!C�{铊��N��͐��ԅ""X��D�L���h]ǩ�r2L	^-72�犓�2οd��8Ղ�J�N�8�X�H��m\ ��~�*l�;O��f]B	8GLgV#K9��q3�g(Bp`�셈q��cBKk7 +�9��7�������{���Ԙ] �?8���Y����
'���Ѫ���+~��L����KR� �-��bj�N{;-"��B�Mky����!wv�݌R��?pie/��h�%�(-�}m�',����}�V`L�bY�k�� )/�G'[�ܡݲr{3��{�=@VE�`5I�q+e2[�V^���j�Dio|�tQv�ҭ����; ��XK���=��������9�_��Z\�C	F����>f5�¨�E��`y��!��qi��65�X�9Ze�
9���I 5���/��+����_C	�tP-�%�0ʐ��6ǀ����% ���B���I}��x=��I�%Tm���>Hӧۉ�;ᒣ�����-b݌k�����@��~*��dJN@J�B��0��d�x�o����i[��� �C�Џ�Ό�Zwy+��[$/~��E_�a��$ͳJ޴ͧ+��en9R��.�y^�V~��M�Ӫ��_�y���U���w��#s����L/�\�a�|ݮO�����+��u�����2�y!od����dV]��#m��:�
 �����8'�Z0N!.`���t"p�V��zS�u��(��/��`��W�:��j�I&B�bx秼�z���(�$j�zJ�3��V�{��@�R��JyoĞ�>J���_$�O ��]��AZ���{a��$#���r�)G�Ī"	O�q�����`?/��]07�y���b�*�V��KN��{�t��.��GJ<��j��%G�4�ʥ(
{�da��S`�j�a帚��j��~�	��Ì�=~V�:�S-j�wD��U*آ�yE�W6�Swq��I��@T6��r��=5��QqO-��M�*�:�T;��ۘW������uo�����~n��BR�z���}qj�:$0�rnH1�d���}S�jOb��]m��D�Rޙ��q�҉l^��ĺ�>�C��/0jA���P Mi���͈��/pܭ �����])�=ԥ�u�D���a�ң$�,"�!�_z`�U��`����ʪ9����f�
��jP�����&�j�N4_S�6��7�U�io�/;�9:��`�C��c͑|X�hh���a!�����\1��G����4�u-N1U����v0��P�3��������H�i[I�Hu��.���fE�D^u]u %Ԡn���]�?����i&l��������3�)
�w����p "����~@�A��}0 U��y��n����;#%�wQ�/e$���������g�ej���{�.>�d�j�If���|�Ma�I��ھ���nd�,��)G
=���.���s�夘���%�\n�W�v	��QG���Ueëɴ��_>7Юl1����4��WLP��-����B�o����1��x�9�c��nZ���
pe7&V������mh���ٟ�	�)a��vdJ�&��O�U��Ӈ��V2�.��N��C������7�HjF��1��چ����Z��*Q:Ƿe�hS~��4	�% ����3|{e� ����i�lʐn��� �AD�tzl�Μ��Aɬf�#lG[�wy��u�f��R�͟�mē�O��:Ȋ��W����Rs(�9�Ĥ�Ds䑑�O��=6�vHIȾ���u���5p�V;����M
���<�`A��RR��y�i��@s�.B���l�&��<��1<h?�0��Bʄ�U�dk�l\[�2�V2�����P�&V$�A6ܡr-U���E�dnP�u���WM���-v+�8��ڿ|\m) �i�y��:L���=�3ג1˝PF#7����H29�F+a�|�Th����E,
�8��������l���f����J!���$��Nl���d�<\&�����8]�G����h�Oz��X�&����"8�:�܄�Oq�L�����Q@�X�¢ �T�`u���<[=H����uZE���&�����̦�^�$͙Ɠ�ذ��J�)OR����H����<6��?�0X��0s&|�]��y��.I3��>'�A2o#bO�l���/�!d���x@̾!z��B��Am�3 �XL�6*)���I\�,>bT�C�e0�sC+�3�F&��!�)�9MMw�����M������xz-���-�'eem��������Y Mm���}IK�h-p1���jMo���{��HÜ9��0˙x���^�3c!��+�W�p��y�SP2(�L3�Hf������4-ӌ����i
0 ν=�FLM������=��d��X}���VE"P����G?�o0A��w�r�H�'�?.�6O���rR�]%���I0mt��J�^ۢǶ_��K�x�fD����6)(׌��-t���OW��Ү�����G���$�~tZ��uX�_B�T`؃V�!�	�zɞ3�ZLې~5ȵ25gx�̛�ȕ;+k9�����H���ڇ�g}jELso&|����X��EM�poq�h��r�a��h,�_�OY��'>r�B�e���ܗ�y�:��Z�|=�F\n���(����U3�9���90Q�(v�Cx�����\����Mqe�=��y�u_���@d��p5��+M��Q�'��h���i�S�o�h- dhX��D4
XO��* r����z�7� ��Y	S���E}�7P��W�Y�?����W�J��ҽXS����e� ߜ�*�2n�8W�+{ �p*# ���_�M
N1SбG��@+(P>^�\`ӷ42ڪuhVN7�w��ʃ�(��;�3<���0�ـX�آ��J�\j���!��͋��~�h���us�奟�1G���(��ܜ��+[��m��^V%{�rpVù<�NՏ8���cz��=r������B?3�f?yn�=נ=�vĦ�,l�,�#աh+�0��R�g���a7V&��y������ 3	&�?I�Bp�����xR�*MѺ���z͵�ക�-�[�D���bj��b�*���dڋD��]M3%'״������� J��/�q��8��`������2n�S���ї�AT�I̾n���ҩ>^���4��!!Gh�b�Y��B�r��)��^=�B<
'*"��!�����A���sK,�hH|��-��i�D�2Wqkg���_��Η�ı�Md�Ec��ݍ��CX�d&�#���)���|�ܧR�WH˳�1���I��g�?)(E��� �����i�.$"Æg�����o��t?!�KHG�E��ՠ�soi&�}c� �� �FD�w�=��7^G9�!����܂��3� �'����#?i[���}R���	c��k 4��y|��䛊�'�?-t�"���ja��'���GvLx��eAɦ��x�.X#�
�����]��2r�$�p���48�7�^����~b�S�^�4A��lu���@.�����3jb������F�I���
i�K�7�����H�Oy��[j���εk�S��S����?�rY��d�J�/��҂��NP���]H,�@C��j)��F�@��?�9)�3�;\'D6(�e�8���((���ߡ�}(D�q�'����?.uY�cd�k���\gL�
��)�t>Fq?�l�H�$U�<R�m*lR��ƃ��Kn���K[4��n� j՗� ��Z�%: W�@#"w���`�-a��}6��� ��������U��ʅ�4���E@�M9�ER�U5s��5��(5����,4�����d}̣f��*7Y�9L��V����"		������i�L;�:���,�X�?3�IhD��X�1�N@'C�pr�̱&k��NPM��V,V��~���CE>�H��Y	���y+u��aGtk�|�ɢ���y��v���;Z�&�������gi	�ݙT%�y��Ϭ��]���BrH�l��#Um��l���q/9Fő	6Ӣ�����W����ː�u�|;���JI/<X���zS�d�c��K����Š�g���Mr%���N5 �O�2�|4鷔�!�`{V��1��oEBąe��'�b�V�f�R�K�ī�����+�P�P��5�α���P�z��e �
N}[����TDj�B	��Z���r�����J~��\�T�<m��lg�-�>��Dٲ�6F��yFʯ!刭����?��B��i^�>���1�g���>��PʮL��,�?}p-�*�`������:���L�_�����o|hi��]E�x \�&�h�lL	��E��^���DdJ��e<�ݟ�T�������K��X�_���/Tͦ.E��*2Z�XN�闢7���:ԗd=�K��R����- М���T�B�foI���W�]���]�����7�++	�ì�;�UGs�Vo��N���w�MEre�<l���\܍�����Uz��T�GS��ε�&C[>�0�$9YV粖��y�Taڋ=�n�[5��X@"�wQ�a��{e"��fAj�T�i+��d�=\�Bk��y6&���p�'�����F0r��Qm��:B'��X��7�[*����$$�9�X���P��y�|J`�G-��&��\�벦�@����l���c���P �	�S~�6r�6ڪ�p!}��}��`�`Ck�k��Ş"�48`\���I�a��<l�Y�b��2���x���=��s������0��X�Sn��Vv�j^�K-�����yՇ%��J?�,����8�
�Q����U�R"!���\�5�ip
�\�g�O@1d]�뫉.i%�Q����{c��p6xxq�YAg��gI���>��-�6��얅��1?-�M,[Z������=�-���﵅�+�_�W�qi���������65�\>;�H"���xd���|�ݰq[P���ANA(�$�i��}MK�X��a�%�R�g�}�ҽuoUT�x��߇[�y ��_p�(�Ԝzc}��mB�)3$cN�62o��$��j�:D�Ohe-�P�Grde��X㹍�9�V������Z6�7��QE��j!1�#;���pE�8����^r$kz���@:�4H��G�������
�X�+�P0^���p��ڻ=NY���i�2JX�'�,\^���^�3���v��S���n]/�]��)U���R��f�F+Ś ���9�Y��dm~]'��򤇇����\ ��On���F�d���QD���C9x��B�N��:���zp.b�o�ڃ�#�0�A}���)wUm���������^�[����E�W�f�;�z�qLYʸ��3i�]'k����84w��X'���\]�1�)!���ֲ��,�h�����:����{I����4��]�&g��\��sV��=A4#n�׊��2�)@���:�Y��b�m�&�+�ˣDV0��>�����'L?�������a[�3��o��weT엄ĕY�1%�f�%��l愧��p�)l6bp����Ĩ�#P�l��͏Q�ֆ|%(e���Q�Yb ŋQ����jW`����5��l�q���9KĂ�'�M�d���qP�3�P��c �Ѻ���@tk69:��W��lzug_�%��?#��4!�sw��EK�D���
.N�g�U�@s���5KN�~��j�
i�B����2`2�ͯ���[��gc�um�`����=cB��ެz�ʓDpɇO�C��۫%8��F�t��5�)g�Xh��-���CL��[�mRtY� Bo���ZШ�4���+ˮ3�.��J�'ǥZ0J�5��W-ݖ�[�*  <#���D�32�|����?o��O���Tk�-t�������]^8��ӥ;?K�q��B:#�D��5LMaA�A��:(�(�"�
�:@
��"@=���V8�u�c�)��&��u��࣫�y��W�$H!,(�O��9�z�<�Wo=*��@�[�_1�.�X�ڢ4w�C�@�EA�yX��g�(�S]P��ay^��d���NA���[^#
/�rܜ�=~6؏^�E������SA����NC�6:_�P���ѿO��������SP�Oك�k~4�\�RS�1��L�Ұ	��?���	�����	��(xL8�����bw���E�[f�h�aK{iNpk���1h&6'&��v�}����$�mD ң7�����K������䋲�",ihZyQHӔ�7��3k;9l�	^�����XyY��6K��CGm�K� ��8��(��
���N��X|�Q��
�9[]4B��$�ސ��F��a|b$�M�|��y,F �g.}�.��|���^-{��4�<d������6XU%j�x�!���Q,��S��_<���G�fM/m���ݙY|�?]� LB�m�ܕk��`"@8�#�Iwq:|���Kz��6L��V�ob�t��Aq����"���j;���w~mKM��H6�=��;��@b�q�	^W������i�R0��8ṫ�[t�J�\����4�'��!�MmkL����U�s�)}�3�A&ZFa��Pd 6\�
t+�ݹ=42ǁ��9Fפ3�E�ѝ������L�4��rB*l$����YZV]��GR4��#
ӥW���٢��a��� ��T�a�A�>���o��o`2<�v�����J�o�28]u�LWM���+�d6͖E\���s���U��D6m�.�D�_lFA��m��Y��=�t�����?��SeM��������_�Fz(pN�y#{��3�B�RT ŻP�\�����	�ׯ.I����둃BlIޘ�E������X֌�ͽ2�9q:����b+m��%,�IY��!���UH��S�S��t��*ݵTn��5�K�/��MB����o�Xto���Ω���O�����6��q]VY`P���
�4�N����%/Mt�1���?gw��&@���U���X��w��&q���;h��9����"�o�>�Mfy���c�����E�2I�㛍d�>�C�T���U��e�g	�M�*k�X�EV�&����t����t��L���f�>*�F���8�v���"��S�J���k@Ma�:H4s／��RN>j�W6!�8=�'�5�n�7���T��|r�������C��[/�-HO��o�,��]�_Zo���]��ޔ�|�ےC�+���Y5��{T���#�4V.\(�����ß�34�pi"-���O�Ћ~#�;?ǎϲ��\"��v��Xp[��W�rxR�X'/V��ЏQ�T=���"a^��B���zi�#~��q\�}t}�,1��)K��6h����>��I�5��}��!����͙#�{�5�X�<�IM^����
tY��W(�57�*����޲b݉�Ꝅ��>ԶL\	�W�������k?�̯&����Q_�������C��sI�{N�db't;����m�/���:wUW�,=\��%�:�Tͪ\��[p�|��B����^�
k�U�Hf���[���vc zeX)X7؞��/D�A�lk$�=3r�.�u��Uw���Q*��>.tZ�2Ҩ�(�'��9��Ql��nu�����rv�f�>P�%Kң�d�(c�]RP&�a^:&5��X89�y����v�����_�������{L�<��1+w^я�k������-g����F7R�%�� ��'��l�g@��n�93����S%�wf�Q�9/1V��C
-ꫪ�i�9�85���<乜I��b9�@�ጡ�^*ye͕f��IEL��ዋ���"h��ʛ
��H�T�';��{�����`+L3���
�N��i�.�xMQ��;�F,?x�G^��S�C��3�.�����M"�E�R�L��]�ݜ>�x���eG���C��\��!�,N�j�3K �q���Y�:d���S�/bh6���LO�l���/%����eo���)�VA�q	�콯�ZU�/:�*�%`�|��6��t�N?���.ZnA�(�e�O)ܽ^�Hg��f�����B��ڔߍ@ݨ�u�lM��k�yã�{����x�V�Jō��g���� l����\fE��� W
����c�Ti���ڛ� Dw�$��:�����u>�g;�1)M&[��UB��Il�WB$u� "�P%w�L�/k>��>7���7qN��1�����ܮY'��ps�t����<{�XN1G_�oT���n{'��,����]M�,�(��E�s�iZ.�.u���ڃ���c4��y���X���ɦ���Z�C�6���fg]�9_Ɠ�M�f0����,LC�-��d����O�d;�\WX�B�^]L&q��dcּK�ut�T_͍�~�C�3t	b�`(~^gԯ2��UbE��A�|��BYYO��#W^����m������E�}<���3@a0V�W�!S�S��j�䡰�|~�h�F��,�m��Xm�(�9T<�J�˯��M�7�8�]͇�;wg��u�  ����[�g�=�g�o�b��에�-~{Ϥ�<߆�;	�E��F���\�5�3�@BHܤ(3d��#b��&-�S u�6T����O'��+)е��ڴ���/N�ʀξ����P��(����ި�i;�w�ΐ�LG���6؊0��hRmZVZ�� ��ӭ,p�
F�Tu3^�ų�7Yp�6�@b���8?70˺ �n4���H�p�P�fo-�cJP����Š��aK�2�_~����}�Q0N�ѩ�PDVàK���Gv�%�R���.��l���}]+�������.��u4�^Q����h؀�k����+�-15�񂆬R�Z�3r��I���Jݿ`OWEi6�f&�ei���lM��>��Σ��W�!����$y$b���HLU����S��,����#}�G���g���f���F��l��0�[�Ue?]���'�?��\��ar�\M(�>-%�f�2ARQ�gH���$sst��0�5^SFQ,K��;l�����2G��-	���PP�5��
�4Bwˣ�#Ո�_�pػ��ZF��ng���Y��4:縹j;H�P`�w8;��
Й�-� |=���ʕ@��_��б :Y�%HC�q�����w����,��X�/){}f�����,�M�J�"x��SB�c������ŧX�f(}�~�H��*�(t멆����jj�=�Ť�H��F����Ŕ?�~�
R~#Rzϔv�$�)���՞_�I鬏�yHz���+^B�v�ꭇҔ8���$����
R��Vo����p0�N��h�:^ ��<)�E�Y[�jź4ǭ��E(����������8�_�:z����1��G���k�3>�e������nb�]�P<�=�*eOz������՟��xD2I�:�z^�@�4���X�7�Kݵ疰B�_/N�1L+�kyD��μ׆��	5UY��T�B@��@�NM��\�T���5�z �쉔����I{�W��q��a�w
�����"]��j�V\����'G��/4AQk��xc��ΐ����Y`N�1���K�G88QWٹm\�1�b�]��f�;8!S���٦� '��?�\�rG�1&q�0P��4P���s�G
v%�'2�|�X��O_Ȭ���Χ1�~Zr kK@�3��[� ]�����9A�Ib'ڪV�<��1b�3f���iC͜K���ڍ�q�2�|\-���7��z̒W�f��٤p�h2�N'�=��� +~r�f��� #ݼ�O�j��G�p��\�ӻ��7<?�v�g�e�q�!'Ok��$����)�O��DҦ^x�I�/S�	���I����%�gpҮ�m�4U���a�
�w���1�6v�"��2��K�����?G)Sc�y�Uh4����-��!�#�7@F�@w�}����<K�D��yB�����6�_�	��ĵ����z�ѵ�=��j��@���B�=_yp��~Cq�Wz Oz����?�T��(�Q����`'�!Џ���KzO|%����"���a'��Ib/ j�'}6����[a�/���X�K.5jD΁J����y�)�~�v;,[����=v��7h���N��� #�R8��?�=6�����!6n�G�3��Lb����]�I��R�7�Ok�S����kI)̤�?�G�b��)�"��u[�&���g�S܀�
�����ڨ��Q\{g��G=(���쳀��%�M�OD�x?�|�^y|s�� ,n�x� ��t�u�Ͽr���t=`��v�(邯����Tl�)�b����ӎ�!�޼�_(`��rhj����}i�6�@e=N8)	��٦���&2�	]$����ϛ���?�{�e>�5	�J|�ת�ґ8��ɒ�y�9~Ŷ��k�g:�U� ��0*���|_��'���H/������ɺ{ȃqNh��l�� Vp���N&�h<[���h�40i�c�9�׊aΔ��P�|���354�buF�e�:%�lxk��2֜�%�B�!,Pr����5��rJ�rn��'h�\_����:,�>Հ�H��&�ɒ�s;^�Aq�+6�k+WG�/yϏr�,S�u�d	.�^O4u6Ρ" o���-r��k&���[�C�\��兏͠�i�������D>����P7(q�M��� 79H=��"���LL���٘�!�[%4��7��^�"���Z����fqڃ���R�;�9���h԰F_ �9�!O�������'?XK�3	>v�m�����c�o@FO��V���,��(L�?öY@���|���\���C$]�3�����g�l<�㉴*���@�"l?'U�'<��#1�<׬���{����P��'#��zC<BK��@�ӭ�%Oh��$�
��Em�����k93�|�A�S��ZKaG���7^�m���M������E��F�Xn+|���.I�x��D��<3J�SJ%�N�̇�<��1�ȕќ%=������}���ܮ�ͨx��U�u�;�a�$��G�jT�ڦ��m+���_�NI��E�����1�]ar8��-	��9��V��5�-�9�y�S���Nv��(f���nX,�#>��̡��bw������3\/����_�����7W��;m��?N*l1Q��ͿK��/�G�N1.8�ʡ.k[�xW�=��6h�ANzl���A�1�T���?�N��������K��DhG�H��q�'o��({��e��;�|$HV�N?M�\��Q|Y����=A��1.暚���1�ް��S�m�a�+%�%�5m;���~�G[�$�錭�4���[��S¿Qi��N���I�%�C}�E3	���z��۷��*������.�`8�W��w��̉w���;�H���XV0�Z�����1ǅR`��:��+&qQ�H��%��T�����{^�U�|��`U���lFS���?`Dza���V@(�MF��.b��ӭ�:�:���`�C�Iǹ�Hs�^k�)��1�,ǧz�*
��I�fJ?woF��
�q,3�v�~ݭ�$M���O�����ۚ�y�UY��n���<_���D�bYj!�
m��*��=�ߑ�!!����"�E�֎y�tu�_au���}���_�u�i�l���~�ѥ�?*T}�B�\��u5�/�զ�Ɋe��inMr�'aC@T7��U�:�PO�&���p��bW�4��)8�H�L]\!&�;+�n��w*A2��DF�9�+	�,����@f�wk����$/0o3Q�@/א�����RO<�����4�q����.�\Ol%P\u�t�}##Pz˦G�a��Z��@��z@�}!�x��a�~�IoC�0�ys����yj��6�JI�;�r3ye�������"п	��+�O��5�XA�������EjU~�E�.�ܹhK��� d�J����i��2aR>j_� Gk4Ms�U��O".3���"0oҔ"��nc�R�)��B�$�����9�7D�Q'	8�9.��ˮ]i����ek����}�A݅A����B}\�P&y's��?+3��b���.�z�N��0��er!�����OӅ}�_�j�k3�J3o����ݙn]/��3'�Vn��tc�:e�o�9v�)<
oȚh�'7���A*��W�ı��n�����x��3�h�K�f���3i�zȇQ�|��F$�~��C�8?z���i*.�n�F�9[�{zu?eĥ���k��;{��*s���eQ�'#��!�=����mʽ;�аd|�s�J�2�/�ؤ�8[�����'Rk�1g[�g����Ǉ5��
�^[���B�@>2�=�x�Xy� uTZ���G�H�n��/��kK]|��|������<�l{��^�/�-�����¼�J�����P:K�ز���@��f�9�M����Sy�nE��ݯ��ڍmɪNƠ�)�?$J�֬��\'(.R�R�I+����������hs���+1Z[�� ��M��D� ��(hGƭj��!��V�8ĺ*JT��O`��9	��,B���ז��?
��.��'�(I5͹�6�@O"��NߦL�'���$��)��X��ra�j�OP�T�O�"SU��̾�v|�|���S�hh�^��^Ј�%f�j� �Q�>b8Th�����&gR�YV�(�^���K}��H/!�'$O��VTMX^1̅��|�)�#k��*{���CI�8�~f��DLTn=:Lo�t)g�-�Y��8N���l�l�M-�x>��amI�>J�= ���5�=�T�^��r��E�7�T��,�OpvZ�A��[�N���GSn48{�Yd�b�)�y>O��WT�Ue?����K�ݾ�eG�-�I�&��5�[����{��ح�д�w���9��l����&��މ3��}oᰌ0y3k�+3�L�?�u7��&� �r��\a���Y�
ہ���,��$
{5&�_-���n����2ϪcN@h,���݅t��=�ošv���?����E���G�R�}d����������=K��>8�6Y����@o�H�ûWL�d���d�:W��%+y՝����U���`��ǻp�9o�E��[$U�I�DN�D��2@'���.�AY��	���� ��M;�S)B�̆�"`�"��;�?����k��LR� �(q���ez\ݔJ��i�p�go`o����Jg븱�Q��L�j�e�4�r��,��H� �Xj�8��Y]z�)h A_C�7��:�y�h�7�v��o��K����8N?n?�Y��D��W��09�)��][;�XR�[s�f0D&im��N�՜EY�E�f7����������D���e�j�i9�����v�Ă���q�`�lɶ�$,��j�����64�t
�	}�,���)3�q%���i�����Ơ���qȗi�0��5/>�[p+x���Y��A]�+�r�l�_7�T�c'_l�뱰��S5�@��<U䙡E�p�I+A,nK�.�Q���y� ���L8�ږ9��R׹4QȾ�n˰m�o	�]+߈"�QVf��u�eZ��}8cr�W������#Y�rx����i��U�!p��-.��f.��5��7�F�O�uWb�{BZ��:��vJx��XT��#f����"6��qb]&W���d�2ou�U�?u��Y��Z#E��J�*?M����U��|/�2���f#x�{� �}�����t�$J/���RC��8{n�����܆�5:��8D��R��=������t��Zm1�g�0 h��>�!�zb�X�J�/��J�$!|���e���������Y��}�v��6���V�i�*6͛L���_憃�k�a\q��F��t$<:L�!��xw p��gy�g�È����	�������=]e"�zCQ>s�<�]P���wf�L�NӘ��k	
��P9��	�5Q�L�}�O�\Xj��8�pa���#�e���QB��
̊1��r3��T�6bw���u0ڦT6ô�fZ���ٔU�tP�Q��B0�=���x���~�����Z�(��RY
:[��d�ub�u��٨�ǲ����Gl�H��OD�/)=@�xF��3 dT���iCD�����zs����Y>�v��3���6���1���G���V�i_���� 5��p���z��1|'{�2F�o(���h�kx�Z�T���� �Ur,�]��U��2�� E����b��x �5��@W��\�j�����X�>ޏ�ո�9�}`�6�6�LXdn�b�c���
=).�7n2�޿��T5���o��Y��dUmI�W����`�z�����Փ��q�u��{��<]����+��i�$�!����Z��uﾍ��h�TZ��l`�ƷRN�QD)��D�Cy�W\�Ru�}��D��~�I�E=T���@��+zx��,��X5*��u^ox�~�-Oj�|k�+�Ȧ��
�o��+����%��V��x��<��Pl�w�߁�?6�t��iY��5�)@ף\0NuY�_��N�R̒�	L�o~�#E���=�H[($cߜ[>�)��x���=bl���(؃^[�<�Agw-�F��*�#�'F�����͝�ʸ��W��]~!n��}4���|���u˖ �%`�}����:�/ v}1�����J['�U����""�{����e�<a����I#�T4n��AUn\J�m(��p�1L�W�n��G/�3��u�I@<X>��v��
�:\i���j��:Bz�+�ȸ�cvZbI^����@(����GV�}?��U̘w��F��A?��@�:����5����"�f�u/DC%� ����)� ���A�&�"xVe�oNН�-��3��F�6c��,�vOgu��z����������ς�4�WE�@����L)m��T����/��s�Eͱ�;���"Z�G��Щ�r�ٺ�� �홺������b]�����uV��$�r��̸�*�ťoߑ�5��)�����ь|^��2�������%�/r�����&����LA/K}��m�	/��[X�oĶ�I?x�}vh��Z%�BJUW��7^���=�2�W���M�	*��Z�T��*�s�C}m"�衸�AS����`�	<��A=���A��k��"�|�y�u�N�����z/����!��mg@���8��/�e�
"4�㻸��VN��l�I]rTy/��ξN�I(6�rָkȮ���L� QF��Ī
N��'�5��D��=�|�@{\�lN�8L巨�{L������5�xqɮrp�9�&��U�>T�r+��UB���O��N�~X�R�����%R�����U7WY�ו'"[���F%����#wfh.��`�Ht��p�uY��Y������-�e�4�$�D��f^	��e�j�A�@�vU��'#3�ݝK�j�����-��j�k�z��N>�C��:s{?���2�D(T��9�I6��;���ލ8�^�NQZ�:��%s��.S^�vZ�6k]�����V�-�t�!��N;���'$��7���h�A�8�O�5���=,���I��/�%����  ^(Sf9����sgzi�%R��	HQ�3ۻ=-7<�&W����@�qE��h � N�Yf����/���7r9���3���@o�*	;�f�	�$ͩ�Vb�o��J�����-.�$}�dD���9��	#��v�2�N� �Hg�si�-'8QS���É��e�}��]��%f^GH�KA�Ӛ�FL��@D�'(ȃD�kإ���s�o�[�f���S���� ��2���doZ�z"᝹����@4�N�ɜ`/�2��FF�;�VL���\@��A4��Ĭy������