��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A'xin�XO�v⨺��sZA�R4��g�psXdm"�d��Q� N�_��b��(�O@���k��-��w��ûD�׭�<l�'�b��++�|��}�]Qh����)P`*W����X�Z7�^! M��d����>�wE��G�i9;Rך���Y���{Ӏ���m����V����E$A�4n�a�(��w:K�g �R������+�aa�h84����eV�袆\:���Ji-
xAf�zS��eT	����e�R��Q/��%��B���j��y`#��	��d�6��Z�;sy����Cg{G2��D�;EF1���#���[Ι�i(�72�I�à�* ���G��6-��-4�bS�g���}���e��'��kQ^�L�oK{%�eV��ӎ4bD��&�/�L%L���� ?��f ��K�f�e��y�_M�������^\x�vz1���pq9��C�vZ=�����
e��'܉�`#٢��\���/O�#p�!�1�)��(Q�6�4�z�� �0��:o����S�
��o�9	����Ӗm�*gt� �� ��pt�T�]�n_�f�2�AS*�x׸���R6�Q�i�XQ������U�{�^�����D��1	�u�O��x3}�O�����Xd
�/�V�����CL�z�(R��y�D����i�i�wC��|+��Τ�	��,��������W��vc�k_�2��Y���B�l����-� )��k���U���q�E=�:8`pD�a�2'�G���� ���8��Mw;C����Z���+���\Fp�5p��������t�OK�����b���fa�ɖ��g�T�8��V��?%�U>��FvFCQ8Xx�t>7r�l݅�B���S�*ꂕ,��9rc��]�����vaw�# �-�<<!f��U�tu���3�/������5�i���L;�x#�'D�Bk��/�f��$�2
/l�n�=M6��,�0'�e ���yZl����9A�Ǯ^o�>in��xz�R����\�?W�uY;q&I��jj�G������:�H��C� 7�m���W/��xH�⭘W7�~�Ak!���-+��	�b�A �9����h�R��׭�iA��cT�έt�<>+�a�7Hi�^�!:E<�b@��(h7��H����[k���BNk
_�i����H� �u7U��sE�/�o��U~�?��N�j�֖�A�+1D�O�Z�d���7�6юb"
�1�x(<���Db�a[�Jc�wN[yH�!��,@cg�����}�/����÷��G�U�`g�4(��@��Ա�,I��Q�Ҵ��Ϊ�|��x>V�R�^�sF��y�%G#M�6�fj���}��T�6�o����~��wTx��$���Va�GZ��Z9�!�sn�Nt��<���x�dAy��������DP�
��%��!�#+�I��_̂���قE"ґb����[)��#M�6Z���������W� :�'�h�4$N�G��c~�sſ�k�'ɕ�O)�H�$�~C�+��m���E��/��[���R�