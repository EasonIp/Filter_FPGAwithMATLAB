��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|e����M`p��ّ���Ұ�Y��&�^�y�w������\�Hz���Xp;r8}�9���6�v�ZJ��k�j(�uK `x������#�C��2��2� �j)�8l����%�MQJ*%/�z9�w� ���:����̖Nݳ�N`|�?L2�\.�2
���sN܃r)�������l������f�K^6��+��spz�2�l~1G�=�=�~��a���t��q�@���~Zfv����{��� �,���q�jM��n�;�����׆M���ɰ��ㅖ�8=>�CB���0���h�	A�_�Ϛ����W8�Ƹ6�Y�R���x��o$E�C�������;����e�CI��(&�r�E& ����^�O�o���p��]>m��$Y_+�_p�����
Գ?KpʣE�������V:�ia�;�)2 3��3U�"���hz:qc��0�T�{��n�V�i�\w@����f�S�YŸ�p^|�u��������e$T77���g����*�e�ԩ�}P�\'a�d��4�a�p��O�a��|���ƃ�r����Ed�rC���f��k�dAH�I�26as��ӟr�)e���(q��Г��n@��<��F��znK��򌇵��\�h�|J��7oH�o�Ou|)}�l�~F���,Mi��DSǨf���>�2r��s��kgn�_��fb�?�^pZ+\���� �Y�8��I;��^R��p�)�i���<0�U�f��L8\7%=�@�rZH��8�앨��%�hdǦǺzA�K@ğE a�͞'X�\����1�Y���NvV� S������w57���WY՟h�'4���Kq��~���fn	=��G��F�-ل�-��7��M��ݟ�-�������]UJ�5����.?{�bMX�<�NO�֟�� �O��a�#��d�۹> �xJlv���|�`>쳤�*Ӧh���k�6w�;Cѐ�����Y;GOp�4a�nf������]��Np�-��9s�C�o#�����R�ª1|��j�*J˞�!��|��s�Ρ�j�B콶ۡV���ŝ�$P�$������u�o:�������t�d"�c��#���������~[�Ju�%f���ɕ��`<�^���	�i�0�&>ڥ���\qK43�=���Ů�!ԇA=����S�n��{\wyBoG��K~ӑ�ty���j������1�-_-03C���6r��)���	Fk��k��Wx��������ɑ�������$H5�G�p�FN���AsH�����0� �Ç�x�b�#	��c@���p���X��G�o\�ԗ��)�S8 n� A����� �o�-�&д�Ƭ�g��&˄���)���Ɋ��G�a����[v#�̐��w�Ǖ�
��O\�H�x�NG�墻����J�m:�2t�M�}X/A�[�Ģ>�.��Z}u�0��]}�1��43�>ܧ^�ޅ��SsLe�U��Z������MȯBm
"&�"Ą8�a9|�;͈�U�d�}��DX,J�ƽ���U}�$4p�ҥM�����j#<e:��"g<pǦ���T@3�B�v7Ơ7��C�N�����������u _��`JP��*t8�T�z��#'3�X�����t��߆�0h�'r �k�Y`���r���8L��4���.�"��t�K���A�&f~ק�v}.�bK�#�i��B����w��n����� 4�k�h� N(�OO�� �'�FF�N�dn��@�"��N�ׄ+�}h���I���*ߨ��"��>V��,��ɘ9q +��9_a;��u�=f�^
�.B��tf�ft�@�_t��n͘�#	o���K�5�4�XBS.C���o�o(�.u��m�/r�����f��j:å����	/4 /�8ko��ukF�T;cĔ�ʨ�b��9^�%����&E����7��v�Gm�	�&�t�����='��T�,�'�b^�YMС)�}Q���E(�v����?"ӬոFC~�`���$��+��j�l��-�O���Sf�H�r��Jd�J������u��
����w�(�&BuG�_P�u�_��{-��r8�8�� �b` ���mӈ!������֟��d��SGE$u�9v�DA�-��K%7�����O�_�齢�b64���b��}.!�N�<����?�7t��1���^]�6�_���;�n����'4c��*�j�XY���e��I�i�ޯ�6`��k~h_�
���Nl~��{I��yGȊ]�]F:u�l�� �ǫ\��Iu�C�2�v|'X�궗︴���s@:�ƕ"T��P�{�}HCG�8�Go>o7���ho1r)B��S� P"ص�I�8��ly�^C���#P�<)�&������xP���b�Ts����[��@]�O��t�ד�,�y�q����Ǯ�������,�n6�Tq�v��M�U.�������H��`n��X(��mϗ}��B�C=��óivI��W���b��b�j#�l�#�g)��No2�,�O5��|HN�	 h�y���킊�mc��a����������d�re@��Ob�p�V�G�.40��k+#
�pg�!���U.薃���l�U5( �ì{�=�I� �"��>p^����G��o�Uso/ҁ�#4�֘@�_���b���5@�;��)A�{�g��ɝ�`<d�o"��+:�V4`:3�Z��*��idC�'���ˮ�[39���_�YC�IL=�;����㫫�`į��䮌��	:�	վJ�ɔ�$ֽ��ш$������_�zp�4W\��(���}� uWk�y;=��[TJ��v��κH��܍H�'��3)B�z�ܹK�o��Δ�����7lq�G����A����!p��T;�^�Y�?o�p���^���c��]��su��R�3���(u<5ؽv���h�`�=�^WrPt�p�d47���UO�X��Lr�2X�a>��#ѥ�<�J'�݃�Q}���yQ�J_�����筨5�z.�/Z��/ �џ�sj�L�eG�$C
�v|�l~�3�VKV���5����5aw8)��(��B&����BcǬ� �щC7��m�����6u�uV�ڃ�����-V�(י�Z $��깋�o��������2�<C�{�H�W��rđB��ύ�6'S����O��k�O�!j�K�A89�1|���e/ 0�F|.��㤖rgu���uzL��l �~�uCM�����$'ڴB�2ґ.�3-YQ���l|N�O0@S����ҤR@, Jt))�OL�7����ts��zG4�c�<2!������K&G��!����SI�iDO�v���3�# "����,�D]O�-A]�c�*�L��J���l�aX1��y``v9�-tw�����m��6��#fL{]pm �C�E[E�L�m��d�j�� ����tKZ��G�&�z��\�*�DV�i�/��ywx�z�`�]`��F�\���U�Yu]��h��ͣ!�LQa�:M_~�/p��"��˒G��� .-y�-�Y]�^_.n�)u��o㝙�S�3L�c�O�rA8.����Em��IB���,ت��m*�dl2��D�*�K����R#G��E�e�Y��p���F��q<��3m�ի�*�ZBPe����g_;Ӷ�g<�4�~�� ~dk�m�����ϋ,=�ڱ�kܫi��`(�6������K����:��t����U��Dn=$
V�yJT�ˠ���� ��½��4��d�΂�R2��=
�����YM*���ܛ<�:}B$;�}�'m�S�_������Au��3��77��$�خ�'������M����Ywr�l��1[7�|it�=���A ��>�M눞ث�'�,���7�I�c�K�`
I�{W�,�o��p���Kμ�%f�C[�SI���������OZ��xM����)��Kd�%������r"�f�aS��,�+����rD���fPK��!ը@���z���W�hv����'q�<
u��e��sQj�
d[��(e}MXI�ʆPȐZ�7*ذδG!��%�b�|V�(K������ki���N�n����I2�F'ύN2lvSis{ֆxF���T��� `a���J	��XZEn�DFL�2�埨��(K[*���O3+�A�T4��H��sf�U>���9��?����o7�*��������8;��D̤-g�i����Fwn۟�=y�&z�m=�)�^��H�H��co*�J�$��8�`�G�����8~�R��;nXy\�X���Zo��%-��*�ym��<�҆&��X��������m����pl$F��a1XO�E��N˞)�Lo���؉K�a��sv+j*߉ߴ��`�1ک�6�2r�2`�V`:�k� p!i9d��A�Xڱk��s���pF���0"h<f���&��T��&����A����ֹL����b�����D��{�
.:�&%;ȯ)�k��}��L�l�㲛u@�� �B��Ǡ>J}�7:�;o��mv������Fu���+\�R<�K�Z'��M*����ja�:J����	oUQ��>e3�nZ�s/�7φs�@�+'%Wp<{'�}�ꁓ'��B�3��Cs���*9X5l�_#@!\�Z�,�+VWGC��Hr���z')���>ѿ7��I��r+^͙_�|]�&?�PS��m�p~�X���>Po�d���3�ps,܁��48v���b����ӻp�J���2P�!��C�7`�?z��;R��/��6��y��4�a�j ����'i�?4���&V|ݹ�1zΘd]��D�?I}�P�`��.KĉFJ��6�sS��F����[�r[�Sw)���~�`]Ŧ���
Gz���4'�*�h�;�m�eg0k��l������~"�O1�4n�%�Q�<!����BF��WS7���|����D��"�=�09�5e}J� �|��~zo���:�[�}S����>FaEdu��k�>���[�4���y�����Y����AAZ�[��~E��;���^���	�����v�p�~V4X��+��B���&�Z<����x p���lTy`.c��ooXxڰ��!L���hOT6{���v��-��L ��m��Z�/1�XGW��D��'NM׷2��3���AL��;2=���**g_��	���!�J��V��$/Cݻׯ>��6�2$ ���ڞ�B�)ZA�����_�x�N�@Ry��`����~!�8���M�"�t��w��G�J��	}��1�))8+�||㪷W��:߿,�N�9ׁE���FG�Xg3[)��XvC"�ǐ�,C;,dZu۬8!ݰoI�e�f����1�u"h�}M'���>X�_�zư�Z;fF	Ͳ��<������QHM�`r�.}'�E��$-�O�������k�}�݆��*$O�b2r�[To�6�\�mp��G�<���J�@򙣔���ݨoR���";B Tu��Gl�Gӣ<a?{��RdKL�ś�óT/��1}�@���(�K�WQY�3��<��lx�{���Q��n��V��rT���SH�T#�(�3��.lR�w�a/�هB��V�>������Gt.,H���6��:dz����S]؃<.���[��DF��]�:���E�QB8��$����3��ʖ���g
��D��Ya�T'�o�>�G"��L�Z��8�B�M)�c�r��7��Hm��<��,,�[ѹ�K\�}-��|w]��y���&�H�:D��2��<���Ja������%���`�Ɏ���ol6��X��ԗng�#$����b]u�W���TNjB�7v��Ľ�~z:�iǥ���"��f���IZ����\�*��.�D�4$�߰��Nn#�tU��K��c��_ nC/&Ƿ�f����4�����JYR�U	�'�93�Z�4L���B�zd��I��.*�gee���J��t>~��0O�h:�.��8]ʠ{� +��d�ھ^���;��;���9}�I�c����I�iP�mltI�<'g�ʣ�Vk0za'mD��cL�_����Þ��Ӄ7�]���,z,:F�a�p�>�$��w1������L�_�y.Bfg�Q�S��ӑ��=��X 	Ol��aԕB���&��@.t\�?��m�{7kP��)4pd!S���j�d��#�(����������:������� �^��X�(��a�aO,�B%�
UD���H���Ǔn;'��,1,�IJ[v�V?u�7�V`����0u&�9bq��$���I��<��u�i4ag�j�t��Z��A� ��оc���%R�LW���o��X_�"�	D�/�
�y5Q�����/)Z��2C�d2� ���u��_O1:�qّk��qe����]ʍ�"D$_�@Ry��"�doG?�)���]M{��ʧm< �׹��T��� �{�[�A��e����<��?v�O��:+@U2`�f���^m*���M��T��h�'�oq�������~_��l8~���R'9��[aYprS@���
�J�P66<[8���G�`b��r��mI:��7<�YGex�Y$��"����3���Q�}��*l	��/F�Q���ϘU<�@�D���{�R�Z�~� 2]���y��{�=�l���.x �@.��U�n���R�OU�Q�*9C����2g�A�V-x��@hLU���~��6B�&�J(	pq�g��6	�l`h�"�Il��weG�iͅ�l�*���h9���ζR�������ñ�m�Q�f5��z)y\�Y�c<Hs�K�y���ɑ����}{�o��7'ޖ�k�A8��I��s6��v7��������FA�O��T8�س��v�r۞���P<�r�Cnr�`���nTgT�V�f�wUYH <oP���0Ypp���!��E:e�]�ڱ�71xƩ{%9�aD_l��8�lʋ<�����m'�~ob}��EĆ�Q��n��j��u�s��v{�G=���t�~OL2T����H�&#w<�;�/-X���(��3Y�ϊ�!X$}�q��!	F��ޘ�Ax@�N�>ʂch�5gԒ9�@�G��(�#_~�EtQ����a-�{@"o�#`��L1�-MJ��������YW���Qu�界�T��#��F0�0b�Kj͌�(�c�bwÈ���^�� �"�ǐ֊4��:[���k+�hV|2���k��U�1������Fo��0���adF�����*/�ؚ6�k�y� ��y�>`�77���T�xA�X�i&~�M`���:�Ǿv �DP^ɠ~�3\/�'��R;͂OK�7; ���d���h�w�h�hДPt
�ʚ��#H�d4j2Xo�'��da��ڼ��aLM���&�q4��L�y���J�#�>$F��V)&������Z�
�H�A��h3L�����B����=_=*7��)ep٭W`${�A�� Ju�،/H�2�i�eh�q��L?�af=4o\I����>8# خ|b?l`��2+������܄��H��>���`��l++��^N���|e�a[$��H��0���%��`�4��&��7��-+�	]�9���+n�ʻ�@�9���˖��2�5�N��&�tM~0���*#��W)�
�Wڦ�B�4�&j2���y�֞"�{p�l�!ۗ֩���ݧ|�8���3��9*�O�Ÿ�C�$��)�6$�_�ո�PU����W�{8@?���rU��Q���Q�5y 	O+䉸�;���L%�7z�c�����D���y�����&�8�Mz��M)��%+��A���~;(춷|X��-�!Mx���S# ���3���$�1�=�I��ѳ���g�8 �XưKU�d����V�Ga��N�H���Ѿ��\���LN���r7����߮�}���ToC���m7��KE>w�F��@y,&�6��3 �I	�q��(�"�(Z�_0먍��*�vA'�x��O�t���Y����xֈ&���e"�g8�̾�@<�!�8XU\e�Ҷ&Aܻ���j�~�C�=C��>���|t���g�a��'�� �t[����Y���j�$º qo xE�k��ύā�
�d�V��㨮v]|(.�b�]������﵀��.�m'��+�x� �0`Z� �P�\>�ړu���[I:��F��x)��	�>o)Y��z��`�{"�_��+�K(u�Q�z�N��!L+T�ח3H�ޫ����]�7M�j�$cR���,�[y88*��e�$��N�c����M%�����h10S�h����L#���~8;��-JR�K��O�p��5�Bȝ��dǕ)���ڵg,*����I�2�L���N�MG~b�p���BE$���Zñ���؆����D� �̒�<���K�} l��?ϟ9��$q��18�˚:��Z�Dc��w�|xBo}�����	�Z	��3v�
��S�見�21Ym���U�*=?2�n���z�-�q�q�:#�	<�{�^e��?i7�f��j�X:�ɂ��_>����6�?����-��&�����[��4��e|
�a��&2�AU�sK�+��lY���K�D��Sj� "c�~� ��yi/X @X��e��S:p�&�Xf��Z����*�h�[K-�,�V$�W���A�{��@X���{����_��iH0@�ju�Ső%%}�?��,lV�_�^�kj�J�ڎ��?�����]h.f�76��;���-�♐F����񶜴R�����&E]xw��6����^@_�?���.�*��J%������m]	\�@�����#���/��_: ���% mj��썎�%��]&���?�X8��ڿ��c�-m�ac��{\����v��:�{�d���(��݈�_��������{bXO^ W���2GJ��E׹�����]jދ�S�W��1D��J}������K�3�l�8��K�(�2i����{x��?_�ʃ#K�Z�NF���B�Q��Qr0�xb$y)�yF���>#�H��p�l´h�:>z�n*y5��䬞Da��*�����Y�0X�=S[�\��Q6-	��[�]N-����'�:�8��G��.���LMv�8U���1����oT���w(ېy����/�5����� �uٚI��<a[�m��@yG^�>��������N��Hʀ�v��)����I\|��Iy_�ɗ3��BT*������](Q�g�X]Ss���ǅ'r�p;���\����k\샺� Z�����P�v_��3�Ņ���B��oFt�Z��^��դ¥�o(s���c4�??Q{��k�)(*�3ė������$q�����h8y 임6�6�Ä�Ms�``����3�O	=X�=-�\q@�f�I]��t�Ǭ@7�rh�pVA�:��fk����d~�gMwp�����#S��(���W@���A�����O��$,����MEJM��~�t�MP5�FDko��dl�Xo�6�C���#s��0�`���ΈH��@� B�}��߀F��Wt��k̍�"�P�3��$WPo��/����;��ݞw�C�שּׁ?����zrL?Ao7��O,i��!&�pb�o$���م�mS�뇜�|�(R3��}�\j��2�F������\�m������ߞ�cU��� ��| )�&�n�6$��z�59pí�� �*Ϯ<o���ͱ�X�Cz�����a'�5�7��r5,��?o���DHmy�[U<q�y��Ls�B|l.ӆ8g7�(���<9��O�	��w���sź�s%��-�7�Y��/X�m�h:T��R�(?,7��$R�8��U���E�b��*�$�3ʨ�O�$�ևF��(��/wL@V(��?¿�мt��kI��� ��sU������֔8s.H�{�_ouy��檋G|�P3�)�\?������U�v4
V���`�߂N�.	���a�㔛�<y�����wnC����ɕ��)��h�ų�����'����M��~p/4�w�=��z�|8��a�Bh[l�Xs<GN�����	����I�4�W@ ��L�t��o�d�0D��k%���z%Xe�	6sx/���9y�W�u\�|bW�<,��*�]��}�zE��]�4�5	��`�ܪ��
��c�M`���y���p:�D�����$$W\�У�[���51�,��j�=LH�����f��b�__�D/�ʊ�mgȿ��N�^����S3ɜ��H����~4���V�g��}
�˿��Jxh^,MQ�Nw�疛�'�F��E�v���������,X�qrQ&���N`'����IlW���y4U�Y L�y�;^����4��9�?��r������)�{Ϸ�R>U8{:\N����%Y�i�g:��XH�����˪70��T�ޒ�2�L{��2{�1�*���O2������"
'W�+�w$B��	1��i�?s�N)A�'��\��w��Z��!��+�N^#�����+dWrtm���Ӏ�'י+"+�)���ůV�`�[m�~�f����`i��1>��(1n��M�� ��̪kh�db&#��X1�x���HD�V�A$�T�etq����ā�v"X�����	'j�p9V��3Zރo!��&w�U�g�F��h,��Te���׳�8���_�x��n��<���ڪ�L�jz8��+�������9�5����yܚ���\��x�r���?6�Z�;�����|ԓƀ^e3��~4��	ck�͸�B���iOof����r[;}�nJ����7:����d�'ۅ"��U�A�#ne8������5�ѤZ"�eT�P�i��2���he���a]��d���xjS ڔ��x��O~�vjH�fl%̞�w�d�+�љ4~@u��:�8F�P����wA�nu�3E�O�q�)1S�LM��:O��ø���;�
��_q�=3��0yf�CA�îcKU�A}��+�:J����-4^U��Z�1'g�Vd�_}a�2�=*��d��kX�2^��m$YW����a+�G'H�A�����i�ȼ.}�(sMѾ�n��h�\Lp5Q�������%�T`L�Ql0	i���~�D��(X�1�pe�,sFeE�c.�H�OX��τ[�����p��jۯ��;��k���h��ZI���#J�.m��g�G%4v	0��8��/���>�E�S���M�]�ʴi+�0���+E9�]?((�q��S���L�f�8�}!���>�iL�ɂ�[���X�qe�
�Kð`~0M.��&�t�Qruz�k��f���M�l�y$x-�9�{vjԟ�u��ا=���C�xB�����̹��f��x����'�wH�Fʑ:�:x��5�K�2�~��/���0���r�e��$έ��3C"�XYX|O���/4c�a�"Sx�o�D��[� ����ƛ-�w�B�-���<G�{�6v�T��U�
�p5�I�P�'�]����4��)�A�y� "� ����Ù�I���v/�a@�K�q�d�!u�ɖ�@+R��ɛI�"F%�d�'��ۭ����,���eYZ�Tu�0SB���#���w.���	���崖}�����!�wfm��\Jҩ䧆L�W�szH6��&����&>i�H��[����-/�|�w^r��K@��G�����{sQ� ��V]�a��Ym��p��"�^`�L�`]=r<����2r%��`�|�_ O4��>ε����v���@��i�R� �Fr�F�m���G�%��PXHU����]��XK��]D�I��y��V�nE!��K|���C�w~y�S�2pP~Fn�<~�@� ��|�6s�W\9]��`mI�?%�������!g0�mx��3XM9�C�O#��;e�/�&���#n3������M���Y�mr,��TGjy\=�s-������,�{r����4~"bzu��X����Hhs�d���&�nz�K-&6��ѫBUyP������'��h���/�JX�=�ܧ��
R�DeJO�m=*�ˇ�'E��)�f¶�ȉ����,�_Q1�Nj0�Bma�1K�l��^!�a]H��:��}�N��_ԦS!���#	��C�M�Z0:��sp��2ٚ���-���,�{t�r�ah�n�|	 JC����dy���c��u~�����\a�RBF9R2(���Æ��-#�?7������a������aiJ4���5�(��ޙh�����E��:sKg9)�G����m�IT�a �S����`�}c�Ը� g�4�Y^�\5���� z<��� {tiތ���A�PJn�2F�Q=h�L��[�s1���wB�)����3䙲#�)E�n���T�
��I ��6��ѧ��ո��WF���-NS�D�~�6�i�N�����o�:��I��ŗ�꿭��0K�l��4��'/�A�`�D��#�YMq�[i�z���5Tqx��q �� =���k���&o���^Fc�3����N�v�	�m�e՗��+�'��6��2�"�: 82}Y���Sݝ`���0���,���'��V;���N���xXhc��=xl�N�ay�N D���p��޴�c�m�^JS�_Q�Y���i{tP�é�:.6�]�s����9���5�r���S!����ٳ��,���'�R�FH���9y-{�+�-����n{�jHZ�y�~n���W,��b�9�ɻ�?�����\�m�:Ǉa�!���m�ASG��0a���1�6�&���ه�߽���G�\����H�Fk�2Ѡ&:��j�o-�*��G�f� y�x��X��<|0���>�E��eB��8�i���4����җZw�������P�3vg@���=1�""�Dz�G�����=2	8�S �.�pu'|�� �؆mh�����!�e���If+�B��z��fH˔���
r<Ü�Ւ��&��6Lb3�NL.��RM�� 1όx���x �ֶ��P>L�//ϟq���]����,o�x��˧�9tx	xk�4�Vf��=Cl����h�f)���gK-s�ML!Ҋ�͆p\8 �����sS��JnZ��$(�.�p�P�!��Bޱ��8`my�o'�|�&7�xh!����׎���󠥽����:��C�ic�=��g驅u@��K/o;*�7��X�@��q��auPX#-��r�N�0M��n�*�YO�J��Tg��2Ϊi�[Ac�2:����f��ߋ�RT�]H�D�혫f�4��ǩ���7��K6���o%��!�b��`�" E����p���ƛwQקwe]yC9�C?������H�3�7��$�_n
���*�6c�#��5**��ct��X���U����0E��8���H���������U_�&1�� ��b��
H�1g�; �]��U���jx!�[�GN�e������-4�"�w��[��:hxg�g������j�>s�V���q��Sy����Q�^��@>�*WIp:j���d&T�hy-#�Z0�_ܝ�3>	�Pl;:E���9�ă�g0"q@�3�/�ڙ/Z!n֓Ξ{͗�� 'o�	9i�3邛�*σvF�Ue�@�Iű�Y�H���2��p�O��7�����!����hL�7S�z�`�i:S;�J��]l��p�V$�?*q��/0��R�Q��ħx��v:�<op �/�M&�M��8Xx��;�}����m���*��͋t�-����(ｷ��K���e�{��-�G�ఐ�{�G�xm*(��J��-���s���Қ�HB�+�Ȅ���Q��$���&�a��V�r�WM�.�e�]7s`���uR��.��\�#��)��8�����u��9W��g�۝Π�����r<�#o��J��X�_��t��z��W��}�#2
]�4��n���uh�#�*�7�"��a�yG�q��.�٫V5�Kp#�v�٧X�,IL���
_������.M��s� =R�ALs�����P�Rߌ�v�^{NfB���8����x�U�
m���s�3n�,���;r& S��Iw\?ʽ��=C&fy��db3�������_m.w���5>�������XG��1�E@�(�����V,��x�@l���Q]���j��hjq0��ѿݔ���r�B3���n�|�ڬ�y�E�*���H��I���]��
g�XБ#�=^gaݳF��'�����3x�%��H"�v�1����E��Kf1L���睼o��g�)���PEOG�k�^��t�iooR:F#3�Z���ʎ>>ﾌ����c2掑������x[�a��|�ʎ�����`���FS��饰س�f�N���\cv���|q���|a�l��:W��!(��W���~���4���J�|�܍);�-J(��'*��~|r%j���p�C�c�bZ;�̎�\V[D�Ə7pR_�quHT��B�v����^yEq�b��_��T.g�̥`�&�/�21��s��K_���3SPrߔ�'�OP6;XO�5e�fnFN���a��l�������h��6�^��B���(?,¾��ĳ�����
�R���Ցv�Y�7�<	Q��7�=����b��U�������D�6����i�����.�QҮ쩎8�+��$�|��v|GA�L(���s��5�N�\��#OzP���\3
s�/JM{Akd��LW���oaT�GI��j�[]����g���.�a.�C�-�&	HHN��a�<�7�]�
�k=�x�78���:�K�����wx��F��r
�ʓ�%�$#�����zy���C��JS�p� J~��p���Q	��/^�oXj(����~"�H�Š۴8�i\��P�in�+���_&s���x-��s�k�;~}�!]3����m�);�:]�)�4�[l���ڨF����hD��t�y��u��y���.��D�-b���LG;�����}|H��
%���.	i+ge.���K�g�o�ۍ��g��گw�_��{�2���~S�����ёׄs�ٝ0Q�o߬�i�ʤ� Ӻ͕]a1�E`g�����_!�n���*}������{^$�OUZ���t�9$ O�Uk	������#��~G�f��{V(�O�Ȓ؝i#������Hxl��H��1%�n�ڦ*���
U[�W��\��~O.o%Q�� �ؘ�����[�f��Sj����F�>�[�ݠ�s�3�f
y���k0�a��˻Cآ�^Am�Xy�֊�.i�
9t��)\U�<Tg1��w�+l�u�����)��䦴W�Z����^�4�z�r���.�!��0�XT�I/��M���'�qLJK1�jg��g�H(�;S���|�oC �,D�"�K���t�Y�:�FoA��V���6�*��F�c�ZS��1�b ��/�*� �D�a��cnT26�ޗ�$p
���S�N�a�KT��P��6p���8O�\�l0m���Ge�$-ɾ��_��}\������O_���r���׏���faV,��U˾�HG�N׋�}2��
,�ɔ�@9[/�̪i=�u蜋0��[�(�e�R��օZ1�?={���5�f\���P��.��h1K��RXLVPf@x;���Nm2�}$sPTӝ!��)��� �f�G ]�~��1159ϐ=���l�O7����\�r\�u�^<i�),=�aHU
"����<��ҳ�� �ѓ��W��r�+mR���Z6�k�^�rF�5�*M=�wY�����x?]�A���#��ܹI��jL7�Ĕ3�̈je�eL��!Ntk/���&�:?�P}E��<�\����tl u�(�0���.-��Κ4Э���8䆾�#iS&����o=�:Z\��,�,}�7��t�(������S�e���W��8-$�a�*�E�S��VO����1�a��_�'2��q9�~�+��t����3罘�Y�B��b��p"��m�D�3/R�9���E�pQY%���t����Gh�(�;A�{�mQ��F�;s�__7�o�!�����s��!/�O���I(Oʹ~�Clv�՞�@C�!�b�7d�\�ƌ
C��m��o�7��/>��:��h�% �6i�F��c���Q!۵�^>�r[ʝ|��$ds|�xAZ�/l�����HhX;����cH���5\bH�|�}��A)�,v����'�������?h��h��q.�7�O�4g��PǞZ����LĪe�bnk����#%���6����'�Dڷ��M�}��=���'�|j�bl���1k�iH���ĕȥ,d�Z}�D�Dܥ�	�`����(W�م�?��{LT� Qg*y�n ��ԙpv�û�,j*���������j�vR9�~��z��GP-LN����t���<�*j��?�5�U�ꚶ���o����dz�r,����TE�Rnl?�����t\.пӥư��ׂYs{��ÃÈ!�.��>\�[zAΉx��S�e|T"SO�`�|`����D��B�T���Z����YƯx��u�hf��+��	�ϭe����L�@>P�UI��k �҄v/x�'���QE��ݨ.���,U߸��~Yy�O��V�:S�	-χ�)�����Ouo�Z�����lM�2��Q��4���C_iS�0��O��y씮���q��Đ�l>�L��,ܖG� u�d�dz�:�h�{7��)�L�d��0�8�	nI�o�tɭ֓�G$�bB�Qڀ*�:�Xk�-���t�����9��>��kZ^ިh������3vZ/Pow�	��b,�QY�}��G���߄,n��3G�f_2�u.D�hJ]�q��e���Z}����L��&����گuZ]\@�jS���#%�T��D���n;��7��5�*��`��$Z�S�T�vv[����cbq�:�|�����e"@F^�=t�P-����BYR�ՔXqYF��P`�d�J�6Eq��b0^��{�қj�H���2� I78%��k��I���YN���s�^����/�\���M��)z��N�R���>#�Ƙ�j�N[#���l!�V �0w��Ǯ������<Jez�,�ʙ��U�s:d��'Cqي������w`X�ϴ�A��`3�̥]�'������^����O+�����3C����L�s�؍|�̶�|5�C j�CZK���K����u�>��e�=w�7Un�'�,��]ꗄ~�4&��gu����O�-�����bnf�n� �ܮ�dSřv_	���{�G:�l��~EUZgxX�yp�G�)tw� 8eh!zF�ݬ*��O�GK��q��xl�ؿ��C�@3P�G�×£Y+�o��D��D�r�e̓3������ˊV7�XB�����t�/E鴓�j������z9����/8]�@n�i��A?���>��*�xp��{-	��S4&����ZU}HxtN��ɖ*L��M�߹^-_���低�#�8ƖR�ܬ&s7�#���>��vǪ�PgM��M�t�ׯ�K��*з����Oyh�f_�$&V�AHc��.��/�4�^u��,�������<GW)9m�2\+ $˰�E�@`K�F3�p�CS��'F�0(Û�U�:��c#O�*j>����T�$;��	�I�� Y��	����*9�\��mŏ`��� ��1KH%Q3 /`�LcG[�0G`\SlV����pp@gxc�KH��'�%��. �ۏ�-Jy�OJ�Qx�D�w��Pǹ�/����*���c�*E��d��S��&��K(�xG�,�\�����	�3]���M��>,j@ͪ����VwO"*�<���u�㙍UR�,����0G�Q�/�N[z����		�|ۧo�W�	�)�s���`E�C��MJPV�N1S������-��9�w'�USR��C��p���p�Db�b8�C�1Xo���)fѠ��������})	r��4㿥�B��>p'��%��B{���:��.&�!f-<����8�x�p�8!I[�5o ?�P����
�mW��e���EZ⛰�g��>BfYW����)"7x�q���`�*�-�ܧ[6>G����URuI�4%��d	�a�v"�-]��R��Иw���d���l)��澁�4�lO11���H�O"&I
���B�Ҩ��`�����y�u�h�l�aL���4��')�X��|��S�0���|\�����r{��L^��� qj=c!�SU�����r��"+5�5B��u�9@���թ��j!%T�rkS���m��s��
�,�M��C��-O��������J~�*���X���i=R	��~RD����K�qJe%�d�ǝ�]���}p�e�mN������I��UW�����3��t�2�'�C�ΐ���m�ￅZ��a�:���������8����f����ž�;���a�}6JT�����S<����ՇS3R��!+��&Z%7��+@ܝ�Ռ{7�>��� 3��d�MjౌWU����oŦ'�ծ�����>8�U�C�$�1��v�x^��������t�o��~d�i(=���@��J�KGl�A�ោ�OF�z��-�,p�R�A�K�^A�{�S�`�z�Ko�7�da_��~.��F��e����_%OmK��L�!�lH23�膺��:-<(9=���Zr�m�6Z΀ރ*>�5-����P�~��R�j$���f���ח����>�D��F�x�!X[B��Nܩx)�
��ԃ;7����#E䕛�k�gq��ly���+�%t�v��&�M:��Y��e�	`�/��X�GUL�~* ���o}�,���7��,�"��~�I��9�\�H�Lѫ��e�'��K�����C���%��'=������?�i�c0����&)ډ��W����t�����y��C�!յ�~�놡�{�I�L	z��d�k��^�8 ��%?�[b�9��v�S�K���pp�_���X���K�s�m�}5S�8�lz���}�ܘ�ۻz%̿�Ju>P��S��M���M>��E$9^m��Ɉ���Gܔ���RG���_x��L��@���U�R��������o2憤��-����G��[��W�p��|{u�N̲Q��#�T's֪N ���Nk�pGO��V+]tWD�D�)���/��_7�/s�f@m�����}R�w���<#��F���
=�ݪ�|����'gpeҒq�E���%��]>��P	�؆'o�ܑ����6�*���N��%=dw+�
�/����k�%��O�K�� �zU��a�羏�����6�ǋ�|YfIMe.�z���=_�忯�k�TCF���L����?�����pYF��b��Z��o�����t}�.����qJT5m#
��j7��1D�����2p<N!�u4A�^��6i41d���Nn�X#�mh=	�3!���YV8X��- @���/��#�5x�G�:�mS´H��s� ,�2ϰ��W�2`%I��A��Xu��p��Y<s̉�Ow��&�g91���ާ��*'���u��;n��Ɯ�� vp�HVl�Z���[�E�q,A�޸��և�r#7H�������M��?�0l3 6:=(�95�E)�f"G�O�&N�^*m`n��ځ"�aV7��l���꧶"�3	y���!���c���ѢR �dv�3���cH�Vs�l7����P��h{���:��K'�q�z6�g6"s���]�py��&ro$Sjk�֯��"��c�S�5Ӽ�㗜�-W���k2MQ;��&+�H�:�B��¶��@d�Y�a�{fa�W ��u4����ڭz���$�6FȜ�	��v0|���*ʜ���^���z�����N�6�b�k�Qd����_�����6x��I.���N�F�7�a�b��hYw!*|ԊwsֈH�.9O�d��i[+�H������s��{����&�?�Ri�ɭOȣ��,R��\��.v���}i����)�+��
�ɂޅU&w�W��T��5����\n����W��m�i"��d&���)ߩ�H֛��dH����:���4�B!�o����M�4hǿ�_
�̓��¨2}�if�
������zn���ԓ��tTr�%��S��]���5�"HR%S�0�ʅ�ʽ��>�Z�ϙ����;��D�z-��!�LyD@
}�����v
����{}$�?��Q���򿗜�\���r����٬aF'ˏQ��vIC��׬�߬d
�VF��PƹD�4�k���a^�j�	��e^�W&,���*��������(
�$��#��F��0Ͳ�e�ki���5�a3k4������1`qկp�90#յ�v��@��Oؠ0��cT�D�pe au��}�HG̻A��9��ni�)����J��P n��.�'q�ٍx���
��D=%K�U����3؈�����NGI)&=^��j<K$׫S,V.���R��/q�P�/����D͇��2�Z4D�t���R�皙u8���sشvj����Tǒ���.��]S������fbE_pŖ�EfD	Z{^V�g���Z�Q%R-1���Kޱd�IV��]�ڕ�r�F*���/��ed9%y����� ��%ԝ���>y��[=	���1���t`�ey%�lK�"n�pU��)���Ny��rඞ3�3�6�'�9��.���}Se �^q+�!�Jס�@K�s�-��$��Z/G��	��/.LYd��<P-�^BR�?��b�ʸ������>��f����{��lj��L#n� QU}�^�ߢ/���;�pb��)9�E�BXq7��&�{�F���`g��W�E�qwr�;���p���9/�+�9��T7!Wz���eqD����X*uE��ʈ5��I�6~Y"�n�v �LV����PJ���n�G��6��M�>��i������f�����Z��7�����s¥F�"�	螡;l0Q�v0掏�~�L6��$[��G���lٖ�2�8m6�Q��v>����x,�"�\G3�x�9N�,T��X(��#yƈdןc�z��Z%J�H��h]w������������������&�[A$�{�5��O���}���r�W�G-�Y�# ���/l<�b=�G���MsgL�==Ps�\��gdI�"��P�U�-��٧x	�p���F3�4i>��W�����4 �F���_���SUAz��2�����z����l�a��g�%. +�0M���r���)~�n���I� ��p�%�eO�f?zX֩�Y,�#YꡕQ���w��C<���9!>߬�~W���,a��q��ެ�}���Z�]�����V�
����B���` �3(W_|Ԏ	G��2p��}8�I���+ؐ���|��L-u�f}�C&.��p�X5;X���"|��~�VO�<W��D��yXX��Aռz��q�)�/˝�X�g��̍ҘT�/L�ͺ�m@�<s��={L��q(W�Ql9"����U���Wqt�ڛ%�����E�?�`A�݋|����~Ğً gD�h�ծ;gh�[h�t&O�陾�����5����C��@Y��ҏؽc<��<�>ذ�.�9��
�B_p�s�;�� �����>�b�.�kс�ue� e��O����`3���|N���*�k�ЮS�8[Pw�ۯ����"���5��
<1�j�!�څ	�� �Y�Y%tIj��%1�aF���q����� �,E��;���;� ~Sȡ����#/ԌK4�frV�Z�9gX��3焖�Tl���hsHr/ L� �m�$�tґ���{��R@�G,ՙ����ӷ:����r`6�݆�0!�@g�v����w1��5���~=VL�֜��4H?h�]�?�Hм[�-b��C�xr�=�S̒�6�C����Q�1&�l'���V�����`�N�d+�|��Ks$:z�q�l� ���NUig�/��)��)�@�����V6_r"��$0��B7d��i�J.�l�~%�?� R���8$(�Pn�����J�F��4��D�gJgJ�1ء8�0���V��/��;bHN�=F�����p���%Q9i�=� �ٷ���h�ڳ��2�n��M�Z�gr�[�\{��a��΀�#�J+�n<��[����s��&�&TBZsx��M5��q�~IݙD���r�v0����N�������5��:@���C�j<.0]#�99��W�8<��ͬ+�����/Ǟ�i#$D����I;G����E���]�yw����ȯ�e£�jd�ҧ�^�l�IH���S�\�s%�e�Y6��$oD����ƹ���»��J657�}��kv�w���K�rԡp�p:�y!H��vp���4m�p/����3�)��X��?��ɥ3�m�Oc<8�s�;�%�$��<QT�d��͞E�NX�ڼ�j��W|��xO�gT&�Ŕ��#a�v�c�;�*f��|8 LCO#.��r�\�+��~��4��CZ���sŘ���t�`��]�t��dR�={y���-���}$U�����vyu9����Ȫ��nM�h��I��3��5+��נ�``E^F��?�a*ʩ�w6���ƽ����樫qۃ��Z�]Y8��6�sW}-�d����X�Is�(@�V(��b������e�~����&��r�n)�y��"	��u�_:�����{�ܽC�s�R,3����@�E �^)zTj������i����wWk9��<֊BM�&�эMj ��Z����d��ٔ.�e���6uw��PI���Vx�}�@)
����6�J��R��f�ɗ1��!�wF�ɱ��G����x4�Q�Os����a��MHۆ;�18o�C��q������<~2���Խ�*�hu��`H�/������Π��]��I	�y@:�K4|�W���+���?wLq���DY%��|�=W�V��E	çT�[�P���O�"L�q>���KTC"c����� �n|b��[��iȈ���K7Dݔ�NsЊa���)춯��s���3���,��v���u�����&޼��xuh��2`;o!�5m7����U�	c+��ix�s2��n��=\�xd�|��j�6|�o.G��b!�޾{�W!݋�D�4,o���������O����_,O�Q]�Ty���H��=�������UU\�O*�I��UE��oSŽ�����A�0+��.	N�$2�mg�?
ڊ	D
��n��5t�R��!�;#.̈́��t�q$��E�B3=������8�*�����F�	�ʏ����"�'�I�\�&�	6<]��yF��$Ӌ��>3W��1��^	m0��$R7?�(	��H؅�S9��&밠X�r���t��F^xB��eซ��xI�I
)�F��l���:��Β����S�hއ5Tțs8����T���H�j��x��rku��Ws�����p-���v	���1���U<	�E��:l2ō��6o�1�8VN`�i��Y������v�q�C�M��<dMű��ƈ�ي�!:=��a��V�U��O��w��E�(8�$1���+�a[�����t"��N�C�ef�X�,����W|�)L|%�$,<���O-S�@�T^��:�̀�lɟ0��<��zd�`�xu*�i�$���d!~1hh��Dژ�ހ�Y2AW����7����[zjʚ?���SMM��J�U͙b�nd���*<|�,i�񶞡�z@D����=����w��l�=�#�DFX�&^�@��A��
ب��d��״��֏�.���C�u�!	3�8I=��,.���0���;]���`n�ɺ�=ϑak�)Zd�Y���e�o�ы�|�0�f")=*{>B�%�f�з�ݒY`o�/IC��t��w��&�������K�A�~M���φ��,�,Zn�G�-����[.��T�5 �jsG5���>�%i!Jb�1t�-Jg� l��dh{dN������LP��/��걜��Jȫ~��������n�<0���rG�j3J��`
Q[�d���j������/2��OhI�%������ ��7�hh�V����� i��tϫ���Ն(�{�G���-0��� ����t�� �s��� ~{���wh��F��C8��Yh�W�1k�m~K;5,A��35�;�,u(D�x�G�OۣE*5�d3f��,�p=m%E�wV�X9��k*��/�r�S�����E� }�����g��"�����Ѵ_�ς9F�[�_3�z� E�(��Y�Y�ip{�?Oq �+��H������*.�i���v{�!�s�Bc6��)�J�\߶�%���spȟ�}w�lZ(�I�V'���4N9��-���q�q��83b�n��Hģ@_�"Gw�k��E�\�[�Q8�VP�ݨ���%TT'F�`3��.|�j��%�Ik��f�_��g��u`j`7	�����L���Z� ����~�1�(��f���Y� ��R�"=�:RE�B6��V\k���I��g_��j�qpm��KG�`x�yV��c</�^��eD��m���3_�3x����P�,��#���dA[�Ϧ���{�J�mVj�ʗ��!��$0F3-TZSu-w��u����=�
2�ئ����{�[�!ۤ��Ԥ{�7�IHv|�����d!����B��h���=����c��́�@���"��7`�6�/N��Fe�[2��D�&�=,|��T
韘����Sd�_xiN�����!� �F�8.vkI��=�z8��K�����=%�!R�x��|��V����
銜�=N��tI��rJ�үiR��Ro|!�#`?�>U:D6�}y94WwҸ4���=w�d����W3�?�33W?��i.�!]��'��s?׸��X��_bg=E����Լ�X���w<���lH��̉a���E1�6KV����Rp��-c��1.��=�TO�X��X�����:�s���5'3����㩾/��� }�FQ0�t����ŷ�6��Iˆ�v?R0��X�=Cv�~��J���
�g�p��n����`x���aO��7{����`O�b�� �n��/���d����y�@#	�o��������1e3�q������1�壚m�n0�m�2.�>F6�R�$Y�"�!?]�L�/�w�xA_oT�GUJ�)���6�y^�� s��jC��C�&7�J���������1���;2�q�wui��W�ɹ�/@�9�v�<t�����	�XF#mɺv���!a&��"����5��Y����7�k��Ci��_ )C��oE�`lPb3�P�=���B��JobۭOh�`�<�/
[�m�ٞ��) Y��ż��!ӠEF�mo95)�+@���Y�K�0|
�.1C���&�z����u��Wp)�'89�|�B�Q��!}b��_7�y����$�K9��Sׯ��X�^���.Ƿi�*�t=�Om�^�̥i�����Ĕ�c3�
���z�u��dw���
�i�!r)C��/Z�H��Lя
q=��,9��r��0�a���"5�2R�ir��G�%�H�
�/�S�G�b%��Yw�U���uvjQ��2{.z5�5��{N�@?f�U�<H��3�e.�O]s�#��X�~EA��&‴ fN��v�M�^:!..=>#c��3�!�y��C8�������S�࣫\Lm�cb!�9�Vr��*�)��?�7��+7��P� ���'����o�6eqh�v����?���Z�Mv��_Z��4K�=�����Y|����*U��R��L	�BP;l �.b�gF���P����c!�'U�|�a���
���m�6�m�C��8|Ž�σ��d�J����ǌ���ҝ]���8���"�]�~����