��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$�ʣi3N����ޘEWَ%�R(Շϓ�l��:=���CW_ь"z$|�~u;?z�]�Z�8����j��޲73L�`5���ehM���m[���
{={��7�M� �Ɯ�g���=�T~g�✓A�ߗh.����S��Eap6l=��e]�S��ZI�q��*f�}�Ʌ�s�X�"kJ�
��<x{6�҈���C��ʷ��eO&i�V˗K��.b�c�\E�;/����1W`��03�֒���
�=M"��}6��6E����W_R��wB�b��Fh� %������N`;ч�%|,W�顤&�ϙ)��1�ˊ�-���`��	����| 0������
�l4M�W'��ȇ`$�M�Eu��ݡ<��9F����.S��Q�A���� �e��ЎU@��ʋ-�Q��>���G fD.��۰���U�9Ҏ[�N��b/�ضhwk�X	���o�� �^O��x@�æ�>�p"��\��2!��14�45�r�	��JWzn1�R����F�=����Va���켏�c9�o劔�y/Z����F�G�'�ϸ�i�yX�/a�6����i$"�`��^�D�ӂq�!��&<
�
�6��X��8�]C��������#�f
��� d"F����B0��|�uj=W��s)E:�EL�X�\�n�%��ݷ̇|_"��9�^��F
.���SQ|5�T�j�M��Se������{�֡�+�*��Ӂx��G�Y�}���<S��0օqu�q8ӥ��H�#�:��c�)���f��g	�ۦcW3����gkȯ��JPc���)
�`q�	(�t�T7�{iu"݌6T�"4)-�t�c���r�x�s����E�!�@J��"k���������~�6^��H��!���X�HHQ���S-�۹z��`n橅�W���T�E�z����s�v�7��O�K�|���gR�^�1ݽ�<2D[l���pF��f�)0n/�rUϿ�늪�t�rVy��[����9�.�+wٷ�b��[#\�x���B��:��`�2?8�����Fw$�!zl;\�\�,7��1�{���Om,����k 5����-;U��
�DG�٭�?�/��ǀ�\������+���(�&ұ��u�NK~�ё���4Q�h-��h�8���������s@G�8^�� I�x�Y<9&.�>���Ðg�}��`���ڵ�MF���,y�<��2;*�1��@0�h~��Kp"ã�f>u�hC$W�����[w�
룊�t�F�OShA�3݁M�KQ*���i�H��!n����Kْ#�"JNQ���h�!����#�	V�]-�C�4:ֻ�O��Lc��5HF�V��(r��%z��r]u��\_g�+"�� ��/�.� "�����ـ_���oL�Oø4�h�%���b�;Z�� *"e�>�Cǣ�գ�K��o���Wڰ��y?�����Rv�����A)��vɣ�r伺��݂K����V@��Z.�6X^l����)Y�y����JeS��0�J0�n��V��\i��Ă>2ȱ�a�C�*Lq/NŮ��T���?Ɨ�2K+�xjDp+\�4�c���I�ς�L�+������p�H���&�P�B��ȿ>��+�|!ғئ��r���p�'}��޲�bX�" ��F⫲�
MiAp"� ����V�	�GF�,�Ƙ{c�J�Q�N踞bU��^�ݺ-���u:.m�/,��}��o�ڧ�Xǋc�����t����d�]rn�4��R��phYh.
uz��C��Y����n�s�LR�r/B�T�M����1s����A��k�M��]�)C�����ǮR���|�"�g�F��J�*�hyOWЗ�D��KK�k�r�m@��t�P0_%w�֊e���%E�ٍo8��_�6 p$_w���t��E��z�UAaH2��ܩ�'i��LO�����/�C�<�=<�ߙW���&����.Ilx��ZLa`K���)e&�"/7{y3��6�Ĥ�~�^䀌܆����k�T�\WP�*�#�O����#?���W�
��w1�T۞����I��_�zW ׷�\!`j���L��,����[EՄ�8[>9\5�К�[J��Q��mR�O|�X��1'���%8(=��lϹ~��TϢ�"lZ�H&���@m����>��++8(��uǗ��C���@�3]��gO�����2e'?_c��"��[40�癦�f�<�=e����>��#�y8���n���@�-��1$\���ߏ���!�?�,p{w�3��hBu��D���te�6��}BpM���U���B���Q��q��~���Q'~?���J׆�/A�\}��Sn�Tg�9��Qs��2�t�[R��K��	 AΩp�^岷���+���`�s�p���@>ǐðQ��9nF@�j�'���|����|Q��Ԗ����,Öf*�&V}/L�Դ���I!�HVZ����(���C��Mv�_1���'�]a([�N�:�3��$�����y���&���5�I� t9�/+��+�!��]Z�9�(�J��g}���&����⁜:���� >�(og���5���a\⽿YB���T�BY�@�='���R|3wR���-��в#��Z�P-�ĜXհFh]?����`��ܑy��ƻ��"��q�E�}h=sW� �[RAu�sqx�H�l��X��B��y�ߗp{���H�s��v�~�4k�h��i��s��1�tD�ʹ�{�n� �B2*��)/������	�d����oۥ�v�A�����w����|�W�*��4��	z*�{-���L�߁�{�204i�n�T�J�ަ?>0�� �l��s&p	h!ߨtO���W0uDe�	�l7B��JS&�H�-�4�PJ�Mߞĩ&Z^o3��K��(] ��i�{��M�\������h��cѭ9H��Pxp���ZZ_�>�芈��%����K�����vQ{����=��SX�����_���"罄���>m�wr���R�a.�=y������{g�D���U�ઌc����~<i���rw[�X9��{�h���zV���.��0�C+k�-������u��nzj�����_&�E�R!�E|�!.꧅����.�`��T�<���s�4|yC�7f�Y��L�&�l%�f��"MJ'�+ޯ�R�3s�~aT�9Q��A;�F�| 
�Z���o8��!��X��z��B0�����Y̤�^�;B��-��zl2Y�6��"�#�B��o���5g)��`B��Һ�8��4�4��A�FY�<^Ϲ�ðB�ӥپ�Ӕ<.V���=���6��%�m��me��_�H�.����Z[�Y�iQl%��"w� ��Z���V:�A`�P������'��m5�`lG՝��<W���n��|�S���v���$��&t�����M�t�(�;x�-r���AR}"^+~|8�'�����h'z�Z�֟��8������Սb�#훠�m�&}��RC��`���'0�+h�]7/	��>:��{{T�A��|�k�1��DI���D��+�`�������z��)U̱a��q�y#[��z�Pk:�.sP�*�f��<��o!柜�Y������S�Ti0��Ā���:��L~�������4�Ã��0��+R�".�>��$"���6h\��+��	`�]�QԒ#:a��6tx#`�E3Z�%����ļw)�*���8����C2ǱG/�>�-~E/��KZf������z9g:L�;-J3i�����ۓbB�8��ލU�O��W�E�F���^���V�T�a�ƅkW��b�n<x�Q>� ����Q V�`7y���P�/��#VF��t�t&�|!�́I$M�/�-�<�>�u��p0������NY�`\��ӄYU| �`t-�.��"�5 MF����MΈ��=��D�'�!5�?#����
�+���f�4�������z���¢QE	F_B�4܀���hi��y�^a�>}]���*b�Cg(��Vy��X���������0�4*����OR�7lˍ�5���uTx/7L��7��������8f�ͳ��7��<j�S��prK 9��ȕ �A������_ڟM�@���_HKF�H?��[�
�y��a����'��M�mm��,��z��\}|�kd��݉z1"���B���U�#^����b��s����VS8�!�+�E�~��$��ʚ�� j8�s� �JBs�	�S�=�"�} 9(�z}���\�E�v�j\���)�*��C���CH)��i��}��8�
R/���Q�g�~����N� N��|3�p�"�P�M9�^�sf	��βo$��d_�V|�2=�����	�+��h�Q]Q<�������p��;�qK��T�wO�d�����m�.-G�7�m�Ű��}�BJ�ԄC������vx|P��U��3���㼑xC9�RL����A@!�zS�[�B.��:a�D	�����o��ܥ�0h1&xT�,��Q�֊�;���m���[�RA��t�N
U��=,,����D��	E%�3�m�y�8�t~֮�3$�I�reg5��C;�.jI�u1H�x�Uc��{��E�8�^~��]�k���O0�z�c�t����f	�˞��&ϧ�W�4��0[��du�^�H�z��C�%�*�~�>��,��'^~|Ȥ�:Tz�I��"i�{��X�fK�����!�r��lR�����߫�E̀L��U`��Й��S<�D�%ۦ"�kr�]�����is��6���n����ʧn�G,6�*ɐ����54�UuOZ]ᩃq��
H� �U�e�̖�_�sDk	�r�J�%�R�n�G��$.����Fj�a��{@ju�٤k�~#�K����]/�lR�:[XO'���|v�G�iR���z���<\�*���
�
�?�[�X���U&��-�������C��ɦ���@1��Oa�>�{���S,�?y�g�i�,�POٮq��Yo�
Q�:�9�����? ���;���T ��F��s�^��g��̌P<KՍ�������E��>�j����\|����]�a��+:[��$��{�B��u��͸s����?���r��@���bW��e�j��x���F�"�k��b�