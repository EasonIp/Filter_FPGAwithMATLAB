��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A&Q>�Mx�E��K֎�>v"wTD)3�2C�
!h׮X�L��,�]�c�:��]�D�ߢX��xs�YW9�=�	]��Y�����&����	����_�͚����܆s��.��F�5@e��1���b�ͻ{Uz�2���Ƀ��������[�����} ��T
9<븇��b�ѹ΀��z�7:C�"{��K���T"����P{AKM���c���,�3{u�?��L͕(0�,W�m?;�b]�Os���!]i�� ��OXc1�Ky���Ш�u+�8��`�=M5'@Bqx�2�Rc��,��=ѣU��2��o����s#s����p�[��M��	���kE<�b�|l���iH���;`�ΰx��e�@�)���tyW�[+�a��Ω*t���R�(����)n�,�X��ɨ�z�[т��a��I�t�3f�'��Bzf��mt"x ��|7M��NJ�p`��hzq���W���]�i�Fƍ�p��i�ߗ.g������"qf��ǂ 5���ԓ����Iq�6�s�2L0�>��D��w$��cM��w�:c�u�_|��xԇ�^i(����):b����RR�[@FQ��f����
 7��J�C��bؾ�vW+?���*���#Z�*�Ҁ�`Y��)L*�E�h=9U�/��oeh�Q��q@�Q���.�r-|�� �]�i�$�`xZ�i?�
�� �t�4��@"ܙ��I�?z�1 �*'�*��"�'�H�2�-܆G'H���@�}�k���@�oc���q��,�����FM}?�!c~�͎�����' �p��uT�#����A	+&f�K�6�VM��v�>�,�{����O�jg��0��|�NN������.U7�h?���q7��Kg�^ �)�Ig&s����0K����`�J�HS=�3��S�AJ������z p4nqd8fb�~N��q�e,�oZY�'�Ғ���`�!DԳ[ڱ�<�c���7ck@�����q�������ؒ��;�Y͸@&��z��&]�Xs���CT�Tq�ar�2��DT���O�n�-}jF*<Q�����"^ﳊ��5��_
�$N����iM����dPZB�i�^٢ �#"��L���m6����@L� �L�+9��J�w��x��\����"H����$���8��~��R2��r�S{ZI���R
�fF��C}�`�J$2�B����?�&W���&DϮ�A�/�N_�vg���w��u��p3@4�u\�<]*���Q�oK�wو�,�N2��L�`J����K���t��j!0H�^�e��d�D7�F�]��E�Y1`�=���gϖ`�`���qƴ��hT�S��� \�T_>K6���h�'���	���H.�+��x}��]J��d�+��׊.�IB��eGʝ�[�؍c�a%F�ba�a�W���p��w��(��������"�3��xo��\T)�
�1O<"���ϯ