��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>	��։�������7��*`�ԇ��h��U
�~�a�������.H��N��Y9Ύ�2��3�MT�������-8]#�X̵���lV``�^��k(C6˞��w��7�w�T]U:⡇J?��\f�խ�@��R@���>I6�Y������N9�F�N�)���S��
VJ�R�hw�@hf��Ko��J:� Ȣ8�j�^c�AʊAl<H��I����k[����г~�f���E��ت� c�yz}�WY�ﵕ�jΫ��P��.	9��t�o�r\^����b-�@�	��0�Α��?>xT÷�ln��$8������8���$�����A�����]�R��������%�)�X���H�=�F}s�_ӽ�S�&�� Ӂ=��HD����6iF��a҅�$��ܻ��h��'�d��qc{8��2�=���&��b ���U<��R�}��Ra��|�YDq禽f���z�Í�h=<�'��]w,��8ws�nq�o��I�{���i��3)c�sPU�=𠣪p��s��稢�$d�%w�}_�\��Xl˖��o�*���6���1��PKV?����7`~��?�3
"߫��g��~���?i �+�;c�gX2/���_m4ݫ1}Ņj��_%wf[͜�/�>��2���Z�-�9�\{�K)�+��!T����X~�p��kn> ��-AH���GB�7��VQx sd���&�;xݷ�vj�v�ޘDOw�R��f�u>ɔ\ծJ۽J0��jq���"���ޠ�v�0�2"@C��S�ڰƵ�^��XR����B���w���N���D`'	^��*��I���d����p�6�D�dr�p H0o�X��;9e��(��üt'��28��pM�@:�W/��1ĄF�m�fj��:h�N�z-�C1��;���]!C�'p"2��)�g���aE��ϓ7>�B�_&2��B�ţ���\���|��9���piR��n��dR�jS �!`#�QI��"�&~�ʖ�մ# #��/�r�J�U�7.Z�ϭ�`YS։��V#���	=4�<�8&z��V���{� ���a?n������C..*�C}-�g�����؋G^��㔫���ҷ��=�@��i�cیV������Y�U^LyÆyl��3e��o�Π�9(W$�*���g��9�:t<����F����u�_��4ڜN�����ň[��\����fJz82'�����pg:���Q��b�L�e�l};���4�=�Y�sG
i�{��?�h��w���k�c����s���X�$5��^
��nYŭ�3�=˒��eSY����]�0��m9u#�Q�|��#0L��6�M�:ce�e�Q�J!��C@�jE,�7$�L�S�vč��3\ �^e�g���:�_c�1���@)2��/$�)��)�,̕Tb^�2rJ�x��CG�+������v�B������%�oOL․�"����8N��Q'����ܥ��Ƒ�V�G���xZ�!9�؂�F�2�g��(�ʢ���^�a'S�y|���v��0 ����ΣjlQb�P�*"�m���ֺK�f<��H���Q����0)�x��
d��N�"#���.�Ǘ��ma�Q]r;�}�(K��M�+�����̲3���.E�g�vy���׾�&���e���,��S��|���{}��A��M$Dh�J�Lr�c�I��T-ʔT�{�M+��_���,��,�ѥ��ı�̻a�4�/���\7��8"���>1�nd<?�y_{��u"�jXj-J��鵥#,��X�{�����9r1ϙMAĊAǜ�U��:��^��Ԗڛ]!������5�4����0S|���*̌�#焨��A�/�b�U��I���?�J�m�����xQ)D���$h ���aI%u��=�%�D��<�����)����kލ��x�M�����}9��B�
zȱ�������Uz�X�C7CzU&^�����5XqM�j�g$�ꐂ� ��bQx��[�rs�Ylˌ֨㊨�[I{5h�>=IP_*Ж����{&@���J��-�U�e:��g��a�%y�,'���N�%�bt0NQKY�yde�6�_?}�p.���Y2n+�A�.A� A�HX�㈧����.�	F!�����KŌ�yM�cm}�lkU�гQ�f������$Y������KgR#o����2�s�Õ�����?�ȝ,Hp��N�1ܿ`�Eb��C0�Z�=�f�64���H��n��m|ԛ'MTn��(j>*Ue�,ܘw��3���t�.?���@�Ӑg���b�z�'5�%�	6��!=����L�2��wu�'T��L�U��@1^�� �x�n�Z<���!�Q`ɘ����~=9�F��d�%�
�‌�Δ]Py�9:��8�=����r�������
*�{A��B�km�d)�O��࣪�'������[J�vA�2��]<II)��ђ����aD�	�0t��#�O�J���=���b]���b+0�%��@&���x��*o�>kt��F�_�Ǆ�}K���q��^i�7ɦ�3�Aͳ�c�7ڜrAq5�nY���sϔ�����QL���gő������ ByȈ>��<�K�ٍ��cx��<$+
�d�hW �z��n������>(l��fv.f���dy�>5��x$ͦ�JD찏�O*�	��t=D�;���gu��Ƚ���)�ՂƄ$�CN�7�e�8ݤ�No�_9�b�q�af;��·�&��@΂�q�j�	#��/�����dE�����K�͟��t1�gQ����v?р�k7�9&�l��Gn4bj������Ե�>�L�0u�N�v��ʥT�c�f�j�;��/%#��+-���Z�bZ�TC�'Xh
��x���0����"k�pB���F���R��H�DZ�
�b��2�ޘ�O�\���⻺�%ܝE��ȭ?A>l�Ӻ�r
3>ƽ�%m6��:CZ�`�*��&fח���s���D���������y�aA�f־o1�������}iӵ,��ͩ,�{��VJ�F�|A��tx��_�юa~m�!r8l��Pa�ޞD�wu��W���!s��i��] � +��� �8?r��.�RO�)���7ō\�'�
Q�=�8��\�\�P��M�y7��e˺��!�3��I���'M��'���Y�!�
 <5����e�l�a���������*S��la+r�c�f�c��r��#�A�WG�˥�(�t~r<ejH��ѕu�K���f�iϤ�;��`�R�;�?�3��x��L�ҧ~�Y� �|e���D��W��^�@]�?�e�ke�!����x����ѯ�@�g7�j`v[���1LU��Q�C�����Ú�|H���2��IV�7���/��݌��d���4	�κ`��� �����㤒�y��h�S�5�nE6��[��(���� �m��!8�M�!�ݞӱTab����.^�"���$��;m�V9��[��8�%-۔��;*={���q�qD��5�=�u�L�$����oĨ��P�0\=�sQҁ�3��Q�%ڦj�r��c�m�
���P���LYo�A ���2K �;��VrW���(�̄��e2�b9R.4#,G�Gn�z�9D;�Kd�M���Ƕz����-g�4�Hr��#��A�A���}��&��X�X/�d
?M)�2i����m��)�+O�|2��_>V�-�ڲY�˟�j�j=��>�mO��~1�/��`y$h�=�{�wk{L�������b����2���nM�c�7�����=�̥���N~����e(�}d`16ъC�� y� c�3{MK�׳6���Vv�N�K�1 ��y\L����H.�p���b�Y���~���b�ap�r3k��G��s�,�e��޴6=�V�g�.������4XC���I^��RR���[dPm���u���~�,���8�"I�R�W������6�c�=�Y�hy�B�Y�������~� ���k��/0۶�F|4�s�4�!5u��c�rG����kM����w�B��+I�d�XK���C��t�A��@TK�{+#�$1�H˰L��h��wQ��_���A��'$������<�}�bFl@B�x�Me(p�Q��i5�}���~I+ ���ڤ^�ʋ���5pXL�T����<�ߍ�*ȗ������=���ـ�a@*e1�Y��@�N )��b
�d�n�`���͋����ey���,����~ėf�VU���gfK�e��fRS�����/ٮ"ȵ��+�([&_��N��w�^�@��~&9��]�@�~_�P���(��
�A�h���_6��5H$�6,طfvA��]ɓ[�3� �`<�{�c��B�Rf�i+W�n&�o�3\��I���yΗ"�_v��\��*Fe�[=��Hs�L/Bm!�WVl��6"�����&��^�`U��F������o
ؿUݚV���9�3�W�i+5����z4����%�S	9��b�f"@��s�M�9[���N��ư �@ծ���������M���+��^j��aP�!s�(A�� ��n��6�W����4N�o]���t�.R�b�/C���h����xNy��_����Nqm�����'9�?��j �A�}kw�V��W�x�����a?���r�ܫ���-��s�l�_T�Z�	#���Fm]��K B��3t9 FXP��I��jf�֖���Gp�~��ǽ���CH[XN�,-�#�T#�f"q�\@�"�1�xm�M�m��bo<�E���C�a�QI�5H�l10@-5m�t^�� D��θ�+Y�q�<�¡������.`~H�؆d2�ʳ�:�֋�i/� ���<S��Vu$F?��'����E��HF����u��z��X6m����r�vn^��C<�F��<��t���i�w��jn�H\�o��2�@�?�Z#��bF%����7�h3{���*�<G3K��qS\9��X�v#}��R����.1�dƵ�n��%�ML���"�i:��Bl���}�D�Qaێ0�zڞ'�K�J�%�$����#��;Rþ9E�!��;�Y{�=V�
�XTh<���"����E��rH����D��W���Y^j���c蟻x˕C�A~�[i��SF��#��&��`�u�y+}���@��5��{?�LU�J��/P(C�����ǖ ��o6[��f�t���'�^ھ�f��*�ys�Ͻ����;Ƞ���ao�ɕ��@c��N���I摚��}�:~���B0}{�-ńFZm�.��/~�>���O�|�2�u#��������e	�S=n)�ҿ��+BX̳ر�jN�Ё� �8ݛ�{��.����9h&o��e��� �F�SN���(�[������h�IE�a=sѠayN8eq̟t�NZ���w�"Dr�F~�
O�T�Z{�;��j���j�9fwf
��8~�>�gT�LHF�"}�fmƯ&�����-$S��a�vܸ>��ca[P�� ��y�Cf�
U�$X�����eeO3"7��]n갿т"��%n-��?�!Z?MIS���n3j��s��̶#��7�'U��NJ�FX����K�K��Y�G:��c�����!H�țd������0�ow��h��z�ag�?��sc���.��.NRA���R���?����Y�Ֆϝ6J�ï�Et$z��4O�c+�1�I��G��ɸK���Q���0��+����dn3��|�lV+��E�BHD�f� ���o%�v�2d��d�dH#R�]�J]�6����'��_��5����NWUn��J�3�x�Ig�Ͼ���¸��q�U^��`l�β�����z_p��6��-'ġ����j���_ڗ��=
�����q��Q�a���r�嚳by��֧];�}-�}E��&Nˠ��8�ѻ�E���=2e2_�)~��Ir$��%��)dji$���j���[���n]|;�g~��0�kCQ�S����<���a�l0?x���� r�j���Ql��I�ME��G~�I�y8=A�(��1ܬ;�/����K���	Sí?���=�����0�F�L��jz������y�z���lf�d�~q�wi{58 bR��D7̫>4��%��"f(!6IƇ��5�dNu�[�4����1>���k��m�����,�clυ2���F�Zr\�e�K�*������wYdn��&�!���S[��,r)���^c�8Št�&-��;���^u՘�J���njvNW��������x~F�&������G�"�:(�}�	��9��N��,M,�ќ �Uli���~.>�Cϻ���>o�omÕo�z��l&����V���6�M[sf����Y�(�ͼ�=���
'�Zѓ(�8q&_ �B��*I��ě�lC!��1?�s|D����%a�d�����eO��h?�Rp�k6���.�T�%�G 4k���נ��I��T�a\�B������;�~o�:
LZ�٘Ɠ�B�>�:���[�q�����{BOz�tmh-��Cq��׾!���6l�l��V���D�g}3�;�f!����R��]�g�5�B0�[ �3[��gWL6��)�Of~^��%OK�(�&�	�jؽ-�?�
l�#�D pe,�	g��<�_xj��/��o�m�9�_����Hx1�3%Td��Ќ����ۃ�Q�s~Y;1试�e�b�0vQ��ȫcZ���j�y� �)�X��*�!���������Ix������+l=S�NX�m��@���2A�3K� ��:�L&k�j�8�#��{x�^��-��ȏ��D�\�f�i��$��� ��Oͤ���<H�Nx���4n��I_P�]����\�m����Mm���Þ1��݃���'�t�5. a"&�ߐ<�3wO�a��y�
%��ה!Jn|ThU!=�c�G��%�U�W�]���t~�Yy��Sי�9��Բ-<����J���>��r{lI�8U�s4�,l�0� �#'����]|����8!�n��\����m,��eK?�RЈ�4��}��]��� y�4Y����zUJ&��"�w(���~f*
��:B