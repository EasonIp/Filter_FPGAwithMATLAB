��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>hs�*�U��Q�����vXH���p�+ׁ4/3��T�?#�ھ�ь�RT����u�Y�����/�Ti�歀R�O��5��s��
�rOK%t�R�QT�� �>���Pr�
������:h�����"��I���*�P�ne��M�O�	r@�/0�,/���Ro����SI������޶��B����`o��~~��n��ߐU��$喠)�� q�L/�����q�E6#b<�h�\�����m���"�`��
d��3�j��G\���O�@o-"����-�&�3Gt�@͊]5�{�0�FP�L���Db�������>ti�.܃�ER9�賿%�o��/DI)hc�E5{ _��CF��>)��)�N����ؗ����H���iyBB��*��!U�������e�g�^Ug�*��ß�ρ5$V sw��+��F|vΩ�����
��83�L�SY���ҏT*}�u𳰳a��6p�)�]��Qw_�m@�X�iz[,f쿡[�X~L'�����Ǭ;0=#�`��K@�S4 ;�3�)�Qk�����r�~�̴���%Ѭ����q���v>�k��A,�$��W�_���3�����.r�nW{�.LQ���st�������W�v��5�T^d�����6u�h5���x*�&��o����
�q�fN߼ܝ���.�'�/Y���(Z2��k�p��ʪ�� G��W��!|�i"2�"br�l��䣙�:��#�lAW!0��R�WS�\AbYV�\}Ep	�[��8�֔]楼$<FK�^�����йY�A/���� ����Po�m�!�c��SRAP(�~�����7	��
ߑ� �3픆�l���q��@��=:8ӎ���o�������qc�
Ԭ�y=D�� l4����u���ω���<Vu�pE����
Zq]���aB�	4�zNqŷ\�)���(9�j+K ���f��#�E�j$���"����zufo�\eZ^�|�i�n4#&w��k �����ԑ�>���O�H6��#AG�҇���(��\�	z��3Z{�� ��EF�%��h<�c�9����S~�B��'�*Q��`x���{LP���ޚ��I��A�7���Y]j��$�[�%����*�f�c/O�s�V�
���	^�A�h�k2���Ȃt��1L�|��"g��
��7��$����5��&��tƄ|�.���}�qh�:j�P=څ`.'�������Qމ��"�W���� ��h<��H�匠7E�F�񭔤�+1�f2�~�q4\-���w�]Z���ȱZ�m���)5u���n�>��{�^�%�k��d�X;S�n9�O47�5�07��c�vW(��-Z�	N���N���%�łF���6|��(T.�bEJ��ϱ�Q[�!�p~��}P~sOWϮS4��qI,�U^�9���DH��cE<��~�G��df\�V�C�T���m��~���9��^:Ѯ����I�L���ݫ�$��-��ZTt���Tt���h��w���z#��z�$A�ϭC���m�vvB��I�ڃ�9
 �e���3�_h=��O�c���h�L,u���v�L5��1��z,y�.bV���.f�?���rF���ı���͞Qvt�Ug�a�ű䎢j�������n�i��4��6���(�+�V�fz���X}�����]����eA��&��H����Jaӂ\ċ��3��'n�%T���#(A��HdH��Kӎ���|X�z��`�1��;�6�J���MO���8V�c�#<W�FZ��sv�n�x��q��q�IN�� tk1�o�P6M�?�2ue6t�5��©������@j�m��Wk��;�c��&t�c�G5e��J��F��x) n8�]��x:D�Aؤ1���)(6�"��B���$�c 5��,5��
�ܵ�zU�f�^���n�(�3v��M�=Tq D���䋞����7Vz�VJ�9���r��$Qpd�����@��{=6��[.s)�z�]���2�����ۢA�h{��͹lx�v%�7�����q;������ޥ`�8���d�́b*�ֶ�.�U�ZpjJ��gF[�(�I�$�騩��q*Sh UG���1�[��ZK�6��@���y^3��F$U����*$ik���O����ɺ�@ǇN���83w>�{�!���w�%m|�OR���N1�"Y�W��G��^�9��Ȭ�%�=���w5���S ��F��)�j��Qc��� �=e�d�=�Y��g~��w6:x�vh�DC��O��[&B�a�g)���6�{p�E�t�`M�7�n
՘u]�+l1���_��l'"K�Rub��V���̚��|�@�Qy���bx*���5e_J�L����Ǽ�'�-ڋ�{�u�z�杁�a��Ƭ�_B��JO[�j��0�wRx�]��+m�l�����F�wW'˩����[�}�/��39�����X�ܚ_�U��2����R6�ld��_T��Ň��c��;N�_�eX�ND�>����E�	��pFA"�박�9+F�?�o���)ꝲ^>�6�۱<��!r4Ҳ#<ɤ)X��|��kg�&i�T7�\'�������X:lb`♺���^bN<fxG�<�m�?�鱳��k�;<i���nI�G�<���J���a��޹K�L�tCOk���"��Vp)��֋�6�]R�X��t�[(l]���c��oy��{#�����Q5�j���6r�M��m]:H\~ľ����ѹ�I]�G��'��d8mN�E�o��R�Z���t��"���5K���+�
)�s� �S��j��Գ����'�w�ZD�]����;@����F�ʡu�jν���AL�E��Ga��-5{��E���{՜���к�Y]x���}.��-����:'��LQ���4�\�m���F��få�lS�^�n���/�ܔL)�R�_�~�v�)�M��U�&�9��D�=�d�L�@�o�)Д�5�Z����5����ɢZ<�z�#ӯ,f����Ӑ�(�8o�+P��hT���8��R�s4��B�=,�>�ꀿ����*
�Pb����I=��13�o��n�>`}���U�'
�.h�vO2�cǽRE�Y�x�~���?󮷘� ]�T&�N��Ȼ���~cC���N{>�l)5觪�uG�k�+@`E����˓�8�^�c��FЯ��E2�DE���x} ?��L��x��S��'�-*u�O/i]��{k�Z:��C�B$�Vqh~A�<#���!�S�ϸþN~&0���>3�O���$j�8��G�c�0�B��0#H�h��4��URwEe�P5à�t6�>�vDz��K4�u�:���*�DJ�"&<4� �7���>����Ƿß��X@
�Kn�V��������<��zF17�:Ԯ�G��d�^�{tŀ�G������CKR�Q�=�
Db�e--P�@�z�/���pohdd��BOL�O"$H�]�R�TU@���L.���W���5�H:M��9#v+u��G������q�4�ɒ(=S�\���ۦ����cA�jǪQ���]r�h$e��|���M܃�'(Z�S�iɐȚ��ܵ ��X5uQv�u#p�{�I��jk�����5���	t�)/����l��]�T�y��i�A����z!������oG�޳���ײ~P�1U���/D�5)l�/Ӏ}�[*��m��*i��V�k�AN���R$dI��S๢/l��i	�G�5�aL�&O�i}�Q�l8�|�Ȭo]�+ۉ�[��e�n�M���u}�ɹ�a�"�oK�m��X��(��� �I������t���G~�X�I���mQ^5�����7����n�&W$0�*'J�4�mv��q�eqx6؏`Q�C��N�?ya�����W]_��Zɛ�n����Յ{�Uf�IN�E����Pee���1���cn$��x݌퀌�-nm��;y�޻����
lG����Iy�	�DŲ��}Al����� D3ɯ@A~�D���Y���]=A�C�m�6?�@i�U}/���^'X���;�0)Z���ES6�dDn�3Q�:2֊�Eʸ��֖�2ۆp��e�в��k�_����������d�x>*a��1�k=5�<H���/���R�B,�+����m�MA������.2w�J=�'���9���M]* ��l�X(����dY����ڼ-�$��S��^Q���8&A�2×�����P�z$$�<�1����-�E��j�7�	i���ۛ�u6c�B��$s1�]G��*G�ڪJ��(�U��c7��GҸU�q�%��Es��;L�g����ʡaӓ$U�R�6QA�ĥ�!��g�0��n�L�zo�57�ǁ`��?�\�9��m��X�jq�q����*C��5����+��n�c��}��t_�t5�L~H����a��S��ǞADΣpUwT�3A����o��	��z>��y����E����U
,��h�ir �����,��F�����4���G����LQ�1�r+�E��J�(ϴ�@x����1r*��ԍ�&�%����%�2�FȈ~��څ"
 �1I	��g���X22�}�}�ŵQ-B��U��s;��6�C{N>�>���=��<����Ɂ0�J����[��ηcIZ�ˠ�VF�͔�:
|��1��'��^-9C�¼�>4�?_C�� w�ƞ�t�ι�*H`�9�/���
�	��;N�ɲ1)�]H^�?�Ⱦ���4C��e��~�� 4��@��G˖�ޜ�ZG$2�k��l��_X��,)�_,�!מL;~I���fCu�$������A�ۮ=�;���80{��b�X�Ȉ��>�jX�������^�*5����H�D��}���:��nn��1�2%"�Z��y�촢eʉ!�B���E��i7�Ol,��@y���'i�����uy��櫠����B�Rg�Q3��Z�,gN6j��"�X_շ�{���Q2�g�8�K��,��Y^���&u�՗R`�1��C�2ă�k����32VV�߂R��^����S��<GN�J������r����
�(={�#�7;���T`DYNXH4)
dr��Z7'	&=n]�������x����:�с)]�%����nd#��������b�/�}зoX>�,HE�f�0BŸ��	&���p�c�PC���;�D����B0$G�b�	������zE３<@O"G,@&p~�آL���a]J�z:8�P���~�oў�'��ᓑ$ቬ��q���e���7�T�7S!�!�V�TҩB�����y#Z�[�Ұ�[��<_����j?�[��_�V�V�C�|䜥%ʹ��H��&ow/�=5f#I�d���(+,5�e��<m8��Ek!0���*�>�v�,x����koFӧñ�+��X��os�<��a>sP$5����0УL:�LFM+F{�]x%B&���0ҳ2፰e���?g��ĵ!���
��z�mӌ�0 &�aON�Gkv�>�/��W�|i�������nJi����O���Hb�<iKIX`T�
E9Ȝ��v2�+ߍE*�,�|J�!<�9	�Њ�2\�r�q�ni���X0� gс���E��U�˘ˋ�e܍)x>��T���=���n�����=y��"���-2�`�5�	h`�8��V��/��MP�Y�@�M5t��ː���8q�KEj��x�ek�tե>�������k�n��Gw6v�~c���0��d�\^Ű��o��ie�ж8���w�WL�۰��;.��̢ �JY�Ѱ-v1�=�N�K`n�'���D6A�تO� ��l�8R�sA�k'���'����9H2��qa�e�g����'�V����m9�ц�xr���o�f�D����[>��8
o*���2��۹�
���]��L_�l�_w������Tّ	����7������ I=n}ϊY��{q��Fy����ɢ
�SP�=Rn�ɽ/{5�����"�b�����r1\m�@��J|`��1�W��O�+E�y���)�*6� �L�3���"���E3o�ʍ��_FiE�]L= suFp���g�ܷ�S�������L�����,���7��w^�q�k%}mT���#m�ml��In%��D��TґTl��|)���HJ�¥yC����Y
�)�*\e�,�J&�MIQ����B֟�?� �v�xP��vYb�Sq�ĩ�R��B�@����U<9f�&I�MH��`=�O,k9�d)w���;�[nu�h+�Pg���X��6���9-ڟ迹z}rB�Θ>��^�#
�{�F�v�r)�����>Kyʊ�O���^����W�MS/3n�	����#�c�<_% i"�*�KB�#t~��ž긃��>w���2¯
˰��GFDҬ����d����V'>��3�����A!0�S�hFڏ���®Ws��.��L:�`,�+�a���^�A��_.nJ����O�}��X�9��iC�T~x
�	^~�Ô'��O���@,�?+��pnӢ�Ml<ʯ~	�57]�[�N�a7yB�]�#|t�}�	�`���r����9ɎQ,���).+���M �Ҍ��M�˸3���q3u��q3��a�1ܝM�^:y�+��dl0��}�}�I�Q�nw���l��Y�E�m�M���_�C(,��@0k�@��P/8�<66�LEdA%[G����4����ڂ
#J;�ƿ�����5��e�`ru�����^�M� �C���P�ˡ�'*h�8���\C���u� \w"�HҏX���q��i�Os>D�WZRt�CĮÒ~O���5�]���7=4Q�YkJ�C`�1������[8*��?~D�	i�`�_�wЇ��P�&�Z�/g�^����I����c�Y}�,A~O�,Zc�~ ���`��ͼ�2�Ϡ�}y�J��$����׺�KO�_�|�EA��l�0�=;���'�5=��ل9D�"I��X�$�LYBR���1t[i�8E����w#7��=+v9��]����d\���;���Ĥ�h�ޣ\��Y���]ذ������W�����ꡧ�S_�r�p����["Xq&�qŝ�PM�`*��臇�9#�hϹ���lb��-iEqZB�Bej�&�/6�	��E�����^���ߔ���w�|uh(s������,��5����L�,�v��J2�؜W����rQ�\�՚`�lI@���}ۿ�Ri��5�����{y�:{����R�f���G#N�0����B�ے�����Ԅ�RRka��]N������|�$x8Uu���'9�H<:�58�[z��Ҿ1�&��k�)����	���12�����Ւ>^ <;n��]*�,����C�!�v����\Z�z�A���޹O����d]z�)#�J�R���8;qx�I�6	>�l(�C��~�����?� H3[fm,I�ūIśX��9���hx#��@G��<p�fe���,��&D&j��y��rjj��E� hz�����4�*A�
QS)����@�Q띢v[�٢���}��{�8W���%�*�������tPf�*"W��r��A����b��7�g6_�ӱx����~�����.�Z,��$��/l$/ӇxU(�i��6���*7�7�uGS�i'���7�7Hc�c