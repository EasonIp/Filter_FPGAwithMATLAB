��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$�ʩ&6� t%�L�HC��*+�?:��n:��Ӆ���V��U�!�����J	��[T�r�rb�M*�gy^�t7�O���vU����߼�~�7{�7)*I0����[�ƦR�/|�5U���w��N���7E�3��T��f������:��hO� aȞ��e�E�s{@��Y0���+RA�,�Nup�+��@3�Ѧ��b}���^�z���>5�wG<���b�	���	��Hs}v�d hp����'?A�̊���~�-�9�����@�n<���g���Pv��֔
����ޙ	�A�9W�O����׬C��vy,8�d����G�RL�_v'����+=U�B�y��6�_����Bt�f�l�^(����miM���o>��.���m�s�)W/o��	G��Z<k�����X�~>��� �h/ϯ����-����Y���mz#�V�A�Z����A 1>�4ww�(�yV��5����=)y�V���%I�޶���k�Yc,���u� �둯<w�s�����z�|�R��Oy��%�/-1Q�q{I��[�z���u-��"�pz����+q��P�(��Y�*1Bw#˂�뚝�k�&���-ֹ�FQzސ��S��+�n��A�
��!���,��5�/�"���V������J��y&�_���;x^V�ʉA���j�p[e�:���mUŹ\�q>����Ɗ����5!���Z�)Z���+��b0۳v�9���f��+�Ĝ��ɉ��6�{lQ;����{�ǆ�xcB]��p#������F�,��g�V����[
Zk5o+*s�`�����)1-� Ŷ�(���b��m��5:�D�u�=h�)L�8F _X��F�d�ע=���=��z�G+'r7��u������C���t#��[)CD�e0�g�kt:`�u�Bz}���5�%�r���礥E�X��+8p��Q���In���1����&�A��.���h4����tO�BD���r�U��o{o2lz�{���"ӧ�$���_����r�҇�i���6�ta#�%�����hBŬ�l|�_�X'��w��d��cض����Gf$�!��	f��Ѓ�=��ʸf�ҡ�-�0L�s.#���\,�m�A��"�ןA�!]�)�=��-7��A�؅A��KT������Ɖ_���2�ˋ�}C{?�����K��`8�}pd�R&iE^܅j��y�?[ɾ^��9X������*pF���H�_-z��pZ�L@g<��E����L��f���Q��$ִE�O���X��ڧ.��]G�R�����H����C���eP�u���`=Qײ�,�M�ᘝ�K	�\�g��V=��i��(���3�T9;�Sd8��h������!-wT�D�X���v��k�FΚ������xW�Ӻ ˛77�5��Pڙz��� 
���'�CsF<X]ԍ�u;ڇ�,�
�F����4�����#e1ydKЪ��(�}M$K��}fX3�EB��UG��&�!�Fl�����q6�@�`�K|(H�~N�x0 *�2f� d�z{>����jGQ�����@�[D�M?�~���c4�\�AO�>�{8���w&15�+����hj�on�׺�$	Qz8k�|@Uڴfx`Vk�&����\&��4I�y� �h5��D*}�Of!�h�88�b}�t���E�L\���!��_[��r���#�����@�M�~�Q���쳜��Ʈo�2�d0h��P�Ȋ�����1�z��pM�A�V�A@3��R�7c򽎷�����m�Q%u%(z^샢��z��(�V���+h)�Ą�n�՟��/�#1����2���ۍ_�xC,��qhBܰ4=)��y�ݝv_�K]� 	M�U�9��\\峲Sǜ�?t@M��p�q��L?��uO,�n!�����J�.h�\'_I(!�$�)�guF}|%R��.�S|;�y(88��ܓG3z���0�)6�Q1���2TOf<E>6��s���ʂ�)�*�F��C+����$;o+;���hΑAp�~<1`�AIn�O��<�H
����̾y�����U�}}Jtjd0��D;����qS����i����SqX�ak:��~`�g��'d����O#c'���������iqhȘl)?Ӣ��å�I}�a��h��+R}凉�IΒ��cWL�Q2MX9��HY���q����՘�r�l����_\���Ӑ4� �dB���C�DP}`�;5�1�iA�I8�<���� E[�U�x<~y�,�(�=�(��o��Me$si-��n�Z�����E���(I�5W߯�7��A���:I�0@B���o>�[�9��[�@�Q+�q�4A��F�����'#�;=�@�APF���i�{�1��6��j-�Ջ�cX�1b�����g L`��R�^8�ME3l��m1��j+>Q``/ι��
���1F����A�1�׾�|f�O�H�;�{0NE�+n�Ac����l���4סT���2"_y:t�ͳ�,��*x^�Aȅ�a����al�d�2�V��lE�C�L�>j��.�`*�A���y.O�&�jV,��_Z\��
�6��Do���s���Z��#b�]��M�0
�G�[	V�M9��7�Ii�?0xŭ���;�i�]�-]�sII���u�ʳv�d�a�az�#nL�SlZo��cA���d���qt��T���7�>�7E��0"�{t�M�r�-��{ �C���X0�iC���&qiȲBb��0����v��q�F	љZ��F�.'az���4���OJ���l�S��ho�4(]�\ y�s�'���;L��� uD|�e���9!6�!I�g�3�)������VX.{�P��NB�6�\��s} 3uBF�k#@�{�y���T���!w�rѵ�ދ���7G�w'z8Y�(?�������k^�-z:eݜPJ��r�_y-9G�-!�P�:�ɖ��F�H�CwR���<v��#}G�u���~ ���P��|w;�$X%��f�����%m*��'��z�FA�jb�pQ�<Ό�AB[3j���F�>a�P�_�
����38E# ���ͫT!�[s��;%���h��	1I^����ش�~n�G���M6�(|%c�1K0��_v�Z�6"�wG�?�5��8(Dd4x#��QI���ђlR�f�]>��ݾK~�:�.��Jr0�Q�K�NC��R�BT�[x��y��ы�Ј��5���+� �\�E���P���e���b)�k�:�;n�'ܵ�L��_L�e��܌q����HI��c�f���1���N㞬�A����X�����M����)�%Q�-��e�[��²�8���G۟6E&2��0��ؕ�� M�&���k���a�>3�Ik�}i���B�>�+�P�G�R	� ����!��_�I+R�"�I�v��C̗H�QqkLWIUqi��O�rH���`�,��v��2hb��qv��tE��.����#������&�N�ZT�[X��i��sa�����GZ�/�S�Xn��м`&5���U ͫ,���cE]��&'�򰰎���@}K��KP�D�g.��b�oS�vO�����Q+��JA.2G��Tn��{fia�#}=-�'b.�i^�ed����8���y'�&W�B_�}�6�Z�}��A�p�[);��xī���Y�b��-����k-B���m��Ad�g*.�?�4򖹠Ѡ��#���\��`���r�p�8�<��G�A�G��y���RX���`�*>0��w�jI���O��|7!�a����/]_���h�^ ���������s���-4�  +Σ	�sy�<ZV�B�Kk�#�F+��eQ�:�R��%D���~Z
W	�AW�����A�13'Z�ὃ��?�x}TaTAB}3�X�fNr�~�����v�\}��E�e/����g�8$2��f���H��oo7ȃ��Aj�ņ;Di�!��Ф�y優��xu}	$l�ov�c�(���u�f�܈�u��5��-��I�,_��En�������V��q����jId�j
���|�C��4�Ǥ�K<�Vz(<�!o�0(�E�}3���F�5�Hz�luoF�e�.�cܙ�z+�z�~я#�9� ���3����ܧ�1���^W��>�	������f�}�XRܘ��Av���x|f%�S��$V�Z�q)�L7�n%�ZAɪ|�W�L�����R����2<�r���/�	�f��jE��m����4��;^�V�l޴N�����D��@�I+-Nʭ����m�/�%���%B$9�0 �Y�.�ɖ�UP�G�/���PF��!�uW$v⑆'M;�~��oY��	Xd�x.l��ࡪLs�&#�b��6��%���l
4-l�K[
�6U0���Oi�sf��sx�8�9�B�Ґu��H��;��;t�:nL�>�/�;�W�1�����S��v�V��m
�r�]��/k�Q<}3Z*�����R3��hJ���p7��X$@�̬\\7u���>���p=*�m��������^�j�HK˩���5��MLH݋\���NG�^;��#�A��,��M'��R�w��d��6h4p�iQ=n�s�0��J#c�%<|��Ҋ~HQ�	�FG���.c�fA@��+�����ɩYQ��Kb��4�DX$ӳ�-4���v��4J�;�S۴ϋ�S�{]�kǋ�c� �Y�_mf����.�{�ŗXԺ�i��tg�"HU���L���i3��x��_��6��X2تY�=z���B�v,�ՆY$r��Sِ?��->F�l}1fO#^Б�E���tQ��r�w�Yh 5"�"s_�?�}r���`XIF�Ů��(�w�����j0����1waOT�}���뜄i\i��5�H��w���������#3�?lw�����`0��"{D��ąJ�W�8�}?�ӥ�ϣ�Ț��՝p��Zk
�����qfa �ĽџЦ��b^"�ٜoc��e��V����k�=u��z,���Sݜ���?߅HXC����1��Ar����f^n�(!DQ+���ѿ�ql��P����K��X�E?�.X��`��D0RE}�G}�9�sd�Ѥ	h�a1)N��@I��HὉ��I~DȠс(��g1�^���*,ծxY�lB�[j�V�ϓ�X'��>��-����T�0z��K����?�*k~Y^���#������+c{E����Q~���g��V<�~��ZI�fA�t~����ߘ~\	Kp��"$��ɬ�D�v&q3@u~�=�~mpȆ]8�Ө���IQ�m9�8�(E���_�^|�i�p9h����͢ΕY��<:u�:k�BM?�Vu@�'��3����L'��g?E�(�ʚ�5X�nr��<�����E:"b9��aZ���\%`����v�F̒*[��V�0�v��,$Z$�l9��y��,pi?��} K�� <5Zq�8<��3�HW&h25�f�M���$�D�d�_��r1���)��q�e�h�ʽ2���JѓS/�H�e��:QS�w�[�H�_{���������`��7pm��-;��>�q�X�v��+�Y�D�Γ\t�������&զ�Y�G��M��W�����/s�AҒۢ�r�+���i2p̳88���}�[�Ѧ�b�b�o�և��2���2���]���n j~�����r>�ܯ�mT�]Dx���4���\?�����/��ؼ�X���ů��	|7�q�'?L���֕�<���%	����^�8�}$5a�y]�-d�(&��	(��h��Ux]�2)X��O�:�d�g����3�^�l�e����1�ب6���`J��;ˏ|�4����֋�;�_4��y$�a�T�q�en
��^|nV���� �Tť�6o�#�n����⸂6[8g������߹ǥ(��P�58�U��$K��M%��+��$���3.�>�iuL����aWT`��A�Ƈ"_m�<F�r�DՇ��n��!c>!���s�qOC6� �7)��a�K�=(��#SR-ġ׎@�d�ۀ��|�J�8�㉑��M�7��C�?�B���� ��lH}_idE*�E٦W�	[�'R�+��tb!M�چdu����A�=t�*�i�:��x������b3��>pƤ��tN���m'#�l��Ē�_��b��^H�%�A����e��-�cQ��w�̝P����]��$,���]�α�v&��i0��?�V����j�5S��KW0Q��9�:��a�M���&yݸ�\՚����H��Ra�O�2�G�=y!�'�M�E��:r�]Üz\��/�Ow7�z��)�$�Xp�,�,���O�V�n�6 *;#��h�j>��S^k�|����Ğ�w-�tx������#Ӈ���L'񽉗�U^��CwD	F�����M��-�m5�o2l�_|q��5�F�U�ޙ���V�Maa�Np��D��LZx����jIr��!����5��J�����w<��V�'�If!k�BBA��P������j�@��1<���Ԋ�Yp�[��Q��ϕ��}��dLP�*�V���?��9f%Z�8�'ױ���\wjQ��r>H�xڑXb�ld�<�>2�	��@h�%kt�ʟB'��<��u�g����w�#��sR��>d!!�EʂCNŲ�7�ޓ ����`� ���w\���ٽ�Ys��i��CJ/L�Q9tF��=�}a+��X	��=l���4\���c�.�����b�ǽ.��ܢ)#o�C@�i��@-M��ȶ��&�P�_P������E���ۖ�Zey��N�Cxi�@L�x��ˢɜmsptL�Bkf����S�trV���E������!�����(� 7[:�T|���pvc�ù��\�#䇷�]h��7��Aߢ��?�~�ӵ���9K ��K"R(���:���E�.�<`�e	�ܳ�C���]����i�1[S��FL��aZS�" ������ce�:P��Cr��	ڻ_=��P���y���4�ו���p2D.�+.8�����d:�4�=��k#���ᠺ�z� gϵ��+����Rz���l^���(��65��dw���:����}��:K/�-H멤�\�����i���<#��q�>nq��n�d��U}y�S�ReC,2���j��+^��������~�3j�v�� ��?��fq�G�ߟ�B0���g ,Yc@�]�$�L,~��R��[�c(�f��p�"�����1*9r��
����xZ�Ϧ�6(�}Y/&D�aw��/[��D���ѓ$�	,��n�$��[Ɂs�L?eh��^�t�w���II�Aҿ%s��g�zd7S�����ݵ!���K���+��l��d`v�eB�R���w� W0.��<���߹��P�JK%pW*�'��Z�J�6G�Yx��J����϶R�hgd�X�/f���X�@y��YB���q�s"s�.0��ȓh%#ps���k�����$�\�w7@�h��M���)Ũ�h�XQOя�t15ܡ�
��9�l��5�����8��|IyY�P�P_]-�P���p{�h�L32�ƃ͛���΍�Q�uե�Չ�8]�ū�,�?�"���4��+��[�X�i����.��Hڧ�5�ԙ���jt�3�-	Ǎ�/���t�ߒx_��:���
���m�~�K}RG�w��9 �����<(jw��Z��[vhr�Z��j�ip�D�yr�|]�0Y�{�E��6%yl��n����5��D
IIh ��%���͐.(&��~�|+��V7gZ <P@8�y��e����ڞ�r_���Z���jO��왋f�ه�H�#"�(����Q1v��a"uHǎ�wx�|�����^a�95�삶���e������|.o}pa:X�`��,g]�V�@��6U�G�xn3��]�W��!����ȋxV��E��e�r���g^�����K�[�Qan���:�qJ|���
�P��B
p�,�I/���D|Һ��)�8 q����>Ǚ����sg��n��d�Rvn�e���Jwќ��k����@T0��;51#��Ӑ7� ��4���*������i���ɂ\{���8D(�q�tGh���G�;|���k�Y���f+Q�J�0g��zg�V�⯻�̍0,�k�g�Ӷ�Γ��x��/�=�����
c���Ħ/pn`5�F���3V`� B��w,�AV��<�^�f�GM4<�F�b�|�8�V{6[�]��7���fz�~R����<�K����,m���a~�ǜ6�H��>c�ip�9�૯Ĳl���~
�KBt����Z4Kwl�Q��23"פ����FAl %��Qb�p��/G���[�o���.��0�����|�+�d瑪_Q"Z1]bT�)��6w6����9�cG���,)'O��� B�`{� �.ZU�2����b�Q-">zȶoM���M�7������vz�4#˄����\�gJ��1��r�x��!4ipT>t�L��m&��,������#����K9���X�S)�9g�ǦV��2��HFR��iG�^�j��/���|�?d���)Ϯ�x�<N�a���ƚ��c)��<~;��j�|ď.}4�������t�E%���ҍQZ@�H��b�������KCf�0U��D(,k����f�i�����!�2W)���t{����L�p�ӏ���r$6Wa%�G�B�g�L�n��'X]�)T�b�5��(��'k��������R)��ח'��,�W4Z�m��c�7�Z�~Q#�L�Ox5����k��5��_��{w�1"�` ��ۛ!HYMĂe��=)D�]G��EՄ���o)���F6?�#r��])�t�t��������q$R�@�c�e��ɝL����R���@QG�~d�ʹ<x,r??@ߦ��C���ua_8�q|EdYG�@�nG������u�_�cv���b�cR�P���U3ky�#�ɕO�)�(��~��NHn�0��ѫF%B��N:rK�8*��:WEBhU���*I$��S��!���%��\�=K�/n��|�����I	 ��!$��o���:��1߼�Y"�oh@�Ԝ�d�AnJ�'�?�������c��*>z��+��k���iv�h�� 8��=��r1���_�d�	��Ϳc|MM#��O�[b��t!{E�:[]�@m	E2B$��%'��3!Ğ|�������JHm�^�`���3����Z��1������6��@
� C��~��t����.K�/C��$�S'���]Fa�X���5B���
� ���/�jPƖ�6�����:���NGI��*n���A�©k���*2��;�}f&�5n7��N�2������B栃������"o0�~�n�UJ}t��W��������|�J��ҖxY���_,��0-\������ae��0�Z��rJ����ο�x����y$�1u5��o���F���av'��3��U���t���^L��dLU�  ���� ٭��z'��t
�m����`�h��D�V��Q0���q��}�C�j�s�Z��_��7�q$	0U,�K��7�VN�q��߇<g$n_W�N��R��7�Vy���K7�w1��R���Yҍ]A�y�H
�+�sʗ�Iކ���/)�b�_2Ϩw�&����|�^ ����ZN�#�P]����:�Hz/V�ʙʡ�t4�Zm7�����	�/i= ���$�y�M����7���Y���饾��g�ɽ ��):��]�������h��u�#�G���)A4i,b3Á�A|<˶>� ����+`�.�����G�4�qy�� �{��}�g`��Dj:��1�C����fâ�¬��<͔ʇܝ��"������y7����&�+_�Ht��`<Jm�̩�e1��g��%^�#�to���I�柱IdiT0'ѳX���E�LkM&(����O�y��(��+ G=��V�8R1�N�K�Ǟ-�x ��]��
ۈlK�e�e�fB@EeP��v:H2u7���A�˙��]���?�YC���k�|�F�ѝR���8���؜ �\�2u�Ѫ���8�@'����:@��M|R�}���N� 6h��a>΍��JT��;���ag�D3}6��������|v8q����T�l]�Z�BUf��];e��m��/-�3�,���P��}�G3j�5q'P���\N���*�2�B�r8.ݹ���6�&m���~��Q �mي.,oS���M7�a��?hڕx�V�]Y�#9H�;R�����?���w6����\I�#�<^�¦�7~-(��k7��1S��g�)Ew��x�W�$
5�jll�h��N1 ���]�p$��m�5S����s,ޯ���5�3�DP(=���S[��������]�ʶ��=0��7=��A߯�G��uN�Uă�ى)���%�)uTe�� �1/g��rR9"lS�cU3�:�W��׮�^�� ��@��|<?�:�G� ��J�Kl��sw�������\& syn�^�~Y�T�w��}6Xe ��;�_��X�}b��H��.�)���eL<?� ��
gIz�˖�u�'�Q������V{Tןm:/�T�V-%vF\��1�/ʣ�F4���|�k��r`!/���K��ա_��⠪��2�F|�)N��t�i\ ���AULҐ"\S�t�C�Ͼ�;Ɵç�0�����ظ��]���~����t. ��֬۬9��>MF�QR�|�iG�����Ic���m.k�;�ӕ�4�{[����^����'�SH��^����J��>¢C18$�}]�`�G�"���Vj��>��<�G0Nh�����"�s.�#�P�b��I��эw]�o��&_��(u�Ro�Ո�d\<�����м���*�R�?մ�������^0NdedpT�3���+<!��'�I�xߺq��������+����r����}�&��&��aM�R��ױ�����/�ȩ�6.�OF��b^�EցUƤ�m�e:rcgU�~���]�Qe���"/�y*'ˠ�(o�_�I���Ү��r���f�]T���=�܉*N<.�n�4�.q�I�����W�a}��������G����)����~P�VM�VrO�n�1�`�4�r�9�g�����+
Sԙ�%O#���a���C�^���AϘ/�fp,����L��Lud�'�d�eq��2m�:����Z�H��t��8�A�h[�fcF(���[y�����Ѕ��#ڝ��A��B�a����!��*YV���4;���M|Q+�R3 ��:�p���_GIԶ5��~ȧ���,�ۉ�����_�h���QL�֨jm���«v��D�����vm*<�:j�O5�1�87]yV�n�zG�vHP�zҘ�V&X*}/�i�y�������h-#@�C�zC�O�����c���xpVoy0Q`o&w[�c���]@�T(%{,@\%:���|t9@�ܾ�S�I�Q)=d�6+@m���� B|�� kL/�y� �֛�Blʦ`�\At��G�Uy����dNY$��j
�0���)}�B����A�k�[>���e�j�U'�bO�ibx�����A���~�. ����;̌���FSޕH�{ƺTII;#�(W"��gTD��׽ym>@��:'�g�����׶#�3ػO����F��F6m�c�}��5.� ����nD�|��K�	d�	��1�TK�� �& A�ݹ��1��X�diW�
{N.��I�~`�<���"5:�K=�Ž�yz�3����E��)�-����|3浥��S�u��/��~7N��\1U�[����~{s��5�T��'���&�m�qM
�2�
ע	[��t
���r��������������4N�{�8e��h'��`p�AN�y��QO&���J���FX�C���#un��7Je4>�|�6Sd��9�1f�LW^��6��UE��^g��N쓚Rn�X�N6)icʃ��<�����rU[�퓣mib�ą$Љd���\l����nM\�����9�h�8W�4�ci���h&�c��r�r
`���ve���W�2'<�Q�Rn5o�D={(�DJ�ҿA�7Ξ�|)Hg�,�~w@�fy#g�JŊg]���R;��EI7.���#W[�z�x��^�.� ���I?DBi�2W"K]j�P�߈!��u�w�N��恭E���VĞ���V>=
I��ac<�o�R����O���7�rd��f��0���Ɖ�$�x��U*����$0'�}ݛ>�.#��!������)#ٞO�ҡ6DG��p��g��3�(ߦ�*����q���4��'i+~(��������"ܐĹ�_��8�*#�LG�MP�Fs��7㹉Cc��`b�©�I��B����ev��"2�[q.���e��T-ڲ�e�I}{���9M�$��*��*�X��rC��,y)����~_��K�DᤞeE��'
��P_�_����F"c��}�{�����)�A�������4��1˯�A�N�<����~�+'u�($�S �'`��
�"��u�&�a���y�!�3U�C���:uj_ �仇�eX:�l:��G�����Hpk���)�-���N�{S{ɧ�w�j"I���MWy~�k��Ȓ�ϔ����%�|�d�-�x���L#���X ~��C��g�$[�^��)K����]�4j�Y<�5��c�wo������o0��I�ۼ�I*BQ\G4ȇo�S(%���}��E~Q��93��y	$N�]@�.����|�]T���H��:��3��t J��)C:�a�@k����X�	�7�Z`��S(��k��Q�<�G��d����
�tZ߱�jy��#%S���qR��O����זe!,��
�.Ś��&����Ĭ� K�1�ܵ'y��:W)�/щ*�~#����v[S�+^�C���m�Z�����	���-k��d�3>
 -�S6é l$�ْ�*sw�� d�V����	��Ʌή=X�����1��Ka�E/ȶ̚�N�~�K�s��v/�Uw#��n�k��d��})(�����Dn��"��z%�
؋~0�c�#�+5"�����&�\1Y�wb�,5��"���3��I�x��F�i�0��^��LC���X����@��o���Yk��W�;NE����󚖦n3b�@��]u�M����i'�?l᎞�r7i?Q?���	�B=���_���f�i*���R�jB06N�/�\��Lk�'"��I�1�~ <�T�t%WE�-nP�$��>8�2L���	D�R��TR�.$�V� ��7��ڙ'����~~$�z8B��i�k�e��3^[�����)'m�٦g����J�k�x��j0���k{Q��ގ� <�J��B����/$M:��(w�ou1�������y[��A�ũl�s����2�
�ƶ�ϥ�_��p������&l͈��a��!:JS~zB6-�(tK��9���6_k�蕁�"+��)v�KwhﳮJ��������+�W���r���tF����m#��X���I^��$ۻ��-
�E�H{ٶ�o�0X�Һ���{��
����C�G��v�e��P8]���`�K4�$l'-v0vCh/�_w~;8����7#U������Pod����=�
��?�71�Y�y�wﵛ6����k;҄>
�:vp���6���r& �ɞ09f	8��y<��G��7ZL0��+?뤿�áYM�'8�H���i�qs���K"�K"�1��6ʴ�G"� 0P�oG��T>!ƉC�����/^C=݊�'�HJD�X��H�4�;�����#����
?��'�-��o�^u��*;^�<
��ׄOj9Y����!�4�y����o���Q�lm��xJg����u���BJ�L���LW��,�[��7f-!^>˖_ە�O���@`E�o�9� H���B��S���R�B�耵��x|�����"����]�	���-]�(��b�G��0�"��%O���:-���*n���9�2���W0�_���mB�E��mU�������,��݇����c�BƮ$t2��cޱ���(E��cM�q���\��e�3���L3��g�X���&Hf�� -�KN�;� VytF<��b�Ft�	*���������8EaJo]��\^zYj@%K���=�7�j��^��[v������ЌF[֡�:����"�U�`Y*Z.�F��7l�tD���������$���V�P�#�
����Щ����%�LҶ�;���{�XX���g�507�f)�����}���H�x��.9��o"�z�Z��NNϽ(	o	�	�V4�t�M�3m��Q��wܻR�+��H4�GIˠq~ζ�+��ԉoa��8��o�����sєb��Gt���,\��\_�h!���7cKG�Q�h�=Q�&b�ۚ��L@	���Q�,��@>͑Ƨ�0ex�Z7þ7��(��P$�Ѡ�|�#ru�� �H���됣����UZ�3Lc�����]��,��z�g������i�k{M��igs.�Y�:$J�t��+ث a�����o�����Eϼ����So������1s��I;`d�c�⊟sj�V��q���j�O��f6U�b���".�m��1�i�`���9J�H�(\��!��;�A4'9�s ��kh���rT����!Q+�E�͔H��@9�bW}U�.�B�T�`,���|���]`��6y�Epl]T�[����h�~��aP,�Ux�!��e�ÀR, ���2w�|�ȇ���s�v��>৺n�X����1�\O��q ��ڕr��B1/���U3����5��N����4Q0�l'�sN��+Bk�ʬRۊ��T<������"��M*��.�]�nh�Q��wo�(�m��V���*�E삏���TyȭM8)����T����Ih$ZIu��F��4W�
�dg��g;rC�&^o�;��m�3��wn%s�A͢
l�^1p��C����2R����,��7[�c���d"Zx�%d��<��m�O�<VT2HC��\�i_+���y��3���o����s��a�d�_�,r��2�����W���w8�f^-��k#z9��d�zO �V�kZTD���=��kH�+�"!��p ��bN�Hb(������u����;���h�6�t�Z��Í:Ω�
ɘ����7����bR������M�]�;���G�"�=o��V��q�&�����[߽����(�<'�r;"U���a�\po�g�g��oA�m��R4�o�������s�y��Xg��+�{��(?�9-��,O)%B
����b���lBP��!��� ̔�z��T�k�H�a���:�7J�B��;��ASe7�p�c�8D�O�Ser��&�CHY�㊠w��^�wu3��R�G�̀�Q�k`=u���5~N���?�~�-2���O��9��4��Q6�Q��k�9]4&�D-ph}8푿8�[:ф�m��e	V�}_:l+�!a��\�p�!�X�t�Z�b-6��R�#>I�Y�ݗ0|�|�cI�D�FQ[�e'��zd�YE����׏�Y'v�體44�v��H
��Z���T�z���c&副Ƶ�Kfv]M�۴��4�F�cW�@\l76�m�(����m�7g���%�n�a+8k��^��]h�]�Swͱ���K*��6!������0h
�HQ�6}�-͜�^=�)�n�>�(֟�������f����/�f���Z�,�:���y���k�;G^�t)}t4�ůT�l2�I:ll�zF;��B�c�f����w�3Yy)��R|��+�[Dh$��.h9w��"zEM�'|�WF]CPe��Lw�@I)�j�.)\��T�?@�$;�H
g���f����Z����'$t2����w��������8�
�Կ�8����4�<:6MOB���h�G�Ho1_��bKc.�w�8Ap��*�)r���!�bl;��,ҵɘ��n�yV�^�%
�u��!�|x��]Y���3��^i=�!��Ax��𦴔n�!c(W!뮕�m�h43\�><
��^�	��k��ˤ��ɵ:���7"�A�Y����P"J_�Oyx1k3R�64��� �����蠺)��H�'I�� dZΘ�LiDMv�����0T�%A�'_-��2��x��6niz���7�nEN���z��zC�T-3�oփjO�p�����N�T�	9��=)U<�?�	`�&���3�r�@�פj��֊��$�2��B
D~h�v�8��ަS��N�k�ᾳHܿd4bP�`���~��	v4�Q��L�<-�S=��8���5�#S�'�=�QC��]�_�o$%�v���ӓÖ���w��Kig`?[�&��qA!On6�}%��R��G��Ű}wX��]�7�=���������Y�E��G��:��Qi%�0�k)��{\�W�rh�L��9� �~�f�]�/;���Y���n"U7�.C^��;�*�"�!�z����8LZ�R����C8
Wsڔ���	�>�x��a���y����az�Io�%��Iӗ\yXxI��|ƮW����%9�./乢9lfT(U(�cu� ���u��_�U�G��Ud�2L�}I0\�*+P��mh6z�m�9��-]Z�I�@��Ƒw	$3�-�o�Ȗn0�n����`M��^9��6�!	5����������1�R8��:��zZt�.s��p��~�_V2�Kh�z���Y8�"�6��>t=��(�M:�5Fp"�OS�{�(�9:@IB�Жz�]�>�w
�u��P�N�����R��5�+�o��ч���ӂP�}`z}sR����ܼw���i��iˇO|��b	x�]It���B�Nx0���.E3[��ڡc��_���2'�塏^*a�a"k�,�' `���ϥ��o}�n	:�#�7�+Q ��g5-��]yG@.$�P��ځ���_}�*�+����q}�NY���+U�ҵ�����@�B�d:�t�4;�LhXa\�(9�.���x��[?�s�@ks���ς�H�S��H ����透<�9�����X���P�Zʪ<���9��"���`"�'�=h�g<��.�2"@6噖!��Ö��=8^[oP4`�/n��q[�����L2���%�7&IEO�6)7�=�t6��S�!�n��7���=��2��%W�kԜ~��'(ל�pWqF�=ؔ����_��	� �2=�ܔo?�jH���i{_d�nI�YaQ��j>�s�\A��2�U�Q���<������4>:�Eժ��V0��Z��[F��J�..ZքD��=�u��%)�=��Ut��N���S�ܛ9���ӳ�_ʖeA$�������w4�(�g2�DICt��bA�e�5;(����vh�u�!��R�-/�i�09�I��_p��ND����N��f�X��|��X�}a2�O54jV-@q���8��B�n+�fDj���~N�뀣f8�K���^Rt_f�L}>��po��{��xt��)�2#&i����D�N��#D�h����u�I�߰��s��Q��#�Ka�\Q��@�v����ns��Y���ǝ�2�v�ZjTPi�S��y��i�[eZ�1�1s���Ɖ*ھ������������?�iVR�P�Dݗm��a��Llٹ�@�䆏�e^�����5�#,>��:�Ԟ-�^))滕�b�~*+n�?�熋ssm����+^&O/��6f�%��@ VE9E��9�T���'��s���`LA����\s��3Bēu�)U�b�[E�	�O Bq7��/�F\���@3����Q̦?dH�ڵ\�n�F�_),~���/���."���l�5��-@�(��àF��NM��?c�t�`nR�!B��6��fx��xҟ?`����S||P���������ʽ�N�γZ簣F׋é�d�A*ߙ3��miS��Y4�Fpqb￧���my�&B �f����U.��+��&x�q��rp}xu�;�l�A��Gm[�7��+���:��T-�iׅ��d�7-�x���k3�}�}�q�'��0�9���c4%s��e�ikR��Q3����;�4���r��`>X2E��wve	{��M�A���Q(�hI��<q7F���Ver�A��){9 B<g��f��{�&�,�'z�v�t� <�w斺��K�@:�7F�� ���OéU�T�0�̣O�f���*#��l�=1M|�����:��ӫW�� �ɐ6�?�$Q	Q�	���8�F�o�I��n�b�dC
ݓ+QN��h@"�f���r�q������iʐ�3�N��&�J�JV�0{��9*�*�+���ܡu�)�aE<Q����~����f́ 
XFkP�Ȍ>�n�_�H��� ������
;�*���J����!ȥ2�gK���/��-$�K��0r�3V�f���ѕ�A%53�:k���0����B�n�Ʋ�ve�a#�:�c��Uu�D�`XE��9ar�Vxi��f��d�ANˍw��o�����cB�$N��� ��B�}�$����7~�N��ր(=��.�kB��a�&Ά���H�10tF�jb���B&�	��9+{�4{�������.Pvq� ���gC�&3���~3�$TQf	Tm�>?,�ť�<B5o�t���2	qJD�b�����+nJBȐS���UH�`6w�\�E�[;�d]?�q�n݊���|�~�e���8��Tà�G���4�����e���S���\���i�E6�O�c���KX������_�*0�GB�� ��@`��]_; 7�^���&�3�8��]���0,ͭg�S�:`�d�|Rt!�,qB�8�ìO��#3Ρ5'�t��1����lE
�ڃn��8��h> I��AZ<�ձW[�+R!8�!�p��IQ�����)<c���
{��z�́M����iG�1�I=!��La�g�8EmqL�G�y jt2�瀨�;,"�4zg{�|=�8�l��pZa�r7v^��RCv��#��+t�QMnҽ������	�E��FT�z���?��B��@���9R�6�]�-�߆��O����h��}��-ź��{-e;v>��yq����|ח������Z�T�_O�و&�ND�ᶩ�"���p�пd���u�Z@5�iH��F����2��3C>�j4��p���ݧ��v���;��9�[�۸y6�'��y�����o��f�K�ޱ��ӌ
�� �/�#��7����#��*��࿲P�V�s���ʌ�%_u�<]E�OM��s5��oO��,2^���G���
��ZIN�Cb�����54# �k=�:R�\������������R�9�,Uݞ�pW�rF~Q���O>�({�̿-J#�6ϓ������]/�������y�t�ς�9�,|ץk�J��?x��F@����ɖ���`5�ڦ>��jDH�>�4���Ai�Ձ�ݳO��$�ٓYB� .�� <��ސ>x��f����c�LR�S淌�Q�:eqVʽ�N�Rq�am.� �����i*;^���	�3�6�8IHwx��5���Kp.y�}h$�֨�og�V�D�7� [e3TSz�㸓��zm>�MUl"���ኰqR�Q�D��h�����m�]���A��[�z�1������l}>�6x�{$:ɍ�u�޸�t��gh�d\���Fc���t��PZ�� ��dĒ�@P� �ZϻU⵩]�����ϕ*��d�$Ӭ������㷣�d	� f (*�I����>6?/z�qA�e�:�2����~O��֠����05a���������DLVL�}��pa���q�j9��i�/��ٍw3�V�P1y*}Q^��o·�݈���i!P�[n5���G5j��͘��A>�0�ط\g��ug�+OQ@m�ÜB,w�!������<fh돰+\#�p��$���h��Q��y�ʹ���ktK����Q��d�*M,"�n)U���P��K�^CŘ�Z{�A��i�����S�j�f��jU�D�k[�k����Wc�:^�a�囦�	�� R��4�Sb!�/�[�Ѧ�?o�~?4�#
�%�LƃF�	�ʑ��#��Á(U��ўe��^�J�{ yY�E�B-�ٟ��3�!�c��?V�-�njy��A�1���n53 �r���d��<�t+(�G�l��F��H�%�lh�|�����iQ�:�p1a��ߣ�����c�·��W�dItK
�r(yӓzۏ�j�,��v~���)����7�F<�ガ���@�Ѓ�u aQ�Z@�Z���\ ��|1��)0��=���r�0�Ź�3����RS��Y��p��8y2��W��@])���;ǁ�X��%&�v�7��*<������(�}���Ʊ[��s��hh�� ���~�,=T��y����:B�#�?02�]��RJ�t������CՅ#��Tq?b>����8��]~~��I�y�&Y<_�˨�O�� �xw�pb�V+�;!�3����
B�L��F�.d ���qg�%��^�$�*e�}�NZTF>�=�w*��JE1_+SC���G��L3B* ��IPn��o�\.��$i�т��us~�rAeR;�U��޶�$؍��=j$�
�M�7v������:����烺��|�&��j��7�&oT�S@U=�1��c���s0@$ǜ�����a�������P���*�_��*Z=m�G�i���	���&���o�1���
T�f��	���[H:�ږ���u�.<TVӣ1�~����[�v?��=h-|X
���Ze`%#z	�@a������D�;I�\�^$W�J�WW�8�ߋ���.���4L5E@ƺ�g�R�C�����ɽ��8b� {�m�����ת�/�Lk�fi�tK�zT�R�D�)թ�ycߧ�Jݫ��=[�@�C�8hWTqn� U���� A0ڰa������v��-�ޞ2҉9��4D�������h�X`�	�6��O�l*�`@}q%�v�]NS��b/1�{��>��}�LRH�P��eKߴ��X���۶.&�SZ��P&�!A�9�e�_��L����_��,��p��X��}FG=��:�t��*��Ԏ��`X>�p%�s�3#(�)Hg��+�E=E�'+��'2��zw�ϼ���I��s�N9JC��	z\�%����U�PN�
��d���Q~���4>"�+��V?$E�f"B������}*���IqD��?�odt/8�b�0#�"�?h�8������V�cW��<��;+o��
+���H���ҫ�g���?�y�<�]��=�D��i"f'�K���7\�O��d�V|�X
�!�J�S6�2�Vw�vBQ;�a��~E֚�?]�W�N��!�<�����׾E����!wq+\�!U�
2Vwk�1MQ|?�Ĉ�.�l�HOn�K�#�����;�yQM�`|�A<4=!�A3�ïv�&�p֐qn�/Z��,��V�������w�ا�<��^��};�*vx챋��R{%0��χy-b�n�� ���s�2}ι��#�_���\�O��5�Uw����f����s�B[��Q��DE3&�����T֒"����D�Bm_��d�Dh3��j��&����5�o�Gq���"�m���(3��'�{��$7Z�����Z�Ñf6�Ȼ5��XLl���A�t�Bk�C�����B|R�G[ A���&=z|��nՙ[L���v�1�6�����	�\� Փ:5��`%�Ț:�*����_*�h��]��6	���w#}u���3A��!#�bX�]u�M�a������Zםi[i��yK�[C3�[pG��z���1fqЄ"N��GT�7��^�$aX#A�]��Z��됌ȱU0���mas�~�i���h���х�����-u��T�So��*����1�F�[r|`%�4%;�U�z���g���v|]�~T���¸$��a�/ܛ�YU�R�@�z�1� %s"����{��a�m'BU�ac�97�y3on�9��th�]#�_�ٹ�����1�4
|G�J�`-�!Gk�T�>�� ��0��K	@�_��?���jK��W�ǽc���z��U�۴�&U�О��|5S)0`��.'����r����ޓ��sDrE�y��ꭐʀGcv:�Tj��t�VZje�]�r���au����4�����;�6�eD��,�ԡt��J�p�M��*�p=��%\��g�/L��t�^��|�א�^��"-��y�|J%ۄ;��[Z��������Q	�7,]�B*86Q�!�S�W����p+^49^��<ۀ�߭2�w�J�kc����+�n�I��%.�e3"bUX&�*B[lP���8����=[U��:Bo���]���C��m��;xy�J�w\`�j���5٢rs�{�C8��!_-'�/�}���^=!��?n���gY22/%��-Rb�ڥ8R��UT��̲��5��O;T�?>i�oo~�{u�^�x�������Ut@��e��i��%{���ɾ:CZt}j�p:ͣ�NU�O]]��s�Q_a��ѹ��JV���Ak����00���M"l�.":[b��,-�mcՋ���U+a��)���h�z���$z)PO��4��|[P�[�P>��:�ެ[2tGu<����P�j:"�I.��6g	�Y0n�/̞Iv�}L�4��brK��;/Pl�ޢcZ1[f~�"������(��x����d�V�N�'NN���>k3��攞�U��K1�56���6�����'zD�n+=����X��D���/�v�E���$�EQ�� *��3=��7-�nͶȶ3>���o(��.G ��|f�W��P��纄��]��%��8b��m�cS|�3�y�8V	���8�c���M�"n�|t����f�a�BT� -A�����������Q����f��?���E��� -��pe&�u�\���4�1u���q@kԛ�tŎ�K2$��������c���jy�o�Ki���z�m��/F�Y.�յr���B�_�F��j1�1��C��=P��Ǭ	�KB�u�iuo��J�X3��vs�W	b&�:�4ӏ_u�!�$��4��s�=�~��)*F�j&�-?y��d>���T�T�ۄ�{��Gm�;��`Co�<6�'�3�Oq_�G�-�e�f�ߔB%����%���'��MD���z8����e�0��;���0��hD*I���P��|���o5S�\�����V��ۥ�ʙp����_6�Ra�ap14��ty`�%�_�Q��ei����'�SC�?'�}K�W�h!3�0^�+Ầ��s��X��b�t��yߣX�ښ�ױ7t��:8KI$[��9�����Bc�R��F���r彞G����ѕ��~�qy�X�4�f!�Q]��ܦ�K�ۯ���>�H(D�����劔1�&�t��no�	�W�7��B�k.� �����w/�tF�W�=]3��n`h���#༣�%y0���� �ke�CZ��( ���u����G�ж`,-H�������STym��U2�?��]�W(L(�ϮW��U��S?��S�a����5Ez��؏���+<B����
u���4�<X�vk��,w�n�Q,	��dژy���N��מ�wFߝ4��}p(n$(ӒFZ���I|�Q]��E���aDuEr�E��ؕ��M�N�P9H-�Ӷ���"!o}�� ���!��@�3��%6� ZۆQ$��y3�є�s�ڨ}���c�i"��E&,���P������ ��n匂��]�7��ZSFo�5z��r-��L+ɘ�;��;(U��iY(au���@r���˘�bLI##�k���i7�T-���,ͤ������������E�9�u��^�JVN�C'|�ڋr~��*Z�z:'n=k(k0=@t�v�B��[^/-ƁP���b�/�A��g��)�f����g�U�$5_�вW��>��ݦ���Z��0H����rњ���MY�o%n�b� Y�'a�e��u����5<���M* ��o ���f����!��K�`r�@nq9T��
᥅�
�Y�O���揾m�a*��m����d8��i_j�~��퓚"���@�R������m��*�5���ն����$��578W�E1�Ά�qB��w�.PN0���}̈́��43�%Ț��3�g���_�DN�����[�3Q�E5��k�0j|}I�H��T`�A[���-3�\�߅!���o���<u��Ll�T��[&|ui�~��ly6*Ɍ-/�vά��X��k�־ ���%f�&����ŒƵܑ�>ʸڐ�7vR��(6�����uE�VL�҉���9�S�I������=b}��+�WtczrEj�k��
������A�QW���l�-�{^��=Y�{sY^16�=��	@Z� ߄?�V��)n��'�1Z����ف?�5R�O~��[�`�����@K �m|��lct�n~�Bz���/ۼ��g1 43��V��"��R��_��}{zdU�6�P����#M.��I�6�ǳ�y�[ Vo�&+
lN��7�D����%L4bE�bϼ��Lצ����k��ɶ�)�
dZ=�2+�=GA�y@˳��ul�£��s�����%�u���*��|�+��k
Zp�� }q"UD��$�j"u��%�/�R���,�i���$�a'�P����n$��xZ)��J���6����=����d�)��{`��߾,�o�_��Q���ۢMd�f?Dc�b���m�%�����I���e� �"��#�G`�G۩@�z8.r��
1�>!{"Ͳ�v��ǩ�q�Ƒb��	��{��Y`�L��&��2[��.���7Cq�ߠjP̄�X1�B5�v�KW�$f��Ѽ�3o��?����?��aMu�T�O��� +ſ9��E�c����l��XyU�jn*u[�/��zۑ�ũ|�ž������bo>��KfO9\Җ!���@��{�rݴ�ԃ��QE�cf�G|�vQSP@9����a�l��4^���-�����!@�-O��au{lu)H� uq�Sœ̈�g��
��l7�Q[.W1$<�>��D*�H7*W!�߲�͵m3_�'�y�MV�y��'jY��l��i�zWK
�-j�
�H�	�)������GP��|��U��]�ڻ��{�w���|A��,�Dd��t9+�4gP�滅�w��#�4�q�|���4����+q�nv�Ѭ�!�+�V���9ҟ�5t����W�X�����"�d���pb��� 勡��a�5��a#D *���ćZ4k�T?]�@_7����sܳ�*�9��j]U��n�^�R�:4���_�������V�!9�^P�$�o*�Og1��UsR��LӦTզ Dd�+�%�a�dP�҃t�*|L��́r�Գ�2�/��~�2X�P�ܾ e���V��KB�]Z��^�SeɁ��2�'�'����N2n<1�( �=<J�0�XM�S۪���Ja����ԝ��i�h�-"��ٗ8¬�!ǖAr����J"�`en(z���A�0���/�^���y0�e0$��Յ��N����o�(�~�fj��ݘd��7��gÒ�(��y�1Lh�1�a��*�R��x�q�%+2�S�7������=Oc_]�c0�0�>቎��y!R����H��Q]��w�� �E��A�����6��$���1�|q��ѴF�tޫkPP�P1P���]K}�7y���+G�i1�P���,�d�?8��/Ak���@借�ܝ�P��h��f��x�e�q�UN��t�3ջǠ�^�}^Ej�暃W̓,�c��]޹��_�a��X�S��@�LF�}������EJ�{���~O�U/���=�1l�L��c�#h��vu�.���y�����6χ0'�_���Q+�+2ȪW�|\�:��BA�v���J�5��<�; p�9����X�n���o�i������0nF���	���׋�Ø�\;��8�ڂ���O�
�;0����jE:��r�T������9���Gc����f�4"��g<uYt�]�,�}�-16EՅ_�/L(�0����񪼜��W��C����P!��K�B����R��'z�:l���B����I�xͻ7&i=�t��Glb�4y�T=@�ޣ��`;Zp�W���!X�'�Y������.��	Ǔ(�^�� �4�[�6������;#�\Q�6nQKb]�W�1쀳�7C�y}�u�uS�˟�&׺� Sn�O��g�X:�eԂ�i؃�gN\�I�rʦbS�:�G�}8.(`�����l�H;�����䲢9��bn�aR-!��u����XTa�=N���:�>�?!y�a��~��ݓb�]�ِ�xH����Y�~j��R�ސ髛Z]o��\p��Km7�N���C����z�o�k����8�<R ^�t��}��K*��z�/�L�Tr��h���O(	S�{V��dk��[^�HT�j�t�Gc��<� VG �'.z��ѫGS�t���#�'�P�c��hB6�wK�o ���O|�<#���aw����8��R���H� e�1�{V��
���䴰A��FmH	*�PPi�K�u���x��������o��A�i�]*�	4#��'B
!e��3�TH���=
쏩�^K	;XU/t���Ɔ��^R�ǟ�_���� f"�|��a�`"�� �0��mѰ&s��؈�z� Ù�����C]�1N%]
���r4S���,~�3�����<|�Y�W���&������8�a�O��8ڻ칲�	��y���02��?07�fK��q������ӵa8�����r6� �7-E[8g_$������M���7�/���W����>�ءF[��m��b�`�y@��Zs`�!�<�e�*�>!(k2�?G��C�b����M�-S��6�`n�ږ��iֻv�� �PH#�a��Ԑ���4f�o�nTk��r��]�\k�X�Jw����(������-�����M�p&㝧kҦ!O΂����GvT�	6�v?�|���{BË��<� ��o�/-��G��#��Ε�����Ŕ�����E��%��L8�(;�]HY�[>SЇ�H�S��(\�߭��$<:ib�x ��6���T]����-I�����qGP���-��t�V�^}B�	H��ذK�h�d�]U`������S;���S>)f�Go��-���v��*)~��#��i�	Ҵ׈��WM���oV\,�|���-�����1���Kհ�f�;jF*�l�3ȝ	�ǻ1)��CT֑p�hſ�&�&@��&w��>&Bl�5Ay���@��dإ�"�ԕ*U8,'KKW�z|U�ub��5$���V��� `�wz0��X୮�FGo*���t-6O��R��z�=�Lj>�i� K^����qh�+E��WO�#�xWv8l�󘏑�w|{�nV���|��]!�;S=�CO��=Tn:f�6��	
�$-��~�YD�s9��[�B�]�8�S��Hg������+i#8�|����8g�`��c��"�B���O�a� ���/l���@Ei=�Ѐ����<��� ��T08���\�Ì�ů�°����2�VL YV�_����E[����U�Ăt��uSC�7��vz�X��%�|P֮�v��%Q�K�[���K:E���RbT��/"��	�X�`c"VًxY�6֭ʾ�&W���Q3����i�:�!�� Q��`���gix��_WҋD�����'	��[^G��,�c�T���!Ϲ�Q4�HT��EBY�>��xLD9�4�=)�	x�@�a��]RJ�Z��1�v�c;�m���m�\]�l�C����ʁ��Fo����iEb��]�<�E���y������NO�g��&)DV� 9�ѱ�]5�Ėq�E��K9Ylj��έX�M6y��#Q����#��8 �n�����[L�n`�Uކ�� �0	��Qq���XA���!~��Q�4�F�=|�6kY����,�f�����֊X�%�I�dU2�K�Q��9�xŧ�n��HOP��I��y��E��|L�	BXkT�#t6��fzCA$�fpl�}�C�� �b#zl�(��j�`�6�q#�kI�ga�2�Ql�ګ�k��|�C�yD�MY�|�W(�����3W<c�Ŵd|E ��Db�y$����L�*�2w:���Ȋٍͥ	YbL�[�j���G؍=P�ҡ�:������nLfG�������s����O�Nƞ2@Sw�'�Z�����C�zh�y,9*����3[�_࿶H�I��<�z�k�yк�����qi0�q�G�ZT��`�rZ[���8���1\����O���i�|J����H:<�.��.!fg�6l!X8�9`7B���h� �π5����j>��B���i�7%V�i�9��<4�zsҀ�m�y�ӿ�0j"�	⺈�:y$���^��.�u�]tXK>b*��c{"Ϡ&��i�#��l{�D�]f,�i/�OJ7�^����P�f�e��-Q��d��XJ�K1J��H�����
��ȑ��؟��?������ٓ�o�� �*�vWE�*B�H�-mJ'�(�g��'7�bTo�i��J��}�b�ה����QP�#��0B�J)<��R?{�Gy8��]�Z�f�oiU���@vYǋ5���||�n��K��޻'G��r��{�%*<���c) 8m�|��r�4n&=.�F���S���O�7���0��h�~�|	iw���!ܙ���?is�լd6z��+���0�RVEq�������9�P��N���~�@��+NY�����q��]c��D��d-����|�9�$F�L*e��PT�m�z�4�b.���8|_^�|~��RIJ/�c�G\
�
?I��
��`���(M& �rPa�]&yҟ
A��S�g�Ψ.�N��k��:�j�;=�)�6k����Q�U�F����%$G�a�{��$�kP\J1�cuL�|Ύ���D�E���H��j���͚P��d�2�������?�4��▇,}�nt��^Jw���L�4J�Mu�X�)2�U��u$��HZ��Y���JQ��gړ�`��\6c��t�T�pW&����!d��a�C���G��.&ڎi^��˯dq�6���iZf�}f_�Fם��L0&>�Xy!��{(o�,-dґ+���c�QAn�)������U D�Ga��?NUm�FO����1r\o�����7=2��~�c�\lKs����|�7�+O�� ��;m���	6yn[=/� IS���/�\3���_��]Hz#�ᑊ��)Af�_��d���r%� H��U8��j����ǦHN�K����C�����\]D�a�k�#��`�0�g5!Sr�#����\��1�/q����c���j��+�8Z>��RuJE���Iq`uy�h���AR���f�z�FD�HfC�u��/�gbf���_��:K��n���Y5��kҀ�p;_���5G�c���$�v��r��ni�<q�2��EĶ�YƤb�娷hmAB���xh_+�a���=r۰���
�G�r���u�V��ݭg��䃻������TKv㯞����'�e���G�9�\{���X|
�,�� ����18<KY�����
h�X˵&:��lXީ*�M��f֞��k�Z�!��Bz�Z�1r	[ϭ)y�YCDf!J�����:�nc�U�a���lc���W�~��^R�����e
��6OS��@HC�-7���'UA8�_z��ֲ'�'���;O�7�cc�Ȍ�F�y��U���9nn�IW��8=>��Hb��G��[�1�Ĳ�׭���?���-g`A3T!����NLKо��Φ՞<%Eg�u�oe�K���ƕbB-Ma����s)�n6� LZU@	�CHL�����m)g��y����rY����� O�ŕ݀u.� ѭ���(R.�����M}j�z�)ܼύ�Q����^�Cí��u��+!.�@�l`��ڴ�����P��ڃ��F�)�y��\ÒiH��\{ܨm@���~
�'z q�Ţ�������)�#-e=�5|�`|u|!������,FnVbE���&Y�o��fC܉�B,����C�$E>p}�tt�j��
(�E�1��K_�_i
(	K
ݱT��J$�g�o��������(�ܼ8Y�s?(�g�eξZ�C����g���Z �Y��)n��`&��'S��^t�j���W:�xE���%�إ���_�wW�hs�K(]���6�+�B�ز$A��W(�|������u狴�;u	���D�s�z����X7�rW�]6�脄���?A��]R�o^U�����i�����w�5m�`�4��N��%n`;,Wp�ŏLV�\���2h�{�V�a�G�YО��<�b����S�FoX�;�XT������f�������&ʪ$!	΂J'g"4��E����]�M�
�yX�r\n4�I�%;���F�j���k���eE�!�1%j`uq��@Q�>�(����/[�05��9�<�f��cz�n��;��H�%Ms�~e,�d�Yr�z�w��D����K��K[|AN~��S�����\�L����o�R[�#���Mx��S[�������r�!�A��e�{�q�X)<v�jңF��-
��hJ��^�s�y\J�.�,cι���n��6ۻ�s�sΑF��~FWY��sUR��g\TL��]�V<�?s�F�p���L�?Y�pz�����K��pq�FYN�Rl�6Z5��E�~X�[�����t|/��2wc�V0]�[�n݊+�jH7�B �4~}��w*@ ��9��8hY�\��&�$
GS}79��4�*2��ԆP�/[�~�������DΏþl����H����	z%o�˰,;$;����d��>F&�P��ȉrZ�}៘I��
	����X��Hq�L�E�!'T4�n���Pe�x&���omOX��+�z$3Q�w��CH#�[�골P�s~p8�5�n 2i��zW'��:-��'�w���> ��K~���ܣ�~Pa����[�� ECq�w�X���Bu6ə5 �_�C��F)�^'d�2�ǖ�'3�"�?�,��֖X7�M)���B 2��A�%��j���!��uN;j��`b�%�3 o�Z�[9�牠`�=�2t�,���c��z�..���kǁ�٬�=(*Eޥ�gW���Ő��**���¤%�<ݶ(�t �����e>�TOF�ܣ܄�!�H@/q���cך��gVV`s�^�����в����(�L�,������������v뫠��I*�č�ϸΈTݎʽ,�J��5&#E�y��`*���`n���G������~^E �����_ۘ?�Y�k�n�6y�>ĭ�*mG�#�W�R��4*n6��p[���3�?�
�en�u5w�%�m����4dv��Sbv�`J��>3��bK?���;,�	�վI��Cɔ�A����[�Fo�0\�A��h|KYA ?g$�����,n�V�ٯۑx@��=8 �%h#Y4>o�V��y�����V�\����bw�ﱴ���Y=���A��w�,7U�I1*�O�N[n��U*	R���[GI��O0!$<z�yp�A/�5VY���GP���^J����ߘI;��d�sr���*�C5���X��8��6��4ھ�����ȕJ���������u[u�s�g(Z�
�?G���C����BU�E���I��(qx`��p�#H+n�x�E^ 6��Y+�����f��nr��Gh�#$������R�fh��7�����g]@Rn%%�8lҷv�0�p��YƊ�>���
-��������G�>$��;�a��^�/yt
f]��yb��C���"�P(��4�ʚ�(je��j�W�媐�ſrL�ܸ���k�0Ξg�ۭD���K���0>`JD�o�+3�"�9!�N�V����g�0���i�������	�)*>y�v��?�^�Ϧ�%���h����F���'�8�!f�ꥯ�<�j~ad�W�2��y]�Q��U����Ѡi�0�M�!��5�L���b\�9(|�ˡ*|�w6���R2���ث���C�����ٛ��/�6���~%+��6ξ��Y��;�&I������ө�O��_��A/ɒ����=��ꔖ��:rEm�h��#���ŋ<�0��FĴ���%/��L$C#Vn<Q���۬<�Q��vl*�C �����\��\�Z�f��WbIR9�2�������!�����Y	B���Gfߘe�;�[;����)�ZO'�
[3�>�q.�p}e��PoAVnT�s.��q:����#v��J�?o��!%����������'���龨���;�kE�j�磿�ׅ���~�%��ϲِ�[��G�Y��1��2��a�ͺ��M�&����fx{��9�%V	J�!��~�d��tWm�7^���h��*�
�������R�\<��-D�ŷ��Ld[p�v?�"����+�e�/�Z0g�>�1���U�36D��,+��rr XVV�Zc��s4���i4jQ��_��tZ2�qZ��EtX��%��l�T�H�hJ��V���q:�S[p�M�kџ)�k>)Bf�cG!N5${������q�:�;�-=�-��!�t�@���wwR�6�Ώ٥�:'mU��D�v�-f6+������/�x��R�؅�}��Ei4N�������n�^��m����8÷��EEn�?�
��Q�
�4�]؅��L{�ӌk��-(�%�z@�BX����&�$�q�~�a�suz��vd�מt@5�4zX�~�Ѡg`;7ܥb����'Qej��LP.�5��!�h��ֆe�Ϗ�#:�X�r��e$���U{�`�HV��L��g ���ʹ�J�;rP��[��̦�]����_><>%�C�皫���FY��jVZv��.�E��f�̝�j]��<6�ͽ��,�^��Z���޿Q�L]hɚ�j�x��7�W[���A�#�՟K���D�l��n�T�&��{:�H_�c|�s[�)z�<Q�O���%�+@�BxZ�62wX���������(�B�jjd�L��<{��70����*��Dƙ�m����ؠ�"n��#L���|��'qKX� �kx�Q`�P�� ��t�]X��q�M"�3�t��iH�5��Vφ5��a��Tn~�eW^��=f�,-F�MZ�X/����C�7�ϑ��
s��B�k��,k����{�:&C����W�^��7���}�����c����@�8��XEE:�(]��dJ�m�M�N��M�=��ӿ������8*�Q�A�ʬ�s_h��/�SiP��$�/�e܄��z�=��r��w�i��|�J���c%tr|�ej���hH�N�a֗�i��z�"����,δ:\�e�N�k��&@pͧ܎�������J�p�k��b]����7Z�_G���V�������F�������n}*}�PUf�J�[�Y����!�ga�e��W�y�m^��W"��A�'5{=�W]S���{�X�\d�^�i��_����䵠lF��pV����_��vH�I�z��Q�/}���:Le�E��8�\��VHK�a��_�/@A�O������a���IS�¤�EK7���1���퇑'�s��ϭ�*Ɯ��V ��1�k�v�0���Kʟ�A���zo%Tn�R�Yυ�i�_r(c��\�wЇ�avf�!�R%��V�1ɟ���k2a�LU��҃�ۘwv�6������ɃB��]r�E�ҸNR,��=ݞq(�0��=Z艴���F�m!˺��7ۥK�*T����J`���6��m�#b"O7�ӆ+�ȶ�{E�̧x\P2E����X�H|�"	Ƴ�\J˴�	����%{��c3l�s�rnÖټH~�%�Ɂ�6&��|�!�@���k~��R1g�"X�Aj��m�"�X��e�ۻ
�5��D�-òÍ"���t�GZ��j9_Ȗ�@N���	"ls:!�{�+�����G��
�<�
K~��Lgx q���#���M7�b�f}6l�^�>8�EHb%�������BQ��A��n8{�����x���	_�_���]�ڽ_�0NW�d^
�iѻZ�R�>,�6�%
�ö�D���ͶpQ��C8%(*6�!z�$�WQ�����Z,0G)B���d]<�^�*���|�:�Lh/2Ϯ6Ζ9�1�)��u���W�*�M���"��Ld��:}���ƣ��ڹ�l��#��k�5�����6�����S��3����i[sg��E�o�m�mx@�'�yC	n4�so�k��T1�|N��o�,�p/�����	0�q+i�O	�^X��J뮻�"�m6ɱ:��f��^�?Il�E��m6�W��ɶX�=t���˹�ś�������3�a[xf,,oH�<�e7��E�UG��%|�>Ev�[ rC�Ȁ�1k�V1�+���#ӪI���i#����EOo�Fm�t�Ӹ�������n��ϥ擡���ĵ_zʻ�3��3�I	�/�6Y��'�q���p�G��t���P�W�W.+���wdkrĄԇ�ݯ�u���<�t��SF��z��UN���nbʈy �ƅ;O�!1SHK�ÊY���f�\5*:��`���J�1�}s.�+We^��_k�eQ���`��t�a���=S(E�C�P�e��\��PH��fxw�I"�Y��)�YQ)�r�D0~�aY�!.����R� $;���4�j̔�����Szû4	��%U�w��#���c��ݔF:�8ug�_�Fy����Ɉ��)�@��s�	h��A��m�`�Q�tjt-��}j���ڋ��{�>�:w�yLn�l�䤸_@sɑ5�IvE��&��qx+�b�IP�X�;uب���_ޒ�y38|)8���|�LX6+¯�&����%��E8+����'��w���*_�&��(����8�����ľk�o(.��^+(.Pk�*���X��+nr�Ol�<K�r3Pi�8�� �,��=x�᫥����ܰ>F�q��\�>բZ/y�9g*HO�r���0�����|�:C
�,��p�h���'V��g:��&�������{��]B�������.-�g�|L�C���+@c��`_���X�z���y�cƾ��#_�~̛�/��������L^���C�u##q���ڗF�Oq6a�n_�dN��YsSH/"倁� n*9?5�Z�q'��[��2�d�|7�ل�9�� 2����}�����Jب�mK���+Es�sΉ"��9ʆ�S�I�w2��T��?<{����KC�Vdv(O7)�?��s��C
����e��,�Y�o��w���͖S<�_����yљ,���S�Ȉo茎H_U��etR������=�]��a%K�.,/�c6�U1��E����y�f�JX����Ӛu�a�@��n>�<�:�Mc�P��v�~#�,��������>����q(=��jU8��H߄謩7���0�`P'g�nVv?_�tܐe�}��F�ȦgC,�ֻ�}J�N|gqlrȰy�I��/�e�ȱ@<�ܒF�8����o^�lI����p���[�1��NK@��CY^�*���w���!�;f�7�3ѿf ��Ll��D��Ъ�� ��!@��W�F+�?N+�����/]�b��JGX�-�U[���5_3��ȃ�.놱��3-�`m�O�3#��y���K�1ө �b�l��4A���>Zf!�Ԓ�7��Ir���ߤqe/���Ӫ�TZ~X�
]�Ŕ�t'��(k��C=7Z"����Z�>���#�N������{d6b?�-�f�4Kz�aF���ٶe\Jl�l�N��7�+���lіn&��W��=^� �L�5e�<�����x'�D��y^�� -�:����r��L����^�Y�̲�e�	\��
?`���7Ϩ��xb9g7��+����'��JS�KOT��w�z��c�a�)�ix�#��P�-�R8B$�o��Gjq �p�r�I��&MܾО\D�{PY�b�z+l�^�t}0&�"kL܆�k�ڜ������oɄ�^8��0���?�7O��8_�z�}��'�.��wI� �q�SV��7���/�V�����m	*D���_��{J�,��8�>�Z�ă�d�ث͎�j��pe�p�e�@ߜ�]z^�����eS�ق��ԩ�PZm�E&O����)'��Aut�|sF=ΜX?lڐ�����������`�Ue@[f�I����Vݤ*7YL�E ��F��D�*>�J.q_��{.�:5��Gg�X�&/6GLb�ڬ�7 -��&\����m�3�p"�4yS�Gc���yY��saY���홏.%�2zo�]R�D�Z�\���D��pa�l��4�6��"F��=�F<n/{�4�"S�=�����������"UM*B%L�r9�AQ\·n6Y׀!�2.st)�� �*|��k-���&�2&O�(y�1�s�-��Wa�����I��;[������/5&��_i�h/6M��˖~�}�0��xK�Õ�ܼ鏢�����"�4�����<�ؗ]�Y@�'o��W��4k|��#�_�vڨ���3����_��fMS-z�:���܌�#vH�U�'u�P1�4�R�9�<BGH��+a�W��,Gb����OK���"z������k�����+<CeQz���*���Ϭ����j.+r8m�^������i�P��������B��!	?�]�!��ǮycDN�����F�~˺�({$��H�tN��o�~�	V�|o�h��p���|��'��E`��	���َ��x��i뽔����#TZ�kMɌO�D�y�ψE�I�5��" @[���Q���n@������T�Q7�4rƑ�tEc������y
y��9�<���+��pft��ʶE������ϛ�X)x0c��^���/S9��[xN���$.(Y�@]�j�D�D�n>l��ۮEkg���jd|wV����)�K��YI�~Qm���L�<