��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�rQ��7%gN���i��v1��(���:m�>���D'Ͷ���tur)���!^���p�NW���^��I<:�E����Gd ��L�y�V�����`�N�_-#�ì9y��^�+e�I�Xɐ�b�oѯ&ioY,��z���ͺe8��l_H3ud����C �V�����5q������Jv�Zr}��pj��5X_����a��H��|���6+��g��T_p:��X��I�o��C��pz?�*��)# ��TMq�҇ �~�-�(�Ͻ��3W���n��-ҀW�J7�j�����@��:�s�6�%~��X��%�dk���C;r�؊�7���	�@�΍���x�Fc�pZ����8�E�HNQ`��X�{?�V�)"��ӑ��+:G�#�A��Q���5�hw(@^��\VD�`LQ���@e���d�B5�T!�@�P�k��*�˻1x*�[
���A�4����Z*!q�X�� @�٢�j��� ���V�m@�1�P<&�d��+�S3����G����^g�ˊ:DJ QEw����%{
��1�MQ^ﳗ �D��A�W
i��q�}�e �c�ӻ�5��Rt�e��9m-k�d��Az[�,9�4PWh ]��sy3x9M�����Vn#��0�>�'�f�i��7Z���^Xh
%P�2~]�mS$�c�w�X�0�|r��	�|��95�z���k���$g�HX�Ζ��̧�*��H�.ϟ�
���b��-h��M���mW�n�e%hm%�; �!@��X���ٛE�C�+�y�ʊ����Y���3���>*�.w]	�pV�g�u��>�|l��l�5�Q���21�wo��,���5���j���o��$��l2u#a�Es�8�^�0J�$�f��61��zҒ��Q���7��N*��#g�sCC����В�O��|�VTlp~�Le��3��P���/��͵�7����C�Q�]X�2�b]����9s�cH:��ϟuls��B��f������ff�p+V���D����K!N�f�:�h���}a1wC���s�����9_.&���L��_�vg�[4<od7���XN�y�"�r���[w\��wp�Z��P',]�s���Bk�*'X m�E#Rǳ��3jh��}4́[�47�E���G�\���M>N)��{Z+&�z���HWͨ�c5!��H�J8���y�̰h�6�1��L
Oe�I+!���ԏ�Cj.Om� ?c��BII�P?Cq�
S=4��f��߽��'���m2
9�d�<���'ŧ�[k�����Ul��h9��l+�EI�J��\�	ٗ(as_������˾O�`Me���Թ����+_���-��m���ZU����u�����{>M��$�0hw{��(N�k�5��sR�3�d�.%�N�}џ��6���&Q���쀍�!J����-����񪱅� I�!*1��o����m]����?On��5��&Ʉ�1ZH�Xm��a�x��f(���\��t�g��	䐺��L=�0z��K�_#.��	��'����q&VX��t!�d�A��*	2c�������u!��'��q����q��Z���_e)�1ȋ��	��ኖ�}K}wKe��\���y�it����lډ�̦�*��N�h�8���i-�"C���-����!.f����}��U�7K!j*�!�}�<s���#2rȖ��us��\	�f��Ǜ$�9����϶ر[�@:V� �P׶/�+�ox��	5e�jXGܲtLr@bC���"�
o}��@	@��@)�T��Mk�6s[ҥo:ߐ��t�P:h��8�]�0�W��?6/�3MnN%v�F�IO�:�������ޚ�K��dR�εX�Ω/����qʗ3U�O2gԯ3K��)wW�(�[���-���xܱ���!h���%�����|R����2��dŬ�Ty.CX���|�.E��HP}�c4W�I���b0�x3_+�)�Hv�ƨ�q ��,%Mt|L�����q�!-w��F��J��9�mt0c-�$����Q���W��I,e�ˋ���@ί���qv$ʾ)�Q��g��C�f})��}�{��ͩ�/���x�EՌ��n�[S8�N.]#�l5T��9���%���pq�]k�ݯ"<	�԰�j]���3P�cU���}������������r�@�ɫ�4��V��$L��ͩ?}V����Lik: �ib�Fy�Ť�l<ɀ:ǰCk�,Y�.��5 ob����[�L��;D��2nɱ}����.�-����0x�'g2($6W������W�RU�^� rx"}ڡ�R��쎫7@�ٷ����4�^/�5p�1/�<9�5˷coI���fFۙ+�]^�w�6k�&9r�9H��o���1���>�O�i%�Q/�=I�DT�c��1�~��Y�%�ԜȚsDO�{tY��8�"���e����o��|N���ƙ=�@ü��������}�����!�0���qCx綷^\!лG|.�Yp8\�VA�q`�U���{o����K��Țؙy( e�j4����Qe����ڤ�!�J�V)m"��fJ�\�P�y���W����XR场Le��¶�����M��������;�Z7!^ۼ��zyQ����&mr��%�k<]���fd���[>�+�t�2�Ӧi�����pO�s+�GI�9Ee��� A���Y�/Q<�WQ�'��̽g��:�S��9p"RѝpP����
3Ǧ���N�SB��/��[a@Y��Ä|�.@+bT��V�����6����Zю�b�klkFv��p�9��)m�Fo�3�x��9r(u�r)�p_X���.�����]�ZQG�|�������[FP��% �֓R7e!ۘY����<�u˨+b�V{tiS��1�P(��$�H 3Z9؅FL��%�%U��C��ў�����]܅�agZ�?������b���9����&@:��b�E/)F��򍗧��Z���V�Y��{����I����e�����?4+$�6J�� �����ȧ}�r^!�:��ǻ�3�;��	"M}~О�g�1r���$����=>Z�7��0��R�iD�Wti�/�:e��KQ�y�<�JPDKBe�ڰţ����Ȓ<��;/��8o�t�S�O�c�t�/m���7����֛ �NO��{J�k_�+.���x�qs�}3z ���<p+�?2W�³�����������&��H�Ͳu�ָ�+)�k��/���Q����Ϭ�F�h�\u�����wdƕp�s�q/��[?s{�y�����	� m ��q��b�E�#�=�ϙ%S���0X���0�v����u�K�a��s�K���Z}�������2�Y=�&�^��%c���.����S���Rl�B�75/�e��Z2�R�s_k�E���Wpԯ�d�痐�'id��z��"���z��',��t��]~����%��v�br�t�\i�+6陜���Hio��l��n>s��~S���;c��; �::O���aIQ�
�^�>ۏpP!�PjeJ{�B?\���-])@eY�hU��?0�j����.c⛅7D�D��읖�+��ET���/���%[.��o*#���-?0�~�����"j�p�V���J��d�	�3�W
��_�<��@GHC�^S��@��`/�y�!�z��O���p��W��,��"�<���HW3����jm!2���.���Z�4�.>֮ѣ
�����2�7�Ww���a�;�|�����\=��Xެ5@�*������ߖ=B�'�&�����_�/o�}��i�YӲ��*�{�\_�N��׳-����јY�
����@f��;�C�Qm ��6o�1/k���2p��)�j�SZ����!&ϋ}�$?r���d�i���O�#�Π0	��7��ݵ��;��!}2(�V��)6Ϥ� �1�`�K2��j�ǧ{��.���=�u����x%�x�=�R+�Y	�o���W�kΈ�����2O_��3�y��4�=��;��D:S�Y�)�\��'\k�K��Ȧr^ g�A��q5ҞdPI���^7�-WNVq0��D��t{��h�D�M��~ȓ�H�4���k�Io�=�y����M&�Ac�.��Q��~Q�7K���0 ���0��Y/�1 Ğ
	���EW���ڒ��.���'^�t Q}�y�<�]��==]���l<��;��b7ǣYH�#s��SJ�?�S��G�/쪆Y���
,�[J����d�H����5�x�|f�x��`Ӊ�5֭L-�������N,Βxt��ޢ�g��K���A���$���1�1Ӷ�^(^!�[8�+����:�$$�*���VP�l�ϭ�x������M3�#��>���R�g;������~שׁq-������h��pŷ�ȵ�&�k�C��5ɳր�z�[�b?|D�_���.N5q����v�"�0�:6�\�*�@9r��K�M��mܝO�+�aG��T�������
�	���=�������ʿ����LV_x�\�8{��Z�ޣ��4�Wc+�T�kȍyS��r����!�+o�Vw�����쌥Ȯ"����:��3��A:�]���KǊ�XA�;`u{�xv�8O�"+�=6�x�4�X�UJV\������ ��@���^�mm9���P{C�����Tqݱ�4J�|��E�#��f���)�&�_��ϓ��c��/�G�&'��f�_��S��*@۽\�n��_/b�6��S��~���^���:�J&��zžo[� 0�In�%���GW�0Z��M"`��9>D:��IC��.e�ZĬx�2-��$n,~,v&�R�_RP������2���ӡ�y�������E�i��)̤��oՖ��.���nh�a�+>��j��
|-����=V�G롹#�l��� �-|e��P���2�g��
��h���m�����A�4ܱ�s����r?g �\8�"��=���)�{����?r� �g�^�Lv�2�����T&w͌�Wq.�1��9�$,<��Z�Ri%�8,�(������ɥϚ�E^��9\,B�����u�]8mm>��=�/ȥ��Q��}.޽�XҼo@�k�?�d;9��ht�kR���U�n<eh'�2oWf@զ��+A�U�m�����bqb��$B�� ��� ��1�*�o_Qki����:�)���W���I�H��!�ȷ�%õ�Af
"3�i�ׯ���{|~`�`e���IE����Su�r�'�cY�!?+� �;���;N���������O9L��仳cY�n���7^2>p<����V���ڹ�&T��3��ebͰ�H��u?i,��rJ~7��We�m�=�/�5t2-�2��e%r+�6���A��+��.��r�"�cԠ�x'����B�n,=��eF@�}_�u�!"LM�1�mY���94�f���!�o��*>�=xz�� ��c��28:��	���S��x9�����z�T�7C�L�3�.���M8�;�/'7:ô�c����:�<PEF ����I�'Xo����Ъ�����\���WQ2���h�hw��SD�H"�|O0�U3(�+*h�"�2ב�ĥ� n�6 ���~�ڡ�|�_�w=N�$:��$%u��=L.sF�8i�DeF���+yS!����Hd�<X�0N��x�sz���G��`��r�'T�\՟�{��yepZ�Jz>~P�i��u�B��aLA��!3?`u㖙V��
}=�@.g�bǆ	�[apr��#|��4{��w�"���1��&���Ҳ�E��_��9��J�VW#x] �"�n�7�q �,Wm3X���F�2T:
I���t�Gaމ�(X��L7p����IeR#^�+�Xr}B�|Ĥ
&1���/bp���c����ٍ�oΡ*Jk��R��C��pV������'�c`O��+"�1�y>t.�ݙJ-��G�]x��h56=�� ��}��϶�G|{a���K8���?�ؕ�ќ�4h��e�?O(�1�Ķw�&�������?��V]�٧O&�ui}t�2�"0k����4��tc|�k�5�usNS(�dc��ЇHv�|��5�<b���laʎ�U��r&�}��{Z*�$���R��n��4�ሶM�S�oT��ڛ�p��|������f;��R^�J�Rt:��Qrı:J����Nh�'�= V��e Q��"�n��Y� SɁ�Y�U!�Ȋ�M	�Dh�"'I���qСx�e���o�C��&o��p��jW<0W�0=�{���>9�Xs�:��|N[�}��N2�^�_�6O�h��'j���ZKƖ��t��L���9؍�g��R;C$�U�@B�(�1�����Y@)Xά�?p�2V���p�����M+���!���|�3Rl�73?���~���9�3����Șf��]��( Ǵ��~ްmDFK1�5S��1舯�_�ܢ�p�����g�0ssi�sv�q������'���ȴ>EMT4ub���d�@�M��� �P)Qr!{�&c?mu#O'�訞�Yj�WɉЀɩ��P'���a57\�מ��N#��
R������F�%X.Jv�Hԥm*Nc3+
�=�o�#BT��g�(��IZJ1�&K���驠s�8|v���s�{��V}��������$e�(}ֹ�y�X�L���;_�d�n�r�d�����#��M����f�������@ �0��M��.�}�z��N
�;s啣��qVnjE�<�:����������~���١��'�.ĵ0����ӻ��1��9��{����|��
������3;��~$e5V�=��	w\��@׉������޽�u�	kҤi�����g���HGh�&O|�;l�h�8Ɯq�7�iQ"����9�2�X�!�n	��3�b����'�.�n1F���"cDq�������R��
�k&8�QJV\餟�q��(_DO���M��gk�}on��kX%�FH�chS=��������/�.|.`"��*�9䜞P9��v>8�O�?����q]db����Z�����Ϳ`h�$2�s1U�����9����z���xo��\Ȍ��X�8��
n��#Z>�������Ž��2�H0J�!�����_�]wS�^l՞ٓU�иrۄh$�}?ݪ�`�&� /x�b���~��-K���[�>���h��sm��P�_ ouy��1�ze_[>����kVq���@�ˉ�y��a�p�mYߐj5<�@�8���2������I�s÷�u�A{s��p��q�w���%�"� J��UTH�O�%F�C� �L��%0�/�g=:�3��������k��B�D~ �0^��g�~�z~���d$����;���l�qG)Mܙ��WPK#���BM���$JT��]�E�G%*��*ON ����L��/M���A��O�d�1rE�!�:a�o��K�\����ʁ�>����L7�͑Q��Wܥ���=�ܪU�K1��2����SX�f��k�&�<��z�c�_�g- �����a�ԧR ��"NB�ڈ0c��$*V:�AЧ�ǌ��V�����U�g��RN�{?��1#Ls4��~tD�`�G�k�5YM�c���p8]���'ب�S�4�����9�e�\SUi����7�m#1}��"+v�ivOMds�^6蚉��(>�t�?��|:�MT�49H��*���^̆qz�p��M�"EW:�&�E���mlB I���C�~�ӊ����7��iÁY$G�������=2�iD�PQ3�R�@���⸎|�,@y���=�ŗ�u�	�x֘1H���_�B;��[YݹCBcqR��Q0C�cQ�+;���T'�ا��_���po/sG�Ӄ�ŝ�}-ht�^�D�=M����I�<�0ʒ�g/��$3#��8�{�2�}�ߛ��Ǡz��0�2��R�Q�u*L<����GqY��09�
K��枨�[���%1*�lԹ��7ұW�G��ݙÒ��*of��kXB���Dz�6�pјTr<_<ַT6X~¾?H3��RL��xh݀�����Oh=�ʟ��g�Q�81w��0$N�\{/���{���/���˩��,�G�"4��!�!OD��p[�-b"�*��L �����mjЇ�BېAnצ\�j�Z,n���2w��'c������M��Eʇ-�R߼�x��>=����ˮ#�#��١�
i�  6ZxkL{�����\R�Io!�a�Y>���D`�U.�g���t�5`c<Z[m1
7�5zM!��݁�,c������,i;
/��~�I�˺+����N�_��?`��/N� �`�\KE&�K��ϷB:��EY��C_��8k97�sK���p$�������2pȵ�H�K��}p�Sk)G�O�x�~'A�W�	 =&�Ʈk4�=i`�����ȕEŵ�CY5HE'�>��8�M��E4j���f>��]jm�B�ݚ���CU�f���@�]Z������;V�4��f��2�0��o�>$�9��,��b�a��K�O<PԸw���>&(j~'֥/����z9碀O��\:�[ѫ A���Q�M@���{_%ٳ�ߋ����"پ��t�
-��0J��>�O���7��M):�:JL�,"%Lw-��'Z�� y�+����CG�+�8���
�վ �S��/��B?|��bV���RXI����Vl��M���R�QgӀ��YD���!J��M7��'��>QKǷ|n�4[1F�ݽca3b+*�_�uѝ��q2Z)��I�$J����	g���E�8��>q�R��� cpN����S���L��A�B����\8����D��-�0v�mW)
_ʶU-*�{^�c�^��ݹ@���1\4Ǖ�S�O��?��wv����b(��)���s���rF]]P���iX~S̱��i�FZ�h����g��<^
\�8��[�*��H�F��%Y�N�0�/���"��ւ2�/���c8���r-1t��Căݴ*&������6!�6Q�Cp&�)��ы��; ��5�J��V�s��V�GL�^��,x������Yp�t��Is�ߌ��ER�͐W?�7j-�,�������z-�Jp�`&������>".}#�����b|��Vb��.����x��+K�F�>4����3v��ѻ���Aw������dwu4���"ͫ5<Q��=�G�⩖h���3�����`�c�y�`QXD��Y���LP���K�}�e�̓�b�N�����:U$���
ښB�qt�i���$�E��u���(��h�3BXĀ�N	�Ƭ��WO�����������C��v���lm���|^O-�8|�1Z�/�Gɳ�>�9M=��DV�;e�BO]xY��:�7�~����k��1�-���$:8�nTq��?�T��a�-�^� ���ב�yX��I����meןd���O ��v��6\¤����t�"��d=�o=o^���F0by���
����+�އqKWe#R�x,r���j�8(H �N�p
S�X_�����Ik$�lx^]곴v�H���,��z|I2`G�ֺ%��+����G!��d�c3���B�&���4oc��dAE}��O���#����@Щ츏^_�Tǳ8�_���Cs��V�$��C�4֞�x�գy��֘� ��F^�r��ֺz��	Q����<k����N1�퍈�J���LP���%,PA�Ӡ%�䒬��D����W�*��Y�|Ht�Ƙ�bg�u{B�(�2���E�c>�*0��ױ��iB�o00x�a*��PC�x���z���|:�w�W����b�k�X>��>a�[�gas��	�B�0Գ�	.ҧ.`?);�T�*�5[@֬Ou�1G�%'���e>�rƢ�Փ�C��(c_���V%�#p�돊���I5���m��2�=�Q	�έ\q�c�ʩ�cMM�;tg�Qѡ�騀�Ị��@�8C/�%�_����1�	��{�������%:��Wч�����"Ulbu�lZ�)��9&�RU%���=8[�y��z`4��+Q��()��G9@0|^5��uu܏�8kط�x �x�ԹekU��9�0��+���!l��RW���y���|��U��CXQ�/�[��<1������Pe��@�n1w$V�x[k�0-�#�.�<|�g�<�_D��0�|��ٚ�xoʹ��qq����ַ�{!����.4�.�.=�'L� y�̉^�b�8�%hQ�X<�N��?�lW����v���ț��.I���k�[,Y`Ng[h'x���:�,�t^�*i�:U\�5�D�N(� �YC��!��DtA"����P��W-��U�S�>5dP|�$��E�#r��
쿹��x��ThM娐��	�鼪_����;�YWNw˘0��D�Е8z4�RG(P�"��=�dLdASU2�ˌ��TPI�~��^c*!2�-�=+�ze�%�Hլפ�G�f�a��,�����<b@�2O�R�	�0��<07�η���RX����g)�Et7�m�NLk���'n���e �Dwq0�!��E<;Z��3�r�d�jnVH������b��Ί9-�����WA�H"�	I�����̤�Y_�WST���+=����<���0�����b��Vد����<�?�7U��u��=���c�#Rh�
�%{x�'|����a04F��K�'�@�ӑ$�}��c�-��ݑ��Z��j&�R��s& ��6Ղw�#��C�Ƚ|[�S`Fgy�����G�ªG�ȧU�ZV��G{�n�+��QW��@�>�Ԣӂ����CTu>�:�9*��o+�^Y�;���-[�J��� �J�Z��fs��_��)x����ިH_���x #sŅ��$4��Q���cS��Jǝ`�[ �C�q�zg}G�@N5��%f���E�9Χ��ETJ7�jsb�({�8Ce`�����A��`��8��pD%�ўQ�)��j,���S=�E+�k�]�X���H�ZLT6L_�2�	�Mk�L�� r��:���q,���}�o�����@�B�"�qW��Ic5�z�R�M%��I[9�f�-�x�h�y佔���(�@�����7����a��*׿�&v��;'�&�\�0��(\�WJ�8�5����3~LG.�b�'��]��B��[���W�ǌ�K�����&�Uu�Z�`���v��<�x���J�Ҝ�a�n�s�j'���S�`C�*�_��
���M�c�ԸU��jԂzz��CM���E��z�U��?[��`����5~K?�V�����2�Cv�__{4G�Dѐ��̀�iZ+�ϓ �C�A*��`ιa��ǌ�mF	-�6���-�N�@o9������ǡd�!Kb�4Q�{xt蹢�@��Qos0�FQ�ݘ��Y���������c�u�p6�ѕ���/
�D�bV1P"�е�n�,1k����g\�{p�C[;�r����K�^�V���x�iD)B�X��"3�K�Do
�l]���`k@J"7��Z��J�������c�{���'C$ѱ�q)!��t ����x�L�@{M_�[�|(5���+����<��T{�Wm�I�h�=�N�F�L�#Ls��ҙ�g7��i�4�V��{�dS�*��:*&p��W �g�����"*��M[��q7��.�UT����PNN^�f����~�;��I��9.�?>&��e�J@v�X~��oի�u�ׄak��`K����2�%�{6��9I���li�]]�/y¡����֜&,e x\h������8�٫$�]���H8��~x{������A�,����M�L��`�k%��l��e�� �{�Jz�*�80�x>6��|�G�O.���_�-s2!�UZ� �O�O_U5ߘ�1B'ju5����U9><l*2fsF[Ĺ;��؇.J���g(��-g��+Q�ml˹z�/�Ӿ������J�����6B�?e�;%&�3c�]\U�g��z�8�|���pᮍK��+?�#�F�?=�.]th6�u'�-���gi~�I�kJ��3��@� j��x�Z��\d���I-�wY��v f$�z	�����$2�<��+��~�r���j)��੎z>8��'x#�ЛU����2,���$����d�0f�(