��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�J��"4�=�7(�T�JѺ�ő��,\��s���ӣ�F�؏�#��ѣ��4
�j2Y�!������/�9:Rf�-���v�b���Yɼ,��̞�SRp�kW�gk�VވT3��$�ƞCY�C��<�Д{�i
E�./ =�Ir�Sa1r ��W��|�Q���]٪��ݞV$��\�|���K��)�6[�~�oz�o��q��(�P�9�A�zHq�Ԃ��"&7��SI�"��l����y	��)��V�h�J�����gOԽ8����SF�q��xO[@O��'�sj��xX;�=��{w/#��U1�@s�J\_�rh�����L�fg���5�%�#(��t�,��ҭAnf��yV�kN4�T���'��z� 2����Xp ����ٗi�^���-�k���Ȅ��c�A�' ���ڮa���)�f�<o�J�C�ܮ�jfXWb6G.�!ck��7��vb����]D��ւ�}c2vP[�cOŏ��"��7pG�G��]���ϰ�Cx��r��>r�H�G��#�]��|O�jQ{\���2���?���;D�`���d��Ģ�m���Y��X9�;���dh��_wO���"���e1�DW��QX�	V��`Vִ���0�WYw2�ٹ�+(<]�0M?��"�����Oj������^�v��.GsA�X�W̅.c���*V�R�8[�nU�ЎCɈ$�j$p�q@�S�8��R�0U��p#z^�X��ո�����=�g�qK1a� ~ʹt�����a��B3��r0Ɖ�+ݟ,kH��Df���o���v3.J�순�]u�w���Juuդ��"����Y`W�p��3���=0��B�b���jʻ��Z"�!&O}��5���r�<kI���`����3%H��^T6�ѻ����l*G�Ð$� �RGGU-�B���,:r�$��
Z��|� ���ϭ��;Y�r�J��pt�?�+aMC�)Q��R���Z\��ݏQ�:YJN7��]���BY���n5�S�^Tޒx~�/��с���3WU����cHt�ĺ8���_ 	W�('�R{��Wj�o���oBW����z^�,1.)�X੔$;LQ�.j�x����ݾ;���}>�yy[ �)�z~_Xa
ž���
���~��4�f�ޱ��3&N���R�~�D�4�FE�p�/� ��C����؅f�Sz�rI�d����!�A���`�d��@�r���hw\i+_�_��v������:�6�s���3fS��	�u���W�se�1
����f�6b�[�5�'&q}H���8�P\n���4��������hQ�Ø�௾l �/|������_Ҽ�z-r���m���OSتg�Zg���F7��X6'��'λ�� ���!���\�,>�Q���zmY�q`F��s.U�x��o��P���NxȄ�/��`%P�Ë������0Q��V��b�oVzQ�P��a�i|���){��� �Pˎ���B�U�;ۃ�Z$A17ܭ�XN:�O.���,]�m�\�F�2��gd ��V��tp2���P`���}��y]
����8nfU�7Rr9eOS���z��()�3-Ҭ�d�t*�e��HG�C<��4p�������>ID�E�O�߫?<=N�$�-КC�Ŏ���8�Y��"�C4��_13��q�a��̀��&���kS+��xaz�	���Z�F�b:,�Y��&"���[*t%��|շ;�?�Z��a-r:�N%�bs��Px>'�2l	t�I��y��鍮HL"�%R����+ߵ)�}i�Cx�N.��Ea�h��w�m�}��~?x�ط�	�\�¾p�����;=�Ns�ߕ��[���zg��׵�[�a.f*�R�9���B��1�)��"HT�;'�B�?wFi�P���1�Ue�>Jɮ��H<Im�/ݨ)�� �n���[a����t5�S��"�~��y ���D�N��/4<�~��
ғikf*MSwR�U��ZV�����|ŒU�7~��8|؂q�&�%yas���U��P��qQ�N$��-�6�2�mnRec�Ɍ��s��E�ܢ]ĭ���
+Tc��ZL���\���ws�9�0�OP-�cw�����%Kx7^������b�"�W���/VD^Qa�c���M���#-�n.z(]�%�8����-}�!��l��ͻ��0
���� ����uF�@���y/I�����~�/�!�`���a7CE/
b��k��n�$���P����u��P �1��FW�$|5 �_*ڙ v�CL:%4ss]��d9oA��f��{/��V(�M9�?8G��C��$���uQ���CF�E�h��WH7�}��H���A���y��2��^t�ڲ�oWkD`��]�JH�S�`�{9ѧ�"+�u���]�}��X�g��*���g�^#�P^�}d�+��w�W��U	�������o��i��?9�W~➺b.<7XQ9�-���ׅ�!3�+X�FT���b�Z�Q~�4���S�B���<�e�OW��O#n����P���;"��9<��h_�-IKX�5��<����!^�X4|>5�M�{�t��/ɖB\|)��ž؏y^���[:������db$P�W�=��Ϸ���M��!�x��i�"��T)�7�
E8J��I�d�ch0|�/���Ԅ2w>�8d�Խ�̫���XCmP��Pvؖ�m\���4#��_����x����)<C��5����<Na�����G%dy��ɣ%��*. Y�(_@�H��yB�y�dL���a����q�I�� )0`����{�n�k�}a��U��au;^��k�B�Da��C�J�����\��)���/&�`��HՎ��{S�ݞ�P��3���]z/c;�EU�r2��FH����T{!�(&�!q�0�:3����}u�6~5��$�'6_���4s����X.8 &vNHmV�?Θ�߰Uo�����Q������xo(KZ��X\~���.`�/`c���dj�A�L<��������R��G8m��6hje��N�ͤX�gO�.tp�8ZY�<�#��ï���,�?	*�c�J­������]!:{�1�\`�I>�Q`�n����3m�<��4��^gh+zv�\>'`�\'hg�����	J��+���'��M4X�2��d���<��
Dd�o&�G��q#���Z��\�+�7�+�k
��"�h����{FOZL�T5��B��f!��:֯1(�Abrb~�W�]�V֣@;6���bA�QZ�I�7�*�(�Zф%ԲTc�dhK�4��DQ�\���G��®l�����䬳�p��GE$
���	 �o2��\Z����RH⍧�;��ɏ��@�ż��Fŋ�s~�м]?ȶRp~j;0�H��v K}5��_N�������3~�2�5k�����D�x:@6*g��&�ƉOW]n�����Sb^M��y"I�ɾ�|�gBe�xݪr�V�
�Z�����2YS�D�^�����֞9�ћ�o}�"�P�l]�e3*q�����R�S���<�d7�+�䯙\���M���qw���j�>��+�W� �BA�$����v>���^�����@h�8�I�rϮR?�Bw�I��03���I��2<wr]��ܸa�W��HmzL�HeЗpM�\��b`��#���5���s�qj8�K�X�σ��n ��"���j�3p����E�/��l�K�[������ �=j��,S5��.�8C���D.nQ���p�� S+��ʙÜW����]9���ajE��bc[[�uA�o�^Ǝ�P�Z�Y'���� �~I˛�fl��U~Ƈ�Я�sE�\�:J���.l=�JViV�@�������+9�Go%>l����fТ��^N�w��y����I�Ao�$׭��X�H�:��Di�\�p�ޫZ�����1�Á�y{� �[J�����Y��^�0e^���~<�F'��t�&*`��=5���N��w�W"��$TE��NΖ��(���H'�{�*�4�(X+��{��7�zy
��9�� ��߶�a˜*m��SF�e��@,���a�L����.��� ��T�j7�][@g����	��:�3(#G�ڏ?t�^�b���s��S�;��J�erگ�5� y���L�I?�n�sF�q��W����h�P�cԧP]�@w����6�D.��GdaH��<�)��\-�'AM`bb8Lv��*�/t�#ÎhՇ�%�r�)_I��p�������.0��SͮD-�:�Eΰ�U��aڨ�l����*�b@0�a.s��B=(�����%��L&)�Jm	@ˢ߷w�eU��HW�L:������s �Z��J�E$���L�r����<w��K#������~���t�}5���زH9�S�֦W����/A�0>Б��x���H� u����3\f���AA����{Sy.��[�ObJ��o|��W-��J?��ٴ�V
:��}z�`|~j6]�9_���ɟ��úq��W�1���"1NYR�<�u��趎ו������= ;��S�Z����c�=#��= �J(1ۙ�s�(�<���z�-�j�B����l�N���>��R�"-�#R������w��5S�^R7X�.�2�[G�+N?n�O{q#�H��bD͚�rRz4A���ey��\��y��r
�RIA�d�8�5����!��ak�%O��=q���:9ԉ���5H��8�o���mG����);�!������Iűҵg��ג��`��s7C�*��4�(�H�����6��щOe�a����{A���G9f�l�FV%y{Q�oъ�y�6�\�����̸G0�f�nMwIq����#��$3�����v9�Ou��8X2��$���aӭ���;��͋�u�WWO~B���w�"0P�!kz@r�\�o]�1���T�Q㑚!�q�T� �B��}�2�r��'Ê}I@�Zv��'�R,+���.ϥK��3���ߓ����{Nc���
.���3��{ج���ig-!��m��;�3!�:���[tjx�C�0��ܯ���C )�;	�?��#|��n�$	����_C��?��)B�Y��ߕ�>��ߴ9��A\W�g����P:o�gу)��Y��lc1�랶ᴌ��{EEf7a&t������1����"b	B�ۇGS�G%:׳��c֜��m������3����<���{�ަ&�L�إ"Ҏx��ymX,$�	F�j��w���'=P��C�N��<�q�Z���t�Kb�����xuoV��i���Q�Nz�hiQ}V�
rӭT�_İ�R0
�i:^��:�9Y�P���i����ն�\Y���L$ɲ*���LVh1[�_�~������4�t�j�Q�1����c����PQ[Ѧ�S��ɶQ�X��0��׿I+��ȩ�l�y�dc�ءɜB��c��ec��̽f��$�@�џi��z�R�i7�J������!��or��T����]�ô��*l����q����HF���/������6S���m/��9����	������n��J�/4�%�\�i��R��O�]��hZ�Tr��0_���ع �ZD�� �~�)��jH��q5̠�P�KZ5��G="N����ϩ}���W�.�u��v�Jy_�bz���RN"��=!s�E�R�N1���
<o]B,�%g�~�q�y����*�í��q�2��Šd��G1��v����;S._F��{rh��)��2����TƵfVw8�};8��\�ڥ��B+ɑ~�{Xٵ�M���{%�n�b.�w��Eg%�������$��K����]�C�q	�	H�9�M\nb!��W{�o�k�K(sĨ�{|ꥂ�1jt>�T�V���������V�N�n�o�>�ӚFh��+�O��He���fp�p��LIq7M?����y
N����<U���Yq���z���R�h������^�X�A?�5Tx���6J-u�/C
��\���W%����[�� Y=���n}w�?�al,��J	�>�H���"��_ףּ*lm��I>�A��@)T�C=<�w���*lfm��1V�