��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|>�qT��>��*�0P��]�*��W��l].UDY[q����<��;0��ꂂ?��Q~ͩ?E�Ûݾڝ������"2k���[�մ 2�c�Ü��N?܌�7�;�~y��}�Fv�J��)m���v�t��s"4~#��e�w��O��,���o,?�1g����;�)�!���oFZ���9�ޮu��}y5����o>�`�^O�&ʯ2	e섧�Ҧ�kct �ZT��n�t�� �5E	'�R4U�Q�$�4G������;�b2*'���
�D!��L�b=5���Cȱ��������^O���_F�����=)H0\T�sR�A
q�� �~�yo�k]>\tv��N�i�G!����!��}���T��m��|8�v(B�a澲`�?��ӻ���<�4�7�K�K^!��V���d��7r�E7��% ���]#5!#F��5&������4nڭ�z���^2(E�0����E?�KRh9�y����ϗا�,�� ��n?:btB]�K�X���V{1Z�F2��{I	�Wb�D�e[3�Z�NIJ]�t�4��|�04�*:�?͎kzi=�vZI�F�����G�'�{�QA���w���:i���-o%`v�6>�?[���2�Zd����|��&A�O��o~9��!.���yb9��O����d�WC�e���td�����l^��8ޚoW{���@��&�;�9
�0��S�R�{�븡	Smu����Vx�����y�ڎVl�S��8�
��3���߷�>�N�߻g�m�_8�.�җ�~W��Փ���M? �q�ho�O6�bwGg/��,������� yG���:�>��dLn_*8�	�C���E���VmK�	"�:|v���O2�/�?��Hֈ�Y+_���^�*�t�:��H�t��SK_ >�7ߔ�k���.��%�1��VN���|�˸��)��X؋.�p�@}�Ib�����&��G���9~Τ�F�oLϦ^����&���HX�I|�6J���FLI�T� �yD�M�૵!���������F�*R���v=�� �lҡ��&��/	�KΝ�T|v���f� �}�lhed,�S��t9�<��K��P�	Z]B�I�tnBy�D���AOt,\��:v����k�A���h�yd��+2����&�^�M������������q�F�dYP�>���[�)�V�anbm4��=e��.'f�P��3y����My�j���@�sU�0H>��Ã������rZ��d@$iǑ��E*?�&�9�x#y���s�a�^d�@����
/�L ��..�f����ͿVQ��fj��]�@�b�h^֟���v}U#�	G��_�J�����SN�x�7�=X�y�\���5�
�A�wgԃț�Eܲ�/�'�v��k��Ƶ��{++L��y��q̌�������j1� ����p-T)]u�Cʢd��NQ˻@L��CB��+����(����!�k���=���^Rk]>ȩQã��8�={g=Op��9,�_����>D;�_�|���[q�Lj.�#��.MO\~R��z���*OZ����!���t�G�d녗�d!�����G
�y�R"î�d����7�21{+\��0�}�%���b-�"�dp�	RZ��_}q ���l�˝���g
)5��.���	��>���L���^p��R %6n$?d���t���$(���	'�1��)��o����P�O��0M�S H�����i���r�^=E>�A������#����9�\�c��l���G� 2[�,Tpx�z`� %���	�+�o|I'���pϠ���tjx��^I~� 3\�QsP��Iq_��J3|_V�b@]���lvJ��,�EMS�'�\� �o�u���@7�Jy
,`2D�Y �Q䝟fk�4�z&Y&�&��IT��Q��cU�G���_'������
��:|ov�gHup�,�ˠ��"�z%�	֗4���V�Fgh� ���n���I0Q�(Бu�6cWG�џ�q�>�|U�:�dI�p���Ru�%�!�	`y�)��{a��ܜs�MW��/գ+}iqs��M@�>ۛ���]r�R�Y��a�����}'W�0 <���Vꃋ��b��XO@�$��B��6Y�
��4�9w�ҋ�)�E��>��']�!��W��&�:,��>���nn G�zO$�[zmO˾�P�2�A�(�^�+@Y���o��*ұ�~(
n�����5A�a<LR3v��$��U(���L���2kZ<�[(��|�ڃ~d�:eYߊj[���䖓�����o���+���T���c��rխ�y���c�"�ri����=`�E%���KY��c5⩕���U�8�"�����������j�ީj��C�\H����@��/}ѓ%��QnGl	:����$й��*�����4"~HAq� q�9
�h���`�������	/|�J5�M�"����t����I5jI���5��Z����P�3):YƟB5��(�0EF�\�ۦ,h��w�Gj9:{s�G ��3"�a�YI��æ%BM�<E
��G%��	M쾨�VF���Œ$(ލ^\z=ܲ�� ;M뵀����DYr�d�k��8� Ɉ��mA�x��ܗ�z1d�n��q(!m�Z��h�8PuیU�����
�N+}�H,~l �o{���_��>����B��1GEm��:Fw2JTJL�&���$X��������c/!
��"rk�.����qZ<�сW\��yי(a���β=��F-3�K�ր���r�Z�E�Fl+��%8��/2��aQP'R�|ͩ���2��c��|&!f����E{�����	�ւ+$��'og�RQk��h�}eJ�m'�(����d�9�znv��]���9�忧xD�s�������`��$���h/��r����hŜp��; ��O>�s� ��������GJ��P�m�(��-����$@s�ݶ�D?Caa�^�.����z&`y�7�Ɖy4�>�J 2��:?��2���a��/�����I��f�&v�ɵ��������-K�|�`I=IR�&�+ɹ�5��w��RB���*��@ �r/�����_]^zp�����t��c
ܫi�)��͸x���!.qh�(���˩������K��%{�NB��f�����cJ����BB�޲�棆�{W�!�>|��(���{a�_-��i��擱�%�-�h "�6_�H+{������	t"�ũ��zƇ�9�{<�	���t7�V�C�NV��x��	b?_Q��1F�c����-z�z�݀�����
�M�������ɻ
\A��'�^T�ù0�$����`�-ݰ�H"����ߌ�Ӧ�eD
����P���d��]���?��;�_5�<]/`/�kkrq0��Mj�Q�@�5��M�����!:�|r��6\�D-�zˋ�B��~���#p�#��~\�[k�S�*�I$�g�I�����fs����C�	x;�^ޟ�|��_w'� y�̮I}��ʿ�{���	[y� z=��&�������A�
"/`�|L�M����̢	�r�2�Dm�q��C���tT#���\�6�
U%�Zm�H~5�n�~X��%|�-у+3;̿Ø�
"���m�0�T��BH��ѣ����6��v�=�(Q����A�f��I�ro������LP�G�Y��}�1�}����'�~�P`
 ����� 3�x��B#�V#��[n��>�57�,5[XJ�K�8բZf�^����x���