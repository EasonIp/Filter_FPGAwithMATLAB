��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$����Ѻ�`�ue�Ú\�Ϧ�9%["h��ft����@a�����w6������D����x��'�S��=�ד�@���Z�S��-J�x�a��e�䱯*V�!wGe~�uߡ��BKo@͘~�d.R�y�(�Ls}�X�i(5��U|�~��P�r!{�(����E��v|�k;"٢�ޏ|K֐,|>���W��/$�{����Q!aq�\ĭW������/���gй��NGԮJ�� u&���P<����$�� F���G��c�$�C����6��=��2r�S�NpKb��[U��$Y`6�*��a����\�"t��� 9;<"2Mv��x��9��_�=�l=g�~Z�0*ü  ޣ�Y���aM��fKRbة�qH�����v�;~ֿ���l���Ou�Rn��[1�`{%�#OHj�2�Ϧ�QWa����ૹ���U0 �e���T��lP��s��W��;�ڙ�5�j����3�>�S�|}@�Eəp�+'f�5FEnZ0�?\+(�0&�8�����_��;H��P�&�	B��4����|�,�rT�'�x��X�{ST1�G�Ԅ����%+"�Խ��\�⟚5����Un�ȥ��<��FH�v�k���P��M�W�=R�"Y\�1���M	]����-�Z�)�1K�}�4��TP��g��o��f�-`{�3�����|�W%���r�ݙJ��3|��z���F17�����rX=�d0�/��c�SkE�Wc!2c��sv�<�k��"�d��~%�m#���ٚ���Uv��F����.}���W�W�j����i��L����aw$�Y�x��� ���lI.H��)��dF���L7Ƌ:��/��ʷ�k�aJ*0S?\�j�^i�3/���e;p�-�:?o|�C{�V�kF��*����TN����9��zh��iS#]^|�m��)-�h"qmA����� Dâ𗰸�V�f4>mZ߄���ݡF�#���9i/a�Q-y��,{��q`��ʏ�\�Ʒ:Ҏ�_����R����Y�ƺ�<�  ���#�LN���ӥ�oQ-Y1-0u�#7���1��;��>�_e����>eN��*z�y�/H�Q9}	��a�����j ����)�)��J+���u)[�5&��[RY����G�Yг�k�W�đȜP{���V��6�m���$�T�B��<�ԙ���k���O�+kL|�ʲ%��uV���7F��d�ϳ����O\���b���~��A)�Q��#i;q�Z?~�u6k��������8��A�8{�BI_�n5I�[��|o2K`$ ��R����i����w����>U�SF��'�@�����jY���_�Y[b�6q1��X���$���8�&�j��j��	nbtH�`��x=&i S��9�^vЈ�2'Ex֜U���O4�NbK�$0�^���B}i8'ʬ�}�6��<z� c!�8S ��{�y)�{�)F ����q����C�x�F"כ>e��4�N������C	�­☝D�!{V��Z�x8�4��P!~K�>X��#\�
���,A�CE�?!��G�^Ť���
#
�(����k���|�3��%�W/��X].J2�ڣ��b�����j��R�q�6�0���]4B[�D�7;�FP��_�����>���&l���/#�G�D)҂�JCH]߼ ضP�h�Ak���n��:�u*����o0���DJs�_N�ڜ㒊�.�U�7��t��=��SCĶǖX�O��KY�0�f��^4�?���a\�^䃫�'i�l��Ţ��An��w�Wč�6�����3��EeAX?݄�а�b�n5��p1D���Q~G�R�$Gt��,��p���Dro����+:XP�ݨ�Tst@���B&�`)�o�\:���U���^~�������7b Sn7r�/�BD(������_�f+a,��>����<
��B��T�l�)!����A��	��Z��b6[7���O܂��1�E�գ�9�^�7���r+��l�w�S&����4�s~#�s�G�U��	!�,r�̩Ր�g���(���K��y��uk%{S^�N
���Q�p���%<y'0m6%EZy�b����B��7)��-"�M��E��0��bDY���Y��F�W��lx�b�8�,�-;0�GT�n��9�}�*|*}Ê�c�@�m����|X/����bNZ��ăCs�f��=Hv�d�����k8�Xq�-��?ɾ�Y�@��	������۾j�{����+h�w�t��It�^��h9��8$�ˎ��hs���P����T)�\U�8	;�����o9�����-��㘗B$�sK�aȖ����>..�y��C��� ��&-�n�*�{������Md.8!bpq���1uA�F��vzd��@�1ZB�eJ�kJg���9�p���PE�Li�'�y$��%,oOp�O�uU;�9G������G�o��gR[>�7�U�Oʡ�Mj�?�⋒�(����e��ֻQ��v�P� \Sy����=��,q���/ �:L�!�ޤ�O�c�ξ ��~� ��gr�"�%�Op~���5���T��Nhb�SۘK
Y� �2ԣ�NUK��J�6k�`ѡ��pQ�u�a��oUV�ʟ�Bֵ4�Ù7��
8������`�-rq���6��Y�Go�gx��(C(�|��վ��(M!Z!���5� �d�9 ���M���Q9B��=L�ÚmFK��ٙ�� a��a��g�G���B8��{�(��..+\g	T�_�;G����^��\�y5#>�S$�q�
�6��/��D;�Z5tM�MI��{G�e����@��F¾�� �5-��W�p���%�kU�.,(���[H
���N��F|��f"��5�qAuf�׬�`MSoT�o���m���;��Lӳ%���S�)���00�Kz�����SԐ��-M^,@��pU���p��/�SX]�(�C��U��]�TIe�����E�έ�ee��\;��2�_�Q�阡�JAU�s�������&�\"�&��
쪂�,��_�i���o��9�&�v�W ��1�;׆Y����ao���ju'B�'�^b�m��Z��`�^�����ZY�i�3ˤW�Te���u��=_�.���_'9�:��(��Rs�6�����>� fB|��2��TP���fj�+��0���(�����\�kM�>�TAg?}�f�; ��}d���YPgL[�����C���Kw
Y��K�3�}V+�*"�f�h"Jҕ#�����-�g�.߈Qy�;�7�m��8\h�	�V���\W��ˠ���x�3g�Y�`�&xX�;���ڣ�S�����o��݊�������HY���ȺIl^kR�J����[ۍ���uu�՗&�nιw�b�BX��:�QݣOlǝ�eMxz(Lc!b���ׯ�W+n8��Y�|L�o�ع����+o�tJ���W�EQ���M�`�!R�j솠��f����/�l�@*���{K3���U���(��-[�U	ꝓ$ �HR���X�1A8����g��p��Tun�T��v��Rǽ�6QV��d�kp]5T�g=��4Ha��$� ?��V�8ǓU0��|�T5l���Wy���|�E��~Ӻf =YZ�ΐ�{�6c6�	�8GGF���A��ٟ�.�����(�W|�g��I�#m��Q�6�F`�|�K�/��jgvI�g�Mݮ�H(�nɹ����'���U��1=l��ճL�c�!rw�x˲�8Ll/��[xэG���SŚ.��$QYQ2��t������i�����C��w�9��61�*a�Mm���(��=��/nbu���'Vc|E���z��QAR7�"K��YQ�1�;w��:H�I�v[���!�ŹQ�y���Sm1@�$%�@���l1�;��D퉜#������yD��p�cU�/����ق��_qo�?� �kN��窾��#��=~I���g}a��|���Bb��Dݷ;���@���,MK��ŶqmB*�+��V�:�=3>ٔ�ʨ,�d&h-%��Ҿ2� �� ls�<����4R�g��.,��Ir�l���A[lDK�?����Yj�d���ݚ��k���rV���)Xŀ�Û
��_��̉'�$5<�~�q��K�1�2��i��mB��|t���4�}sړ��(��Fpu�<������R]�Y�X`]�a�m"�̝�pEd�'n�WB/�DD�Zw#���|Y�u����|��2ө
����;��_�;/;W�w� �\g��
���������o��>̌蚱��7Brq���^5X�@����č�
�p>ׇЂ��0-y@W�Cue�������Vq@��A���Qu��ê�2Bk�?I'�E������x-����|μ�R�3�0�Mb��N+H
,���;��6A�'�f���0�Z��T�~�p�_CU
��+h��G:,�D528�� �gϲ
G�
M.�T�f_� ���FJ��Ĝ>����)�A�/�Ph�k�ۇ_�b87dL��T�0��W��"���@u��yv���C��t�P�lW0�'pw-:�b)��E?�s:��.#4ϕ�R,,i)�b�#��39�b�ne����z�RP`�J����Ns��
��:�͆�p#��V�Ʒ��\K
G�S돏�4�p�e����po;�*yw̓�����O<��9�jX ���`e�A�b^�!DW�.D6B!���Fo��P�G�w�J�Mc f&cZ&��W�o|)��Q0��$~�N'��/�L��;2��j�=e�[�d?����&DO��yP�^���\m���9�dEH#��5����.
�jYpɃ'lnv�8�Ks��7W���}H�*�*|L��"�ګ��IZY���e�d ���T!�����Ԟ�?��P�{M�.! �*0�o�MFgɓ��T�e/��⭟�]�4�_��_�Fq)%�3�%����X�*?��Mtȡ!�5�S=�%�~ɚ�l�OZ�y*8qln
\Saa��{��F�ơ�"�1����!����U�AT��R�1��L%�;`1�hG�;��xjLa� �,����I�z��*B^��?�-�+@����š��u�T�9\R�Gpq�H q��~��Y_�[[�4�sh����A6_��$�Cg��M|�x���F� �~6 mn�&|��O��������w�r"un#�k� ��Nҩ�	��S�� �`:Ί�_$۞�$��ؓ�T���{����5�!���72�J�?��Y��}��9`��}�/`}y�%
�o+���Wj�Qy<��vkv1]�d'��;1�
�ޝ=J���F�uT�j@t���\9A8�s���G�!}-.'Tj37�<X~V�Y4$�u����=����jzE�{+ZS�r#���Y>�!�-��c�B ���W�~��N�PO��]�_M�6S�Ģ �g�;q�'�(�2��9=��M�H�1(4YNgK,¤	vSL4��_�+`M3=��;�{cx��]Y7
���$�S;V��"�;Z���	K�Y|��"��e�)rdYl��2Dz_2�m����G�]�4d�J�!�*�뼬Z�y |��P.�V�n���Ϫ􂱱�K��J���^��UK�����(W���#q�m�۫���b���5����9�D���?��l;�����XXn�5	R�j��@���,�?�^��`��G�v{�G:&��i�N�����M��`zOT���j�������F�xg�ӣ�O<�o�+w�d�C���M3�t��עՖ�2��O�
C��!�_1�u�͘�UN����=o��0�G�ZDL��İ�v.����{�'o���(2rQ��S4��
�H���0N�i�1)��6���E?fЂ'Ab�e�Ԋ|��T#��IŎ��}��b�H
A�>`}VG<�X�V^v�X_���p��'���h�<"�k��
a���.?P������R�LnK/�!�ƞ��ǘ	�J�\���nn��f�	nf9I (����&U�_Г��*�Vv�i��D+���p��m���\�n��2ba�\- w�Hh�����c�~�/]�K_�.�@w��&��N�\���?�wׯ�:��s���tcPn�wN�J8���WHTz?Z�V�&�c�jE>i��b���4�s��n��D�Q_��AvRi���0|�fƁ8V��0cG3\�sw^���rˆ��7���2�u�A%�,q�/��'Kc�Շ�i�?�
���g��E�J���X�!��G]����y�$�s@�2��Ф��m"��}W����M�dMX��F�� LG}g�أj�R�w`���6�Fv�u�<�n�SXL�_I�4�|Q6���^ծl�S��	�����	�!���� ���qX򻉯A�7���Lζ�>8a0�3#߲0�5���)?�\��{�W��NT7�+F����MP�m�6��Ȕ�gW5��ӎ!���q��u�C� w��ӨY�5����e���cyyЮ�Z� Fcr�2qVw���P��@HW�_�Oq���8����Tw�����[�����Qx���)J�p�dG �b�b!b��1w���v�ʡ�.C�Y�*ƥ�"�v�N�O��r݋�n[5TRx� l~�
�J<��7��p|p���7��0�0m�#����T|�A���/�����<*={Ggp�q�j��6��7B8����N����G[�7s���2��ޯ&��2T���:@O��44L�(d|��z֑'\���`�-/-��U����_h�z�Ekpp���D�ԗ{U����iK���|��a,����	;�S�������&3�~����W��$�i������mxi.�U�ʁ6��-"�	'~V�y��,�����zm3B���h�9$��Tج��+��e�^Z�L�ct�/���^��"a�>�0��)�gّQ�R�5�m���vl!�/��Jѯ,r�^i�?�U��:ԝ�\�P<���׾���䱶���H�F�ް/d�9��o�)7g]�}1',����%�ߝ�9�v�ؙ}��u����p͵�E����?����AF����g�a^?���"�����e0w��[�ݗ��5�F���7�B_���|)K��HIT@�La�h�Sq���q�҃_�8#�hq<P�d��R��B1�XK����|�=�j��@C���~���$��d%�{�)6���I���8.F	�SXu���U�����^��%��ˡ2Mi�o�-(55��� ڻ��ie�Ͳ��ʖE=c"5�yBp�2�M)_�����u����7?�����e������	��E砞)��JM{�pZu�CB�҄D����$8UL ������?.��!�Ξ`aߖ��)(���u ?��%��]������;�s�|���QƑ�N�֮�������Q�i�#��[���f��O��uö�s��TG��gF�6u���l�9����DH��ۧ2�6�¿9^� �QtiX���ET�v����J%ZJ�č$ޥ����r�Ϛ��7���A)���>�y��X�5�a�T*��N�Qև<�b�c+ᶝ���5��cD���B8�v2�q���<]�r#��+t��mN�~�fE;�|$_��a�H����1�WL�!7����O���¹ LNpQ(��4�b��ę�k��y-�>�Y" Z�����}Cx]�;@at�i���H���iL��>����Kщ����9|h��&�y�[����B9T!�>��eѯn���NW���8ΜP�7Ι8[���Ƌ�X�������*��f�3!�<y*Aϡ��vu�L���+���2�}�ꑥ|'���)=/�~��b����i���![�D��]�J"�갔�Y��_@9��(�F�1�eA�� ���P��}�?B�%2�NPm��hB;��	#�p]�衡�@�b���x�w�{�A�&���F�D��І�"?"�BF��2��ą��t,��H���Y���HC1TA���刄� �	��rnc0/7��I��p6Js�oN���Pد �T��� ��2��o��`�|���/�M����yL�{C��K�9�wB_>��_�*{���m4�7�L��A1dr��B�\���b;���g�ڀ~9+8��XN��@c�;��N-a����^�e�ڛ�Xnmӏyl)=��w�Sn�Ι��B���PK3@�,�Q�}Z*�y�:��L�?蹧`ԡ;%I��v�5���ja�*���R�M�l��+�����l#}%hg�Ba��&�+��9׃����X.��_�a'b�J����ΐ/_�X)潖��#nWܳZ�]�з	����)}��=��ɟ��3�Ӓb�[դ�la�eR6�
y�R�WdC�vA�E��f3e����w���
{� �i�_�4��%?%�w���a�y����	�# 	��2C,LvyJ_mx)���(=T6��O��9VHH!��L��p����slU�w!��^��]?c�	G(^���p8�qphy�$V���~�͡_���l5S'��;z�4L��]r�\z�$����^TF���p��ǁh�D�/��hnϪ���sBV�pj�B�C��-��{���G�V:�0���[�	I9�L0.�!��J���N�ૉ��O]����Z3GG+c �FF�Jmsp(>���P"���a_ۜ�hϚi˦V.��|i�u� ��Ã�O�I��C"��bK�\�&sb~�!��R�,{B ����p�Y <1V�N�{a:��= ���7��2��V�I���@�%�W��c���f�������EP)�!l'o1�N7�}b��Ag�k]��J���Ã����M ��zP>p����qq�.�4�37=�Q7Ԡ�JH�^��Y��b�j#q	�!L����m��&�`<�o:x5t Ä��;��S<���%}��x�k��m�1�]���:����1)�Ҹ� �O�".��{����(����@s'�(!+�U	��
S�dGK�'U6.S�é%�?�'�"_E�(���S,�eGs��̹��q�\�W�OK�����U4R�7�zUzQ@{���o׸A�R���\cH&��h�s�t�Z �E�^mSI�B�s�Dri� �\B�Lb��L���v˗IQtV����V+��8�/W���[�jiT�;�ܒ�T�/Wդ�.F��Û6����A(Qec���-�fG�Ao�N��ݽB����m'_���IH�ꡉ��� R7�3�R�q7��n :H��?���R�_-F�[��3��O��y�6W��5��\�S��fc<���.͂�#J`�*��;
-WB����I��p=�&��m-w��-�BO:��7���"��_(�O]��h���Sn��P�c���r���O�N
��m�	_?c̘��!�>hꎐ-�HIܩ�5��JB��})�#CZ�԰�EU�r�d��d
Z��If�^_ؔ,E"G0 ��fN,X��ӽ���ʗ"|IH�_-����_��;n�%�CB*����3?M�s�b��
ݜ��j�=}X�įV��� �����D�/���]D=w�#��&�ʻ:���=|�����EB}N����T�	��^���:��'�z\�j��=ԇq�@�s�(���j7"x��������
�ue�Ԉ��|*���IR& F�:�$�@%����A3�\^�Kx]1���A��e�����3U|[���W�`症�z�G�|���	k�X`���g�����2%��|I�=�'�����dE�?���O�0$wo�5�|�R��Wƹ����ª�h���a.S��1h�N�.luض煵uy�SJa
QE�i���ˉxE�-��xk"���+`o�����9�����M00�p�i�5Xi2Q���u���Wp:�z�RB&�K���+�t��r��D�d]hÞ�H���l���1�a<��~+Ќ�T}� kQ�-,�AJ�ަ2�^�a�Y�R�>w�<c�����/gĸ�L�6f�#WW��~�XU2ܦw����ښy��ި$ :r3����D���2ڔDh�nXK����"��t���P>?��e�? X[��S��jo>0*��y���o�S�ط���)tY���D�Tr�sUۀ�6���&�����R_�~�eLk��߻k�Z��ֳW�����8�/!:�v�Dr�Q�&�������j�ݽI����Z[��
�x�H8꣆�Z$�;M&��͇ZAS�Ht�jD��O��c���s�Ƣ��	Yj/+����jr��T
��`*�O�f��]�w�P%-��N�aMc:ծ&'��uz]{Ǘ��)�z�zB�
�6ɘ�z�N��v�`
��B��W�fĝ���K�Lk�~M+B3����-T����_��8�=�~����/q\ܥ��J|�Mݥ ����&^� �W}?!V���?&mR�4�R��A� ���Q�ݑ���CՇ�:�LmM@I�`��?rg�Z�q��!���w�@0�G}d���Ӳ��'xb�=�` ן̨/Y"0�EL�c�g ��)��X��߻> �Ua����p��PYJX/��e$r ��QC���ݑ�h���?J���d#z��-L�w<JrU36
��ՙ�|q��VҼY������:�C�x[�ċ�R4�ckH���'��x�Ҳ�vd�%d�&�f��,�G�~=-�%V�i�Md�p�O�ݥ��$�tƫ-}΀���� WC�H���
I�����g����fO���@���b�$�e�������pUg_���_z��t-
_�U�Q?#���-�_��)▍���ϋ4爹=^������\�]�\V'��"�
Q�l.� �O4�TIR�&�)BQ�m�¶+��������ai1/=��#2�^bQ��ɟf�e��ꪋ�L�0���#�^�;.�5Ke�W��f�fUt���#{� ,�@��Ezl��-l�����5����}�)Ư.�<����iv��m�uK� ��Y~��H�S��C2�({�a�;�c��b���8��q0f)ݖ���1
�V����VE�_�ŝr�"T�i3I�PGrx��%��`��FrŢ�}Kl���޲�X%��.��♶sd�;ةw^9� ����e
�� ����&,�7�*i��mPrAd�g��-�v�S��-�n����Sx��+�������i�v� ����{/����V|/U.A nU�7L��g�y]qF�i��䇻�!��x9D���JR��(��E��s��<
x�e9���������:RD��<���0\{�C���������C\�@�B���7�{�l�t��[�hn0喻ț�t3`�����'�4�W��a��d:<������,.n�(��gB�+������	��T{��h]#s{���[J��J��
3�SFA�@�y�E��~�YO@�봋	�V�q!�x^[��œR?+Q���\�US�k��J�P!b{�h30Ƒ*H�@ᬮ�q�tC�l�Y��'������iՕÉǨ�S;\����=aʁ��uw.���>�W���0�b���˄."T������l����O�g�Q� �
��#��FR���ь�cne^?$h�A��?D����)�6�l%��,93�D��Fp�dʩ6���w5T"�%���EL���]3s��M�6�r�I�l��-겖v�W=������kRY6ڭrc}j��X�5E�:(0���S�t�@,H�3���A�ڔ�=�H
�=�h��8�B&��u��8k	�
�(̱�u�gס������H{;xbg�ݜɿ`�2"���3���vI���lL����!��ć!2ʅ�Y��0�%�Գ�O��O��$\��h�3�x6mJ�خ�9��M�Ć, W�����:���p��Ld���We� V����R��)��A�ƽw.Ĉ��t���񃴇֍��)�l���-��1�������W7��qx(��"��N��{�)S�'R7E�p,�r���$��t ��;�rG��>$�f��7�|ƍ(�װ��K��q���'�&�2�"�V��/l�C@�X�������ֿK�n�rԿ�F��*����ߧж��E�y�)�)=�i5���,dBZe�/v�9C;�i�;a蘆����oisQ�4R/*�B��%+���拠{HY6p����/jڤ�Þ���y"��:�?���7���"�\�0@Z����R)��k���&����ip��FA�A1	�
C�E-{��O��j��C�U�R7�j��d� ��A�K8�����i�VsY�*uQ�=@@�0/ܢNd)뮾��R���D���-K��s���PU��:�Y��;~��5�� 7c���9�Z��r�}S�m��bq��I�4H>Sw��m�ll���9��n_G��yn���c;|
y+��O�
������}����4��h��	ǭ�	�S@(�J�5���[`P�a����¦jX�������̴��eC
�2�_���.����W���1�L��R�R`��~aR�5��;y�����v�`NuA )�
\tY��0��x�B�Փ�t�*��_F+T n���}�#��v��/h�{S��Vl˭���IБ�.�8o��wиl�(@��y��%��ȥjqC�K�}�?�V�c������2G�yN�a�Y12�؟]p0Pv�	�@�%��b�	3��.�ӣ��-��R��sd������5c����d-˨���*�J��-��}�bT�ok;9t��%{�N��tݚ���'R�A�����X���j���:�E�rÁ�uyzJ�g��:q2汞Ю��Y�`}ʀ���9"�'�\![�07�����L�o4��؇�ا#��9�X����ձ�}�*�+b��؄:_Y�Z�N���3L��Sg��)�����q�	�:�ω���XfP���3�}܊Z��v�˙PzL#F���|�9	n��G��G�Ք�ݩ���Ut�l�wi�D�+�l{MJL
�3a���iO�+�U�ouE|�.!���@�r��#��D�2�I�n��ݶޥiK-y3	v����+���2���(�ۄ�+�������W��>�aXz1�8Ԯj|�t�)��<=� �T�����d���M.N�*
U����1�5iʈ��	y�.�m�n081��/5�Djh�����# e&�qT�T��9ꚫ�HlaB0�b�B�eU�,��!s��/s��Ȋ�%�X�$"8i�{�'����~��������&UG����;�Q̉�K$"P�]w�U���2����zѲRK���ӭV��c"P�Ҵ@vM�bU�]��PS1gyD�M	��짔����Q><��>����y1���AM�ʓ�U4n������l�z���^��d�g�pP�/�>Pe�-�f�����eMUε{8�	qac#��m����~b�r�K�
Y{E�T������=a0ECL��ep���9���s�5Db���{u����azw�|���(�J��F��
>yJ���-"���	`[Oq�@Q�:u�.lu|4��L�)�#��bU"�z��( ���9�D�=��WcaΖ���x�.�*��	D2r�#	<��EɃ�0!0,��s^��X?�h.p��"�8�0-�a�$�*q�Gt��@���pv���yJM�M8",�B�E����;��~7��2!�(�p5�>��m�����x.)���"o�X��t��T�)A��\�̷�1�s��<~��IZ��O�ȯ����<Ȉ?#�J7���[.lw?y͗H^�oH{+���H����{��E�@��wH�h?i�j��q�B7`;�=n���C:��u�Aܮ���4���Lf~����:�9�HSK�}C�Vyi���4y��>�ŧ��p���04�_���yji}���khk�DXd�G`��Ff�~�{�Υ���8�����e<�F�b�hP�Pj�A� '_')'7tÊ���p;x#�:g�+-W�yOG2�cb�]�6�IS����Z�_4�H��)|^�3�x���N����	�$9�`o_US����)�B�ɵq:���-�j�Eu�{�=y�k�F-Rd~���~�kx�OGŗ��$(����!�rrI�!{,�[w�&�J_�
TҤ���z�c�}�?l�׈�Д�7:o��G�Z�QAg�x3�n�m�#WH�]��2)"������㠬�g��p�b<����W���">�X���Q�ގ�#��>)������a)R��]`�c�9F�BJ��t�<l�ڄT�M������8�w� �.N�+c�U�T�0�5�������35�Lb�n(+X�橞��.���Y���vHf H�������)$�K33��Nϼ���|طiG�Vt�3tEC�0���?D�Ρ�e���m�}|�b*B��YDm������J<��~�&���9㢘�CwE��:��C�;q�.�O�U&���;����I�H��'g���_���_�p�]�����nn��n	��4��	�G�&/����HNo�U�<\�W�p�6z�&�f֥_��(�-i�0%��[��$Rwg�A�H�g^Kp�M��΍�!?/g��] Y"l����OrqF����a�Y��{��Ĉr1����G���S�v�ꯒ4Q�Q���1|J�w/醓�.�>��t�eu��(��#4�~�������s0�:f�@�W�.��gq���&cL�[n�|;�\��v��6����V>ڞ.2SK�un]Z<GKYE �)/�\�+Q���3�v���Z���s��*"�Y����1<�B�Q�s�ʐ��GGtw��>�����D�w�k���u�'I��H�A/{��/L�2=bx�� ���/���se�^����'
��F='��� Ɣ�t�h�D��c���DK�y��3� c9�R[i5�Y{0'}|���G��p{FՃ�\�IO�}���/�8�����O.y�j/����7��K�6ӧKc��M�O7򘙸�ѷ����ɐ7��ϡg�J�~�Vr�'%Y�j��t����nm��l���VY��xߴ��wa���Q����z���X�bE�&1��%v�Ѵ>���z!�E<�����'�7�.��o�:�|�2�7�N3�u�OwX�!`&8 �Er�P�)}�-rY_� ��̈�^�7�{�
�<<5�Yx��Y�Tw�3���HS���/��4!�p��93�K_��#��$h�?�1�X���}dc	����BpuyąB�\9�T}B��uw�Ԯ����g;x=� �[� �0 XW'6�0D� \�����_�)����Ĩ���ż=��ZRV9 ���|LgP(&��|ָ;�]=s����&CS���x�V;�c�����2�nN�\ez|APu���FF��{��A���F7̼iʾ���Dͱ�	 ��L���"�%��y�,���BV�Bo��k�Ӥ�kS�h2�֐6�G���3H}��`'�໼s̯�z��6�<��H���"��V��*�͈��q/�8^:�q�;�M���ֲ�*�~�m���>���M�iv�>�~���r��5�	����j!!fIS�I)��0%_Hzd�1tBo(i��g��=�:@��]��oV���\)�����`D� ���U��͌��ث��h��+��&�]L�����::��&��ʹ.��s�ˏO�,��r><�T��\��m��q�]J�/ڐHi,!j���j&\�V	�r��n�1��KM腍،�<X���fw�y��*ᘴ	��;_������7�g	�D���4}ȸ����v�~Bȵ�m��*�r�*����D*e�7[c��v�BQ�z�
��>���l?k��pt-AsC�vA\ϡ^ڹ\�r<���D���"<��'����N�)zE��u�ke�
�;�o��y���{r7�v�5k��2]�LB��1)�'�����_'ZlNJ�0�֬�F�s\���è����?��gƫ��g��+R�m�F|�}w &�r�b)I0;�8�Y�t��y�6n�o ���Z�f%$��X0��R(��FSQ�
k�\ ���B#>�V���g:������T�nM�y�0�j�y���u��o�M��3/R�>{������N׋8�\��w��
�/�?y9N�+I�f�H��`-JT1��:t�2���eћ�p�H�0�6�§�Y�>�Y�>�N�������[)�]?��?�x��-������zf�8"����}a/�:����b쥿aP+�&G�����Bm{%(H��;	x��}��������)h~웷3�_D�w�o%s��ܔ�����6�O��^�>�II��D��4 �i���Op�Ymg������J��O��AY|�n{�<��ʉH�=��fU�o�YH2��kr���>r�HQ����0T!0��R����+MpJ	�����HNK�D�U��sC���F�G>�n���P���{�f`e統��S��[Ȣ@�o�j�"I~�NL5����Y�NYSR�F�oӪ�O x��!��ኾ����ⶑU���Ω�.�:I�ʋ���%���(ࡵg܃�{G}�t����*/J��o��B��w���˿��U@�$E5�����\�+�o�����ظG��翽�0��c0o0!N�Դ�3q/uT�:��U���C��{��en0[(
F�]դl�H�Fm�}>L�aLw��
��Ѫb����-�k������Kɯk��j+>>v�}IE� ���N<��cn$��;��3
�}��?�]}h>`&A��&j�1�=x� ������Op! �ԥ&������k
����d��7���O�����T��B8�z�G޲
�	w_Lw�_�5%�
0�.�OZ)?[#�q�Yڞ3��|!P�}�������[_:��`��$Ôs�=�7��3� ��7�C��`BTD�<J��5!��lj�5&�WJ]��60�P*��,%����9R�懬)��'���60Zkt-��61½��Ç������N�!�������}<Z�j��2�P�Z�����&�&��j��H�����J ���K
�.�A���!)��D ��[<��U��N�:3#Θ�V�����s�mM��r�x
�S�7!���tgqD�.&|��jv�6���[�%�#�8�I�`�o��|�p�s��l���x�O��sPX~�X&�}�L����,_%^�m�=O��b+���~���{̩�(�$#S�؇�5�]��`"�(����
j�9���VR����a�M�V���G�M6>u�4��}��J�y�̳��I�v������7B���g̚M��iK�Y���w����Ea��e
=)s!�I�C��ɫ�0I������+J�f{�	a�ӝR��-
u��I;h�8�	�7�հ�"Np����9�e����':w�[�aQ=�I��(�wb,�FU��@��ء��~!!�Q0��в��HfPa�:��y*��fS���+��f���p�]�C��{x�����ώh�RJ����̳�̥�L�
�]2����2s��P끋R��r�s�g�|z-��-F=�]6�}�����|�橆CE�.�tu�O���[�4�zm����XWDY���f-��∲�R��!ᧀ'�{�t�\�i�I�Q��N߱'r2�,NBC~����x��`��U�rH�9KO1F�`����iŞ�)�1��zC:��l�I�˞�$� �#���g:v�I���c��h^3G�ff��N�%@&�����O��n�RҾ�X:�|z7�<WNf��;p����

I�9J���h�A�/kɤ�MA���Ĕ�o&��]bo�gm�����v���Ԭ�đWO&�1� ���3Y��z?��A�O�̅P���t�X��:t�����v0�3��2���j^�/'x0�M�3��D�d ��4� Օ����,J����Q�nͤU2�I��]gT��MG@ʄ�j�Qa. ���W���Y�ls!�`��q1/�<'
X���}xLEw��෶MՐ�
��`���U�0��<�M ���aq�E�S���,����X4��%�������t�w*� �jQbO@�� �%�� :%p<&_�D��B��.M4ud)�i;.p�x��%������k��C�z�qU�>쵚v<��/N�C�g�"�#6}[�������+6t�}�(���f3�`S4�"_;؛4&ݥ�������,��7�Z��7M� �ġ@G$�g>�������b]`�ñq�D�r�ǆw��S�"4���@���u,���4��B^���*"�����@9��R�[�FA��.��.�=FK�����MjUM�Խ�d�m�'G�|�ʵo/��+:2��EQ.��m��hK��#��"J�
�5����R��Q����I�;�����)V@^1ieYk�/
q�0����5��1�q�618�N��!�q׈�-�1���,�|Z�D1����Qj9�9't)�}��Vw���Ρ,9|���-�t5�\�d^+�����σ�Ԟ;@�O��k}��o/�|�rϰ���>�Ϊ_����C� ��g�,�K5>�����g]�WY���⑐���e�S36��0mS��C�N��;�τ=�j	�}��xR�R���A%'�K��tj>�$İ��@�R>�q6��{�6uh��e�B��٘�ߵ2*���Ll?���tgȞ�X�b@�ꝿ��hlȰ��_�����綾�)���ހ����o�9P�-����qO�����_�D����z`'0��V����dcmT�ۺ�$Vpg��mt�0ɶ>���`$-�z趠��p7�E��_���\�>��J��1�5����,V�(5}��:'�ï�}�Ǘ�<�j7n�_���[�1�
I嗾�֬}�����#�ƻ�>�l)0?��S92wd�6��^�|G;���S��Fc��hF.�U�q�l�C���C�S|�?Fk��n��'n��h"@V1��~2�/�	���fs(h���As�@.&A�n��cP�0�~F��n���f5u ������-�w��@3q���>�o�.(�ֵ��Vǔ��tE�gX�08�Fh�:)0�W��5Q�vc?0CK&��n�G�YZh�X�d|�=W46"��F������0tΝ�Y��5��H`�{�@^�N�:���f�L� �(5��;p����O�kq�[;�4('X��!�^��������ҸY ���`|�����o�����n��a��DΉr1m��|��"0�/a��l���;����޷��}��q�3��x�Ȁ���4�but�,�X�����5�]�f1���v�B����=�
t�RQf��좟��x�Z�/����|Z��e�j�smu��w�~�$3�?�M���F�"91﫡�Zcb��*������	_���Ř$���rN|0e��{��Tj��(N�ʀ��g����ӽ�)�vl:�>�lw>����
��ﺯM�] .�8�
�Zz��n ��J��P(����J���Sj*��,D��+s	��<jI�I�u���6�~��/hF0�yν.�/ �?��cP ��|T��`N��߼��� �פ�m�U+�V�D	gA)�]��B�ӱ+���~�=�ѐꛤ"�D^�Փ�6������N�!�q]��EL���=�~Ţ�j�5C������T]UQL�Y�]aT��Z�����*׮K�O�n'����x����n�{Agm^��A9�K\[���I���������*%�i�~��[��s@�{Rؚ�SrM"L�GD��:�5��9$�7 wV�������
݌nJ+Cv��Q������PX��q�i�_��B3��e@��ʱ!@�2U��Pծ�~��0�K^��`Y���D�z_Re�W唺Q2�O��--B>
꧍�[K	���h�.1g.���|FLYHeTO�1L���qT��˹�J���gTBh�>9 e�����q��C��60ެ��2V��Ҥ�7���<�?Yt����ڐ�T�擤�V$�i�hn�����Lp�+�仚r�K/�W��{�핱�di��B���w
�Cj6]�=��Ջ\����]Ң���2�����8>���������s���<'���wdT�H0��PslC�����鳲��Rc����$�l�k�,�8�����*�4{g|�����ͅ1��k��� �t;�v[ޜU̧��|2)���T�w�%��e4=I���i���, ��Bg���+�H���MEo:k�(�.����`eת��tHy�OÅ�G`���ѳ�~"9Ǭ�` ��\(?`7� 4
e_�~GN�*�����(C��I��	�ʫ�jR��b���W�WO�>6jf�'G����u�'dWb�[#x���K���-��--�	Zf��vx�|�d��\O�K�g��lv"�zJ���۝�y�=I� �K0 �V%�/���`��?0V"L\�j׷m(b]k�9�1��fBi�Y A\yJ!I��컛���L޿04�Q��I���Z~��=o�Z�#��ɗ=��QyI{YuI����ߕ���Y@�!j���z��%�ž��N-n��=�8��\�8~/c�+��K��'̓WbJi89���(���а���n��&~��������G����ر�,P�lv%7��?(��P+���:J���*>ه�V��v[�>�|M���s�nP뢬�PԄz��}�H����on!�`����v�*OŤ$&�ڢƚ��:�X����W'�4����3(!�s�H=�HǦq:洣�@(PW�G:>��V�V�P9+?�]������p��HZ�cI�e��v<�ЍWG�q�#Pr�L-o�6�>{������6���by'��� La�+Hi�2n��c��;Wƫ�O�W>���1~�Z0H���A�Q4�{��}�W��䉦Sm�_��ׅ��bF�^ź�[�+6���@Q������G��t%§�h��L����K	q���v8p����9I%\�<bBcyc0\��al�f�H�ٮ�aU\��4���=E�C�ݢp�z#�h��{�E̢;���`�#�?ޓ�6dQ�k�aUM�Ӫ[�Q���Kl��m;`FM�n��I4�9����z��x7���u�b}%2m:�hE����]�x>F����,�#Q��O�z̩�m=ͬ��������B�
�����~J�i۔!+J?H����V�}����#�!�tQ���?A�a���|��uP�5�,���l7q�5���0E��X��*�����~�Pe��̞Z�
���"�,@D��]؞`i,�E��/�;d���_Y��D�9~�{�z�n��<9�[�����A�T�6{l���H?3H+}"6Fz�v��0�'��H�?�6K��"w-M'��IO���80�;��חʟb� ���vt�_�?O;�m�B�AE�̔��V� ݋�� �bD���|���hmcJ;�3sR����]�"9��	p�9]6�yŹ�s���?�<��,�{(f}U�F@~r�@���g�>���F1�Z���qŽ0\[P6�������g�����e݅�ko�C���h5W�t�u����/a��O3��{���7����D���?�)�����o�E^4ڭ�K\7��9�|\��X�X��,��fHnԿw��>��Q�PM�����uj��~��������ڬ�~���"h9�p��4���>��w� A�ammS�(�����Z�o�b�]Kyi�d�Vڎ��r��<j����"�J5w�̾n�<�tp�~�����g��o{���gP�_��2E��n1�>|�n=������: ��Q\K,X�jK&����������e���.q������-B�&?zk�)�ˬ�������Tgm��b��L�)!@�ە*(��}��Q�ՎY����Z�r=o��C�i�z���<�m�!k���|ڌ�{m�;���LHF�H:1ʃ6�����;5�Lg���ţ�&��?�.�3vo��ݭ��<�p�f�v������9��vA�n���9uE��Ү?�^:K"�7�P�ɸ�\ٍ
ͮWa�4S �Ž\�з�j[��	 �+i�MÜ��ɧ$���p+�c���iAh��� V�����ٱ'�p�ҲJ(�� O��;��>!��у����W��Q�L�x��p��:�V���ܮ�/<�(�ɗjs(�%G����3]E�gT~�GU)��I�}������~��guz�6�Y��V���ޚdQ��*3�%����*����ј���u*�C�'c`!b�̰7��`��G_�[��ԩ��7�&�F�gt��A��Dz:BŃې���!.�b��1$���An!j�8i�$´*7�|+�3pc������_}D�m����G�<n���GvqP�K������9�Q�A�;��>�_\��h#JL_�(S0+� mE�n�4l��X1�2P:*�t�TK����A_���g���{2�̝y��P;�q�wF��G����S��4BW^�ή����{ғ�QFA�W�QO��h�ϕ�U�QZ���|G0}��N� .��P�]�z��r�m�#��
�M2W>����������c�:!o��K���v%&���A	���?O��F���/����ɿ��-K)`.��Q�f+��h��ܡ5V��_ȉckmڮ2�y����-�c
� i��u� 2f�tgO�BQ�P�@���F��
o.;I���ڋww��)	O��Ή�P-a�k�3h�����"��Bb�����T��w!k�!g�JM쭸0u8��%�^d^��W#
9��xıJ	��`"�3����Ӊ$��f�f,΄���Q�������^"�xO�l��j����y�}R���T�o�6����L[d>ED5���i�+��j �j�4*�R!�4z�L������%T�V��Dl u�Lr�}s|��� ˭� � I,�}�A�|Oc��Z�1?�	v�:MD�L�^G���,�X�,�0f�����p%(�z��:�g����ޏF�������u{� �������{�<�P��V@P4r�wj�sP�w�����o��8\T
��˽�a'-2���5:T�=`D?Qyl���0u�ܞi�3HcVA3��e�W:�mK���'E����R_��k�VK�8��7䆁��ׁ�0�;�x���o��?A!�q��F�BD���hYw�� ��>�J���\O|�C�|N��!�B��=���N��)��ɭP<����d�΀�si'�0�9�ƅ��ag�DR�s�:�$�G迵��; ߫��7 �B�|V����ϛ��f����[�"^A��ô���(��z.;]�.�H����?uI��Os�(�$������F��HB2�ׁ�~��!e.����/,�Jw�v1"�ze��lX-'�8�3εNy.?�%]�5�^t�+��>h�w�N����l24Q�$�B����8l";�v��d�U~4n}��ؓN��i8�h�|��'��7���e)����#Q�N��E�8��}���r~����?��נ� z�^L�n�j��t�Q�Йs�lǠ
hQ���z��dqx�D�DI��,���A���h�hd
g��n՛��5
(�!n��%�$�va���)�?}w岅�+�A���L/���{z_o��rS���kD�k�1+�.���NS�ĮB�S�-��e8��:b�g�p[�mI_�
�%���5ԛ#�!�-1���^""Jm4���Z��9J�*a��]�8��6��6�$^�I����ۖ:� ��8e�y+��e��Yz��
�@�^�������V_��T��.���J�*Q���y�/��An<=F2R��y�Ug�l�P�T^f1U�l$,�F?�Vdhk��Y���J���]�|&?&�~���kʍ�K��([7���b5N�%���z�
w{t��9z�O�z�g�7xN�e��%@hb�F�y�^崀�&��=����2p�.�n:ΟjzãL�e"r���,�V����'v��N��#����W���w����+��}f��ٽv�Ke
�h S����8���>�w2��i��~yN�F&^�^�S�,ı��w��|L���($:wՕ��DFRw���|���{�������J�D^�y��Bp-���bL�d����!��ii��:���:b�CG�(�6R�~�*�;��2�vąEh�ohŰ�2�}�9qσ�	*��2/`�M%��>��e^tLѓ�P����C�MB��ra^�֧7H�!w�Mv��&yh�浏#�u
�ϑ����$��Bb�4�+='�x�/"X�oD�\�[Z�0�8�jvFQ�[���G=�&��rm�3 l�����ɻdpa�-㆟R�y4KP��$I $��]�]�8�֝�I6F�^h�Z�����4F�& �(���g���t�Z�	�K9g`��F?
��o�z+�C�ēm���/���-��m����B�����f��T�.���d�l�Mb��O�������yn�q�c;�mŪ�0��' ���B؞� �ҕE߷yXF��d������4q�q��)pr6����
<�uq2hc��j����|�.f�
7�z�ÃD�=���VV70=�E7C���Q�\�Y�R���ι������N��|���B�I��8%Hgc��Qf�؇��*O��+�v�3�;�c�k��S7
r��tXr��7,� �_tptS���b忠�����1=�QI���ØC���w]KB�'s5hW�Ε\�)�Fe%}R�K� �o�lbL��п>_�y�&c�&Y�$:������e����O���ИrS�헪j9�b��C�㔩b�|�Q`S�*��fN��&���5hB�E"{iގ�6#���N�	���h1#��ѣ���M�k�`�K7��"n���X�����g��V��UGW��R�G����g!*F�'���
*'�<�c��L'�WX�6� ���8=�i�.��s���� ��j��$��M� >f���+��r94���+�v����2��3��u�5��,] ��h��+���(+7ub
��m�ca{�ȕ�2S��.���#|����^�~�`?�8r`�Pc_H�HE3V�ԏ�sd�B=sڹQ[��������^E����>����p��(���X��I�M��L,�OD�0�Z����B�����!0��ǰ}Tw޸�\����_dJ8����g�ǥ���qx�Im�"K�܅�?�KTc��Z3��{��Ǫ}Ϯ�%r�t�Ճ�z���ְ7�gJ�e�=�P� �����b���o2 �t�2Brv?��R3_ԕB�p�拹x�;�M�η�u��yՠ����f�C�������F��� �=07(�g�=қ\���I�!Q��Eu� �!oT�	&hU�G�V�7���N�9��s[��f�Խۊ�ۛ�+��x����ݒRqu!�������jr��������� ��"mgh?�m-Po'
�F<�4I�	�-d�7����h�gv�&���2A��6�>�z���{��KS�D{�����l!Dkr}k$��Yh�O2!f-9x �Lr�i�[	��8�����U�؂H��o]�={�We�y����"�팵�%��HB8� ����N%¹m��Kr`�H2����D��U���vN���/�	�Ԑ�Ue�S��-�<I�U���^�6��G�4�����Jb��t��u�G߶�_�y�w�dU���\�N$�J����[�P|�V]+� �t�l~��.�� �2�r����A�j{���:��K��c5�>�J�Z0D}�	�Pմn�/~k��&|�c+]���F<�Ԛ)�ש�h��|�/���Q_�υc>[�m� �
��p�$�[�q�ۆ�6fQF#���0�����<�M��D���.Va(a'�#��L�O�ߤ?ww4���;h��?RT�n��X��@6��)z=��N�R}c��߸��g��"]RF(#�eY!��X�Հ@5�n�ֻݦ����Pg�a�ezʥ��r�Yb��5$�:�K��6l�X�R�h��\�ϥ08�� '�	�j�������xP(-ю_������b��<hT�����W�`����Z���D�n�������2` �͜_.u2���BO���н-��sS5� �\�봉�bȷ��#��Z���Eb+wW):�j��n(]��|W�+5�:DdQ��.�[����a���P2�Id-XV֫9��sD�h~X���������6�M����K�[`A�^ۆQ��l�F��W����,Ĥ�� T~���«�n��.U�(d�����*ẸXV��(�Y�����*��tniW¬L�uy�ͮ��7C�-�$�FU����Ĕk�8d
��Q_:C]<�/b�ˣ�S�Ȋ	򧲵��@s.ݐV�0�΁�3ـ�^�B7;`�e�-�̘ ����chS�wP����-&Z4�h"�N��^@�>��Ї\��?���c/i`U���HCd��Ŏ�B� �f�z9B�@T�!���H�I���j q���T�_y�>�7�������9��T�ʚ��k{jk��E���-�Yצ���u��̿t�����8?�p��>��SU���^-�0�y�R6�F��QӰ����o|�WU�8�1UE��Es3�6��9�o����z�T�7w1B�Ͽ|�07]�Vי�/���/�{{ ��ry"
���
=����x�I�w����C� �ܕa�N�qLV��e�]
��C�t?�B'�΁՛���O'B�Y�}n�8���P"7������ǃ�����)q�-�@d6t3ư���\͖�"���# L*��fI�z�R>z6q+�ۤƫW_b6���ǖ	�����N�����׿i�<��V%K�ER��,Q˧E�e��]�P[���lLPc�V8
8�:�� P�l~�}=�`��K���#���Md2�6�Q������|+&$�:����N�2�"w�@}�Z.�8R΁"�`ֵ(�Y�)y��p�i-�(�j��8�XDvº��JjX
l��!<�4s�pp^��6;�b'*Y�wV&/Q��Z�Uq���}�M0�]�k����R��]E��W�r�yO"r �CH��4ѭͦAn9��K�JH1)�aއ/��C�D��C̷H��/
���5"��f@5�71u�G|�E�m��]БAI	*mAY}�#���WN�ن�1�ۡ�eVQ�L�'�\���.$��&��0JN)��lΜ���N�5��7h�fR4��	��aD�%�882���Қ4nOG,����(� !.T����˱l"��;�j3*ܘU�	�y�m��BK���䭇���sл$���R�d��|��!�V����C�l�vZ�,�/ﴐ��Ȁ!�i*Џm���	��a𱽭l��Gᇂ���ｙ�U���B%����	�I;x�Q`�n�۷dȢ������3���/���5,5�Y0T"r���TO�=��jqpB��O�g :4Y�}��ft�!����1�NM�E�^g��G��e�"�w�,7���A�q�͎e���������W�Imh�}J���L�M�ƨ/��nO!�w��C�_'k��]����Vx�u����6z����c�<�5��Z����~���/(q� �ǳ����2�J��d�~��xo~.v�gR΃���_�����τ�$����)�UHv�!�!D��/]��$4Ht�Vi��U?����l�	�_F�3]�5	,U<,�R���y7γ�
�ԋ�[�V:���q��#x~�!�v3�@;�K�ܴ��׉�'ہ�ߛ��QO�v��>C����R��0�kFB���F,��Ce��ɩWX��:�\S�X~p��d���d�2�8�l����D+&�c#�Zu�N�l���=��H"`������8��&9��������.�P�Z)}�`۩,��(�M*�g�.;���ץ�U���/��b����T��"�_|�v�Ho�^s��p��B0$�G��䊜�/�ce�����A"4b�`a��i�����/�#D́�H�ಳhnx�C#�������'+�u�~�D<��l?z,���@��㞝�J��u����B���G���5I�]�Z�+X�*����e[����Ns�Go���Үr�������+�D@k�A�v��/�f�dh%VPh3>��rػ/� b�Gu+^XR
�VI�3+�?�̡�5�X�e0��rm�U'���8���!�]�uB��W�	�����{R�7�B_[֝�r+"�;z*���3G�2�y�� �V^����$����S�Ȉn���&L��,C1��΍��Ix�m�� ���| wD�>��֊�;�͕4�I�h�ޢ�a�Nc�����ե��U�4V)ze���B�W%0/3>�;�"�+0J�n5<�BCl�{rL?�����c5�Yy�o.�5#"fc�4W"�Ma|��բsCO����}TuQ���� 
Zn�w�5��(�Ạ�/	����,A�����T���X��f��|��_[91ORy���>��:��3�\3g�59�[pI��NX�)Y����qMIaV������+3����P�ۺ=�5�(�B�aC$v*N��G��D�F�qJ�T��TB*��u�g�僿��re'�_��P��jy��6��R�	��M����o@l.c�����
T�th��s�s1��;�0k2[_�"�6*�d���e� 4��n7�b�{�N�	���-rb�{6����=�Qs���Hl�'���gh���H`r��J��R�w������k�ip����1!�d3=U�^%d��b]��w��7�>>�����c��G���Ȩ�����of#�e��Av�R����
�*[�s�ѧ����i�27E���%�8�����;}�8���B����Jƨ��\�e�~ك]/Z�tC[X.R1��vr/�3�m��eߑW+�fn=���q��]��a������8Ƅ3�Oo�ɓ@V��{�M�0z���I�o�W�Fٵ��8���;T�s�f�~rbs	Q�Td�e�M}Dp�vU�a�+�����Ȑ'{	�RU0l9E����#8�#�{�A���?���O���s���hE�#���	� ��y��h���S�7-�v޾�f�x4���,qͅ��=*�a���Կ�t��@����y�~�A�zt��1��2r���i 4(�0�dh,m��Nx,���T�E\}��iu&ÞA#�h������� �z���F�,P-g?D�l\!	R��.��<�7�I)h¼�~�"��]�rW�9kS�^�>�8J��\EK��=�(JK���A,���/� ����"���b�.^��2��B���l�I�#i\�k���o���/<��j6�E�sc��ۿd2�B���#}��Y2#9� ���Z.p�~�I�E����<i��<�t�$;XƠ� �JB�8��Q��Pæ��6l����g���n�%���=�.���,��[��~3S��PU��*�V�γ�G�(�XA�|w�� �m�\_+b�_�-���Ԉ�-�^� q�(%�݄)����w������?$?f㼾���		�T	�	��/Db�dm������p��냵p��;���a�ڿc��l�?��[c�=zGbsc�1�T��̻���2�Rm����;�e��6p>���=�����V��*�J6��C�N����!�sn"Ӏ �H�+�z*;��{�k��N:`�U��sH���t���|�34�kei�^y�$ݛ���&�g��^3m���s5%}�����(�:�q�I��${���.E������t_�����?�>�%,��L+�淋�d(�*ݼ3B"�̐��s�r����TU���>cT��FJ�e��Aˡ���ȟ��4c%�1cr'�$ZK���ґ��͐>Ͱ@!t6˺R1�-X�Iŗ�2�kkmh�4f�"V��p��:����Tm���e
��I�-G�	���X�qK`�(�&�8�v�ܪ��� ��g�5�P�����<MVf�T�]K�ѝ�YD>0�B��_|�I\M�P���֠
���8˺�&���i�4�i�aC�	��c�-��f;���	�p���c����d�;<S����[�9����������nsZ#���>�z��a-nc}�{Um+|�Y���T�)-Ѱ���C?��rBN�Ae��
�(�xi�(miu\�d��ݮ�� *��{�Pu�~L�,���(�D�ǹx�el[|0�$�7�0R&�Ъ��@�'�i���|t��߆�?|�d��R��TWZY���z'������dG���K��1o���(���7��d �"\�h\sF�$�}�0�����y 8W���k�x�v�o�&s�=��W
u�� ���$>s�NB��i\s.�#oit�_H��[c����X�>|�[�ȴ��9�U�t�)Lq������T�ɵ������HX-&��C��!'\&O�����x�qP`�%_ ͣ���Kl���d�#*��A���(��wᔚa��s&A��ͅ#�o������qƛ����%p8�MaU���:�`�g=g���&W׹�<i��xP'D
)CV���{Bu�޲[�L����H�D��w�6ze`��1�9rI(5��Z1!Պ��ܾp(�,��Fl�����$x�PT`GuR;���"o�dHAD�;��s&�ۇ;�p�!��q�;]�7 �$���n�����t�2�4�8�q}��;�'2�Ct��Ye��]-�6���P�P�U'h�2�Bf�Ʒ����g p1�d4--9j�`�~C���<�<@Y�
��74&@#>�U"f�;��a���]�}���e�\�E&���5��q��2�òD�� ��ts�A��Ni*f���_�Ei#
��(���z��4���t��=��M'f?8���y)�C8w�E����r���d;G�F�><On�`�%1.���Q��N��ӫb���\�{��F�Y���	]���OU�M�m{F	Y<�[�W�3.o����췉�j��*���k��q��A�x�ó����9�2����2a��!�xL>nud|s��א��0`�T̈́j!�rʾn{�ٰe^.FO,7�!�m��ʫ�Y�L��U�}X��^���kB0j�[�����5R��UU�F�%��Dd��t�U+�,��O����.-����
��%�uF��^5�H��.� P�(#xN��ܜNuϗ�ې�idB�6<	��Β6�r�RA�f�*}$"~_b�a�Q� �fW�\�/��T=ța8����lxj�PiL�6Ɓ�dM��eT� ���J���t�0$*y��U<��O���bL�S�T}\��Or��Ç���刊/})�%��q6a��F~���#o��%Ng�;����D�ԅ���L��g#Jkh Њ/�L(">E��}.�i�a�6�0v�
��H��O4�'~a�������<��:�Dt��O��/�����s��Ve��-����jo�W8��p�a���@��eKeދ�iз��n��Nk�ef?�)�W���G��+�u.r�x_Ʊ�XOC
8�je9�\zG�+�CkQ�`I����{�;�oi�4�ʅ��-~��MS��?T���s��c9{R��O�����E��
BUW�Wr#e[�ETA����^�%�=�"wka:�o��b|��$dH��F�-
����,|2j��Fl�J��,�������6� �}M}9�C�(3�P:4c��R�|: ��Gg8��q?��f�\vJO'��1��5�$�;�X��c��R1�`�"M�zs.�vUR�9�p@�W �<6b�b�����J��Jkty�A�1m��Vڎ*[�nn��:��&U��P�� ��4�kq��:^@���V鼌��ݝï«p-y�ja�W���I�����o�)��f��]]I-B$'!���`Â"]-w(���㰀�n�S�:�r5E+���kW��/eVV�]r�qb�S�1�Q�w�R���t0��&x�TM'CT��ٟ�(����W`1��E6����U�)9�t�;��f�[!P�Xå��f�(��<q��la'��r+���k|�
��;3$��`mc6܉�Y�$&�V/����0�"��V���Ы����/��+�8Oa���n�ncb'��n�0���ːj�D� >u����JR���������+!|�핤@�"�9%y����Lk4w�xΏ1R��X2ŔJ��k�̿��y ���j�nf���s%'����]���y"G]oW�PeqՐ~����x�(G_�9\��ꧠ�D���o����+>�.
�����ڟ\Б�Y_ �/,Z$��=�v	d����=g��,�bh`ź�y�=�'�k9���g'�B S�V	T���S@2Zg|��B.0��2B�����)�twe�ŷ��k�M��W�c��f��8�6-�S�H�	:g��,m�����~��BF�}��f2	�J�����n>��%;d\	t;@?!*A�ſ��QB�d�%J܋���c���Ӫyy��H�uT28���Ƙ�}y=0�X��K%�;��!�%Nߋd>��;>y�,��yт[��Z��ܝ��d��WhT�`$aCU���1b
�����^P����3]��r�J+�z��g�|{:cB�`���$*{
�����"�}c�������ʱ����ɣX9�,���]z��	���W)X����1|ɠE�E�:8P��f��k�Ƚ(ԬT�޸�M���yB�����e\6wId4�S�޲����6L�Yn���R�o������`������S����>%"�-t����&��"����[��ِ���M����З�V���M��������H��\�����M�Pƨ����v">���NBeG������)�Uy reȲ�+����G��6���a��8ڒ�q�6PZ�Et�1�ޣg�ɗ֫�5W��Cm�Gr&}+5�R���,Ki�+�+[�`YF^VS����B������|f=����O�}�d2_5�c��l�{!��b�o��]�m�ۃVy�\��9yg�_��Ⱜ��,s��~2у>�#J
ı��µ�^-E�*����z\���3�x�z�9�X�9�n�{+ރ71-�.5�Ф�����m@-� ��F���Q,�MS5��oc�P�{+����=�o,����+��J�Ri�%-����Jx�O�p����8�����%��=��Ǳ~Em�����?VL)�P��|7��{6��1�������F/)�\��_n�,o�{t�r!��n$������5}� �Z�R'r�ɟ�s�e�����}�~�i����|���}����YKn�z�J]ǨG�AMQT���'���c
�/��Zq��YA��C�l@N�M4��a�D����?H8��Q2N���pQ�QiT�"k'Ӧ��6��~f����kg?.�bNĪ����޴xsd����~!i�+T���( �r9i��1��D:~����ь��8���lO���*8&vΤ���8sFB�f����	ޚs�b�&&�n"�b���|g�x�qM�qv��z����9��/�j-��ce�\Ƙ=�2�M~-=��)SK�s����>�>&G Nא�nC�^�<xG���ί@�}#X Mz�|K�a��D�?Yx�iI/	_t����Q�?���tmǽ3��/[�ʢ��z�xw,~���?�ah0���v N�Њ��f�Y� ���:���0PE�6��wB=Ƴ�k��ju&�c�� ^-LF�MS�.��M`��;�1N��B%���a��Z�(�F��U)��)���L.�\�Un�J����`X@�,R�s�u9�N�����s�~y�(���,��G8��.{u�Z���]��cטd��xn�j^z��3�����.Zl��֜�'�A����W50o�/C�D��Q�!�7�� �PG��vM��V=���)�?ό8�"
��?pÃO�t���-|��Z�r\@�}������������O��k�d�vޯC��2�����﮲���l߇��0�z�w�y�	պ�7C�6�)�6ž.�͙�~��I�ô�J��( s�������V8�p�5���
ی�}�a�T쐍���F05��D���7�j�Lz��DiRf���+��S���io�V[CE?��U��i�8�~Z�,��l��ƏV�M�Tq`�vLQ�-�Y��laS�chj�֬L��Q�̩�F�7�_A�!:�W�K��R�CX.ϙ�X⃈R�ܨ�:��z��z��_��>��ڳ?�?�ƚF�q��(�n�]���Ț��x��q��iYע��9�9��Qnp�aM�/�W	J�s��0!L4D<�#tvwn�X�|9i�'E�y5�#�"�d�*�[��w��#�MWg��zL8�A�#dls����3-��<U(�v�6f��1%�)@Ne�a�JxtF�YW	
>�I
��&�[yT��y`�_������g��c��62����e�\R�u���3���T�ؼ8�Jhg�_D� x��U��l?nwc�lս<�w���Ӡ�ۅY_���`t{���o_�ġY�U�%�C�#�	���	6`�R�d�]b��ɬ��c$���?��� V�ۧ�����d���:�'��n�D�.��v]�8x�pY;�	Ĵ�B�0Ғ]�>�K��~
�;��H(�w��q+� �n_�[�x:����T5��)x�Kz��@�o-�o3WI��n	���`]5?2A�С���'[mu,Q9$��Ǣ2Sɰ����HE��q�����؛iz��	`�%��fSDEx��Tk}���O�5�A_�[��U�M&!����'��P��XFmC�\<�	�]lc���y�v�&��"o����I�)��g�tfC߁��I1Ԩlz�B�v7��e�,�_�IQ������J�Tb�5u�����Eµ������/wD��o+V�S��g�Gm��E�d
m�����+\�Y��&�e�xSB"Fʝf�u���M�i�ր�#�4��G�E�C̕Dw�8���l	R�xe}hY�,��W�� h�n���O�7�ؤ��aA"��2i$$É����>f�b����9�g���Uq�;,���A����YꅗC7v���S��NR���b)�a��*t �E�g��;��oE��Y�18V��F�E7q�{S�Ŕ�F&Wv,�ۮ��Uk��y��)�ëI 2������#E���
�&;I_M� ۵�+�rL��@	G�m5o.�^fZf�����9�=�!\�
|�r�T��j��$�;�N��X��E��Yp��~�?�թ���xT|�_���Q���"<���e�.�}G�]��`G���-�ۜ0H'��o�V9y|�h��sS�	�ZqJH�� a"���@�<|)>^x?~\�wm:����3���2���)����������u��v���k�X.�������ZmI0���s�ԭ� �a��A"ެuv���6����ʆ�ڑJ�řdv�X���䚲���g�B��O4��}	}|�G��-��Wd��W��"��ƌ��w�9�����*$����n�x�l9�V��B��ܩNA��~�����>���zш��:���X���8�3�I���v�m�}~�Ûk�מ0�(X��z	<f��ZT���{\v2Gen��jhD���V���$r�vc�q��O�}&�(�9p�j�,�BŰٕh��\=��֪�����ҪY�<O�>�9X}���Ц߼#�EE�~��0�$�o���J
?��Ȧ$4o
�ѕ�y��wf��΅A�y�n�f.�����nYZ�BwQ��O���NI�1�n��}H:W�_<���_t5�1e������Q&�>�z��$do�v� FP>�����) hqb�֦pZ�f��;f_j���qAE�D�Y�ɚ^�,	�9bs9bN����k/tr�膲��X�#�~��+V����N6����I���U��r��1{hC����� ��muNSk>������;��V_�2[i��k���݃"hyq�uI����ݷI�юU3J*��%鑽���}Z��߼$�W���xΤ�2>�A�E���{A/�� ��nqC?9�"���.��j�՟�׸����(8�sXJ��=�=�|U�Ⱦ��W�� GÐD/-ƾ3)���������V�y�K@�ˍ
-ԛs�wͭp��u��P�w�΁�I�oe:���]p�^םT�ã �޵ߓ���:�=���uf��2�(�����Ӟ(-����{;��a0���S6C��P5��ܰh��6eӥ#CHg��f��wr�i)��$z
�ڊw,nb�<}WC�Z;ݨ����>�_jo6J%U�ͮ��$�'C|�qFd�D�>��D+v�W~^�t��� �Cz[�������E9wh���ϕg��-��K�sRP��'�'?6ՌR-��>3���<����"�l� �5�x�L�f���r3,1$Y��T�X��i~} vL[����\ʂ"R�>�6CD_�
�q~�)�|�Ȑ���<���2)s���1���["��dr�k����I'{[=�x�u�dׇ$E����B+
=b��T��B��P��F��c�隵���u�S��@��'���T�Z+NжY�Ta�%��y�>>�~�D�b��n7d�0K�yh����C���YFь:�B��3�#0_�GY��£��,vYz	O���JV'rnR���=`ѱ髮뷱���$�i-�w.d��@o�]��֜�u�F܍�W��AF��#o�LP�L�z����=�_nnR�?��xs;���`��,�2��u��&�
;��vC�����Fo�"��ܐ|��'�~(��	v�<�X,(c<���{����b���\?v@�l���l��e!N���0>�Rm���9A��oNԼ��[\s
'@�'�� �3��ߩ��!2.����&�ގQ�M�\\fj�#Ƞg`R����ɇ��SK����4|��vr%�_\ �Ʊ_�Ή&%Q�-�P�ˤ+
Il�Y���2��g��cv�%F����7�r�?�V9��4�|�-/ho8Y7dT��dr���
cϠ �����%<_{VȩdI�V2�	���!`L
��wș����t�[�L�H�KfNrY�A�Tc�p��U��x�l���)x��:���'���_Xݛnmy~�Vq�r����s=�V�Y���1�↎��x���d����!��������9���a�f*��9�ssv����|����kp�kZWcR����)<�TF���h�wf�yp��~�ȕqQf��;:9b{��ڞ�9H[��m�FA��{�p�������К�������K�.v�:x���v�-r�~���"���'���w���n�=lC�)ܾH���Cϊ�C��������[A�
����&�����?�;��H��q���i���7\��+[�a�dQ�y�"VdI��S5��@�v�𖉞;^1Wz���f�|�)dϣ%�9�DA#��wJ\�L�[��?~
��d$~WoNаF�����=:��E�䐉���h�v��$�y�����m����gƱE���P$ᒳ��^��s,pL�F���qG�pp
GՄƯ[èg�A1�M~<�H_��ht�9�?�R�Q ��}hd6�_�l�ٻ0
���%�T���'�-��+t�D�%+{��dJ���e��`3B�y6��M]�v0�I�nJMR�ː9Q[7N��@�#�}*Ԇ���q��?�PW�%?ߨ~�k(QE|p���e��1Y���m��%^����y�l�#���}��Vv����n�D�颻�y�abB�1(R�sFV��uq����ٸ��¾����ب���y?�*�̸�6�zʒ����O��;D����-��W9�]��*��f��3ֳ��/+.��5��Q
H��+p���&����+qr�$��>�%�1Q��A�{G4��<�N���h\E�L��B����k��n8�!O>�����<����!�$fmc�='`=[�*tZ^LYq�jVX-Ŏ��}�)�(��4��rA3��k7���u��Y�P+͢Tf��4Aq)���"�@B���L�Ѩ�7�t��嫷h�p���hp�����"2~���dR�k��{w����FG���*�a;<�2g���������KU��v�ZB[�m��gFO��A��@��F+,�֣K��3o��E�h�N��r��BL� T
jh�J�O���G
�p|��-n�<�ZB����X�4�=����<X��N�"�g%>���*cC�Ⱦ(X@+4Q v��������P�3�	��7!YN����4�")#>/��,��+���>��}#��4���&r\!9�:�h�ZX<+���"�;��l�Yk ��V�3h��R��*��*Ǥ9������M?��=Ce�%���C��Ҟ��oI�(��['g��]ѫg�g�b���P�T�<�W!3.��AӢ|�x)�S�Di<k�O�()g�(H�Tg[�u
oal��鐃U@�!��M���H&�Iy+{Tˋ�]��v˭���k�F�Bp8���5x���r x�߃�#��
tw�E9��O�����2����26p�B	8��+��KԱ�d~:�c�Ÿ�ID����QM0+}��_��04��k�}F�"���E�|F"_����϶��=PҰ��ӧ�h�J)�Ore�ZHxK'��������0pc�A
X�}h~��)Q�&CG������Ć�b�t|9��f����Gez�ɗ/j
[�˞�7�����T�Es�0� �sבE7���>��KR��V��j$�+-�
�F�ݿ[r{���'�����TuC�a��y�0�_�<|8$�հ���c٣opn\�'���R�bة|�%!&%W�R�$��>m7E�#�t�Zwf̭��(��Ӕ�Sx,	��$�x,�5�6#���U��=y��6^����s���,Ē�Ղ���\�b�@����kc�r�JZӁ^Acvcl�ǎ�4�46��-%
��\C寐�P��}i�M~ۂpIGl�A�`ݑS�!'�'!JZy3(�q�4X�����:r&6y�9��K_(�j��'G(C-Q|��݉�� 23�V/h��6��tx�E;�d�k:�.�r��8;�pfzP�(Yv�-^�/�ᮖ�nǳ��_���A�
��.)�x�_Z��t��"��]�N2�v�h[G��Eik�'�����#���{���p+Pt��0NgTz^B΋f��2^[�}ѿ�f�^KY�H�;c�eu_�.b�����v!�wGË]�U��ҥy�\(r$'���8�K^	�} �',��KkA�`,b %�?t���!���$���-�w�4�<����H8�rNx��k� 簳&�y��s�v0�j��<eg�M����}>wHms.�≺��E8rœ��:�)�J1:����  Wj�&Y^о@�O����G�"0�z���!��DŅ�L�z^Q����Ds�r��-��J��{�Or�ռ��g�)�2��INѳ�7�~�z{`O.�֖�i�p��ٴ�?��q�����9�:˱��H�M9�(}���,��y��8������o�	�T+�5�O�́��<׼����/-��Ȫ��jH�-��0�������U�Z?�v��W7�=����
(ěq��\1�u6�k�v�E�;�T���ux�W#�O鷨�2̀BΞ1�=<Z 0���(�=��_"}?������iU�#:,���C�G�J���8}7�:�x�7ȕĸ���0`�����jz�6a���C�;4�f�=�U���0���2�EP+�DM8��a��U����R7� �DIJ&�I`#J`��FW@��!�҉v���@9/���C0���`�:���Vĉ5u��j#\��]ت�m�"+�T'1$$3w��w��(Byo����/Ҭ"�s�}i�2 A�0��ܢjpi��3�E�d�hѯ�{?*Z�'F|�X��+Wu���G��[k�F\���U��5��4��û����(a	���,�E�E����p��7L�d˦�`�(̫X'���E�󷎁�u�Zg�����ԉ�R���./:/oQ��T���[J֩�Q,3����uO�����P����ͫ���]�v�u`��$'�;�lr��V-AȨu�s��Z+��滝_�Ľ��Y�#@���jw���H��˺�)}=dy�<������E-	�~?�}y�klR�� &�����Me�D���U�� ��M�1��0�d���0ӭ�'_}�A2���P�Z�%7���\��[VG������0�䀹�"����h��2��)��s�������z��WZ��Q�TX3{5���.jYc�q!�s8S/kXG.�¥�)ٮ���UPn��J�[�{<���>��;��B��L�
�����(�Q��0�!��q�ͭr�Xen�#��[���V�B
���:�1f�����`&���D�� !t~�Q���ŉCr���.�a	��A8����� B�2ʼg8�y��ח�9�z�%�ɢ�Ѫ{��A��	�3�}c1{�0��z�JmEއW��X�t���Xb��x׶Gl�&�"�6�	씮��8d��}�;�<
�����*V�yo>[
CM��Lv�_�e1 a�aY�";�0<�is������1r������_G�ί��l�6BN����k��M�y(R��5��}ڮ~��ږ1�*���`"�
�����ԫA�ޖ�B
���λ����a���T��k5˰�B��0�5w���b;��Iڋg��LT����q����� )�i����:�!k��W/F��$ Ј�Y�<�����"�����6����E>΄��H3j��d�3yŰ/Mx�`��'��]o�$%'�O��U[�Ш��6�P5J���	��p|R�u�[#qBǢ%������FKH� Ԭ p {��q�i>�
n�'�h,��얜�̟�����1:��O{v�+'\^��:�c�ؠ�B� :wMzw�ْ@�� N򝱒
�w�u0��7�T��x5&M�r�8L��ǵ�f��T�QA��� ���TWS�/4���6��0��(�=�6�*�k2a�J
�c��]8�����@O��<N1�c�f|��mh����t+�̖��'$�3.�ƕ��5=	��"��/z:Ӿ0�¾�I�o��:�;���$�ʢYvC��d�U�S�\4�B]ra_�U�9�O���� _~x;��Л@bDGw��)'S+��K⌼wIJ�'	U�{&0�a���iYq�w�y��2�p{[�XR� 4���s�4�X�x׉�Z�_D���Vtz��4�9P7����+���,v��I���
��S�n��`PwtF�WK�At{�ǋ۵�V��N+��v"�[!�|è!0�N��4�$��/!����?S��dS��l���O3�~��k�α�
v�%P>1�
�f7����YDI�:��P,m^�ovˎc��yu#��l�$,�ҕ ���gM��5�39�,�}͐1�(��K��C�uO���צ±a����ho�k�=��sQX��uUq�B��� ?@�E�E�4�w;7�)����@� y}�7��KU@�Ր�� tm?�2תM>I��}a���8�{5�� M�9r�s" @	���Z��p?KD:�[�2iV+���8��u$�Y.�$ ��!��i�(rd���ٜ	ST�p�ſF����E@�jh�+!��r�J�v!;e3fn�q�~���.���]��Twr?�����Z��ˎ���Np��'��W`�>�V_��dn���VY��ޝ~�%q��f���t�|5�r�ѮU�4#�����CQ_d���ٌPr���ٕ�m�*���%|↱������4��Y���a퓤��pD%1��1��p�SGNd
U-��L �C���'+�����l�X�-�>�j8��hh�eF5Y�BTZNbw_�j��I\^ ���C�a�%�N��P�%�o��_�4��KH.��o'��x�^"`���ό>������H-�V�f=�P:�q���c�a(��L�wժ�;4[(�� ��@d��Q�:zu���qG0 �_��>�j/.v��wL�@���IuT)��9!eu����<Ё=FQ�K�`@�b˭�+0*&� �Ť���q��{zm�Y��� �&,o�2v��h*�8�g�[��<0QCIe%�.�!B�v��gG�ԫyҥ���W����r/�i��!?-//����N�6��'D1�Y�H�F#SP�w�tr���פ2���K-�T-,_�%�!��[����S_+��;֔
�+$ ������ ��S6����v�I^���9|�xl��k\�[���Gr�e�d6�SE)sCi+������mf��彟������\�!R) v,L���7��{R�����W�m�?2F�����?1�}H+��AfsT˱�ԫ�!�ܗLU�`�Cc�]ұ:��l�N!oX����|^�^�c"�	1�Ӈt�I��*xT�ܿ[��QѴ ���z��5�J4�Y��Yp���<R菁�]��ڱ'�%�zP�?�i�&���A	�#}���T�AN�:�A4w3o���{NG�#x�n���W�[�@W{v3A��G�	�W!�.��.ŉ�e�y;�Մ��A�C�u����f.�hݴdP����22�˦�I�j�?��{�a�z��1l"�j��vU^SsD+���T�MA2�{��C�-�\�Lk���Y/��ؖ�m�R&�����]L�z��/F�~��Yg���f�Ƅc5bJo����08���X��ײv�Y�̴��Y-���Qt�[�U�1m�.R�|�Jg����t4#�Pd�D5<���|d"���j�]�V�	ЌQ��bEE�t�U����Ϡ�����<����H�ǹpq�?�8�Z��u��b�:�v�"�q&RC��Rz�2S`�j�[���V9�&tc���\���\�4���qM_����t0�kSw������v�^�tJ�!�1��v����9p��4_������%]���ACApa��,(�L���z��������;߈h�pk��� �{�F�'���!W�^"��y%��p��[��H�n�/��t��<�}O�� I��-�i
���N5��,�7H�h��ג�a4�aR�z����^l&�k�|]s/L����������i�@#�:�VG=2}w�+g*C�<EFO���i���Z����3�!j�6���@�A-��fx��WVi�`�^��a��Fh\+SN���㞗���]�Ȼ1��^�+��3 �%�I�碤Mcp�L^m�R�R(��S�#L�l�`3J����������B"�Q��H	���l��;��^��`4ߢ���
����L�GưQ�Yuz,Cc�`p��J�3#�bxZ@�S��lr����W��w��X�y�*x}hq���O�R�d�:��]U�biB��gU`���$;�h?)��#Vl1���Ե������Y�%���I9���U;�zm��"qߒ����o��ސa(̅�L�5v?�t�%����Wȓ�h7��K�5��!���{���y�|��g�fnon��.�r��[��N1&Դ/im�_��;rqˁ}6�Rf�H��	\����[�����+�,1y��v�y5^�=�z"���,�o��CS�W�&0@ov��W��T�h&���z%U�lU�����Q+*�Ͱ^t���y��,�YG��;�s��M�CG�@cY�2��㾫����İw\ ��!r��{���8w�^���B<��\����6��gQjK�@��X.�;��ڍ�� xO����>��nb����LM-:�4��d9֏"��P��g��Y6x/�S�j�,*��g��i����ס G�������+ٱH����t�����){n�&�*��)2̕P�Q���VY	w�J�l��f��N��z�K,#���J)���x(�������z0�ωEed���=�J��T#�H�A��-��j\��m����՗�"Ĺص�����=X���3��D5̾"�+xx��c��1�:R~;�o�_�U����������a���ȉ�Q��5B��7�9^S>^�p��撶$m:bSc����!Ϳ_��.���:�7]��-��xo��Փ�t�b,xL�3�������-�K�X{Pڜ���E�}�K��v�IH��]W��+�j�kɫ�#g�U D�G(!��)��a���8Q�4͈�]��]�j��6Zo�hF��)t,��_�@��?I���m`U�6!UUP�_!�L�����{�K;1�ɕ�]��d�ڤ�:;P�����y*��G��2#0�\���ն�vl�3��F楯�>Ca4�q���ȥ(��q2���� ��u!cH�kw�1�U4�]����{b�Z{~T��J'���䃕�<��
3+&s�#1�h�X��)���Y��qr ,E6|�W����P�k�Gf�w�\>��;�P��+d�T��@�`$���R7�>T�gH��N��hZ$'�$ޢ=�	���z��>��:=����6���YٻG"�3:H�$����h��L�#uKPBi�k�sO65�j^���7l_I򒰯��2��*���ҚPr3�\��S�&�s���1`��F���M%ZZp ��Z1�&�&�n����`��}@��s��@��Um� zՖ���ws�O��u�'�i��9��G�VIu�2e6�3c""�"u�q�/g*�L�c���*����5�J_�A��/6O���l��1�]
	���� -h":��JX�$h0��V��x�$��2�;!�p;t���p�� ���@>�����XM��U��V�`��S���0ɩL��lj�W�eF�[�K�K�������9��:��Vձ48s4V�~Ns�4sF���v		׍4I9F��>�����m�H3sU;q�f��Z8C@p�Fe�C�\���;D��"zr��F+�ߝ�����x��`+����<a%l���B�ߎ�Y����?�|���tr�3�A���AfH�����v�o&z:K[�(z�l������8�X=zU:OT?�U�/<>�
y�Bၠ��e�P^���:��o��wQ�c2�>(���֏e�|�`��d��zS��]���oZ����`&g:��TzsĽB�xk����ҒM��`X��
��@;SM��u����ͪ^bd��NXhH����<)]��1W}��\��A���n��2M�q���\���zv_�{W���ZA\��0Ĳ�&$��O�X��p����g���gK���������.S�1�lxc�܍[Kb���V�M���L�@|ȕz8��i�8y,s/0\�Ў^�5��
+A'5ߓ��ɂ�A1�1��<�A�ׂ������e�D� ��D���48�?u���09�x���:vGa�8	�J���iC���|on[DUc��Ė�")$z\٘ov��k��9�a\A�h�^U�Ry�����6��[��YIm=K7ڹc��y�~&�	�5�\y�i����|����+<l���1���@��n�A,CI4��a����/F��%2h}S0��Ųp�=�.�9�ƍY�B&�J�y�����V���O>IpЙ���~�xPN掾:>sz����$Z�����.6�{(���Zťc��B}��DG)[��I�e�8��!_����>�����C\A��/jS����2�%���F��`���Ǫ/�E�}*$��v�:�*�4L�V�+�hkЭ*A��r���s$Ȳ�Uhj����������yh���貐�@6귓�j`�<˓K�$P'������j�xF��V��D\1$t��݆���bY���N}؅�@���2D���Ja������2�D�ML��'7�2'�R"��$�F߹{�5�\	o��!c��'C��
�#H	��M���G�{;|<#��	i�?��&�b�5-��h>o�0��l0#�.:c�שk_�YLx��T�=�� �O����V�=�2��R�� �
���FGT������[�P=$�t���}O�^��X�A��>s�_��Kn����l����N�e���V�����%�(mV+�8��e��ѣ<)M@ť����U�:FZ�f��;D�|y�9 h_���Xf�3��黰ƍ<ǯ�&��>\�! �{.���#�
�k��5Y��0���� x����j�;���19���魮�Ģ�f�H�{Z�S:�;����B�u�я3���U|zCS����g�е��+y�g@�F�\��c���p>��nieħ2@�e��wc��W[�F����p&����m�R�N�_I�=��k���JQ?f��Ip}D:Pq�q���x�;�r/�v9&z�����D�̡M��Gԡ�8*\8:��fZA.�N&tB�?"jhd��,��%�u�b ڱ������$�vi��Ǭp9s�*�v���=��Y@ɥi�^�Jy��,�VV�
lN��W��e�Q~S{��������8�u�3�6�|y��N�R�#ǫ*2�	�A{�t�a��D& ?�ԥ�E@av�
7���R�BP
PD���'�'�$\���xS .�nwXgF����0�~����%�;���fm��[R*4����.��ī3�=��V�I�k��Ƴ[x��qۀ����<�i]5_y���t쥶�����c���9u���C�`p���Ms!���^^h�R.�fAo��,���|b�l��5yU��M]�Ĝ`u�T�`2�%�;G�W�wڔ�73�LK�6ʘh�u#��0���.a��&��B�gz~:�aY�s#\��@�)e�ȑ��6 \�I�23Ə�t4�bx�j2[e���s��
�4ݞ\��x���>&�C�-0����s�G�"����p�-��X�N)*;R�`�w~�E],�c����*e�ځ�K�����O�ym�(2���]�dVh��&!:��PO��\��������_�O9�X���XR/�����V[fdD��W��s������Z����"B�:�4J�)�4��*ʆ������	LC�4�v��DR�m��'t�ݬ-}ܖ������:b�0�"d���im�m�P�)�	��4��H��t�>���a����� ^0��t��\�z�  e�z4�1$e;�N�1O���Mzn߻���c%���6��Ɔ���Q�:�wZ;⢆Z6zV0j�X��&���k{�U����m�>Rs���?��~�3>p+nC7��,⚚��.j��Q�%ȱyee\�3�J��o�ƕ_U���3Z��"	�X�^���>���������_�:ia\h�Qy�~��x,U�r\�A�tP��#�u����+F���J����� g����Nqȸ�\��?�B���9f.oK�KԬښ��נ��n��0sOT�����"$�a��p!�z8^�A���l@�}�9�)��Z&QԜw ��ނ��Z�[	�,�����Q�jR�u�K�!v�`�PH��o�cIMV��%6M���8Z�2�y�c:�<��*b��/$���%�mr5g���1������#]���g���|���l"Z��:r`չ8�/}�*����Ơ>/-��E��l_nm�(�1Q�f^u<*�y)�>���m�V0W��f�^�ª��ļtz��v��	ks��4��4����	�o���1Fd��;._�@�A�Wo�n�d#�wq��ԸU[8ZW�'���uf�e,2Vu�b��m��#�`b�%
��3�d��&%�8��dPr��v\	���������v�S�g�(������ө��ݍk~�u�o�A�Q���������e3����9�V�3���u����B~�R�<�@�_���C������A���_˓i)O�'1��[�բ����RRd�%��m�ɺ$ݬ73C�H�t�;��Gi�J�ǻ�����̩p-��j@�t6��Ѻe��@p~�	Ze��q�ܰY�W!x3������G��V�?3n:�[��$��ǉƢSA�f*| ����u��@RŻ �s0�,�/�$�Ȓ��#5B_�}$F�e)�G7;�I���������P�̈
��g�A7m�����;�����&�=,�4K}�@��YP?�͑]���=�<?[h��>������bB��)�F��5٨�tU��k�8<_)K���#~�.'�O�&0��~����\,�Ds�HA9���������� �l�E���闋�)T�]``tҡ��F1��
~�����k�D3<r��A-�B�7-@�����Y_!]P��C�r�Y���#Eyh�>�\0�[߶�W��R�֞��'V��*��PEB�Bە��i-~[Z+u�2	�R�ß|3�����{��cA�'*
%�)K���3o��44�~ZA��:u�ȗd��䢛����t�� n�����6|��o���^-:oo�'�ƹ�O��S���;q��0fE}H��*���A#���r�1v��Y.$4F�(��;b g*��Ab (*�i�6���?.�X��ā��8OĴ�Z�{Wl3��0������(��>_�e`c��y��5��j肹O��ind9q��@a�%b�gߵ��g iy�2m�s���}�1Ʈ����qˁ��=��孵4�z)�6T�4�W�S�$t���S������� �U��+�)�R��<��
ב��b@��y��$�0����co=w�"����F� �C�H/���IhN�N�l�^X�{�����M�H����[�[7�� ��m��L�'���{��$[���F��=��[��,։_1��g�b��I�p�h�YD��f����g�������R�̹�՚^`�S1�>=p=J�e�W}�aa]���Ӈ�L< ^��p��{)e��pmZ�XN��>�6H�����R&�u߹�}7lJq����.�0M��:��� ȣ��~սwNi��Q�i��~.wI)�CL�H��7���4"���Y�|���cÏ9̣V��L��(�!�૭��%�d�z�3�;D"��:���Y�ȋ�b�8��2���Jm�RVJ?�\�qG�F���7����6/��g���O�f_��c�3��DQ�t���cg�0E����Gxt��&�%e6��cS��X�ĳA���'���%)ϟg�Z�G�s��p�YϘ� �B��k�'�\�(�������#æ;��Ǌ�Jƀ�=�{�Gj&��)���'�/���?��(�N�2њ�*��/��)���%�:m��4�*���PL��KR��<��]�̌�C��v���L�}���J���C`�Nf�~`�.N�o��Y���[�Zg�p[����0>d
����G#}�E9w���#� �g0���-�I��n�/�N�D=̀���u'�\���_�ȍX�F3��3��~�]�>�:��dGI
uH����E���^uwT�:D@f.]Y-�&��;���Ǚ��O��eim�}�!�ON-�lT��3_v;C�Y��"�x�T�ÏLLs��P�`g��$�	��f�>$� �d's�Fu��������~-�X]��%�2�δ�d ��LVD�6h�)`p��<�H��ۊS6�7�>����\�����,�5*��鎧H��d_FiZ���D�?�RF��8y�rx���Ǉk�P���P���
�4�� ]_[nFQ$|Tm���
yJK�]NDQ��ݠ�_E�K�B�U�"�o���K�u�]\Ynk�IN��LE6m��v�ϧW��C2��>�Z_*�l�n\QX�}���2��s���b�P����So�3�����id�W2�	��8��Y�a�"��!�br�9�Qh��
T9E[�qsn�Z-2b\Wu9�C��n��mGQ�a�,�i�{{��{�ؑKs�me�L�=��6�hG"�X��A�_5��&��K\�Bq�Tky�����3��視c$O4�G	��]8_Q�ġ[��~�a�ܘe�����3lb�Y��e��ѸY@��a
H&'|�wn����sL�E�u��|RJa$O���� ��u9�e�u�#�)!H��gT\��-�g= N��i�8��/�ݟ�ls N39[:��) ����e� �������k9&���E�)2�xA{�l :�0R!�q�\0�]IU%���/�# �Q�=�>���-�~(��n~Sk� ~���q�1yr�.�C�1Z�-yB.]�7Y��M�Qf۝�<��g 9*��k$]����ڔ���=�X��L��s���9��?_���ز���Q�fc�RT����@jB��0��G}����7"���y���Y-��lI{ۻ �su���cč?q��j)$��K���]#M���e}�ڥ���-Z��!�'>0�P�@ݢ�[Y|v���%�uG�3���Ȓ�S�MF�G�4�_?x�_+�T�y���>�ң�jĤD9�2*W��
���Q
�4򥠬�ߢ��UP�M�G �ڭ����֊v`!��!�،%9������>ø�HFؗ���ǅ��]�����V������e"k�q�~�D�R�X���/�a�������-�E��l���D?/����[�6���F��fNŤQ�q��ŞYX�ov�Vul���7��8 ��h�4�r����0�`ɜ�>���c�ȁ(����'�}����9�����-���8Y��ܭ�X����'�O����[`/�Y��K�������YN�����%�ٯF0$R��PPsL>b��m���z�K��x�ZƱD$�N��Ye�n>+mN��W�b��d�C����sQ�\Ԡә�$�9�ޕ"{W�t�/ͣ�>\�x 9�̱����+�к]�ChG?U�on\��52���?Sb�5yBw�*K��Q���o)k�<q�hL��'�>��C���|}\�4X8Ȉ��P��U&��l1oP�>�i	�<�O.ς��"m%�K
��d���:%T��U���ҁΤ�r �I��7�Z7�ԪC��"�|i�Z��'�V�+��"�{��R2sou)s�H��|�)� ��{8�uL&9�����c� ��~��/4�rj9vQ�>W\i+\k�*�yy�!�g���&W��G�:���+�3$p�g��(]K�kR�'+��Z�Ѵ�b��.��}p��{�j�%�Q0	�����<�"+�����X�����9^�+��<�.�F�Yg>����_����P�Pa��k�'Wcn�������2��7 �P2��9�C��@��1���Xl�S��C(i¬0����k�����O-�h��z�V�Ͷ��e��f|���ҩ2��(�<ɳ�S��mC�ݔ^�pG�YC�;��Z���W��2��0PN���q��߾'"�(^�8T|E˘�{��:��E,eO�A��
�-�t���ĥu)��26�˚9&���5��k���(�+|���&z�{�<-�WwC���g4�yh�M`�[�4�EL�_"�� ��0y�5��%K͗4'*]��纩��!�Q}fц JxQ�����i�(L�5�/�o�k��nw�k��� �{Z	������(���[l��k+Y�9� o�6s�����2φ�Vf����]���R!v&E���<@ެ��Cd�1�sK�%�|_q���c5�V�"�))#ӍUg/��Kz�.����q�[(Z&
8TVr3����T���;�8aLm��>���	.y��!�ʋ.4#�������d����2j�ޡ̐d�A���3�!�1�VN7s��$۫Ij4��HLH��Q���!癃L��#�%�=,��֪��g'f��M�Mf�׷�C�d���8��3R �7�@@����oY@\���7�"����@���LғS�i*�"�t�-�f�dY��󀛜��!5��͟g�t��d�#5�<ֺ�3�Ɠ���/��
���=|��~�;�'�������H���F�FL��8%]Tȭ��R=xe��@��a�O��KX�I�'hH������Q�}�3���#�ث����%d�|�������������.x�t�,�=4_*��[��/����6��T�G�ca�A�xh�\Դ�+)XZ��l�9�}7k�,o���H�u�CH�H��3�,�I�ʬ������}*�!g�|2ӌsS�c��F���&) ���Y:���7L>��+%�r̟ظ���@FQd�R���F��Z���5I����)��A\_-q��*X�"�w�������3�9��>�����R���t��h��aL�^��g�� ]~�zb��BN�Y�Z� \�XE!Zp�A���1��`*C�~Y��B��໣�QK��h�v��qG��Ʈ=e�N,�3�m�,�W���x�Q�qwC8�ߋ2�{��z9Z�oL1G}�~������p����t[^	��A飬�u����Y>UP�� ����pMpg@�Z%�����Դ�����d9p�7�QG]>a� ���0S��1�zD��wU�}�K�a����m����L��:���┢�%s��B�^�����u-F�W`�)��\-��O�9�|>�T���Ydx���D�����5���Ff��N�ĥ��&����C�F*�D��=�����Ҷ�Z�A|R��%4�UΘ*֔Ƥ�C~���^�u
�-�k7�b��RXZ�����n���R��ʌ0��j�G5����ФD.�KpC@|n���yY���E���A�Uɹu	]����K_c�r�NУ�>o�a�qK_����:���u��'AAoFig��?���T@q�Z�ޫ�K�J�A3�bFE5���p��+u�ڇ�"(ϣ-�"%T�x�jLNw�������4�8�۾��4�FIy@Ydb�m)��	�y�~!���}
�VHoOP@*��ܵ��ۭ�d�ل��!��s|�up�@M
|�͛����*�ݤe�]�vٱ<A%�x��mf�@�` ��@��@?tyL�y�
��2��uc�uO{�i�����=�h����k9��b94�LOrSؠ�|�E����D_%���9?��;�܂�?�SbA~䈳7��/4�f��J�B��^�!nvP/޹��@��;���F|0"��|�J���$}�B�v���P���,ƛp�>sh4>�Z�pk�,��6Rm�#�|��-DԷ�IC��D�- �C�݆'GD�z-E�?�o �2���o;���~/�+6U��7��M��GK�N2��Ea��	��'76BFYiE�%Z?_��D�"5 ٫)��[�
��uIg��\P~!0�6u�hOwQ�:�_���k�l���OƠ<oZ��TQ�q�]���x��*X�h=�N6����Ղ�C$���9�*Y�J���r�=�+��d3c�USв�O��y������p(^t$Q�;+AM�+%Ot�{ߓ�n8��ʄ4RH���'ڊ8������T< �ȓ�x�+%|K���"�<�g��.Ws;�Z�3��kM��`��1w�D,{O
���W_�2�,.ф�?�M��
�i�J�� ��.?/vF�_�X�B�4��&��d~��3+��.6,2�����ir�@��r��Fg?�,V�tb�X��Y�>�����$!��ՙ��,44{ʉL��VRz���ę�m�_D�<-��׋E5��$�
��,��wrpo�d'��|����7m18־QO�}�wUx�MW�UU���~��EW��oe=~�3��u7cMjR~N^��44��d�����̓~<[�a�`N���)�#�LD��rЪ0�h�xb�j݁�4>���\�}~�	�%3����q17�:�V��n.�p��q)�i�-��?(Ř�Ro�F������4����N��Z$H)�y�џ
��:!_r���!��k��%�fޏ��Y�H6�1���T��Y���7�H�Y��2N|���7�d�cA�,����� 9I&��U�mtiOu�Plg<�݅i
��u2�iщ!�{����f�c�i�����0�0RT����t�e��+���0E�H���{������L~y .Ӂ�
�F�C��]r�	�w ��J$՗~���%E���'��ӳ��آ��@U2s�_����E*:�AѦҫiy7W�H���Oj���S�0^(��w&�xz9���;��fqg��ٌy��{Ǝ��(ha�ڃF�T�������RL�u�Q*u�C���|��/��	R��/=���2�(�Qr�)f�\�p�*�Pҽ�@�M ,��]�f�`̵
��7��`z�qmR��Ώ�s5_��I)i*�����A����3�� V<(�^��ܪ�#�Լ$��(�ȫ�mn��é�+e�P�����@Z���'O�S�S ��ud�|Ð�w�8�v�b�8��Ns�q�x�~n�e%jk���Ldl=c��j9��~��w����3�D"�Ҫʮ����_Փ���)�%��rqV���*��H,ӗ+=�!��YV�|���q���S�ŹT��^�}��`lmB#o<ҭ��+jC��؁�hI����y�����x��FQ��b�us̂��`{��|J�g��03�=�,�y�.q$u��i C�R�e�G}�j��V���d��h�1��-������qxx2��	�خ�3O��h���꒢�^(܃�� jZ
;��kM>�wm:�8;3��B����F4/�8/W�7����7��j��(�IK��Ť�T;�|F�L:�N����"1a%����}$�+$�h�����a�(�+ȫ�)tZ��Q��inRB1M�&�4�s�U�4:J��lc-ءϛ�0��{�2|�-\�3�ƺ��V�ZL|�6�Ƃ�؜w���&�?@#��r�
a�C��FI;�*\��:��+ĩ1��+T��j�|p	�`��m�	vR'���}N�p�ݶA\dz�.~<�ڐ�3��ѕ	��H�!}��5��w�FW���U^�	�w
J�Z�GF;ꗓ��'	"kY��̠�����t˯	\w����s=��q|�k'��X��-d!9��k�ҫ�c�z ]H�)��+s�w��w�>�q�l[��aV���~0���<���ug��8����ډ"}�D@��4���h��o�i�����q�l�72�h��c�
T%8�f�C���4H�ȉ��b�K>�����maD�ff�A]e�D��v�m��M2��Y���
7?(���3C������(<��[B<�D^!x���6GM3TT���;�3-���x�ݧ�Z��G*Ԏ��z��EU���3�3��]�����Xw�|��ݶH������@�K�d� 8Y/}\�i�T�N�O5&�]�#YHNS[ҥ.��]�g&uUw�Y���ary��ȕj�O�KE�P��:��Dl����n��A�]H|���,��� 7Ř#o�ြ�)�pz������!StZ���Nn�\<���2�@�:99�4>���׋�I�L�?~�|J5a��ҍR)��_L[�>���OB[�<���眄�.pX�Ξx�X��ǆ:N�a���q�;n�7��1��C���.Ѧ��$�p=��%������0�i��C��;M���ȻW�o]�*�6I!]+�䆒���?~��àو��ru�׊o3 �E���͒9��L�~r����Vm/;�"���r�%1Bڋz|��{�rr�>�R�{�y�й@[��Pוּ5ս��9�-�=,$�͝Ȟ;��o z�Y���@��I�5+�?�%����еf鶎ݭ��աO���_�4w\���S0v�
��yH��Ǐ5��(S�*��U�:Ƕ�{��X4Rf�B��lJa3�V�����9���)�x�4���<n���)�ҽ���v�u���%�9�cҢ�w�X��ODC��xu�V����<�)�|wt�ц�ނ�mp�0v��\���6g���}�c'�H�pXعD��E�lAK�����c�Bv= �
P�A�������9��� ;
�T��
ı+�5�<�g]�)��^m`��2�͓M،7T]JI�X���bj�)[��Pr�"K�4�A�g���>�4�h�DZ-xo��hP�6�����`��":�4���#^�l�,S��K���V	�'�	���yyMO]��D�,�h���^P�ԸI<������h�V�G}��������,e3���LF(=�4J�C;ÞȢ�xk|Ρ9��o�5^+bU;[�0h�xX$�H�']���̶ �eڭu��u�;�/����mtQ*�����3�e���F��AƯ^=��s����Gf�A�(�Y{�ݗ�q�!�%D���cx�!�n��g}�����Q��,t�j��Q�5�굞��2�3�~xG>�0	Grqzu��{3�]�S)`�Q�쯽�ۤ�dN}��h�p��/�;�g~WÀ��+{�ŧk�~������E��v�s���g�n�ū� �l"�R�9_�@y���P �TA9�rl�Q��R[b+u6��v�Ů5ZN=\�Q����ӟ�9@�>b�s��/g=!!���,��?}Ϸ�e�]��� �� ���p(w5!�?�L�'��V>C�8=!�6Q�R�<�����rN�2�|�����t�R���\��bU��S�o�םV�֐�/���$rq��VH��"D79n�D��2��z&�|��+$[���4F3��鮴&�m�h��}��Qe���ٞ���1��K�u;�p����v[�t]m�����R'�5��e-���rO�	7~��3OZ�*B���듲��Y��C�n���5�O&y��=����3t!�)_	�wj�������W	Q_Yz�3f�n�'��ч��%�R����q�3�V����v��Qk�+ x����T�강�������4]��ƒZ|D�Ֆ�4)Tt��v�ęA%%�9���Zb�c�IV�X5�~�w!�����9f�~i��ң��'9�.Du��~B@�����:3��S��/v��ei�}��ȗ�[(xR����#_}�7���t���V����8���.��,ܥ��r������
�w�k����������`�H�"o�g;�� ��?�.���_���	�x�	�s<#b��٘�_Z����@���Z�&)��D�.�R9ӫzd��`3�)w`7���f����T��-�)[fx>C���G&c8�����~F�Q#���T��C�$v��g��>Uи���$m�#0K�/fu��l������c��㼡n'��B���3Kx7��G�SmVJHT$��4���a�&6N3;�}Oھ�����~�z��*�� �9�L�h �'��p8�,�MA��
CO��R0��;�����7Xb?�NZN��+��~�幓>嗼��3��KK��p$����M��O�)X_��"ņ�3��X������d��YM�
�k��W�c���E�@��ʲ\'���^y�d�y]�Wb?�]�ѫWt��6f:O��;���)d���p)H�jqF�!�ĨK:)��|	*2�V��9E&N@#R��4��7�ڳY}���a�^qSt_�͘�D���j�o�iH�)2�=�!��E��|+5��������#�u��Qe\��P���P<V����fҝ���B%��$��W�=«:�b~�|i,c7��
@�#�jU�(��=�U0j�`�Nf�+ �g�pu4!�C�6}�����\V��_�^u�Q��˪s�5���0,�.�P���!H��,�@J	���^�'�,r�:�t�%^é�Y����K��|�&V�L�	N���а�}��h0a�&�>d[����d�������\�nqB�/Ҵ^�H礟һ�Ra�{q�==U���˜�*�Q���5������xy��1
�n-���gu��b~V��g�M,��T���"��z+�5�U秉n�컈��6=i�k$߿U�l^�'a䔜���u�����I�D�rr(Th����O��$]N�w�)f�l���r��l�r�y�±���tԨ�>:	ZOg�c���(�v��"���7�omh:�!bD���Ϫ�$�ʙî�]�H\�C?k�g����d!M�)�N��i�Ή�Ia7�ԹoM��w�[�,�(ODB�L�ǔw��z����F�e��Ŋ��6 �`�t|�BN�C���Yl;s�i��	;�ֽv]��aol�O���h�_ɡ�FDn�I|���?�������ʆ�*�����yC�A>�M�ugQ,�D��p���G#Y�`9��l�l���-ޠ	�m��0H&����ع�緺��p��Cྞr�t�'�kx�
�A�e�ڂ�_T
�X�-pJ�w������Uez��:�8�㴕��zd9U"�Bk�hv��b6ί5d����=T�"�K�����h�rz��^���e������J����d�z'�O}2���S�8���!�ll�n��2���3�����9�*(�>7�	InVp�X�p�.Eׁ}�I��n��Pj�b�1ҧ���	�ȃ�`��D@V�[r���R�Lt;>�+�����<.�6�x�L
�Fl����s���{��Y��st�l@(�(���?���s���f���q`���G����3Mށ�T����v|x9�m�A��fi�U$�NF&�l!����[B��~%�8Q��ML�����*h#�ud�0��ͳ[Ȋp����U����'�5���Wy�o7��̶��X�@
Y�Y����ƛ��5���'	]�J���⠈�!�� ��/Z���L����8�J�xe�f+s�=	��a����[׮R��� 
�K|����z��\%[��WXix�@3��~^� ���׆I�U�Y���h��,q�r,��|�q��!�FT���֙e�L�M��p/��X��hX�{5�A��L��&nɊ�t>g��o�z� k�P�Zs�@�'U�"g��'���!�(�zt�w�j	,p�𿀇ԃ���Zӵ�W*C���C��a�ŵSH��`)��P�1ҁ�4u�:��c)?$wT�lOr-�H��M��`=�i�6�S�!�"9�O�8˝�����#(}��y�3�ymG�03 ��0�G�g���Z�C�=�F�L� �0b�oG��%��]S >��8*܅��5��Aw�G������
���f�	�O^�^�kz��lF[C���
%r�'N�K�@�1s���T#�]]�@<?d��UD��UϜ���u�@����G�lt���<f�Ta�XеJ��Q�Qk:������ա[H�c
�H#���r�%�w@�Kb!�vײ;�ˮ9��:1c`����*�r|��ۼ����zVͻ8j��)D&Svu`��0��+�A���*zVY�F/�":,���~�Bo�u�$0�ˢYÅ:��R���A�O���-p��s��hE��:�������8�^�dx�A	�庚7�V�|.��Akc}���s���L��v���Bk�-W͋���)���S:"Z<���'� :�(wȘ��W�?�go5�<�&�T
�3�&���BY�f�������*ga�&�i�Ÿt����+U�2�Ƿ�\@�GE�� ���'�c�ϊ����`�b]p�|�B���9�El˧��!�O���qb=ȁ�'�A�)�jO���	��ˠXc��ywc k2K���ޔF���A��tЙXb%$2�?]��&��7}��7�a��s�N��*ޓIM�|�{n��r��Kw�Ǳ��:Lȇ�[���1;s�J���x�'�W�*�ͧ9a��i�@��Z�D	$�ޚ�GN}y�D7յ5���;.I:p�4*���#*LH�!��5╚~�Z�d!�=<�٭x�E
�J���,wJ�u��0,����؛��cG�xF�*�O�����*C����W<u�?r�����#�g�g+��pl~�Y�/�V�f��'��r�-7+�J��ff����E~��H����0PO����-�T�?�2�
8D.�կ�o�l��^��Ťq�`9��ZM�װ�ğ)�fm���	`��t1��.��/na1��IUv\S�ErA4�5x�+��NUX�����3ߎF�0o˩U�9�1gDBJ�q̇Lx�O�ҷ�	�w��WZ����OU�YS����b|�ʶ�R��$���-a�P1��=$��R��e�-�0��x�Z���6��!�`=�`>/p�=H��O�Ġa���}�BV~�!��nsW]N0��ó�I��WɲlB�n}?��.H��Ez��טH�v�WR��	�	����$-�,�1C#����=G�nĔ}��8���:���RW��@������u�y6�+Hqݠ�@���==��w�QJ�-
q��%���2����ЇH���"�hH\*�-S�T
���녠�H���2����b�:a]+�Hm�����tG(�a|��_�_�q�N��v�]��k��0x��p�\QGz��s�x7Rn6:��)V�X�Ɖ��b���WU��L���3��R�g<.��Z�Ɖ�f>;IviiK�?%��@i
d|�W)b֣h�1�w�yc Bt�핆�Y�~�eph+A7��Z;:|B�"2&U���2H��1���h9����{^1Zn�m�6b4�J�94���$�H� ���qk9��V�k� �d���x��H$E�6�(\�T��*V�\`�-�N
ʝ?@\bI�K����@�3�hj�p�>�q��-��\8N1s �D�p#H[����s(3B_��;���~�bT^)`N41��8���yw1.B�G\e��Qc@�c�$}���<Ȩ7+q��_���)�w]7;�kS��3w�%a%�D_֏�.�Q��8�
Z��=��zEJ��{F�}	���!�{�����"�?��+a��)��W�an���b�E"7s6O��o;����l�;&���"&����iã��d�a$`��h��CY��Q��o�
]�?_���G ��NŁ`,n�cH)���^�|7jx�[|a����`���Q�u�O���,)��)ǐ�[	T�0O���Y�����G�>���ҡ���Wh7ϴ��.�6�`�g��Ԏ0�U4��c�j`���W�l���bj��шC���n�O����9&t܏K���Cur�nW��2��D]��C�H����	%���|�[B��j6[��a��w#h�
A�8���5�߾j�xR�Ghi��ŀ�<��{�OK�6�@�
v��+������������{��>9��"y�p�\�wL��'�F��q|7-o�#n_�(�K����Px��	��2��C~G��	�x���t�,���/�5]-R��q��Մ|���J{���߳���Nw
��+�Ot���2;�5I�C��J�1��)�S�^k�U}��!}��W^!<�X�Jl1L����Fa�*�SQҗ<���~����F!�u�
v淦#����B<��Iz�g�s'sC��p8�s=VW�}�R�8?��L%<�EԱ��4#�6(�{���� d9Ad�b�����!����M��ְ�F�~�&���E$W�=Nwڀ_3e���\�z�����8�l��pk-���tG���w(1ɂEa3L�Z�@^��[@&c m�:�W<H����K����~��f�(���*�+�*7�pSLQ��魿����)���X]k�i��4��0�Op��l�LEH��V�o��5��hi�|�WG\訡i�Ұ���L��aܐawF� ����,�������+��$-K��l/v|�u�x��Iw$��U��˵wBbx[y#R�'D�S�{Ӏ�)_�q���D����E�̿��3`
���-��l�,�[D�耑���E�1Q5_�,9������Æ�k����Ι�߽]K��[b��߫�S7�i{oUTZ�g���}��\Pο�
Q���3�@ĸ����� r�uR�F�5�"���G�ap��Cl*�W\\̓=F����j�ˀ��+�X�c^�7�8�(����#�Xu��b�*���$��kz�xb(�)����@G ga�qm��i�i���@�5D������9��^��q��ɓ�&b�|ǰIU�O�O��9�$�R�����["A
2/��#d����y�r�}&`��<R*���)~���}�T8G
B��Y,�C�[hm[YY���9�
�O�kmGf�Sz3���@�sƟ���<@��V,M�� T~��ь�vR��b��\S�+I,����/?tY���dX.��8A���̘)�x�sr�����4^���~J����u0��*?#�S�ly<�10��*���ts ��fԵ;u�S�(	�_��_�l��7 v���Mx���Yɂ�o�%;�S���Ln��U�V��/V�ɳ�Y6m���-G/�� �I���{��W<��?G%:�#'MJ��md�G3d��iz���uH��iH� M�W��vQ�� RC����m�N�Κ"I�.��� T����Oϳn=~r��(��>>�`SF�:�( 1iZ�-:.t���d���=@$��`	�wյ�2fpMV�p=�|7�9�o��IzL���fM4r�Mk��1{�����7}X7��L�0�En$l�p祴�f�o�	�U�⥸����e�A2g��,��b@��ٺc۠���
.��K�MPr����ҶY.���l�Ѣ8݄tUC��(��;Ć�4�Ih��a���`�{>G�����f���[��R����w`P��]�dҗ2��dX&Ul��neV\�p���������^-hv����c�QI����
b��,0Q@�pp�r؛In��DI�6�mڰ�n>�����}C2���>�Дn|2[��1�b$��
"��dt��+)��ip�S-��G�IQ�r��g����jD�6a{�b�l4:A���_�B���� �Osɐ}#���@ۤo���&]�!������ݜ��Ɓ6��Nw=@���"�?^�)����\�:[,6��i��։BFH.�K�y��'��s���P�r��5r([��t�o�w��yy�~�]�a>VϢm*N� m���beMQV�&���v�$�:�D�J���#���גe�Q���7��NuG2+6!�E����Q�����	����������i��Wr��
&|�1�sT�W����\�d00"�ςVy����0�A��׶'�S�ⱂ��K�6a�B�
�M�l�y�#L�u�@Lysx�ͦ8f�F1Q,�����I�$b��#��Fp;V��[5�f�E��Y�7�kšFo�ؚ[�M�p�����R���e�4"i��d���Y���������?ZC�Ӧ���+#�b(?�XN~N�%6?�8�[��]�Y����|�H�`��Zަ�B9�A}]�	��PPH��Vh�����E����?RJI��߬7�~�T����\6�oG���/r�2���	8���NT=F
*#>R���B�%����d�`œ+��Z&`	����2ן�a��&&����$���E���Y�� ��lr�����= ��Ɠ��{��N{���H�\v�h7�r_��xC�q���O)�����yr����+	�x�ʁ��ڡ����H�g������O: M�8JU����a�6"���h�6��ਜ਼ғ���%�x?N��I⡝{%�s���#aFRH�"-���:ٸ������~���/o��}�L���' z����� Wɾ��\2�P����02[6@W�X�;��N ��W�\�P�^�3�ZY-n��D��ƪ����P��C���d�>�q�8x�!��Y6e��#+�S���
�����}�|r�D��� �x�Z����шOs���Ym���PÉ�nd��M|�����(n���.u+�V.�}�<�,*�����Uǹ����L$�f�o[n�f��Cw�u��Q�x��"}m�4"���w�ϊ۰�S�� ��_OOet1������̩�B'�y1y*�u�R3Y�Rc��QN!�N	$���R?\��h�peh��a:ۙĺ�L��%r^}�~��"Jp%^[^�	j^��)���:�
��caK��"�2[��ӉK6$��Fܱ��-��W�{D2������|N��]p�/V8J�cv]	5}d,i{�j����._w~y���z�L�5֓¼��t���7��Ķ���R��5��ؒ6����ǸK#Yho��歋�r�+��J|y�{ ���U^���tD�\�y(����'�?uX��R��W-��D<�֘�N��T'+�~J?�Ϸ��},,�%�L�W%`�t���+�^w?)�k��l=8A#��p*Rm]p|�8O1�y�u�l�pJ<|I�(���c���Q�*¯t��=�5�O���e���t���}E��]��4����Y�pDP��b腦kj�u���#cn�%K���Þ�w����yn"�| ��H����^.T����!�H��p{�4D�gd�0�A�%X�z�(�w������d���T�1t����f}�a0p�pd�7��ȉ���dVVSg[�!ա��@�Y�:� 6��>?���2xْOƭ.f7��E��\�4�v|H��o��顱8U�6��@$ڏ+���=<J�Ù��},���3v��<���e;z���c^Z�d�
����3�kZ�EypÞB��zH�ھ^�a���������Z��-ͳ��w��������s)��άF��5��Q,���)�Z��A>�&1��,LPʗϺ�,�!Ƹ�iap���𳲡�׋Аe��̣u�۶�z�v��Yd�!�@tr�_QQ��Lmts����Jk556�a�<?�� Hq͆Qx]�@r�cUޮ��� ��M�q�bX{�
���ʔ�NZJ�&�����j5�E�S��er����c��ta��2�Ӛj{���M�4���h��Z���!���F۠Y���;F��ؠ$~�����i���$�unt9��'�ߧ�ȣ?���] Ԥ�?�
ǢB?�|�)�|n�� ��n]4n��^J�n�DM)�y��!1fv^l$�����#؉� c�I'V.E.�M�fט�o�)�k��������H��C� �ϛ�P�-�ف�۹#:�3�#�?�m�_$�f�D�35��xX|�_��;�������ỦWt�%.���5�ۭ�F��G�j�6��G�A��g:|���[�#�3dro�2�`[@,W�r��Z�o�~�D�,�Z8褥�-K1���m,R��2\����u���FǗ���Qcf�����$���%a��^H	��v����0�,pAl>��2�:��:FZ��v�T�����Զ"����ˑ�����{�����)1���~z�9�4A\A���h".E�De^S>ɲC�W�p1ܿ��؁4$�;�9y&Xl�o��b��@0�˽T]�(揑���*Ih39�:��d,��	X��� �;��`�|�n8�Dؼ��"��+����`:Z�ƶ������5�Y�?`̱���V�J�}��(F������I�宎�e��x�"�5)X�.6iqYx����^
~��Y!�D��&ҕ���h�y܀q	�����aZ|��������r��g�]_�2�bz����oV ���5�H��@����$��7�#;j�]ګ\v���B��uI�	�Ǔ��3���ñ�V�?<M&�h
=��v������e�!���U��)�����%�e*p���A���u�;�ik��A8)�`�/�R�=��=�-̲�QS��C!i|���T<�9����r?��T��'9 
�)Z �=O�>-Ͷt!Ol�j�1(_)�Զ�=��	�;i��ۉ����/��8E jlInb����H&���
�Cʄ��8�]�tCh_\U%l�w�ʖ����Lp`�¦;����r��/� �n�g<C/����ߚYȒ{�8����ϐܶ������b���E��L�+��pK5Jspp�(j��RoY��Ƽ&�>i*����Ɗ
��I�)]�R�8n&)&n}�:�rA��te0�St� �G�}7`���e魹zs�2<�Ʌ�p��#����;$�bS�^ S!C~h�g�أ�z��eYIW�2`����uk�}��/T�����i�VX~ٵjEՙ�0p��z�ϱ;W)�'_�BC��ӷ����ųg�$Ag?����L��e��A��D�x;�xkّޱu?>P�8_0�N�FBVi����:�A�껨��K�4I{����urT�oT�������R��CBG y]�;��Z�-0B/%ȴ�6q�0F�<ޱ&gg��o�CZ?Bۓ���x��gw�^�|��_q�/s���r����7��l{�	��3@��,�y"�^Db�[!�H�T���y�-���F�\b�ӝ�@gOײ@�;=d�� \ͩ7L�Q�@y��DLW����c�?�b��qù�������bu=&w{��IK�]t�q�`]��5Rr���04�ŀ��PhS���+?0���dP׉��
 
�N���@$!�d�Wx�`c��0�f̎�����V5>�kN��2�;�9�<:�Ӽ�ɡ��ʶ���3��zj�Mbo�<l"h�԰:�d/���N6	e�%��#��&�#�Bd(ݙC9K�'�.�f��NJ��͝5g��Eޚ u�\�4�k�s�/�V.:m^-�+H��w=���ݱ^No+Ӣ1�"t�!231��{pE��l�x-|��`�L0\E��K�S(A��Qŗ��5P�P~�&�Yh��{"����~�oݙ[����� �=CW�[�O2	�ɍ6)P���.�Kl)�3��%��n�\���gI|-\�t�@������=�P����5���Ϙ�~����L��S�KB��֢ݪ���A��8�)��_/uIZQ�����-Se��h,�e�R^Q�cIᎤm�g�^�㵓p����or���kM�W(`;�*\^���"^뱚У�|�-��u� ��Su*7��V�&�O�����B�1~V ��s�/[d	�GN�I.J��Y��`"|�ҜAȢ��H�=�-5T�����V��v�-��_n�P8�g�d��E(���m:?g9 ��q[�V�� �
�\�v��;���u9�y"%��^1a���Bʺ��.lr�د��Ӧ�ǭ᎘�#�E7��
�N�=��#
|�R*$�zH`�Ǌ���]ð<c�s�jm�K�h$:<��*>�*��n�����G��w�9i@d��qc� �d��$�λ�xy�}I²����-��
�#3�ɯ˸�"�D5�	��Ä��+����A`����1��,diO6��H�W��V��4;%�p=�z�7TI�U3����@σu��6�s9N��_fB��ys�3�E��LG"X��RS����g�_��q*��xI�K������#d�V(�<X$X+X��O����=����;F�ShM�W�2�d��ő?����mx����p8"�1GT������%�=��J�^%؅B�2�o���n�c5�ߙR .��yD�����@��$G��RV%�4�~�͒	�N@��jM������ʿt��M�@��`��JG�ˢ)��@�u�;H���F�,��W��f��/o� ��,�>eV���R��/8��:�u��i�ы�_�����r�3���:g�FJ�j�泱�V���\��n�,.W��a�2�2M$,+v����6`ﮒwU�&�pD��J,gDG�(Fe��5/'A�����U���vn��PwW�P��zQ��p�;���*ͬ�� x�_Xo��ni�Ené�B�q�?q%s�\G�OR�{��
�2��C> e&cT�[t�q�r~���g�ȗd_����?��}ҫ�~:��`�?�DʐR;�����.����t�c�ĝ� \�JF>!f�2���*�mx��z���Os*{��?��$��S ��S�I~顣|2�
�=[��0s4hܯy�s�3�����x��ví7�X�`����5 �/��>�k�\�)��7$���X�Jx���G�x?�/��/A.�:�;�e����6E�)?���Gt��z�Qǂ�
�P�#��ٿ�:$����o�_�fd���A�n|�"�)����(G�3��V���qL���`�ηx�A�F�������w��"Q4���:94]W&��tY0Q��t8�:�4HAZ�TG�#�L��?[�=����� ʵW�N�0N�',��z\]�`��'�!�J���%�~�$ c03Em�L��"��0��a�;�M�?n]�isaz�z�����}6���G�������9�9�����l>��c$w�!l $�1jh������D3����룉|�be���n**�a�z�	A��?�y�b�PfE,�9��:��݄����4�׶i-Y.���}�L77-���2T��0л��~E�� �M0z+]���+��@�9k| xyV��s(�X��U�-ΟuA�.�.0U��A 4:�&�1�:A��zC��BLeJ�pc�Z���V��ⴷ;�������q�,د��P:7�7���=�_<|܏��$� �dq���4�e��.��*�{@HC'�n�C�������+ZA�$��{o���5Ɣ��������E�^S�лG$���M{9��I��Z܇����ЖN7�\)'8�[:��� Dda��9�,5Y=ذv7�>�f�N��W�����4�R�b�Y,W]�9q)�ި�B+��)_�H��i6HsЋo��p� �0����<��5S#�!z>����jaK�=��j����X��7"�	<�%K�̣BI�E0��}�64��(�A@�Un��b��g�&��G./%�.��I�w�#���'�W�q�٭�,���r�`��~B<��������i�o�D+���s&���V�祍��gr����{L�*��7c����Nb5�w����P�a����b�4Gn���ݳ��oi�/c�m��!J�	>��ڒn���Dd����z�y��y?9�~s���'���	c��-�[��غ��*�������1Dc������",� ��Q�]�>a�NT�9^���v/�5Q�:��d��'jb��e3��6z�L��Mh	�c ���Av�#��W��L�]����%�,�Xd,1tCɴ�h���/{��O��ETI�����N�e6�58^e�#�k�" ̕�Ȋ^�F j�A���=W��.�*��T�]�F(鍸xɷ.*�zdԣǐ����'��*۳$'h�ǋ����7C����`�P3�9��V��C���ͰpW�l'xoDF?�N��L�D��a�����C�E3�C��߼+B5?Z�����c]SP�����u���S��*qB�����{3٨�c�Z
z�\GC�[/'1ʛ��ʺ��k�������/�wך�FS��M�7w�l�z i�m�,��*���Z��u�V���aǈ�Bã��-gB�'9�UI� J6��2zx⪗%N"1֘��;i\�̅.�윜��{��)0���� l%��J����ƕq�;o/Gȃ�OF��������8�VSJX��C׊DI�l�sqqDn���V��^��U�+�@Q	6�J&�1X�;d���_�ZS5l`f'w�3[n�9��U�(�����HS�P��:�m:6�qE� ��Wӌ;Cf�(���dV^�v���mp��E��=a[# �� h(f�n�`���b��l�`�������a=꯷���t�:��Q��<���3��K<=}���!��=h�)���$r��f��1�(Œ�� ҥ���l��
|���C8R{f�������m".!Qu����*'���7��5�`
s����ۃ�`%�(�JI��N�K}��(�����N���-C���е�|bԗ%�am
��㛒�F��d������ ۟T�&z��ӷ���r��1iPvz��'j�E��}�j��P��[?���������Fᚬ,�������,�k �t˅_.b��q�'�� dՅo��$~z"e�!��aZri�Y�J�K0#b��*V���*�Y�a^[�I�woWN/~pcY���~�b����u�[q^-N�S��ѣ'����r!���"iS3{�{�DՄ5�S;B��?.�b<��=ORε��:��d�# �ػf�)A�g�d�%�cR�)0���G|.��x�c��c�w���Eۭ�W���n�h�,�/�a���̘٨�kJ ��6�U��vDh�*���"���_�;�nv.M�@�&3��_'�T�T�R�ѻ����t�8�;�b��8a���©i6cʜ�r�N�\"m[}ⲏ�=�x�KF��yF��v�8����H���/Q��|WZ���_�|C5�)�B	���=�N��Я@CH���Y�e���%������Q[+l�%�� w?�v��jb�x�����v|\���nn���C'ǚ� ���������˪������~�ZEN�l��H��2VI��-��f{��h�mQ�A1�uj��@��P�Ccz*-�j%��ؓ�Gp��d��I��ؐ"��6��U��8�.^MC��'��A>a��r#� 3c\%o��9.�!��V5�b6���}���͇��MN �K� ���@`�6�1����o��<�s�Ϡ檮4���7���_�;��Z�qn�>N��:R_�$`~�yv����jvU��)~;�G�hN�2Ҷ1R�O׋p:w�|?�[����6����^�����®��g}����qO|�)7\����<���lL�J%��<N�����"A���
}�ܼ�jc����kSں]��� X�vΝ��H��,zV�0��]f�h��аԆ�&��o��ɞ��*���K�	t�r�V��F̢��FIl�da�Gzv�c�B����3ټݣs��Q�Oտ �w�Ak���$3��G���ź�~��[�%���� /��TⅧ�7R�|��J�No����V�!Pp�XUg�H�)b[N��
f~��W����x7��h�O�9��0p�nmMM%Ь�Nq�E\��UA
4o=�2FGiR��º��LwBЂ�l�� M��g��r:�?����B�_î
��<�(u�$���d%��[mwZ��@�K�{k:'z���3i0����yN�2�A�J��)\���ԕ{�*Q�A��X]�����n�V-���R�1�͎.AV�ˈ����b��m��v~nv郇�m�`rI�⍓���ܝל�$L���Դ�j�ET�G�̸gVf,�d�Ε� ���B��q�!=m��7[�Gh�4�	-Զ��#�+éJ�:��7/�����sBr�o�S���\�,�����g�֌S��;���sn��'P�� ��D?٦����0�d0��:� �--jt�|��ҏ4��9A�n����Y��Bp,�j:�F]y�Y�D7�6�
t�X���|VnHO�K�f��(̭}c�Sn����3�D���I�S��h0�u�RL%�� �jv��MՆg�v�o��	f�p�]��z�h�&����5ݸlNZ7L�� �A(>�����kX���o����-����P<l��_��1��9F���%6~��$�CD|��e�X@@���v���[���h_F���F�L�� ]Ē8^XJ�o!�u�eî޹,��'|Ċx���G�Q3��RUB�F�	�8���Ӵ�Y����s�-90L�ٓ�c{g���?����G�������Q,O�9��~��@$�:����=V؞�Am�����w��}H�?C!��g3���5�;���=����	#z�z�g �_��F�7�;�7-�_�"�s$�6<y��4ю"��r<o*9�)Ѷ���2C�R�3�t���yb�&e��+N3_��(�u�
>@۵&l�	i��}�>�QsF�� $�r/.�q$J=�}��k��QOĊ�eb�KǬwLB�]�NɊ�R���� 2��R��7�:���5�Jռ/�f܎D��Tn�Ip�e��x1v1x\�ǿ�ףM�24�_�]BT9���ǂ{g�#����
�xD�|�ݑFz���u�,E�f`n�ޝ4��=ځq�H��˭�kEC�Q̛��N�W��.�mQ,M�o��Q��_O�B����=�M�H�g�M�J'&�O��e�N'�EX99��tfU����9��r���V}���.t
����Fg��$}w�V͏�L��[�I��Q�.��;�;�l"��T$&��IM�P��l�)M�"�`���iL�gP�Φ;oפVq��iN��uk�	_x\7
����2��E�)��4sf5AA[��?�r5b�4��hR5j��=Jl5���I�(V�3i��k���6���5��\�af��7��0Z������b�
qs5��4�}2�M�J�\��<�N��X�!z�!�\�s��G�s>�0��GQm7�?���`#�[����w�(�%"~(�B7#�d����p��P��9A���/{�(��+��4�&��q��=C,\D���[m��7��sK�]7R���Ka#��u�s�N��8���`����A�F��$Xգ|O�Q�d�>-�h"`G��;�B��d�����ý�ޮi{��un%�vQP/
�V�����ߊ�PW�լp���e֩�!0�e,#|A!��.,��g�'�������#:�,)-�i��m�_>���v���r>eʽr�=���VV���ł���U������̶&����(�@�Q�c:� ���;�V�w�R���� �Bi��)tފ^�L���oޱy
�qt�y�*��BPJ���nkwS	�ف�[K ��܆�\tK�"�4Xrزo�!��`�Q3���\�'��)����V��~:`�|6�$q�v��`%S ���n���Y[Y��np����7��s�Z � �TY!J�<� �w���UGl���֑����`GQ�0ی9{l%��^]��K�v ���R����o���Է��ظ������Eڀ�����.�?w�/*�������4����|�8*��ԧ�M���gp�J���sѹa�Jʔ�#p��1U�|�3	m�����u�1͐���Lۯ�/�����v�(�c�����B	��iE5�x�<���M�c01�4����zl�N��?��vN��h���������%���r��s�x��Kw-��{��F%���ls}��q������)IGne��jp�@N�UKQ����m�59|���W��_HtNN�<uP��J�D\�g�޻y�un�a�"��,�[���t�{3�1�)�7W~�Z#W�$&���$ET���/�=Wm��S�)P3�t�F\��V����
�!� �Ѵ)G*���]�L���x�M7A��n��썟W�&d�{����3�ڗ����2�C��>�Ϭf��4؎��E�2�4EP�᧑�η׵�� �r�޾^�gt�����X����y���@d�kV��>�r���� ��k��!�/���c��MY����n)��N��z��r1,J%8�����#獃�r��:�vu��I�{�L��U�ƌ�#+���!!��i�6"�:�V,<z��1�K��z��2���a��!�y�!��F����Eξ��k3�e�呥�js易�f�hBv��ᾃ	$q�zt��\�+z^V��BI�( ʓ�dр�o�:h
�n��i�$�{�!���(?	��z9��E�E���u�h�����&�c���Ja�Ǔ��p��y���0�"�I#@�tD���]�B_B;@��WȶbK춫��ؼ�h=�7�]��J��u��v��Ft0]s��%(�o��W�-� �t�����pr�|��x52P�-��Egb��(DB�Yp**Gm���%�QHN�0D��B�W�&��9�g��Î��&�;��L��0&[�j�y*���;�����Uu!�4^	�M���Ie�@ϰyo-m<Հ���<�X�T�q�y��lv1Vt��B�0���ק��9�/�pZ�Ɗ�:6�h`\x�9�[ޕވ��5�'���0�搐nld�������c�	C.���y��5~s痰�m)&�K���;OSQ�R�Q�u�nֿi��6iN4mnS=��{����8|(���,��=0ʱ>�����+2�f0ҩüH�^��~D�#v��O���ņs��,�%��?Da�{���&��IB�O!|�g6AU�8qU�Py��pr}�lq�_&��4��`ڭ�󂔀̨9�x�_p�x9�;d�χq�e����h�C�/&͂��t�ٔm��ҿ"?���,ۀ�����i�W���,D�@�k!��Ql��5�#��9�k65~������Y����1��]
�$��́|~hm�� @z�=���1�m*^q|��g&lD?����h�*ӳ��+\c���3�NW�WxЉe����iM���Gn~�w���� �^,��>��~���`Z��>:����� H�)��11^^:=�2��H.��C��>�璈�|�v�i���뗻�x����0��Z�"�
y�=x�& a�Vc�y\��q�9�v?�r�}�68�b��[_Z_�ьX�tO�Cw
f*g�Z�[�t=�dp��
a5��uu�z�@���לK�=��r�-� ��.�i�*-.=b���w�wU�F�.[W�E)�[��ə׈ӝ|�=��3\�Y�@,�����`��������ϒ��$��P�ԥ��d�i�Z�X�lK-�`��p4,� ���X������!j�����4�:�-������?`x�B�M�%#Ԅ;i㲊��HNw���%.�3����ø:6<�]x5�9�4X�p����|0����e��Ԋny8���ZS����t9�X�xW�t��>��&���P��9�;oǇ`��iF1���ð��6�8I��O�7`7s^賙î	��M��U��G��j6�S��S������N�j��sɁ���c�n�Ya�yrOUH��)_⚁q�ze/���p��X���l��j��G|~$�;!��0~��vC�a�����6`�S2"���+K tw�L�(��!m�����/&=����YO�b Z��`�������,�����hәc9��Q��K�a���t�֌�}�C�V�'k,Lʠ�h^�|b�g2,�����귬��,�\Y��qKJ�珨놙�skZ`��fdcf���#O�aE#�5�j�M_��8eT!n�'��yCڰz�cL��
r�s�Y�X�����Ә��jG)8�B��.�M�*�п���(��Fڵ!�`Z������ʌFˀ�9������Tnt�A�oˢ�~D�"d�o�<�M�$�Y��fU��Q�`QmF�7��<�Q�W[m*ː�,��V���TJ��KC�5.��)n�M�|��	[��G*Ϧ
?Z��#uK�𮹰]�0	�P7��N)�J�s�×mV��_rLq�O��K_Rff���~:)�Y�l�s~��*I�;?��g�^��`�����u�=p&!u^���E0;D�)a�z4����r��������2.s�+�n� R��n�y�Ò���#�Ͽ���.�0w�H�*�-�Z�X�����J�ο�B%Z�gu~��!��嚆��0FO]�`�Q/�����;�gH�jԆT�b�;���b���1�Db����J�^�/'�9A����%�&�P횗�����d+�*����u�y��2���;�k�⻕쌽���Gb�d����s�"i�7,�\����ZÎ�Lu��EDz��p�o��Ԧ�/w������s�:�$�E:PU��:�7 �Zf'^�J��(Qh��+��0�T<%�����<�bm�p] ,���l�+s+Gy�Ƕ���Y� ��;K
��/�D��V�P�&3I}��~r������^���Ji-���?���g����H0�Կ�� G�6�O�2v_��w&-\�|��˧�0~��H���S?&����۟�����X��Rk��(A�<�F�eڬ{tvWh����N����g�i�k;���1�+l�`~�J9����S�}57�[ ��л�wB8r��H{����&�Y�ԕ��~O���{��E��Ȼ#�#���]���
�B�Aݙ���cI�c�\o��N��PE���%���_Q�-o]'�N������P��$�P��r����DFr@ɝ������}Dѭ���|?��	G�j����"V����ˬ���l] vF�]��j���|}�@�H�����M
l?_K͚��I�s��)q���y5e �:�g� �pK"l�5��)�wgA���GLa���h�T�Ҏ�k7���z}����@N/E�rV�I}8�.�8��&F��M�h���v0f��`?֖���g6_s�_K���-����b��S�� �ɓ��K`a�c1"��3���If���� ��Fay+e�\�׾�@S�������Lp�Nǡ5���~����������F]raB������[K��=��3����G��s���J���o�x�����,�"LGWes���I�~�L~��ܭR�}��z��T$$�2}DPK�lJ�GI���J'!o[�y�{؋-?}���[m�e�YI0�fGE/��kE��Nfp�x-D,ot�0�L�$T+:���r�c�Iq�R�Э�,Vrg�j� �ϭ�V���-��G��?��q_����gKo<��}��&�����Sok��$X���$�H�]�02'����a�C5�)C\J�d=x�:4�Nݤ.0�vDs��0����r�~�h�؜6���/�������I���!�4N�"3Tw+�	0����R��E���j�e��Yeq��m�1YV��Lh��4\�ڂΦ�Q�> |�EFj)Y�mއ�f2�1�h+%1��(�+lZ�0.���7�������x\�DK�iwC0 �ʧ�	�2�`#A0�g�j�B.d�o	K_���]k�q^K�]�y^;�bV6|F����Y�(ɑk�:�9y�M�kҥR��0�Ue��S�_u:yE�,f���O�� i
���\�u�����-��ӌ9T��S!���M.�zP>�aj�µ�]Q���/R�F?@m��,s3x}�զ�<��x3��v�:'�Ɇ�0-�us0"ъ�PB�ﷆ>Ac��QE�����������!��u���&��6��� �7�˘�+��8�>4���PaEC��?�RO߶�\|Rǭ�
�	lFl�H�p x�����K��-5�9��>S�z,�5x�*J6]z�º���a��!# {���)k��mt2K���C�H��U�G���3@�譄n:l�8&��d/[��0���>�-&O���[J���k~B"�m!�P����g���uA����(j{�u�_� �I���~�&c���&6�v�����i��s��5�>�$v.I�<A�wI��Y>��w3�4'��Ş�F ������B�������6S�nn�n��t�jP���)�&�{�MC���fb`1�b�ޅ���+����}�����tȁ^���3t-�}،��Cz�R��t�{ }]��Ҫ��^C�O,�y&�ğ��hJa�t�sh���ݳ~`GЀa���P����h�1Ȁ�gT?5��'K�����x��+����s�f�W tWU�����K��f�3��Ӂ/���-e+lK�QK}B<`��D�̉�7y�&檬�4��IWzڕ�g�����91zB)GF���x�>0�>8LW�o���hA[� ^>��L��>sN��P��Ǣ�>i��i��{�1=nrBe��v�� �s��r�V[���m<�X�g��Ԩ��E�5�v��a�����&��3�ط���� ��s"F���<�3���FB�R�dG�S�gc��@��cR�8*�ú�Lz~�+4��)�s֠�OQ���X'P�vZ浍��Z^&)�_�'��3l-�:O��
�
��)G�y�������s�����0�\�i^���;Q/��*cшn]�&��&��m�'���1�&��H��K�|࠘��>7�J�@Q�	W�N=���v�G�MhI+J~�M�Xv�{h?���h�9�)�Ze�`��T��u\)b���>�󍡆nB+,۱v��Ի��}���`��Tȋs���V�$�&�2�h��_jMj�	�v�ܷ�v��M ���׾�5�L���q�Bq�;��1��/�`
Mo�|P�$9Cʥ�$DԁGˢ�v�^ٕAly�W��d9��܍,����~�6[��[R���+}8O���Z�ML͓�Q��A%P϶�
���x�c��WG�$/u���w(۰�/�z��y�:�.EI	<DYB�}�d(x�e��������](��7G���Qרu���|:�&�M��Qw�����Teu}�]�z��Zա�޼�ށ�A����vKS�5�$�@F���T7eL���,�S�_v�v����D7c_�h��3жh�C�hG��=�o�5����Ԋ)�\�{*$@�����~:���D,F��<sY:�FV�i{.ʏ{�pZ%�k�Kp��t���h9\O���=�<�P��I~Tb�����,��M�vg�]��$�XFQ���iO�����GW'�ޘ�6��sMy���ȁ��������c��m���/�dT%�NL�Xkc~*#n���~/�Sl�)�.G�:���
��W�ը�fh�X�&!��bOB ���>�50�����6Fω�zhaI;T@%�!s��Yb �����O�O�Yo#q�����]ly��IzY7U#�>�#��_�Ja�h��o2j:�a)
���c�y�Fڒ"�@���`���BC�ޭ[LY�M������.7G���M� 
l;�6��h5�������KQn�__$�Ph�Jk�=)�}����a3�C�
�@R����amD�����ˆm���1s�!~�p]-ꁦ��un���m#�}�����TŧF̖D��G|'f@�Ր#3�Ro�8L��en�����*S�7j���:���s��\�ԭ7��ٷ�����<����1}�%Q����S0��U�Ey/
���;�r`Ku��I�u^�2:'�<]�����C�CM���菬�����(�:��Z�H��د�9Zn=�ر2'���_�9}�+R����+vQ�{��.�/!��q�Q)�g�,�5h�!_����D��_���S���Y9TC��jt�J�� ��0�a*��/�p�r;ݘ�&�?=�C�k�J���.ŀ��:0%���Rh`O*R�,�&U��GW��ř�\�����˒S9�(t`���С9�W9����v�g!��A���lݓ��G�i�G:���[a��]���I�+�U���MgC�]�K(_,̞w��;R�tm�(ta�kV��m�uEJPv��82J��p�cX/#��I��,����upC���<��OʩӃ_�&*z�GX��6�����6f����~�\�y?�?���s&��J ��jw]H/o#�l�_�|J����*b����������)�ɶ�vtY@�$%b�W��X��+�6�9���C�R	͘���ۀI��/{��%#�W����r`��$���1_�XZ�7Rk��K(������Rw
D�4
���Ŀv��Z�D��|@n�	Y�?4�4�l�h����7{q�A���:�9шiM�WHtoz���PB}���էr�)�k�\_LL ���3|�ř�&Zi��9^n�׳M%��w��(.%~D��H�(�]������!o������|=�攧t�)��_?��6|G;�A]��:�7k��kY�Ej��t���c��h�o0b��1����$6?���w�o�{H�Sʫ�rU�$?�.!�jb䪎Q�W�^��GE'�`,�LA�̊ĥ�zqe�$H�I��zR^���a]<
S��c��)�� 
��8R��{��JWd�jme�z��`����ޗ�X��� ��M�H�v�r.ߐp�;�����XUh�z�z�`���~�0��i���3�
Y��x���n��nڰ����U���z�
��.z科�W~�6�J�eVA�c/`)/�Y轣Jm8��`�"X�����Hg�:���*]'���s��qߏ>K)Q=�]S��?�Ҁ��لX�e|t��p���q�#��%��1�k�Eށw��vY~���־,
8h�g4��P�~�5A�f��C!��x~$ۑ;G�^��-��8�TJ�]��X��U��+_&�;X�T�Xo�!,W4'��c�Pu�fuY�GX�_d�2ڙ
?3�f�L��.�!�Tp�j�ʛQ)�Έ�E�ɝo�3Ν�X*�X��9�hqK&�.x�kc ��<�j�#u`��Z���G���M�Li���)��!���'�g���M����=��?�n�GÆ��:��i7��}��qNH��1�ڧ�ϡs�BJ�,�����EO{�R��˥R��}������ؓ����E�㭮.�ER�����9�m�c;�#�F���ި@�!���Eh4��;pw�sP*q�?�w-
����繨�h����B�ӨS�քi�-+�roD��F��J�kl|�dp�#��.h��v�ڣ��#�F<�[�H��n\����/��}6����x겴9�1o�s��EZ����噝��VZFU�]
ߟ۞�AX���ç��p/Fz"�����C���΂���\9�1�r:gA�)Y�\���3DIy<%�~	���o�wMw#�����}9o�ȝ���T������a����@���X�[K<u�yhΑ<2���q�m�Y+"��i|�~�)��i�V��Ԉ�p�v9o�����P}�2̴��r��޶	���I!�b
�&K63v��)�C�%�jsl�7k\�
d�[|����[�$i>1�A�����n�}"�`�e����h&_m��nP�;k��k����]���#�*O�B����;�9�x��ɾ���c���;ZU�h�j��Aާq8Pz��4�J}6�K���A}��q���rB?���spY�2�g�S)���3�q��@~��y�s_����78�e<ݭ9�~�U��j�EJ�:�0������L� ���ҡ����e�[�IW�M?\q%r5�L.��hx�Y>b�4�y]��O/��N�l+h�m�2X�2�[�}cKYe%��k<2l��M��Md.�v�+�9����ڨ�P9���D<'�N�ee~���n����p��d��Q�1\����F��1�I�,�ϲ^O5��%7+.��g�:a��_\፫�]\��C
��*��N+�I��:4����%�gH�dHLE�i�y >6nt�F��е�XSDEU�V�e�3�q���<o��}�Z"�sbB���Nͺs����X�������i�����Si����_�⽎�"v8�e_��%��c�/�6I�"����ae��PҢ���u������_ӑ^����C�~� �g�q�<v�q�$��f~>:/���um5͙k:ػ��R�m���fZ����aW�����e�ɀ�X����Q��zi�W�!5团����Rϱ�ݲ�^��Œ	���f�ژt�4�J"Z�]���-�|D�	�hD�Ҧ�k��Q���-C�q��Ҁ����+�wL݀��03�1>��o3�N��X�D$��'8�^6D��Z5���/���|��,�^��t�xU�Vq�7�:N� ��)Ŭ��Ր��ǖ��y��y��Nb�.��?��ҭ<�ʱ����:#�8���q����+��ԟ�Z}��:B��'q`��ª��x������I|��ٌ����Ѵ�Q�sr}ܺ#����2��{~ISA$hٿI���փ�譏�t��pj2�Fa�"���B����a4��HoN����'��S�E�l�q04w�3>v��S�T��9_�G� ��pΞ)JO��'�7S���m�﯇Te���8XJ)�p���
�V�7@�?G�L����sQr��-M'����0"=���f	Di����x��;��b���������؛��n\�>)6���`�ZVP���|�M/�R�h"U�>գj����v�v����R|k)�~~!:혊��/�i)JNτ��Z��/2���ll9B�cQmvB����{�꦳g4��4��8��9�x�k�Çu3!x�f+�3-i�U��FZ�uO\Hn�o�����`�AŇpp�%��CyS�
*bGͪ�TrC�%�H�b��C]5��#]]�
����HQ��;+�0���:����C�YQf7��G#\�t��45�G�P���J�<�����_m�<��I����	�fP�P��ay���1�1�|�p��G:J7���HC�8���]<��7�P{���{�K���1�Z}L����2���Vcq����n-(O%���?����D'�;h����=�:D�Cj�_}��N	�مJO�W'`���K@�w<)�Q���t��{Mb�9��yx��tI���}��*��/�����ƹA|ۏ�!z:�G��cHcj��09{%�R��g/g�7�!�6I�bTTh6�i�A�e�Rt�Ծ�`�����B���ۅ��`�0���K�� �{4FsP�����R�e�Z��
-�*��R���6�m�L���5a�d�.nZ�z� I�H��f?�O��'U1���B�HQ����7����~�T�{Bs��VV��8�?%*�D�!ZD�����V������I��q���FF@�gF�Ç�*���DҠӜe�^{�x$�)#�Ф�N1���nt��ԝ��T�s�+��8P�M�1���e_�����Հrg2��AX�ZZ�U��`������$J�G�'f#��MI.-uz��<ߒ�*8P�$~`e+X �|_��nx���:�\��B]�J�F?���T~+�f��7<�16V�}T,���:"���{j<`���*���ٔ]Y��3a�Һ[�Y�O����+�\��A �્iµV���G;Ծa�eg����ܚ��r�<��,)�V��u��g���*V����v�"K�)!	�dgQg|-+�{mL[�;�-=PK��P�ζ$ch�T!�bL� ����qO�Tu�|n��q^�7����	�]��-����xb�{���J�o��֦I�z�I*F��o�T$�K��ɟ���F�k� -�X��6�-6��n죄������`v�4/��� ����4�� �S�~��?���q��j
����������8�גRA��oCM�鉴���]�����NWB����ɝ!���X��
�e�j.���֒����3��L4�쭢�o1�C7W� m��o��}���s�q����$�x�WBE�|�q�lƢ"�j�r[L�;v�!7��`�5�?<ޚ+d��*_l�3ޟ
q�CHK�@�ݠ�q��tF�}_�ݐ��w���lM&B9T�l<�r�9���q�[j��mqw��2τe��Ė�%;~��'�H��l]�}��CZӮ~��4�8·ov�פ�f�$ޥ;,j��<*տ��$g��Ǿ�}l���j���흴�T9�8m���+��?ݾ��A�5��>�����aLR�QI��6i��>�{&��"����U\[�6���q(Oõ{K�b�Y��yd�~�{�'=�j[���0B�d&'v A�< %)Y�'�x(���J%��<�RJCF��LE/�ײ�u�l����Fh���z>;��I7���c�B���F@'P��z�>%fW�� ��Pk�N{��C�V�u�f/�K�����sl	��Ԋ.��Mi^+��;&xe�x[2"`zK Ԡ�π9`�6��RR̸�S�n�ϡ�,� 4X�j���+nM��Ѿ�P��L��RB�d~�V�9�zNM�� #d���?��Ccg�X6�'b�_�����l[~X��M7ܴ1���d��k�/߁�)�r¥(r��N�v�S5�p��.�#�U�.6𸇁>"A<��A,�����aB��kI/��)�['���u�V�d��R�5�J��?��P~g���BF��=z�l4�HW?�<�>��Y���K-�f�Q�Y�d���3��A����(H��rk�n�IR�a�FTPfD�Tz�V�@�m�;a�u`qN�~�Q��	ܝj�rn��	�2>����E-��Bs�4�ջ:�R��CͶ��iTʆ)me1zd�E�#�d����^*����U07�T Ⱥ���F�|D�#�����$�tG���O�$�<�_���?F�]u���yi��D�6'����9ۄ�4�*7�p�{"j=[t��i�Z��#�0�W��\;T�=}G���\�*wA�\:ӈ������;����Wa���^J2����-�V�˺ �LF]����w�ߩ��-it�2B���^X�*�j2NX��P}"��GŧтZ�(q�ˈx����8h3��&���q�l��Wǂ�wt`�9����$r�Ġ<aХ�ђ��#��F�Lp�K_�&o;�?�k�۸��-r�=�)h�0�Z�`��߈��/|� E^vA�R��ٲ�����7��Hf��|�N��2Oc
�,�)��t��р�/�撛�A[H��U)"�5~��̛�d-����� �)�� в���N��݌�K�!̕��A�X�m,*�S[�����`D�Z1�U��O�D�޳�ce_�v�ш.r�mm�B|�g�"��y�*B���ʿ�n��J�|�ZI��u�=*�c���r���(leN��J�H���w�2+����Wc�0��2���9p�յ�+1�/�;XO�e�e�wE�P����S17q��ǖkb�(춛��""&�O<c&���8�W���w@'��`ҁ ����9�(��%^S��2)��gARc�WZ�SP��vOA�Q����V���{)�	�?��3��Ge �����::t�ߟ�,p"��qq\��n�2�×(�.������gԯ��H>��F"3��k+�9���ŧE��Z�p7��HO� M��Ǔ�,�>�Z\�V�qv3p��{�A��|r�i'�&���_	`�*���iS�3��@���/b���q!���
� ��h蝵~�-�%����VV���+���ڷb����5��6k_�DO�B9��)<���>����͝�d�.�W�1� �#���zz#^勺�)F��¡K�є��-�IX�*j%_�ί�*c�
��������q����E�w�M_v�?<�!-h;��u��C⿦�ᖛ@����٤�n_�t��'΋�.��MZѰ�	$�`18�vnx��aV�(�i�ǆ%�j)݃��K�0�S�Q��Sn��˷,N���S�
0<N[Q�j��d33�� Z�ĺ��0�� ��Bդl�[��1��[�~����
)��X����瀗��}��2���������2�2Q���P�;�z$jP!6r~3k~���?`5����t�=0c�RĪ�m*�Q�P�����t���T�v������׬S6�EG�Lď��V���������)<��U6)�n�����w��,�Ք.��Z��ɒ��Z�.�ߧ���6�0s+9�p܅#W��a�Nۚ�K ���>�2�eW��Wc��p�� ��	o�Z{v��A�� �[�Ω�@]!��=�}��Q��Wr��lQ�������0�7�n>�1�`�� ���o��`���K	b|��.���I����y�Ӧ�䰫�����bX"C�,�r����@]�����NeƜf�MN��頢m�p9��z��/|�޻�|�"�D�[��"��p�o�!�l���9�<NX힡��o�s}7�O?���L��UrΒ2����������RE�����g�%�[�Y^�E��`�O�,�}H_����<X�CO
�~��Y�>�ۉE�7��ap6�(�;EY�S�4�����N�Nw6
h�ƳQ�A:�I1Z0��-l��T�Ub�v�lˁL����̰7a|���f)�S)�z,���κ��c����`�Q2g�Mc����'�,�d��\���]F	=d.@�e��f�H7 X_YrO�ye�C��1�~�A�2�'�gr���^�O�_���,��
���p%�XL�;k;U]�R��05��M��˘����oz����I��������<W��F��5�ce	�v_��t@xc�������lU*<bI�I��4� ~���DUK[��?^�0o�}A��P���j�Z���`Ӭ��q6'���ix3M����n)h �I��XdT�������=l1�\���椯o���i��C�����O�0�5��2�^5����ی�'��1̖w��T��^E��S�uo�6
����lQ<�Ho�y�l�	�O|�wY�/S�a�a�.&�k�ԙ�&�	;X�H�E�t�X���^Y-��������<Z��n׈H뤴�ֽ�<�&P�5'�~X��������
�u˚K֪h��+T9���0����J�nϼ	1#�2���Ƞ���b\�����ULs�Y�F��*��A�5z�H�Ѫ3�� �M��~z��'�y{t8��@���q��c��o<_��ZhŤ����� ���xR�����%�;�+�T5V$U�r���fo���1;�~�x4/�'=�r���b&�L���7�?��f�3R��$B�d��J��"�By*�D:������:������f��3�����3Rq��7�g����#�@��cgl !ߔ[YA.mS��e���@=j-@n�(�}$����WK�OÛWf�T]�=h(Q_7M��b��l歸'2ù5X��*��4?���F� ����F �����u)���� �F�	�Ol�}�4���d�#_���!v�;�@��/..��C�G�����hu$>�y�'�?zFn6a��ZiYgƗ_�%طԔ�p0
�O�J%�w߿�Br?�
4 @�w/���m�$C��At���[!���`��ǡ\�_`\���]X۰�(�5oR�q�r/�=-黶q��S��f^�r��g��k.A�7�^�nߚ4j�)�y�t��DH��V�I�V|C��A�=���Hşx�{o����<�8l��M�ē��/hƚ)a��b��Ӆ��Fma�r�
�\��`����c!�!�c��K��}��;��3�#�^���肻7��/x�i���,]P�k���}�e� o ��t�����vĭ)>
�R����Y=�����<*�[����ԕI��"��
:����&��s,D���u(��,]��W�����;�X��Ϫ�~L���hj�E8�j�A��Dx-rk�A���P˴cRkr>F�y�Y�}>nG�q�� ����.)������P8�`Q���q�j�4�zt�?��+y˄h8zcm˓����oҪM�$����P��Wa��]��zr��2�l�`��Z �bgk� e�/.��XQ���a<]n�\4����+ˀ��3R���0�DO)�`my
�>n��x�TC���T�ߊh$�aV��A�p��oQ`�-�y#��z��"����v�]T��'���3zz��|{u0e��b���S��}Le�:6�&�IP�<&��b-)��&�������"��#�Ħ�2l����R�ea,���,���^,zH��ż,'�i���������F�K`��ɐ|OӤ&����
��l�b�l��������WD�ȣ�]�Z�*n��.H��6Y���nk��Y�� �Q�a��9�{h�~�r����%�7
Ȗ3p4����f�V����@#��PC�D��l�ɋ
Cо��o���L��1Ì&��p�N�T	��� w��E��G7�{��rT�c�y���z�4e�3�B�-Ҙf�\�c���̤��r�J��R��=�8�4&��n̍��C3(e��0!v}�sV΄��Z���(�t��%-c������|/EC�n�^���6�Hw0�TY�N��BE�W)��۰_�L/�"z�J3�������Q~I'�<
i�sø$no�dN���w�����bSs��	ئN�=��V7PGwl)�PL1ܐP�}c2$Od��%�<��k�K�H$���N�
��8�xt��R=Ý3��wڏ��>XPh�ߩ��%+=��u�6��|@ �fFuV�O�,��Y��K���^du.�hu%n\�P'̚�mqdߖ�L�o�gU�������T��� �R�s[i��Zè���Gz�#�;*<C���g���d���2g��b~x���}�A� �|��C���y��=�^�P��eA.�\��*��,��h\W��3��@��a,?�!i��|�ΪO8���DJx,�B���`��Y9 T�l�IV[`W�Y,b����ܸ���uJ��Fm���m/�ձ\��0v�|�\2UPF;��.7�l��W�L(�����+�� ����
��Ѡ��3�}��I�?9~���ʞX�ϋ�X�F���
ܿ��s�漜Ǣ'-�"���z-JA�H%*�4��Jˠf�\��\��VB=	�
�9=�o��}X��@.B@@�tś��~r��F��}�li%�5���(�/�9�uX��Q�ClJg!,Sm�II���
�Σ�[*[���~�aT	"��Ez͡�4���LiU2��f3]M�4����@N�=�}='Z�'�
4}�NRi@��]v'�W�u�?�MO,j��"6ge~�E*�w���_q�^��`�������{����K=�����^9��(\
�L*Bb�J��e�6�.{���.��h���,�l�۴%
qح��`��Gs۶!��E�?�~��k{���3i
T�6E�&.Mp�gX�4I��ֳ3B�^r֣z!]�=wFy��޸̋kzi�W5��<�G�@�T�a�u���'uU\���zH����3p8��~3��9��Ữ��*�
��N�I{��� �2�A����m�����bzl�P�y�R��C���|fm�; �ON!�A���!�W{+v�U���q��|�UKGxé4�~&�O&�H�����9Ai>k��-�/["����¹��j[8��Û�)d��|�@ׯ'�I0��$EցQ#/�.7�AYb�mw5��U+�7\��1�F����I8��Y�����ç����,�.�^��P�$�}��������\�@&�ϣhtXd*J5"����3T��a��	#h�3��P����/!�ׄ�8(835|��1�O;�bB�0m�Z|Д���� w �z+�Z��*�C�:䷘�
�ATA�J�*�j��Q��7`x���+��N�ڭ�;%=�ȣiC>���י�7y�9�dY��g���U^��ɲ���L��p��Z��6,'��ob�����ƴ�J�6D7�ۄJNC)�$:�f4j`��k�W/<�V\*��6KtÅΓ��z��kxm&�HkX�.� K2)�i{��E�n��aH���5,x���ޑ�� ?��·��!W�%�vѫ§Z4���a),�;hei1գp8�0�\�z0	��~�Ɛ�^:)�OF�45n}6�5��w��;��5yjA�����3y]���ZPU@Y�����ع��R�%� u�g���a4B�;ߜC�(�5s���#J�M�E�ԘV\������ȲPޘK�ރ���}H��-����%u�h/��4�ڵ#��!���L���EW����ʩ�t���%5{w������G�Y-kwq�;��xU���A[Id�����kc��T)�㋴	��e����:uR6u����^�|"���T��}AEt�{�%o�#˥�=�9K��@}yN)?��8��dAn����*�mn//�T�
���6�p��X��N�������JjAUm2J��X2��U��b��D��2��p�n���u����ǚ{-���=6��,qF���;	~��)�{��"�\�ҕX�\CA$`�)������{�[��^GDT��NK8��4c���:�5cR��ax���A6�ΌĆ�>�W`���\E�bB�,��@�"���[&�87�]��D����T��3-?J9�o�'�ydh�\���qB� x��cw���׭`(�Jh��$�ֵ;�o��D�����J�H�����ߍ��6���<Z������5���F�"�g��3(6��G�'ݘ���B爙m����N�V1)0.h���>l�ay��e���	�P�t��n�  >��*������YYye̟Ijx�i�Q�Y�</�6�j��0r��|_�0!k��vj��g7o�(�8Q�h�N�7KΐU�T1y�@�&��G칙 ������=�%�Yo6�<)�ZGqŁ�c���MW����a�O��i��*���+FB�lyx"֚�S��H��>6�k��c��
L�.K��|s�cUm�
�АԎv;S�@ھ9m�ڐ�u@6�9�#��e�0��U��Q��3{��0��n�Fz9#߸�tR�)��&jUg�!����)�aU�HhI��Os=�^
�x���-�$��~aԑ�:o��wl��M��&��
#4��A='�܇g���0@�/?����ȼgR�W��z%#C�����5
3)�]��cGR�3Ih�_7���?4�C�3}ި�=	�p���m�]@h$�ZoJ�)����R%�2��9�C|�M�|E>�?{I�9�ښX��e��d�3S&��}�Ӣ����8F�Ǜ�Ab�i�<��۸Z��C6�d9�
i��SƾN4("gk�lElx��P�L�ZR!2ȴ���x)���;�l�J���mĞ��x����"�ފo��j{�_�ު�&�T�5S�'S��8����o��l�x�8��s��jT�	
���d�ְ}n��s�jpE{��9�&�u��C+���p���F��1��1�����t��r� ��%�
R��h�[��a?�4�@�r���=�%6��'{Aɚ���͡�����.����9n���>9\�፜�����A���Ja����S�x�WcI�$_��o���6e�i��MXew9�A!Jww�^���D	�-Y�ϻ�N��1	B�b�x0dm �U��ީ�H�N�17݂��H ��ACgi�f[���D�]�f�5��2�^v����X����v ��h������������5Y4����b��9���Pf+���]�tW>B/�LǤ�x �S120J��ڲ6D �&��%�7�������V'�M!�;��;7yp��@|P�|4mO��8V	���%i��6eC�:{�Hᘓ[��K��ު�B;�[,8�
7�ٝ=eޞ���%�hߵ�l�5L��Q�e�8��=)��G����#o�웤��Hr	Uv�So�-SL�E�y��=	���0|�ΈL��ݯ ��Y�Y��7�X6>-��o�Dpi����A���E�^�#~Q��/�#�L�9�C8��d���>�M�8Sx���)#��F�	"V��,~A?�Qlr�.m��r1�@ycT���iS���2�� [4Q�׋��Ƞβa�צL�� ���w��2_1Hҩz2j>�����i�(�)hn�Z8��J�2�2fj�����H�_lއ#�>�5��6O��6S��:���?ד�� 1X�	��m}��w��N<��������Z}�I�ބ�R63��Xo��M�� �0r0&����0^<���]P�IK�)��܎;ɍ��*�^�B�� 'H:��_�V~�|v�]FhQh�,v3�_ws�%��!�.O
��=�۱���{�3&����B��I�Zi.�j��w��Į�Njk��aO{�wi	��\�������X����~0�`�f'���ԕ�����T���9.+	�$+��w�U>�iU��ۿM�=��EMv�`^����0"�0p,S�����j;ak�$�:
f,|?�wb*��̣}Dz�j6վz�-~R+H���<Le���-�RQ�gLzs��Jv٠T���,���r��s_+Zi��
�Bt��]�:�~�]�im�a#���1t:�!aj�ި[G�y]��В�: ��1��C鋊�t'0��xa:�@��=o�[,:��a�5I��ƲV�O��yc�4B�i6_uƌ�Ț>UѶ!�x/��d!�>�{X$�R��p߷g4�^����� �f�`�R�DV�S��5�f��ޅ`�����G$4e�}o$�����C�0���]�A��$]�������]�Z�xh���n)�dڗ3>�o��H�| �8B�'�t�hrF�K7\Vs\b`�~�\�7yy�_ܰ�r2�A�����]_^4�J��R��};�ێ��O�	G$�����zD�VL���O���ڒ���E��kt����qnؓK������Z�~�_K�S=
������C!V�4e�I�8-�}�l���|���
Q	nn/bN{Vj��I�,��X ���x-9�����]�;�xk������t��	 L-r)�f��uZ~������q�CCW��^l�I�D�o	U���1!%�p���q]�e��Ѽ$�(1"�m���QY6jt��T�|��5�:���ǈ�і�.h�p�a�[��z���	� ��z�n�4\�%P�y�M�q��[t�ʘV�:c,���\Z�I���� ֆ+�jｼŞ��G�~���8��/r�Gd�!R'���x�^!���g����x�u/]�]�˖kp��s?U�)FA��n���d����ψ�m��L��x��HN��g�$?I�t_Ɠ��'Di���Z�V�bz'�P�R0i@77A.k3s��=`ħt(��(�S�<4w	��G궣G��h}��VD��ڃ�l	��p_6�ܪa�͸����sKӁs�3شj�L�����7�{cK�[b��;+gI��H��C���}P�;)�� M��ķ���2�]	{y���+���Q�27SS��{
�����`�=\̙.��mE!�q|ag7N䙥���X�,]x���ې��x��n�Fo~��C�g�Η��ݐ�/��y%"����P�Rj/	C��d𰍲.佐3A��0#�,�! �#u�f'�V��)�]"��]��m0�2��3����o �g0�wV�H�xcQ�,��"7�h������_����w�n����|�D'����r�u|�l0�,Dn
y��8���`�+h�E����qV�8d�;�"���%V����3���Ϸy'�8�4+d#�O_�FF�˙v�A(�V�7b��C�Y]Ζ?pZޯ� fl�#�����v�2������1ۄ# �8�X�ˆ/`�k�[���[�K�*�?�w\�>F]!i�$�~U� Eu��ٌi�;�#�Q+__n����7�їF��LV<d��Rȑ�E�6*(�H�/鴯��h�Y|g%�%��i�cf��X��� ̼Ћ<���v��s�	�D�Zt�y�	�"�̡����.ZfT��Į�7���1��O�k���_����6����=���&Ö
��;g$��?v���%J_�ن�&���f_�S�y`���+����l����7�H�N}�Y#��G0��$����Ჲ��֠1=��p�E�)���8$��W��5UD��f����W�(� L:v��z�8����Ow�#�i���ĕ�2�x1�x]��k(�e)T ڹ�ir2	��\+�������g� ̚Zy�]�v�Y �qG#�7�\1U1�2�Y#��W1����1fp���]�BuN�����k�Ye��v�;p���qu���} p&�g������(��p��hB��I
��q;H��׫�IS��7qe!�fJn#�$�����#���F(4[�=���P������4�д�f>��#��n�o&������Qv��@����3��Y�ߺ��zd$���)�rj��悶oxd�ß���8we�%J���]e�w8�'ԃP�O3R��ߐ8��d��8پ��o���\�R��ϪH /��70���#���� � V�˼�~C0�=wT{�Z)��`�� ���]r羵��9F�RG_����!�Jf0�0oB��O�����q����r��8�-�'ukuXyX<7�2��9�)EpVb�A2��T����V�tp����o�4����@6DtC��y�I������C:Cum�o����[�8p
��>���ٱ��9����~��ԣ�k7))�#Kww��yP�~꤬���/ק�ʯ#m�g	�0��ul����lR����@*�]����R4T��^�Q|��&\i�q(X[��J����pw����;�_�C�Fh�Q@ڎ�jB�s��h� ���)OƘ�e�v_�L�!���K�
�mw�dߊigNW�H�>x��L�<���|pd��/��:�n��9<M ���Ƀ� �����M����Q�w<
�����X:/���N��mle���fA)�ӯ�Tq� �C���ؚTЬk齪9Bh��mdjea����0Mg�����HY8Y]J��B�C�S|�Ct�ə���tXv��}��7.lH!�%o&��H L A�J�-D�8�s�	G �6}S�U�R�84eI���R�L�в�~��"�%�%o�'�j{�ːB��A��\C�v�-3�Z�L��X52tg`'��#�8�'6;`�نђ� c����P�VC�h�����p��X|�����6yx,���ŘM�8���5e�p"})D
� �Z�xޔ6�#D �;���&nttL+�D�r�,��Ǘ�/�}�e27���[�PV��"�Ã�	>��#�/Ͻdw&*WN���Q��kr.��.m�p^j���*p�|n�^��FF��{f���+�V��	�� ù�u��� �:��� ����bu �t��Bf�F��^f�B���U5!y\Rl��b�|�Ft(�q����.��O����E��P}��)b^���&��ah'b�h��7��q�j�rv�>�_����ے�"S�ks*Lk����b}�z�s#��r
�VLͲ��v���]�(���P'\ɼ��>Jh��½z���Os�jL(��B�ИD]=��� � �AB^�b���\V��
{�_P�T��L���e�d�̋�9��Q!��U���9&<_˰{_�;��I3T����*�kB�V�gU��#(T�o|����]ċ�8�_!��Z�A�T��`�`�yHk�6�YS���*|�yn�-�ر�	�T
���7�n��d���]���Qj������5@�Hv�+�အ��v�iS�h/��������:��P( �1
���dMǹ�p�8�];1�Uy�DM	���@��t�,���!�900i�I!�u].������y@*v}�Y�'�T��r�$���W8����=7�����0S튵��J��y5mq:���Y|h��q�����H�n��W�i��z��_C���o'	g�r8�8�֯��l-� �X�`ڳ�Oץ)$�~��b:����3Q��;J"S��C[��`Q^��@{9���hbzR��wJ|s��`�������51��B���YD6�Q�:TŎ��Ω�&4��V�#�kMLr�?�O�c�&�q�ɹ-\h�1^�;��Zv@�v��[t�`C<�Px?���z�Ù0������zy�(�3�V�x]��I'��N,�ߍ���P\�t�m�3zrj:I�<i�V���m�0�j"[J �y�o\"��'���4�癴�$��E=}ᙊ��N.��$�U�_'c�o�n�*�>@:ϲ��Kx�H4i����r�0L���FV Փ�|p�AM�6�g�VR���XXR�c*�l����_� ar�FQUa��D�Cô�*$�J�aӁ�x�6��ه^"���<!6�(�?~BӠ�5}6��+!A���~a,���mw��P;^�b�w��ڢ���Ay仩B�l v3�{y�܄�9�w�����������N�>��9�xs���#u�X�) C�Poa�J��>��,=��^�ͱ�\6�m�'�"�)�%�gQ@^���::�r�&�h-W�����?�6AU�Lf'�Î��Г")�HM>�,S�@���Pw�R��$'$���.	�����wq|�t/�@r�6�_�{�J�*����'��
�+�i�f�ou���rEk!���lY�WAE���ɡ[�fa�v�}�>���������֠nly���C˳yJu��>׃w�Y��zZ+D}�����P�:�)��3��G9���o�Xs��zvL�i,f��L>��$x-kZ�憧˕���_�e�b͘��W�;�z@�;�k����Y;]����g8��y�KsE���*B�X`w�=ҳ�,�!c��n�ݿ�h�J*�x�r��0x:z='�l��PiqQ����=��zJ �����cCA�eSG�;�ϛ>�j{�E�)b�
yD_xO@_�z7��|��;m����z���FB�p�$H70}_#6�b's�Ў �M�U`�j��iv4@�l�JF� �˷IR+5��[I��U���M�&��O,�t�$mX��zy]�Q6�K�U�h�|+).�֔Q��Fp�U��trR^O!�Y|h���<ZfW�c���f�OnD?<y���-�'�U�T*'E����,>l5����-9��8k������}��yL��ʋ��wp�^�cm�6�5~���B,�	0Ȥ�<�<���R��d�2��Le�r.��띸�V��|�>�LK�[Z"�{O���d>k��Fx�,<㮍�YU�GoFI��r�Q����9)s)�Zک����:%'�Q�9��73ooD�N�}��9�Iw&��`HҐl\Fel	n��&葓^ ��s�(<,��a� �o�j����T�ܚ�a���A�7-��!��ܺ��H��e0�^�A�MV\�$�ey7��ܾ�(_���Se�gT��%أ�4YG�{ހ��ɲ <�'K)m��c ()��l��mڝ��͕!ܙ�]�l�|���jU]���a3�[;��>��s[��`���Zr�#N¹V4%�{�r�.��05�k}����#���m��� ��o� �43}X"e<w���J�H�o�ײ~]��2���)o,cOy���n���vC1U��9 ��-�]�懟p��؈�j�PShw��:+���>�s������;�T�n9y��Ρ��t�;ȋ�b�U�u�֟��q)y���fP8�16��ò�wL��I��N^]�t	���SB����łh���xϔ҆�%�:3�j+�mn1�
SE�6�.>����~�{�u���ѡ{xp)���g�M;�ۜؑ�����X�_.J�"�պ �S�f�2���<��F�<�LFv�q5'(
���i0y,����p�Oҕ6��kI�I]�x#�5��55�c���d,?��Ќ.t�&��e��n4<�Q�Oڰ����]�,a �	���	e��z܎�������~_	�T�k[�	�Hjh$&��m�U�A@�Ֆ⎜� ��^V���J�id4G�[׏"_s���2'8>"�7}��]J�2(̿"�4��2��1_�W;Tځ�$�I�?%!� i��ؙ�b���e��݀Wnh""l肥4uv��=�8?^F��j�ʷ+ߐ�D<���ڀ�~�XL�$F	C�ת+H��\�k�z�N��}��e�<�<u/�|'�E���,u�ND�y�'�3s��؄�|n6y'p{�X%_�	z@����R� ���Fr�#.r�2
��ʔ�F�j,ՔQ
�����n�7P��5��e��W�D�e,��v��Ҷi�d�K�*A��׀���Q��z��]k[��h֕1�~�{y	�y��Y�����Cʦ�98�](vY����ε�@�8~�t!!�V�6�D���HP�.C�W�����+�^]wQ	������-'�b}�O,����߆�`��,�'�b��Ka͚�4\6��U��9���V�1�~9����,������x{i�`�N�i2>��[�%��W]SL=���9����}D��v��̳~�谌���ũ���R��_[C���R�L��N��� ���,׾�";�'�!���'|���Ɇ�AEW_�A��Ԥ��j�#_�b��	T>e`�j�������h��O���#����i@y4ŔfgO�
!����5�+�Qz���di5A����6����1\ᡵ�M�㞶h��
˨,��$��|��LJN�p��O\	�K�)A�c�U���N����_�Yu��6���u�Lw�_y3#����t��`����P|=!A�~�����*i֣����"x��}��h �7әd?B��dX:�w��H0�O��{Ι�,F���V���yxu�0�S�����a���H�\n!��x��S�?��8�DF��]J^�Zc�t��0��%�4����O�\I�|U���KO��=(�dv��'q�����º�.Բ���	r���B�x��Mp�'�у���נ����?~�df�O�2
�V(5����T��|MSwĀ҄��y�+6TG��
�x�&['rq$'ą�~�q(����8��!V�d���!L�"eA*?�0Lҿ�0��PTZoW�BMt��w�?&Ё��>)�"�Ҝ�٨}�\xe���11��!qU��n���sދN:R/I��y�c��r&���T��$H�kFN��-@�8�u
����N=7-�޾9�w�:��ޕ[���2���
���*%�m��輨!�7BZ�[8�����Cd�k�����+=�_�t#%�{\�y<߈�v�7yl�CY[�]�Ɨ�{2y<"�##�F��*@����%�
��1w�gu����lA�P[��	Ka�ݮ������/W�?�**�ݲE�o���Y��j���j�+:w��٬��g���UR��{�w�`e\�>Л"�+9�	yN1���g�'2j���?��T;%>�~$\���`��3Tq=*����k_��l�R¶�ˉL���M�{��&#&U�.	T*{d���tH.����H ���	�J��t*��4-��SO[�0lAH��G��[����+)͎! �� ��T",���>��DϡZ��t�<۫�M�^/޲Ef=L5��j~y�Jƴ�\�-u٥*����E���|�LM���?�r��,F\��@6ͬU�O�o8�o��
���͓��S\�lԬg䤮��F��������2_�����: )uC�0�m�p�B.@f��WEK�����,�dP*�p݅���~�����u*�\e�[?t�����׶_�����X��+�C����	�I����.�N��mw�����B]ɕ�.�����R'�<�1Q��w����܍J��gM ��@���'��!���Ko�i��q�ŀ�ޞ�2L�2�����hB��[�r&!0y���y�1����|-����*��弐���D�a9�~��$�`=���grr�"�"��Y��� ��z�C��Kj�#=Tw�*<��G��go��*v��:\�sJ�5�D��ʤ��������`��yBM��k�\��C�4��=����U�5�H�������p�'�Dy2вwc�C�J0|���/p@x���x$��'u���U��y�	&��\S���Iס���Nx�Uye ��?XTM��t!�E�ܒ�,e
�Sp�*ud���H��:|N�#���	�{��+���n�/ay�j�39���[������.T����>� ��m
>
(oө�?����#8Nw����T���5u�p���M�>_U�o�p�Q-��+�Mh{��Np_���/�� L|!Uk���6|�G���V(Jla�����B"�o���˳x���Rm�5\�6c��œ��%+/����q`4#��X0�{Y2��}k>�ե8�����TA��m.��Ǹ��У�;Ddy�S{��i%�+0N(!;���;C�fFG|(�H�_��@ߗ�h��Q^K��v�=^��]��߳G(!�w�Ŷ���,u!$����^�%�nj�전�&n]8C�:��_Z�H!�@�sՃ�=�=~4a��5�Y�G�&�4������7X!���N�u�Θ	�+Șm��0Q�'��<�B"��uP�5x\lB���b��ͩx��,_i�zRG�ro�	��}�Qf��R�9.�j�e�&�nX-z�������l���hC�ƒ����Fzdg Kh��/��9�g��Io���_�6v��%=ϗb�����Z��s�`㏯�c���v7Bh�%�MQI�D'j+[�*[�Ȁ�����k?��R�Q�Ջ���ˬKo�
�{��;��:���)��d�<H�Q)[`�c���7hU���ks*U{�J�_Gw)k��Ą|) �Uv�p���	���,��̃���������-���:QE�����EpX�}�^gqdV���<��T�K*�pI���(�]�, Sl�?us1�?O���c��v�õ������]?5��_c���W����xt�!����w�S���A�UL�Ba*��G����ߚX�Z�=���H��$G *�1"��Ku=����;N�$A�<�¿�d$�fz�R�-w����H�ĝ�cc?r�Z�z]���?��e7}����#w&=e�$� Yǭ��ef���j?Jh|���F	��$h��쎊B��\�ʋ��Ɂ���W���"�M�.~M�܆O�����T��g���bx�A3*�[��s(b���+���Z���];3]'�>�����w��BAsGF�5�U+����tm�f�k�g��2���)�l�`I`��-v��	E@c���ڞ�;(<g����k�!"�'�h�9�}��!aXt��� �bW�(b����"S�)�C��L�޿��f�AT�9����q��9�l��I�"<UC�5r�A{]������5���a8�V�9^"e�+`q�E�Pb� k���Z����mP�}��L�I�����t�[m��+�~M����Ʊ@�C:d��*��6�'P���A��GY�����+Ek�y��ae�FC��d?~�!�&c����l��O�ދ6'�M�� ���Do�+�T
���G��lS\��w��H��z���%�t|/0I�8�/���	�����eX�����I�̟y�y�^�Ao�����#��x���݀s�Z�UJi�b��Y���z������F���p�Y+�������hm�c�tf����RE�S��h���D6��?��q�w�t09�,7��7,'�j�� ��K	<8�%J��w���ׯ���]�JXv���uɫQ�ZjCN=ns��]=0��c�i�oyUQ�A4�LǾ�`��wW[���B:"Z��9Wfd�3) {�3&*��� *�����<��fI��h�N�r�M$������=�,]��#p��l��٘�=6�U�o2.�*gte�:�];`qT)V!~��o�>lx ������% s�C��Wf��̃]�Ԣ��	��F��րԳ�s�j��(c%�Y
�$��e�y���Y�� Jkg��v\�)ӯ��%$Ȋ���G*��h�h>�'��IIem��t���R;2�wxRd�.D�Ó�I�����}w
�'ҏ�ҩ$�{!������qdCl؛PTK��y��<�� *W�1l9��#��A8f�z���AP�V<"3�k�e��I�N()�(z���ég�g�3��	�Hyz��^�X],e���6�L��?C���,�b�>`�)GC���f"aAv�ߌ�p6����¦;���������+*�Y�1�i���׸�e��S�_u��s=�a��:���~���������s[-2��z�J�qL�n5}}-e4����f���qb�&oB��h]"j4%�;�s���W�/��kw��t�|e�u�y\NE}����m��!����<M�/!�I<���γXh�����BzH��;�v���ѼW$�ww��@��y�Ƀ�m��&up�g��n��юʇth7����;���y��O�OeU�ͦ����'Z4Y]�$�ώoMC�	�[��eP}��{{%�wT(�IG	/�%�Z�'�evH���^�E[��z=۸������C�}_�<$�/7��p����s�:���D����Q��`�MM�F�O����f�`�s��z{�Tay(n��S]�#g��R�C�5�gz�8���%������8Ѻ��ΐ�R�h.�-g,��������l�!����Q� �9������	p���%�d��4�:堅�̤��Y+�Zi�~/�SU�Nh�������@ܤ��*���)�ӡ� �}	u�݇m/'Aӧ���o�a��k{W�aŠ\paS�卜��VF��X;�?hK��������V̓���
չ'8�|c��<�lM��K�.\! �m�C^�H��	bi�G��6]�����c��N�uJXIP-�ʠ�QF;�w���1�%����+����]1�69�&��D�$�ã�9��f�1��!�Ն�P���cZ����]u�	�����H���P�y4Ss��2 �︲~��Z�co�F:a�:!Y%��>'���m�˰�!�G�:ǋǕ�-�ȶ�#K��4���5����{��xB�o�܃x�us��V����u�6�P-�s��Ǵ:=ГSe�1 �b��ͤ���0�����t�EGK���p�����6?���X�����UW�Qĉ]�hr�Q�iK�`Ow���/ڽ�mxv��� L�Z�)�&����>Pz�Ϛ��!G`��m�7O���P����������`�ԗ�P�Z��ʡ�;�����\�P,�����ӱ�z����t����R�׵P�֓�! �����|d#�{��6-�����%ξ���k�Mó�e���Ц�kc�Gok=J���X��Z;�q�gN��S5��q �l�~!��r������r��}؇dU.�~}��e $͇!U���$�W(� 7BU��JX�S��N��Y?���: ���NO��A�@�k�Ʀ��9�k	6xL!˽��m��eC�=�2�Y�<S�2�Qo�R<7�.�KH$�����y��R	9�ΰγ�ו�*�̎d��?� �yM�-P������*Rz��^^�4���"*!柁���T�	U��$m]���&fI|:������t�j��`'*{�zL������x��;Ҥ�Xqjݱ8P<LX�@�<��ǧ#56����u�p�TԽ�����;�}'�T:�_W�I�&;w�1���'��5 ����+����՟�1�Z�p��8���n����R1>5Wi��c#�B�Y��*�4~�ǽ��K��H�f��0h?j�$~WT����+�a<g��AldO���^L�����\��v�͛�g��L��OM� ��5�+��^8O���֢��������Gl_�tz�����_lz)�c�x����$���T��JY��<��m� ��4���2̹F�����"��2e*U�#1��Us|���TK"�t�4���y��.-�+:#�,��Q�k����z#q2�Fl�'�9��C(y\⒉�wC����4�ݨ�V��xC��-R{��Ά�<��x��=(�J����	4j��GȒ`(l� k�;Q!�D��{�D,�l�ٟ�6��6⧖����*���$+~���l��r����;���Li�znF�"ǝ?&�I�m��킗 X��������~�Ĵku���н�Rj�+���V��82��vxd���7��e���>���k�a�qvd�f���t��ʹ(,��Yhy�#i��G�$�nxke�����9H�����5�������2����B+�Y�[�f�A��$��8�mi�M��̬��S����h8��L�>��y,i�;i�b�P�w�SW	����H�oܻNXT�A���M$��9�
/�y"��_͛6�咪t�d<���i'ӂcw9�O�V,�(_M���I��0��w�+\�@�1�2�ؿ
QU��9B$���U�'��8+`/u�	�0�+��{�2�������D���*�&��Hq��&6+e��9���`xb�O=��8�D �ޫ�ճ]�ϕ�h�]�H��]�#Ńy�Iu[�� a��U��0��T�;\a�_�# ��=�ɓ����5��4{N�c��2���ӥ6X����8)'�F�w�6���^�ދ<��!T�|��o��^�/�^�L�4��v��+�RdH���v�,U~�>xl�}n����у�������4X9�B�{^`�e�z��ß�'�X7��YzO�n\{M���s��=����8W��vG<��U�B�!�c�'z�/���d�WZ�U%Z���ɼw�����c]haw_H��9�MI��(5Vmx�]�Zi����M��_M�vRX1��/����Bݪ)��env���o���_��W'�Q��f�&��GZc��c�|}ݧ
�xQ�$�{%8Uo�i���"�`ߏD/�f�*d__�
�����&��V�ZJə���k�=�����8���j�I�8֧��n٠H\R[pDD�`���-܋�z����Y��W4����(�����J]�῟8��d��z��>Ǭ��v�;QX�V�[8�����
wY��)������@��b���[��w�)N�y��i+p��p�J=��F��4`&p` ��Sh�Am�^��\JTX�P���)�Ȏ���R>��1���S?(��Y?"�,���M�m��:Ĝ#������FY�S3��F��!S��"+������|Ϣ��������>�`I��$�gƠ�(kg%�K�� �>Ia�:���~}��DQ�'m2�1��o�E��vS�$�A'7�6ø��s� �� S�LCgV�*��dy�)?@�%(�u6���`�\�����>2��˕�����\���~b�������ƕ9� �����k�3�>�Dp�
Q��׆e����؍�P�r�l�6t6X����\斆	c2�!>��SE��b�����=����Ů�#
�����L*��]5��sG&���B�=�9����q���)q/w��jϱ��1QЛ�}s3��	�m������N�#�P	
�$�Qڃ��٪�ۏVu`/]@޷h���u�~/n�5�ŠS�1:s�� 
07t�����j����m��Z��f�� ����#˺�
Pa��b�1(������_����`�%r�Y��n�=n���I��n�?E 
/����mS��j�%�y)21[��̠�*3���ѯ��J@����m�AT��Nu��x|��Η����!�L/"���u��Z�$I!W\�MQ͢�sM�c������`<��zr���&�yՋ��Yq�g���y��A̛�Ǖ/�.7�Qv[eͯ�FI?�����j�n�������v�U,E�V��Ĥ:�7l>�̂j}�f�*p��*���0iX)z[��A���eɛ]���m����a��;V����k�mf=5�����h��DFƹ �P�	����D�(H^^prS�Iǲ��;��ʸF���<P�c���`���n8S*��u�Y|��)YE�V�f:Of���.���{tA�]��x�%��K���]�LC���	?IWH-]�����Ci�#R�H9 hs���[U�t�[?˘)G�.m�J%��u����w�ͣ�qh���p���t!�&�	\M��Ff�ֿ������P�U���{b�����?���g�r�8�G�$���'j�ƪO$cV`T��tj� m��~�ɝU��]�^Ժ�Y��80Ǹ�e���,��^�n��K�����b���n"�;M�uD�~�P��-�=�n���х�q���4��Ng~��2�=��Iw@wo_�?mdӴ��2Ջc���O~������nճ)J$Ǎ����;HI�W�J�/�Q��?=',��l� ��ד0R�{����¨4���.~��>��` t3h�օ�/?{������z��ܫhl���������~�YM�q"J�E<�)T��;;��T�qւ��ߋ�qUU)�v�Z|��z>A��OԮ@�)K|C���zQnz6����^�9�x+��	5��+�yy�6H�a�UdEf��l�
�c��l�w^h!�.�9�&Ε<O�-t�WY8�)�\��Κ�K����R-t+��*�v����'IS�����l�m���	��:�őuo����e�'�h�͗�����5w��3���<K��Zef'�7;�&K�i����3�v���Ns�(I��G�I@�(��q���������j��X���H�=M֑��GM��+'�O�/�!?��@�p�,Ey|�L�K�[��N�SkФ�����S��ef�B$C��M$IB��@+̗��Űak�Ў���'�Q�z�0�t#ٔ�(#���y��Ϸ��IN��\��jE�R@�5��_���-�����u�3���&�/�g�YE�k�&ŋ��@�Q"�m_���5�?���\�H�]���<�(^�P�����L@ �5k��=	B�Y��|#�dz�o�J����4$�<�>�#+&�g>T���.ڻ��"����pS���Q�ft:�������J׏
��s��xhx���gc�>pM#��s'�SA�.P�Ỹdup�LgT<����VQ|��j�#�_�!�Ic�HF?1��d>�H~\��>�.׭�>J�:���Wi,��G��c#��
���dY8��q��ؙۮ�����YG�Np׸�����8����(#�4?i��o�g��&����&�Й���ш�/\�������x�C�J�5��b.[��'�ݘ�:�M�ت5Gd&��-ݢ=�!A��:�����(u�w	�37�BT�d���drG�_����{��4�R�(ձ�0�z\{���͒���qK�;(v함��	�F|�����9����'�6s[��G���*$O���_�Q� ڏ�L�Ѡ�V�h~ q��9��~�k^%du�Bai5<����L�u2��o@sa���O�kI���֔���`��
¾��4x��Ik`���� �^����O�C��sm]����{Yܞ�Oav7�LJ�+�� ���y衐�ڀ�Q̟z�+ђz]{�#8�̺d���s[�\��J��Y���$@�r���.��ib ��f�	������0t1����$��9�x�YMj��N;��u|��D�|g��n"o�9>�R�����B6�B{3�AH���♏>���[q'�E(��mxg���i��GپO�ˑi��d�2q6��]s��S�f�h��x ��<v�փj��kK3�5�i9��!�3s?Hp#��+L��j�F��5c.ć���H-ﺿ���`��
��H)�VXu+���������*z%��
p��X�%R��gHT��e��s&�0�\�B�L��z:�F����CR��#�v?�G��Nk�����y�&Ā���S��jw�f�c
=�����g�:mpz~�YZa�����b�پ��i����_u���:�C�/ʟ3W��]B�a	��=o�ߵ2Y.�
��O�P��jE�djq�5;���Ak 49���˖{F�H�(��Rt-j�v�s�T�7���U�)���5�`�h�%����N�Ӆ��-r<Á�X�+Wid�%P��r��HI�8ά�.�;#���(���l���f��6"s��M)q.?�T�Տd�>������P���(�O�Y9W��>����f��B�l�n�f�g�B!����W���?Rs�}������2�b���^�m� ,]impӤϭh��m%�Q��#�xx�K�aW r�Fy�@�Ś3PzK�A���\������Zg��mȲ��;��R����I
����8lAY�l���\Ri`\F}�S����������9O,N��d��8Ͷ�ιő�����n���s�Ċ/�P����6`��D���/�V�p��{�?�l�gy1yK��V�W��y�b@����Q$H��Ç�
��=/�7�Q�KmA���e��G�n �y�
Q���dF��֫n�����ٿ�h ���q)��|y~POڄ���E�c9��,̣0L*P�mc����^T�:���=ݷ��{��Sz�����.&��Ɠ�9�E=�~μ�W��53�~�kS�Ȣ3XQg��Лh�����N����|@��:� $�!QA�\xQ띥�8
�ny��<������W�Ii9���U�i�Q cGC���M~@�aӮ�)���f;��	W��+�	eFլ�:�
�����v�:��2̈���2�U&Z���G@6n��<�
+D�qB�`�>�8��6r���2�	��D�5x�]dFĨ�3=�G��� ����"/��o.2xK�Zߧou��I v���4�Ӫ�U�������t��{����5hLݥRW�:P��>5곕�0쒟��`�)s�v�H���/()�/�]��X�r�����]�-���h���pkdz6�*|�^_���Wg��=/��v�����me�}z4�\��&�P48W���h&�wN�Aw�7�>t��x��h�*ޣ<D6o��Lp,#���I�	��_�����1��w�^B
�A�m�3�=��aJ:<��m.��{��$��M%���u�BbE�����8G��+�%�����
";���v{{5`J$2���_$t�W�o�zWn��f��G�!?A��S���� ⤐�b�Z�:;?h�ě�f�NB/�ÃPh��x�k)-�[��Ġ�3����p2J���Ը]9󭭭3�'е9X��q_cc��!4\���d��(�	�F%b��J�,t����˒&H�(��,���:�a��Ƞ���L�f@N(���V�R��Dq+��N���Ī}��e~�=k }�P�mi����@��2���	�7b��h	�5C��n��?9�
���y�䲞7�Z�����=e߀��AEAx���)Ψ.ι;�k�Q�{+���{�ο�Q��q��=wԚGX���IvޒV��7:��/;U�b�ٜ��H)^�݀�^�iq�'%���5����� ��jk��U	�3=HU���O�>4�UR��XͿ���ßM6��V�/ʑ�vI ���b��r��z/j>D�h�6���USA��v�*o�N��x��53�"�\�൲i��J�X3X�iss˞BQ>�@����ѹ׸�V��p�k%U�W0#F��
Ѯ���M��솰����,��5���O�v
>��a||Q)��6�'��s
cVC�D4�! ����+�7��GF�{�PxF��k��לbGxV�Blf�1�l}J�zX �K�y�G�7!�W%�8������J��_���ȸ^��#�aQ���#;�qA|��ju��]��O.r����޼�8u�/7r�"y�a��¿W�j��s���TƟ���(�s>{�%sk���1�_|���9�k�>�M%6"�RD��DV�i���ʸƫ>���ϋ��BB�?���3�&������(�ǎ�)A�T��w����,�>=���)3�敖:�ة��̠n�"��q��&���a���^����jhNK�Mb�ML�b[7�\I�LE�K�����q��s� J3��rl!�xxp�-�|>����[�,��w*׈С��hv.��� f."^�4�O�y�E��ࠟ������~,8H)u䈱E��h��9���0��1^�?J�ԭ�{N�%[:D�E�!I ��J�k�0eĳ�������l�[[FG�c��OiZ�S1�-3)������@ɯ��_�t-�T���#p `�(8�,�$��Z��b�|w�^���
���Di�����Ȃ׭$>��d�"mI3�l�&s�v˳�6Lw��F�ܿw��ů�w��M�l>-=C��f/3d��bLq�˲s�����	kA�IaW��/#o�_�#f�]4��LN���,)�;z�~�vX�2?틝�2"�1@��*У���?�e���ȑw�M/����T8����?9��sX��<�'���a:�$|�dU����jc��8:Yj�^$>���a�W^���_��7�ʑ��3��v�2w�[.n�g�Û����kϒ�=?�Z��S��>�G��B�B1d�l�SB?}�H�D�Q�auT��C>73�XM��Ŋ#�
"��&�lh���+�a��f9�8����Lِ�G��S��*�b����L=]~��K!
w��)6�P��F�"�'Kvw��µV
(G��X�{���I6��*K����M{�z��:�LB����0�{I�?E�ݐ�HL�Y��ͥG���m��Eu$��� >�P�Q/)�<;GG�J�pSS|�.�Έ��yٱ��=��p\O�M�&u�;6�}K|Rf�c_��<��~�=|k��.�{NVkϷ�+Z���&��&�,�)��I��@;$�U�0@z�{��ÎI�\b��BB۳�'I��q��J$+�^�U�{Ű�ac	�Xd?x��Qpa���g�^����Z5�}��΅(�0b�4����%m�ß]�=�ǆ���DA'�h��=m�ZGQ� �u�h.��pSc��q_��fn�m�{����k�Z��D+�LNC�{�=��>C����bn��� b,ً��`��
0;��~��H���.鶓�+
�=Lf���V���57]�Y@��a�ÍU�v��Qt�Ry�����"��8���쯰�f	{�Ϋ��vm�Ia����Lq���k�T��"̋ZF����?��#�����7��$�WFCT���49;�{'�kQ��:���UXN80���Ֆᱦ�Y��s���lw����4 ��^��85�/������$Fk�J���>�b5�<kDʅG����V @'{�7��~*O�� ��z�=�p�DR5�3�W�������|��S���S0��)�M�U�Jc���tx��-ӿj��{`�jϴm�9����@]�d)�}��x��Z��7�f�En_2�K��.� ����J�xy|~A4;�)�[��"Z�Ox6��2�c5��C3�ԗɈ!��y�q��Һ��r�����2��*?2��F�/����P;x��t=� �W����$}��D��5wϖvjF���b�A�WHq��M���B_�[Yw������;z5os��B̑'s����0�W}��:��9���8�b&�P��;�lx�r�K�Dn�u���������L��￺*9�j�.WC2X�`3�b�̹dS�rh V d��Y�/��U��^�ݞߊ��+��4�;��	&k[/�q�������Vt�b�cp2�]�V��4X�L��E�i7����֠)`����x�p��K"<�CE�ACkw����A���;�3ٯL�\��)�f�=�+�~/3)�V�U�*�U`�3����Hb�'��ܫc�ʕ4��QR�	�t ���1����+}#z�)N�[��Ll0�y��$�<]_�9�����v�;�,�9�p��jgv��߯�3<�+y�d���ծ��m5c�څ�;��_`�ވI��ҍ��#�H�rc���'�Q�z��=J����� �9��
���d��Li*f��,��7l���	�b�e��G�)7���/��ZKC]���B���n��(�a��4�Z�أ��I�8觧��w0�)s�^��m�_֔�>���I=��k�,aA�Q_��K��*aB�]5w���$��H���tI��L��;q����>-W����N�+��X��1.Pbש���˗@Ӛ��Y"�%&=��؉Rh��݇U+%E۔��Hn�G�����̐�s���:q�ķa���i*��5_�T��)�/ŭCjf��u9���#5w����\Dн!�H�|�ΒZq~�)����kR�g �e7T��<u�׉yBq`m� J"R�q)퐠�bY����KM[S��q쿛�X�[<k!�iα�],���b���9���J](�#���Ĺ�J���$;��������1U�)�ql_�Q��& e�+g~��G�V[��1'������t��T�ǊI1ٙH��bQ,�!'3��e	Dhף7ݼ��Y�Gm�X�����C���u	�� �a
������+mIn�}v��2v�w���,z����	
Dd�#����$�'k�%��{|(�϶��D�0.l��կi�5�.y��P�uOcuG��D�8/8dkf+ȳ�KС�_�O��U��}�(.�|r�㦻T�`]V���ա͆"�[P��`(�|dь!�]h�e����	6��ч�3=�G��뽭y�(�▓W`T>�k�������#L�	��|��/��-��]�ǵ�>����(��g��6.wk	��c(�4pfn�9������8p��qnfy-3��B��j�	Yz�Lۮ��p��f������(��)[�Ʒ��(�@�~�?���H��+ �Ѳ:�_-"	�9�}����$i���=Y,Zpb�%
Y�N`��K�S��5��^0v2_@ط�V�Z�����K�Q+��^�XJ������-�)���kGWa
Hxw]f�"�~�9��g�S�	���`��-F*����ê���:_}�������0a"�����%����i�׾�{KC�qRbۺa�u�I#d�^����;��@M����ؤTÉy,��H�h�)^	/1�7���Գz}2C��ol���S �P�|q9O�´Fq ^SZ<L>/Pа3	UCϞ)��j���^�g:�9Z9�G��qA��E۠�p�خ*�ּ��,B��$,[��m�%J8�`��>eP��l{7�K����o�ёd��v©>	y
n!�"t�����Rx,T/!`���������k��mam��X��Օ�J�V���?&���1�hk���ׁ�M�����>�'��T���KU����<�c���zJ����?�
 ��{�ĥ�2�Rfb�]`L]����m
3�M
�t��D���~j���魺�$�l����n=ʇZ� ��������hC�>��98spy�9 f��Os���(�󉍠��|ˢ��_��޲͕E���d���ಎ֦O�l`�?�5�]�)	����wQ7�G.;.ٮ"R^q���%��ME�>R��Ѻx�:G/%@�;��Q2��<r���l�s���Q�}�C=h����AIs�����g �E%��z�����[��?a����ot�!�߈���{�ŉtY��m-84���-�m2�)]�l/A$Z*b�ِH�!�ZVN��ԧ|NEY��R�$����Oz598u^y%-|uWe�4��*
eIL@����J+}4��T��E����"gВ�� cn/�ޥ�U�e���� ��9+q��Pǧl��z���,�U��x��'����S=/�ٗ��χO=N��R/����*�^-�#�:&&r�|����뗘�<;�Jp.\+�D�7��V���΀��YX��o0����������#ш.��ޖgS7`�|�U\kYJs{kR1sj2��yk%��l�"΀j*iN���-��3����h���c~��D���V�<p<kϥ�rT�QȦ�~#/Ty�w��}�`��X��0i{����p���)���`.�z����tv���8fj�[њ�A!pn5��K���/���5��|w/��H�����ѷ�k�C?��ð�!�@�w��͕���8P��l�!ήnaaǁ*�k��D�q_~���Gf.��?�H~#!��AR�������^�Xk��&����s��hi�	P��K2�8��(�C�M�K� >G!51a��吴��R;�"��
�|�w�C��K�Θ,?B�����&?��,�m�L<�7�O�	��[�(���_��3B���`�`�? ���K�}�%/kH2]�=�^�0�����t�q �1)��N|$�ӆ�ʠ}��*��9���|ܜ�si���n<�ot<G_�<F'�	s>��𯏠L�Y^���5:F��P?�l�u�$Į������ӯ�H8�a>�]g�\��\Ї�Z} voT�*�To������u?Q�1B�^�lW�x�3����]��pU$/�i7��R^\�7o���;�5�D~�~�:������j��!��b��~��p���@w����:�T����,��8��MO�=�f�P��{�t��=��|+1� �WfVPཿ#/랥�m���CC�W]�ģ����b�L��b�b�,w��4Ҫ3��gUK�y���攏�aq�x�Εt����Q��?h���Eݣ
Q_p=6�.
�4'
�Kk��m|�V��`rB�J��&xd1�G��k"|��m�6M�X\CS�M����n�9*�o���h������	��b�i�b�`*��������<Ђ�X	�lxL����Ј��2"ğh�`�l
�����E�,�h������5�nbPk]s �
��!�ʈ-W-���q���?$�=�Q\ڈ�H�Z��By��c(��=����L	H���<��0l��`��L/?�L��ymqgx9�/��m9nۦ�L���kr��uTwH��Gכ�8KX��Y�P�3��j�����Y�`�����m��$/C�X��gK^.L�V�ݢDb5 d=�~����y
��/���%����F��- �B�V��x+�Y�s�EC�!�#����1՟|A�H�5r�>S� �y4X�m�S�IUOl&������K:���8{H?ۉ�<	�Z_֙�>��PWs
1֮w�aB&I��9�\Ծ<i����d�ͤ�xI�I�����()��eР8�4 i]��}�=eYï���b���z5(�"-���>F�}�y�����aK��tI7w�vAM�G�Bc�@��RUjJVRo$��=K�n���P��=!XӜ��UN��N��|��j�����g9��y`�_QT�d��-J�2��@�����[_��iW����۩��R�*�Is�TPUXh�Éq0�ɝ�}=i���@Z'2�@ޑUҤlQݷj|��
O� �!�,&�j��Gy#�/�Ju6��8�<P�Rc��kQ+/���i���b&�z�]Bcj����cY��	�X����初 =as6vۗ��ܯH��^2��R7��`���@�4��da���t3Cfg@SF�R�g���"?ԑxiR�/������Fe�L�&G��mݾ���H�c�	��"��*�>?�宝�1y4�6�;�ݙ����h��g1*G]��PH�4�J�*�y`r���sE��(�N�e�(�0P��-�����-ɖ��s͋���������k&t�"�@���1D# �\ޝ�� ��P������(�s�,�l.��\e�K�����?r:��U�fp2T����t��!�%F��|.��k�qSsjBx(��q��*~��m�q�P4x��hX�_q�/];K�b2�Kf���hޯU�:���O&1�A��?�>xɥ�c�FNK�⥛��0Qsh�24>����3��K����M�A���wj����;8�M�nTT����TZ+M�4!������5��
0O��ue�|d�i�D��S�����+}����7uSA���e���n�.�W&��6Yڶ_Ȃ�C���"$��S���/J��$r����-i�rXX7t�;{����:Rf*��������������촡�����g���{j٭Z3�C5j��f�׼���e�IW}�d�����&
 *�`k68C�����1#f�K�G���WO�D�yhd"��>G�쯉��0r�������wh=Z��y������u+�P�*/��Ӗ�s�<������gS����Q�$>��~[�ؘHlXm5x7����)5�z�]X)���H�.���y2����3�|��W�ٲ5p�^�􀤅[ @f�t%���#R{R�Xձ���^��Q�Ob�R8��}蝢�#�%A-Wۓ`k^,���5Lk�����44Rt�*����'_��O(��7ea�O�t�IFq�jP��lV�	4����ң��{�6{Q���!C,p��ذ��:�Zx�è��=̭�{�4WA�U���߉�9�!���\	 ��K�'Y��k~'n�{rpV���K�{����v�ae��6�go�����w<IPHNWle\e�9�<�֞�/�̨2s����ྒྷޗ�]^E������NI}� ���������o&�T�/7OݬQ�R�ݗ@L�O��+�9����g��-X�k#�9��C�ŵ+-�	�:�Dcu�<Bu�ڙ/k ��;�tMfl�%NA������L���C25�Awk<���P�T_��㋛�ۮ��V<�+;XA��n)W�j�O�ܰ��S�� O0�;	L8rh�/&/E��c��}�S��=�|�,�kΠ��;���Z���˦p�F�O�Xp�L�s5���*�%䢪�4ƌ�ZJ$�#Ι���<~cC��'�E��Q!6���K��q+�k�Q�7���\���-k8Yn�ʫ���my���_�<�I����C��,Dr`8�ڈa�\Ww��Z� th�0	�n%3
�5�'[ж��B����4X�	z)����j��d9���R�Y�^#ڗ�K�+�Гp�[�&�P���KE4��G,0�p!� �������r7~���Yi�-�d�+B�=3��6vq�������	Vo�.��"돘��sbe����CRLu��⡪�MG�h�}�Rs����d�m�2l��]�Ğ�v*��\��a�1٥_�2
`!��|�vɜ@��Ϋ��3�H��s2y��p�29moR7寫��T�e7�`	��wA{�[��|'�6�Ԯ��ڃ{���p=����˹~�.v�J�]Jݢ5��:��63��%��bǦ��`D�浿Ű}n,t�J����W:���{���׏��۶ʼ�E�x�BCW�RUG��"�_�e�����[�k焽{[Pf��hŌO����-�͎��R"�S�]NXQV�����M}����r���"k�(#us9��j7�~��j���%�$�/�\��	����ɶ6��b����8��4fsDS����_�	�[�/���l�W�-�-C`[X�g���t�mĴ^6��uih�������������É���2��P��l�d|��@P����>C��eٱ^��Su�g��ss��C�Ѥq�&�p8|���TW�a?�����&�� �w$��ٟ�h/�����@Lت��!�PtQx�Eo�B�����[���� %M�v��Ϥ��4�#���N������ΐ@$�t�aq�1�&�ׇd�>�-��ހ3?�o�G�2�����3��c֮�0��s��	㦴ꧡ��Y ���h��
�)靈oU����P^"qAߗ$�(�<x�N�l��%xwp ��:��g ��A�u���QELӮC}xmnL�Wv-��"����R��A�������Ȏ�5�<D�����\12���c'�<-L7���:"��� ��_��RP��;л����E@A����)�*��U�I�o�3�"��1�A������oCױ,CT?���j ���������Um<�̀�f�.j��JV�=ua�Í=��R%\�aQت��la3𣻖�_(�k����cfB��gpYzmE���6���I]�G�y�^,�1U�nOVZe5�v�0K2!�<.\H����J��J��-�IG<��'Q����bC�,�:���D.5����ըŰ�����X7�$<qb���w���Z�X��2�U�����'���i��r� ���F0���S��3��96�s4�X+��L{$C�}�5*U��1LW�����j���.�/��x��j�+]&u�m­��8��:t|���ΒUK�?`��U�;�����1���$+���*��#�����ZT}��3�����1	\?��W$70�e�+.<vU/S_��5�.)�s�Y���7���|��}=)�D�VҶ��HO�zv�}sD���Ogsn�є7���}�]�
t�j�䘋�&���S�Y��f#J������4�8$�O��`�l�* �2,\�l.�/�����	r����1�y���o"�n��D;2���-��w]��'Hq�'����&����tY���UQ�OS���i�9�u�{��{% pY�V�H���jBM�;��Y�RnSr���[��|�s�a�K��B_���&o a^��y�Y��'�F]O���T<�2�4��ah�OLJ�~Ώ >�y0�{�h�FhA�)�^B���U
��ό�X���S�?�����b#[�:/����7U���S�PM�0��dL�x��Dkb1ot��t�f�������D�u�����[�#�$]Ɵ����/P���N�);lX�����w���]͛��$AA�+��W�ԧ��W��55����.Q�#��b3�(Z��q�W�Rl%,����	���.r1U�8m����yp�X��gPU���D!(1��H6z�[%%�]	����|A:Q�ؔæ�t�A�c��W�"�9�\��Ȕο�P,���5j�m�}P��&*s@�6���]��~���U�VS� �TS�����ӦJBe���M���%�e{�r�#�W [�lU�ۊ#�)H��C�1�mÄW`#���G� �?�p��4'����#��_�v�x��-3c�59���pQ/q���~XIǵ���x;լ�����Lή�TS�$�P�R+�o�D�E]����DL�:�^��R��dB7��='7)X0 +�Kf S ,���E�����}�#Pdez5�0'fsy�w|�B�쫦l�OE^'c:���H-{��׭���.����h��J쁲�R�n�"�'m��ez>Ca�F��t1���-���zw��7��-��������N�1O��L�]�>8�i>MR�qƃ-7�϶)z�.��t_@u�Me��)��f���3��'q��Co2��[u���O�B���k �+b�/�3�����a���6�W��XŒ�����>/x��ȁ1�O'q���|�b��I,���}49�:f�y�q�}�d�@D�\�˫�=��oqD���<5>�sx���="�l��*|gr�������Qj*<����W7���Ixau���Ah���H���@l���J�Қ�Ɓ��@�!��@[�+���/ ��RQ� $E�CِK<~�)��%T"�D$[f�%�ړB�OC��;)%Ě�����y����ĬO V�ϣ��alp�����'�vL�u&S¯nL�@ON{5�z$���ñ��,Y�lS��;k�D�F� 
!v�A����p�?>�含q�H�u��ÿ��l�ٚ}��ԅƹ�juP5�M9��͜�B�#� l�?\�#!�qX�b�\n@�eZ��uZ̿�v�!��@��Hr!��a����C�Aߌ(Ϩ��o�8����n�*�ѐ4���|����v�@Ds�|_�X ��Ȇ��}&J�|�D��BF�iz�R�,UΎR��T�^��0M{8Ug v4=Ѵ	����A���7���SX�{�P�$�=���⋹M�s��������v5��"�~��5�@�������/� Ƴ�0/f��I�E�ʳ��Ty	��C�aO"�t`��r��L����.o��P���b�⻐�1�7�dH�X�4�[Y�y:��2�FD�
�W���<���V�R�+��4`ȵ3�oY�}�GK?@��8��
�O�����U&Q���� 9�7����o�w�H��CEIP�$B�$���+Z�tli#p �<�S����˄c0�U��7�Q=9�>����TI��RD:��.��,�9(pL ��&����m�ڱ����[�����|�4��ѻ�8/��Rx������x t<7K�!ߎNN���M���>tJo���m�}J��w���u�y[7�,wӣ�+�ѫ�^/����A�߼��J)�x�}T{��|����S�+�p��'_�S�"!��;���,f���&W�Φ7�j<�eֶ�ള�&�_�|�ȶ{l�Ҥ`wm8����qsw��E86��4ݝ�p~*�M��/� �.�3@�	K��]��=�w�9~�s�8��h�b�;����_i�kõ�<n��$Z��u+�c٤��X&P�2nd����	�H(�d��-~���`H�$9~�����.h+%EɊ������n������\��B� @ӣ��|�	m3��x���2#
�"H�un0�ɻ��2��4L9rlE�~j/�����#��EzB���]Y�Q�B

�=�Pw��.���.X���\�h<q�	O�m�� ��A��p!�m�'�E��g��GP�G�c��̀5�w�����i?#J���Q��~��E�
�.�yCE�B�H���v� �A�"H�k'�� ������0�EϲrK�Ifpg�FҪ�=e.WެޮD���_� y�DXk
�:�1�M\O;�m�ۻ
�>�(-�*mF�:�Ȓő�!�lH�W�%��Q��s��.��4��2dѵX�{G��z�+�.g����t�S)G1A6\ӤC��q�:k-a!��HFxz�eX��FD�֫����%<��8bZ7�S䜷�3&�3w�
�����
�)w�F�N��V�*d5���8��q�R� ��	���q��-�_�_��+e��!e��۶Ͼ&X��(�z��GR2�
��EG��f�D?�l謉�'V�_�`/*���F�Q�M�/JvX%�@�ڒ<]������3\3���;%���(q*��8���N����X}ű�����9]�*���UC*�#�P���>�dZ"Ů5%C:\��!��s!y�2�\Us:�2��=�@���ȧ��X*���.쎾�o�A@<�{&��Z1+ c#��Z��M�kNށ�]ؿrN�D��b��Tk��]:��D/L�66KHT��e���!�������$�*N��(���̚�����NW�'�@���J�D1�O�BUoEw��TJO[�e��<i��v��6�� ��I��ȋ��%r�w�J"(����v�<#<"zYOʋ�'_�}4���a����ˮ`�Һ|��VM���5��G|�wK ޣJ?���ؙķZk9O�K�{q;�P�'2�.e �Up��On����e�z�Nߑ���j= �Ma*�Vc=|����X�n�C�̱>/J�(�)wK֠�P`��;�tF�Xo�!�i,b$y֣b�w��y�ͫW=֐�)��s��<����1�s�"�39L[�Ƴq���KJ�+�>�??$m\FI��k��Sxk����6��*�b�*�;�WY��6O��DĈ#q$&��m�_��y�RP��UΡ��&������=��]gvxʭ�z��X�d^E-�#
J����n��G=e�iaj�����6ô�	�K��SUM f���f�/�j�*-I�н��!`��S��R~��Z�ox��DXg�4-�e4�4�*zD��5�)Xq��9���w�d71����D��y����c��w�H�DL�.~7v���J
&��Pml��0:v�@���)�^�k���Ǉ'=o[���L�����Sp4�@n����T:�{ʿT8H�ਬ��k�t0�t_���<�Ǩ�N�2��붿�w�������?�;�;N?7FD3y�nTx�R�8�5��Xf4J? ���yV����G�� $0۔�u�����4�=�l�2Aaz#Z��Z��c7XX*P�� ߈�7:��o�6��˦���;��|a�Ⲷ�>�e�h�?���1u~r=�Vl�E���'y�}�GSE/��`!��QYmNА�:C��?��EtO9Z�'L$�立�/�ǝǷ�I�_�-�QR��^��$���'h�p%��Pk[~�$�CjR�F�Ӆ�A��.+���!��[�)�s���&d��tT��ZzW�ط�9L��qq�8�_4poe)�n���͝�z��d=>���p�k��s8#��8���N��lc:��{��sU�&�7��l<����2�����~J�>�z�W�ڋ
N���t�k�)���H�G�sS�+6	;r��FEsO㢐�d������QC%���՝j�ԥb�����8��挌-//�n�E+`G��Vy�FQ�VJ�����k�g�;�-g��o�9U����3���Qx�^�ܒc����V�۝�s�Y��P�fn��'�Q9z��j��ŕ��!�m�4�9u��_�:��ѧ����@��@v����8����d�o�;P ~\.�,Ad����Hg��O/��;V�^I�\~�2'4"��'J\,i���&��m�^���9��Z�L%i�F�Q�6G#Y�}�����+Ȋ���o������6�������Մ�����G�"b�����sB����%����dK���ڄG�*�Re�` �i�j��{S�4�p�\��Ȃ�(�$V]���a��Ih�'��3�-�B���T�4^pF����?���K\*'*��7��6LBq��L�Vk��E�7'��mCE
�>�m��<�*����Z @n��UPt��L�L ���'��;�C� �W�[���'�k\8b�a�k�E��i�ô��d5�،)��:����F�Q�o�x�����`F;��.O�0���1,������Xq��ƍ3l����%ߗBL�x�-�䘞��b���Z����	�7+R�PW&w�������F�lK��Rv�dl&s5c�]��<��O��7�(����D�d���x�YM
v��=6?������0Vv����i獼n�J����6���Vo?�"��2�a����:G�jj���u�� 5B{�����b����a��h�t��aإ>�q5ڰ��|�6�b��s�[�]��K��<���/��
����c�\�S�|��&��6�>%^�O��4����hE�-H��#U�f�ˇ<������JD�Zp�bW�%�QQ ����xW�K}T�Μ�-I�Q)�?6v%�`�^6����]�J���.2&�џ�b��J�z�ˌ���k���)��!�OZ~��^DF_��3p����"�O�� ����ze.�U�_v�Ά#aX��?�6P2�m�ɃT��e���������銧..����H�_� ڀ[t䡡/��|ކ~�D��LC3%�(��V�qα�o�?�.$�L�{V�ަ*x!���fGq���}�e�T9M�˦��Y����ZTP����zF��䐝������5AU�ֳ��� ؓ{�ky���QT���ߋ��$E�}^��^�.�h���ܸ����Z���s�wPZ&�oL���C���
u~���#�G{wy��K�n�sqpy.a����]o��W$��H�%�[~��+Zgqʝ���r�.\L^��}�j�0�~Q�cܓ�t$��(UƏ�w��+mu�p}�ޤ]?�AVW~!}3 ���;��������6�].��Csb���g~�(е`�{f2��Di��WW���п+-P�w!8� �x�cY�ќ- 2�~�����A�	�D�o��Θ)�A<���s�W���oeM'��O_�9�P��)P�5'�4vS���p	K'"�m�Ê�߈�Xߍ�sR�E�=��ppgr`�K�2STr��\��9=aъ��%ږ� _�}�S��W��b��C'8��˳�s.Ng�>�:oޛP;7�:�!������g�Q���󯸜c��^#Qg���xzBr�@��4�pDw k���=��%��y�<@������P�s���З�9#�D��x��9��5�v��tk^�'�<O�1�J^FctL�	p�d��N�O��zl�?~�&"����T��u<��Y��=����'�ǯ,�r2��dJDBGsk�� ��$�^�γ��ƃ�����B����) ���=#)CB��#�����\����0ܝo�0 Y��sx'p(lu]���U�77���n�ڦ\���ϩ� �g�����#��o�A��K�@����%LH�B�y�@dzl����98w�t�x��(��0m�O���ʘаNI1�Ip�ֱ~Uˢ�8�x�651�|�����v�c�U��ϴ?�lT��)�����o_�p&hT�mD��	�0@6��G`��:N�>nތv���0�g���@�&��:B�q��ܹm����<��I/�¦gt�^���T�&�Đ]������
����efM�fKw�A)!HHδ�C}�[��JD/P��YR��:����9�[���<��C�5Nb76�
)��Zٲk�,wC��KaΊ�Fi���(
�{s�P�
��'�(O��ē�ݘ H"ZI�T�"�Ob��y5���e*(0��Ax.��/�����t]F���ka�D(��s0��g��D���*�'<Q1JSm��eS��sM2Y�f	?YjE��-��罐"���|;�րSrA�Ro�<�~��D*�0YbVM�{G%��F��!���?�<���<�p����C�����N݇�-v��n��-%�\޹�j����M�0s�g���j��D?q~^,�s&y�D簡�o-hG��h!����0�YP��mMa�[������e-TV7���W���1�vs���֕��,_��V�W�~?6]YuY������#Qp/�A�Y���Ūo^bh�{��#BuĄ��
���؟Gr��u���A�b�-OH�G�}b����z���&����������A�����N˶C��f�վ�+���?�V���1/ju_��2�Gű� u�2Lݠ�it��4k/S/M�O��qk�̒��_^�V
2+dv��!�Wp�Ke/cQPDt�>$6$��'����F��Q��D��n v\��2���n$߽�9��C�� lQ{:�N�������4q匒����l���Xޝe���

F�
�Lڕ�mK�[���Y�#�S�o慮8�Ŧ��w�R�}Qy��5�V;��}qb\���"]��m�o �e�R�ᔁ��PJ>��?X�4��A4�+i�|fY�2�G[s����wUd�JO�W�Ȓn[\(f�RWI���/�H8��S /��\�{�D��IPE��VxRꋌx S�v=ѧ��VejX3�|�	�������/ф�ck[^9�zF�Ĺ�c���(׌��(�H���yeQY1�����.ٙ��+���-�w��uUg
,�{��!7&�C�b�}���U�+!���z|r����>:��x'�O��
07��ͼ5]9�j����8��:x��s��\w�e��Up���.�AB��ʇ�.��--���E Oƨ�n���0���hna�~ד�pQxt�r���ܠ��I��H��>\�6��?�ee�i�e!�����nT��lT5��2�V��4Ku=�}�\��Z�Fp@���:Z�_�١P�H3x2u�r�&�~"�)�����GL��T��%w�+���61�l�I�{Z��#���{��%wD����)ܲ�3(3��"Vآ3���1�|����e� �TmN&JV�g�����Ӣ2v&O�ru:�G@�M�ʴ����u���c�#��{dQ���|3�������_�AS�s\�'�2�� 1T���!�x�?�Lxp#�g`E�q�ji���D]8}��'hL�F�5�k���!�f���Ew��������X�»����=��-2�$���zD��H�hu^;��X0Ї�c���Q�������w�ᇝJ�����������1����+0�
Q�ΝUK0U��4s��Jo'|�L�O�¬����9�v F���>(%�
1��h�r������o$�������:��p�=��*��)UGcH��~����1F^���4d������ZV��i8s�ĲA�����dM�V;���T+��h����#y��[|q��VQ��H�y�� xCBb��hͯ�R�gּK�%�KI��1�_
�Vm�5����;������ȗ�b�ma_����H/�$��Zʆ���d�vġo��}�"h��������c[xC�N:��Ɓ��k))�u��鱜���0�<��U H���y;�~���f<!4�nִ�g���j��'�9^i4�4g�>U���VX&_�0\z���7Z�Q��h��J������T�ڈ�k�+U��LǼW��6��ʣ!�	e�Kȷ#ĚDa�+~W&�Pzd�������dҌB|F�k�H6�LIΊ@V�,�?����B�����,K̰�'�Ǡ;�a�yg#��9RE]��A��Sߋ�bi����1hq�\�M�9��Kݛ�ԕ���\W��ӥ΄�D���4\��j�7Uj�.b��5z9Z	$�@���:U��z�p�
�
��9T�,5��M�2��� ��Ð���d5��m��e1
H
��X�I<1%R�;mI�������X���S�!��<�FWz<���al�mچ�]O�p"�d��e�W"0*���N~HƠ(�o��w&j10E+�}B�.��*\YB ���
���|�x�q����b�T�| )�.j݃�U���D{`ޮ� "��	���ZO�L	c��Ӟ�nH�n�\t,>��ϒ�ka�:�̆b7�|@��W?iw_³I0�4�Z��Vas��uV&��k4ݥ�C��u��ЛV�ƿ�Q��}~�t����g��8������1e{��q|;�Â�K1)( !�ӏ�u�t�b�b�A�UAUO��Y�ʟ@����k��I�j�����,�*�V�z7����ږ��\�����+Sz�#�dM�N�TG��:�Qᙿ�]osբ��+ǔ�����R���'vZ�' Ӫ?�~��aQ[dxc�:y1�Du� �Q��j����岳N���!)�iO|�/�H�Ӱ���l`��A0ߤ?KyޞÁ�-܆�����WG3ܧ��EI%�k��ʲٓ��J��F�c!��E�6vcYՁ#�mp����� hq	!���?����[���y�Tu)�r n���h�Z�E��(a�W��㵙U�m���q��mcs*�˚�&�Ư\��>��ߗ�lv ��/�h�[�E9��tX��+5Av��|T��,PnS�b۰m#V�s�f��ߥ����ZT�T|��܆��+���qg�Z��q������$��<Z�3,���L@?��_!�R��*�|�WI���X ;��ܐ�C�&[�f�x�����r��55A���M�))t��pXcU��u�Ȭ��3T�+`�0�d5Urj�`[�]^�Xm{�����D�����en3����	�%^�tb�Ke�L6�	��4��7NP�7�W�+̲�f9�<��Ž}��%��)��F���!����}p�^�/��������4]/ ��v�Q��A#FBhS$V�oRK�$�4��SC�@�F�9��$D�0��F���� �cWO'l=��ݑ*e�R�\`0E9�)��HP�q�A_E,�'�w-r�bsH:�]�{-]������ׂ���e�\*U��Eo�ݯh��Xy"L�I��7h=�?��4;��ot}ǆOJ�������)Ʉ�.O�m��J�XvK�#@� �v��S�z� M<�RE�Qf@u����
�@�nDu�\3M��
42�����2]��uŬ�I�Iq��g AWC�JPx5[@0�/$��d&9���?4�̭�Iy�T�hi&��f�Щlۊʎ�z��e�5t	��W*�
rD�tGu/h=nrN�ix�:�Y�e������OCVC�Q���.�be�Ii;)�d�?J��~8G�m*Y-�AծA�:�OB{"�j��su�(�R�x���̐�fT��A�4乑�i�=�Ĩ!�E!�Rl!��}oL*�&N�*vw��������m�5:vKd�N�I�)WԀ0�e�_�:J[�λ}"���$�n�u�XU�WSc�R��-E,��6��˙��T<96��I$-�+�?P!Qo�G�|5�T���z�^F��?AAVҩ��(,N��4�K�1�� F�m�W'Ƞ�M�Ka(��x��Pw��'��*h��?ze�!Y&�r��n
Un/[��;��%�ʈ�+�9���	��$
ܪ�,t��uBf>!�<E}��CX����q�R�a��;a�(C�a;i[V��>�D�jZ05f'��z	��+�4��eܬ�f�W<�x�y,��rDDh�F+��s�KrD�gs��[�h�8�P��+]�cr���A*��ۚH3�UyI��'��B|����D	�	�AN�on�A*-��y|�!	My1�����<����f*|�ao��6s*j����xk�v�2��Fm�?���=�e.��'���S\ui��/�����@�.P���ˆ�Q�a�Q���^�}�&�L�u5�*�oᅓ��D7-�e<^���?%͕a�^p��ˈ�*4m��d!��c`v3hZp��������!R'�B�����{W*�Cዋ��귱}
��d78�����p	-�(&+�=	^4�_�Z�l	M�P������X�6{c�YhE��, `a!�l+S�m�L������ ��&U#5�`���ܱ�Y���Vc[������&	����LL�u&�c�LN��³i�K����ۋ+��	�	���P�4-4�""���ͮ���rB�d'�
4\�f�ڴPF`*3��swqܑ��ڒ��-��ҵ�9p��j�2븠��]0��!z{�<[M��2����R���i!�+�Z�Ꞓv�E�T���%�fǵ+��f���d��JO^b�f��E�p�B>y�=Q&�r���FQz����}�u��l�H�4>ی 2$�;��K�������o>sż#7�>�jB'��[��j�. �X3�k��ZZ����:��6�ܾ��,EL,\kC��J��Q��yw+W;-O�Y�^G��8m~[�q�(�A���d�i���Ϲ�#�,ʵp�[�y}	���s���A��B�+�ѣ�i�I�����:��m�����wo��*��|���	Z5�[�B�q�p!^�oZ ��S/�]~��#/ػ�C�n^ϘO�~����B��2�����gd*���=�<�@�_���f2�qS� n/�~U�_r�a W��q�p'8�!Ծ�
��a��c\j�e�>D���L�6b*��J�ߓ#���HON6!�&��rMv��G��V
��ȿ�)2.��=���6��D�#�GL��hj�� ��|eTQ���
5۾(�زȞ6����g(�d��	K�P�1 HK/-�?t�<�|����a���!0��C^�>{p����P�X��Dj����J'��m*aȼJ\I%f?_v^����5��Z�����ʄ�NART��Q|��o�~�!c�dvS��;���ɠɌ@� �Z��X�G����m�2���"�9_I�/����(��� Vml��� �T2E�!7'��y�����Y%��c������3���I{����3ZڥFya������k�C��x��|�pNR��9_|����P; ��{�ޘL|��2/eN�E���3�R��_�USX4��eN��7v��"L[�M-f���t�K�kM 
��8ֺ��6�Y���2��w�
���M�d:'p��/��1�(EM�ml��r"El72�s��1izro�:��#���HЬ?Iz�n����J�
�ⵞvA`��+�<�
/^�$1��=�S���$}����^ ŝ�30!s
�Z'��"]���i���,�MD�՛^�*3���k��P��-��R̆s,�/B��*4��?6	�[��<�[�v��Қm;V`*(>�2W�T�ϒ�Cvu�`�'���{���@n�7 }�x��d㯞��{�hN�sD{�3lg����������a���WʗP<���1Sz֟�p��E�e>����S�W�D���/�Z�"�ʵ���|�_�Q`_�9�8��P���5fDֈUuy����t�7(_�L�?-f����`E�c�aJ����*`�R�������a}o��֚ֈ'/���x������j_W�.��&!��MԾ����<#�*�G���^%p�9P�^D��N��MFV}V�XpR�lD@��&a��C�:���6.��2Hcn����C����_����#HA����~�I��GC�П��p����;`%����&(��4H�gb�Ф��qu<�����UwoJ�p�M�P*8��	��'�7 ����.�Y8���J8��:'喂!�p� #s���HlM���α�ۨ�K�nܷ������R���
������b,9�t����>)�g3d�|9�YUX��Ej-����D�Y�,��P�&�M�-o�	 �C\���!y`0�øk�=('��Sީ��x�k�[���\C���U��6���m�����4��K)\��3��q�D�}48��b��p��@�WYÌ��G*}@���nZ���t�wR���_�����If�*�+'�p.�A�ߦZ��5ӣ ���
�=�6	���e��(�!�v�v����3�10�Ag^4�:�9@�-�c�Iī(�R�=����1��_۲t|��GnM�z�S�S����ʄ�V�����`6*�3��C� (�.8�����f�#���Gd���)lxf��D>m�O��9G�%�����E����3��u���`G�I���5�g␘k�b�i}��K�?����x�W�xpy��W��r�v˗#�ݮ.��I76���4�L��M��8� �ϭ�x��m�����	�8Q�,�B?Su$�S\��]̗2�7�_�}rn�X����z�ym���2�l����t�ñ�%�������G�eq��p]� ���WH�,L=�����3��R�&Õv�),}tMa�%0��&՟��T��k�j��(ZE��JO������-B�����ʪ��f�_{�����-ğ���,���'��D�ӣ�`��±��(�G�Cw�~i��F�g@Ӗ�[E����f��nB�V(�k�>*���#t�u���,��H��d8��L�Y8��,���F8�)��[;l�\)����JQO�s�ED���GM��[	���-D��/c��rʃ���2خ�4���T����B_��\�s:*R���2�j
�;��z^�qKA�j";]Bc ����7��K�Ύ�M�jB$�����@���RH��5^T��E~��z�gՙ�)�U2���\��NB&NW�w�9���D3���t4��a��{�����.Fz�������n%:;]ԯ����%s�W0g����7`��{	���%��XXZ�N4)�[Z!n0i{�`��q��� bFi�^�����nH*�**%�r�����ӡC���K��[�;O8l@��q�u��/���9f�T��:����2uf)��Tb:k�ջf����PIG��)w�$&�9��x/r[��������n�#�s��R9�ƀ��a*גw�qr�N��:�%]��viE\� }� i�?��R���'ۜH���^0���y����,��_�'�&�a�K]{D! u���*����Qk�1�ݡ��n��g�Wwq8��o��a��3nĔy����ٛo�lĲ
����A����}[��`��&!��!����_!��-�������$K �N:�/DN'���%��l�!?�����Y���9��!0O�X9mRQef�8�-�U�����V��R.E�|Ɏc�r#��LߔXf�˱^�Ro������a�r�ɑc�a-�6.��|ՒvJ��_���T9�>{D�����G ��|n�A�y�"޷�a�Շ6�`�y؅��jU$�Q'Y�K�� \f1�X]�5^�����%���[�\�*џ������kK��=�)��7e�y�"���ew���*�lwI�WIq_�IJ��܇}!�d��`��/|���L�������5�gq\a`����t�c����6�����aK��#�xb�?��|���[4P��L����x�����/�nzX�v���MtZ)���lw��Q��3&��˶3�]��Y���Z�j���>��ۃ����l������k�S �0����<�$�ȫz����G��_h�3޴t����� ɵ@����/����V랫��3��ҀS�Y��\X.9?�j���1��j�β#7�R�K�&���!$`EW�)�i�������TT���g�Tl���L
���[NAϔxl��\|2��S�%�� 0,�t|�� ��
����1kA-�Œ�aV�Uk���]U#//�=%�1�)	g*P��*a���9
��6�����2�T�[o�-rR�ꊚc5�=�]]~�ǈ�5������������@L�F�q��Y���;F�'�'�.a�	���ω��)$�cX3dZ2n���Wg�~Ll奰*��T�%�<�Eլ떥3{O3}7�7dl�ڞ��gܸ"D�.�����:hȯ�����W�D�@�%����Z�!��G�&��bn����6i�~���C^ms���\쐛������el���_fFelPI�~�{�6�<�[�-CUc���[�f�z���N%w���6�țFU���p���j��M5�ϕ'B�	��F����[�v��͚���5}��i���K4kU^��-$6&�gP=a{$#�;W�7�pJ�q�pfn�+��a��M�mt���R`f����"q�u.���Dx�{��I��w�[N��#��]A����e���猅x�phW�̏t�kI�İ5E�����c��W��5z��ቦI�\>E��j�>��3>����R�<L�f��:���J�+�wܣ���Xy`٢U|���v�$=jX�/���UC��öH;p��D*�P���I�v�s�x��$�����l<u��\�?TƑF;Kb�4��.�7�+����W�F��oZݷN�ko;��%
��������<1g�&~n��P�S<��45�� į�Ǥ]��|��l���$���J�wfD1T���ѯm?�n�7��SuY�Վ�DJ�ff*���7���z��J9#�@�9���˥����H���T�6Q@%����o|YJ8.���A�V��h�A`
�"�{=�g �H��"ʈ������^ p}*·����i]�-� nى��p>QwR����֙����Z�0���WK��N8m T�z����#�|\OE������a�C��\҇]�&�+��c��L��k&�aۚ����h��f32��}��L�%L�	k��}�IU#9,�]t�+���+�b0p���8���` ��R����9?�GY�˄��r��HD��W��s�!�N�̚��a��p������2Q�%�i^B5P�@�21*��H\��	RXC�bf�Z%�&z�n�c8[:"\�Eȸ��k��
pw���?	�&�D����gکԜ5���'c����:���������U�MZE�o�J�	�6��{��k�E�>����[�W�U�
1J<�;؁R�l��ŵ<D�]#"!��y3B�-޴�������a/[+s�L>��C9M��M��z��E���+
`à@�I�Pm�y�-g2�������?�k��_c?��@���t|� �.1q�.]�O�
�t�V���A��m�?�N{�����ek`�]���w�.~�Zc�=k0����:j;np��Q�L�� T9:,Tp�� X0���ku�q��ÛI=��Q��*�
�On֧����������G��D�N��~O�f�d�ռ�oL[7v[* �@$�2uf�r���nﾹFS�f|��bČ�r)���T?����l������楺����B���ei�=cO'��]��T�^c�}���s2�9J�fwP�J2�ȕ������|��I�/�f7^�F���������sɩn���\�����&��-(H��<��f���`j2�sm�5����^�6E"�+q����ŗ��86��ȋ���ꗌ������p�>����H��qe����̀���%2Qb�a�}�6����*)r��<�����1������s+���B~o���!A&X����Q�A�;q�����L��z���Oq��\�fS�(�g,Z��Z�i����/�m�*�5C!�z���&lݸtxe���h��a�*�r>#�f��D�)�QK��a��9h)�O'�Y���1K�{�]��هnE�h����v$=+�exIO
�ҋ{�1��Q��@Z�|g��:��7l��|�?�E��#�j����Q����ߧ�	��IO
w�!bځ,��͉�e\<Z���G�����q��(TFЍ�?I�&Q�R���^Y�h}$���}���a��N�����6Uf�UL*s�}������9�������`�iM�6�0%����5�cdIƯh҉��Ð�)+=��;�F��fD�����:rӲ�Vgi�dt������Ѓ^��q���"�]�[�#��K����y�=)a�'�$|�.ͩ��I%�d�gI�,�%�T�9�%��43�;I�͕N�^�cT�
�7��KLr>Q����%n�y��°1#�h��BJt�kh�!H5��F��|�d5xo��yǷ��lp��#^�;�f��6���0<ͽ����˂������b�@��r�A�x@��k��ҿe�nh6�X���t6�G_�W��,��C���|6��(�� ⢅2�]9�$���Yƴ.*�~�O�q2���0������4��4m��6X?���	��� ����1v��6��ݎ�5u�u�6��k�l�� ����fj �h1	�K���â��g��怦9�@�rh�4)%�iA����X�x�ՊM�D��II��e\y�:���Ê���}>�䡪�NV��e5^�KG�-��x���]8�0�k�d�w�д<>�N�����
�6�f5n�P���c%lߧ�,aFn�Z���X��F'R@�'�q�@���}Wb�J\P)����&s��FCۊgp��V?b܋yl|s5lZ��Р������NSWA�����L̱=W�?}�7�W
1��g)��7��'	]h�����V�/
���H󮾦�ӳ�Rҿ�Б�lBW��l�o��5"bL~����Z-|ݯs�$(���������d[��.~�	��N6��a�^|�����q�4���اd�TP����5궁�y����-Ю����z��:����EAk�y)�8�B��Ћ�Xs��aO�8f�"�Y-9�sy�<��<�d���q4������?>���!��{�|z�*��q3?�P�&.��-����Rz��ʰ�Z�r4���M#)8@iK�����	w4H�h�b �*X��a�-�'�	W��0����3޼��j�'hj���{xf���o�=��BW���l0|���g�A9��2�<�#Ok���!B� |���cW�����E����uZ��J����'y��4�^FA�+��Ǒ���� �F�1m�,�o��b^.0�?�!}���*iA�R8��!x�,�8�x`oj��i}���w;*��bg�?E��������flN�C}N0��׫��5]�W��M�U������ܯ�E⛪FR�w����h����FQ#�"+��趹"�ʴ�|L�F��L���&g��#���K������Bh���L��w�lzaT��Q+f�=�^�)\���>�V��_�=����MV�ʣ(�k'3�4�Wu�V�Ī=��C&ӆ{�.n\��� 6���Ji~h��"�zl�i
:n��&�����u�Z
�h�����DL��2�k���Xdl{���B���;�������F%88�c{���c�$�^ی��: ��+`42'm���{�:��l �4U��=�V��WV��`xӸm"z���Vs_���h��Ɋ-�#{�_e�D][��P�	)�\�c{uN��}J�፱�6�T3xO$�M��	r��QHs�*�2l��ە��7h��H�����)�e����m��;f���z)��*��� �y�O3R\6�d�2��MĞ��f'�N�g�Ɠ�P�M�<�"�{a��v���Ӛ�x���C��<���@}���/��\��z�w5T�t����σ�d@�{ ֻ���.��v*qM#�I/������,����,��s7�ZO���@�����{|O�V%��;�6
f�ʮ؎?��.��	�B|�Y��&c�����r��m7������N�7�L��A�W���*�f� ���$W4�Qs%Q6܁��: oB�Z��s�G߇�{���C���B�[�-L���yV��V�Ya����R8�=Χ�v_�r���Z3I���ī��2u��mCϑ����c4�$�&�J��h�^��'��Zs\z�\z��g	���?�ʓ� �x^G�;M��Ke�4����F��1^��\����b[��(�߃j����u��Ě����\��9�Ww%L<��f@��F��u;	�����T��ӌ����lEy�#��v\rj=ڦphf�|K���Ϩ�����#$'oF�&���kd
IKhltُ��y�3�[�<����=��Rx��CgK���-� hi4U�ϜV��Y7B�bПe: U���qbJ6F�K�ۥ u���X��S��ҕ�Z�$]"�BP�|s���#�!!g�=���S��߄[�_?!�����_�&�Yޔ�u����#���p��)�8���ۗ�E��	`��Y��|?3�����Z�?�M���H�f�&IbU���(��$�$���%ē��Sl��C)3 ��Moxx���DG�&;f��<]��ۆ�U�8�$���1b���c`�T� KС�����M�@�L%�0H�� ,e�33ңLyq(�k��ܺ����L��*H�3ny#��4�U���(O�H#z�⿇���ҷ����u�Ja��&X�����K5/Zvć#���z�cw~շ,(Q�84C'��,�}�b�<�[<FB�{�g�i�� .�	�}�<[����
��;U�з]�m'T]!�2~-��Cl�r�p]?�,.��V�L)�������DT���.����K%ѡ.f�\�ߤ���tww䬅l��;i��̤&�q�9?�$��H;0ki����6){w��h�|PH|u��O��/�,曧�+�+�8RU�Tj?�TM ���|�]
��j�%��K�D���.��N+ˍl;o���cP.=}m&c>�&3������q�ɻ4�k�LP�f�N"$K�h���+r+�x7�������Ht��A��t���M�y׮��gy�xO�H��(��7p,���h�����E���3 �{�����5_�����*u~�ҝ�V�W�z.���jw�x�u��$���J�%G�B*�O�^����(4���^��܌$�#(�L��@�4��v0\�c��]3?�d��e�=�`t|CN|�"^������.woOK��C�K)��}����Da���%=�0�/�����49�r���e��$h�����$e���.ai�'�K����]��h@;�e���!�"/r����<�h�X��
�&���@��w�J`��׀�� �U����DP�Z�{��)Q��z��+����O��d�����o�>�o�'�]6���5lI�&=x�P��}p~B�0~$�:�!�ȔP�	�0��Q�SL� G����]m48���g����qo�w�g��/���9l� \nB��h�>C��]�X}�q
^�*��?|��X'��7����ٷF�E�;�|r�i���ح��=ۏ�b_������5�{|��IQ-O<YIeW"�-�\ʚz���B��^������_��H�历¯�L���k84�܈	�|�{Q�����"g�-d,���['�&Il���DB�?*�nZϱ۳�m���TKHE�F�������Z�Fξ�L���s:�nb���n~6����_ �v���8Z�Pu%+>!�@q��Ā��q��=f��V�7��,�r��r�����v��s���揝6�U+��Κp̒B ����H�蹅J��Ç iUC`9PӰ������z����I�n��IH�X��!ڐ�uZ��K�=S[t�;�/g�7g��{�v�YҦM�
�]U�n���MoJ�V�Y�Ɇ�x�{�6-K](4{�iRa����1�v����/:�v����v�a�HH��u1�M��a�Pz��o<ܼ�0�R.�����!���(}G��{�hE	,��CIL�~[@���7�<FCi�rwa�����BQC>2@�G�+h�w돺І�*���Ć@VY	�P��%KĹ'!f����}0��)�_k��H���I�����dH�taiS�A0��7	C��[��S��=���;�E��3�wQ�|�����9K��ɭ����[��:0�}A��pֱ��y�<��W����ʙ���r'�)���^���v�P�,՞1�t�~�0��� Z9h7�����'�� p%��-ǰcx�¾ZE�b��k
��?�_�A56�7\�5�
�@-��<�
����q:hR�k&H�#���z�'o�x��1s���ґ�D׾���MO���bq��k��2����;�i;�xW���&;�1�,�.���L_���[���"����t���������]�8.���c6��V�ϲ3d$���M�I�����h���PX�K\S@ p��g �Z�<�LǬ���ld����^��_5���փ�k�B%�lqp}`�@殜��Qߝ��G��>��,���dǥ\o�1#9WJ`K��"h���;���.��rW9���԰l��t�h��M�&3�Cw��v����ڲӫ�#�^�S}��xW�˿��]�U�����y9J.&�N���� �Q��h6��"���C���K3;�?%?!C�
v�C�N�݄ibg�I�D x�z[t,Y"o4Ե(uZ��w�|��<%{vX����O�~:$�'U���5V�$���al�"�c���Є^��%ʡ�Z��r��Ƃ�8c(Ƅ�T!�yL�&%ؙ�AM��\�w��W̴��ml�M�m�U-�c�u㫹��%�+�;���
>��%K{p���l"�{)�Zv=�ȐNY�����sⳛ!�D�	�c����6dFƙ耓���g ��t�m���U8�p[v�4qI�*�X����.�,�a �
�v������A^2kZ1���Jg1�? U#�K{Po��^�|`���C��.��;��'y���&�S��
[
� �o�_������{R]@�������3�����8�� ��b�Q]~%�1��w�`��{;�@&ٞ�Es��9��>ؼy�@'�!�?�&�7H�U/�?��G�K��Z�������W�Yh�`�ނk��|;A{l��y�����	W�۱ė��bZ�F�������EOQ����H�Rہ��QKTz)HU�pٴ��"�&-V?����;+� �!���R�&�i�[�+������m���Ox^���E�����������ĲXd?z2��y����h�G��>�-�X�p/F���A�"�UR ���~�n��A��X���|�S��~�����J���j}1�����i���d�Z�ۜ�,a������j���Ud�D,�� �O&*�+���Ixa�&#�Ի,X=Z�S��a�ֿe�c7Y>*��x�~�F��*�TH�I���w���zW�w�Ɔ")$\�?T���Rw_���[����?Q�~ֵQ�ݕԊ�.r�8�T��}%�������JKD���
GO������}i��|�cATr���}��qэ�w�wQ�*SV{3����RזTA��i�Њ��'�0���2��"�t��#�֊�$�w��S���j���DM �n��.B�\����!uI��\���Ϫ;�s���X\���͈����]'����lC����_�^�w�P�}��/l�k/kva=�I�%���m��U\��/�ê�:QMj7l�Gm���wr=T4�V=����wsVF*[E�k�^M���$Y���3��Q���>�v�;Xm����_4�3m|F�d�l_���M�N�(�^t�|=���E�4��AL�?�sB�<6�b�g�<�������ld�$�����c����?�(ߒ��������>�~z0�_��\����h����>����\�Y�����.{���{tp�򄍲�rH*�p��PLPc��og;\A̩4��0z�/����k��$i(�������f�lMT�ir8��&J���*GF��P���$9v8-�u����&�7��0`�ߟ�A����c�Y{Vfs�?^�����}�Y+�T<���8��{�$߶X��U~U���2ZZQT���_�{T԰�O�%�1(#Z>hn��)Dë���%�O�3�C��FdAt.�c��~&R�5[��`��<� �w*����96t��t�����9u$���Un�M��h:	���٬MSHБKd)�����m�r,R��y~ ��۸v�˧�X
����9��M�Swu�l���?�WD4�g�"���T�.��u��:���!��%#{��yɖ���u����?60MNv�`eiF t#P�Z��Q��<I��tt���?y�L�q���>�#��}5��f��H9��־<}!kzs�!�(�ߜ�#`X�o�j�.K\�[�x�2j��c�_H�}r&0y�]`|�U�5�Wf���[%�N�E7��
	�5�q�:<l�Yl=�\A���38C8��Qy?Q�4���a�����m�3��7��/��'�/-�H�_%�9��h��t���R��f���ՔV���7�םn��u�k�4��Y�fTi�V�8*��0ry�,%R�y����Gk&�8���Q�j�� �z�*Lp�Æ*��M�~���Ak���$�%����\D+�:k2>!<�!ʼ������d���p^��⾼O�t�A%jB|B��p�SޙU�O} иzзH���*���oc��:�'���M8�����ʰ�reܡ�-�;�̧�얦�U p��շ�v�!�n`��NDnW����z���	�9����z�Al 隅�'���AS���� ��m\E��r�wה��1�K,�`'T%?{��?�L��*	�rD����Ɯv)u�Fm����>18�p w��҃`IM��G�<"��T���=B�c?�����6.�X`o泫��6�����K<ԩ4pmq�#�����k{.V�7q��&LF�v�w�к���KFe�5Uq|�:�Q��6y�$2�B�~�緊P��$�8��h�8�+eA�g�a�9��w��ɧ�ol��u@7�� rCH:�����v~Qk@����3I��,��]�r�뿉��O�Y���!JFM��&b���g��taW���䠣���VZ��ʠ���j:�&^�6�ӿ���4Ln)e�!���UaH������RSs"�?I�@�af���f- ��*p7��R���1�[3l(�Z�x�{����+��z�(M��c E�r��|�'�W�B��p�9�s������Vt�ZzW�%h!�,E�V0�U���S�o���0r���������}̊�Jg,[�����yg���{��w���N��m�F�=ȷ����u�?��ߟ����WBz���#ڛ/��eA��~Iŀ����U+t
�Bs��ֲ$�?���C,Ͻ^ޔu�H�R��sBK9��R�������؊M�����$�l"��]��(<���$����2gMq�)/!z)����\u5���=�M��tJf��D��-]�ՠA"K�Ȍ�X���0-$B�E'��	vX���wg?�	J���Wj䋛G�Ѵ�t�W�{@LJ���;�_�]�j�*�-������ f�m&�E���4������!�Γ����'����"�J9w� ]�]_�7䱎
�bG���f��d��Dw��2Q��$����t�lIv�z���ȵ�M�=��F�~�o�c�0���{��3ه���Ts�ՕO1"*�i��]Uh��`ʆ�^��(���x�PT�gMjƖh�}7�����\WC�v��9�+:p|�dWZ�.F���ov������S�J��Z頶���@���P��R'�8��m$Nnq}=,H�y�oMU��7<ď_�Maoy�v`a�y2��F�&4��#"S��k�1D��*�D?-w�i�V?�_zEz�ϴ���'��>��l��k�W"����������7eI�llH^o�6�:'_�;[�1'!�"4w��'ɽ�k�.qY���|�i�|�.y����M� ��ml'oPG�w�p�;��E7hnQє���]�Wŏ0*�[�M��:���ӟ`�٪n;k���Dΰ�.E��c����$姗!|ʾ�26�j@�S��c9���k��V*e�k���v>=0Kr�X$i�/p�V@����D����@���3���R���>R���3��%��5�6�%&1�̝��$�*�SR}���� ^��Ż���cO^4g9ֹ�O9|�Y��F�:�q>������b�4C~:���;3�K8Fi�tt%�[�B��τ-�+����"�Ð˘�_�=����f=��Z�3���1#�5E�;�c���k��n��G��c;��
c�Β]�[m�-g�f�O �3�� �?�B����i��W��-��xa�f�ɊƐvJܯ�n�{�i�Z�R_;8M�!@��E��R`�e��1�����<�t�De��>���V h�<��/���;��D}����$�}PZ�a��ۘ�-�!���L�L���@���BZQ}���5;��t{���~,Ձ�����rBO����) ^p�W���Ub��1��x]�\:��DA��J�����bh��(�c����Z��D�=EY�U���5�� ���FM�_5�j���i`
y�E(Z�b�������5�Ď�l$�6�@H�'S�2��҈>i���Z��p�& ��l�]���I{��힟ćԌ1ñ�M}7f�Dգ4�ޯD��A�d�N�w[���~n5��ɯ~<�-K�}M��*�>מ�7�R3�@���N�O*Í�C���50.�S�`��r����v��2�L�8"�fx��-]��Ma�h�1�TT�JH��֣���I���L>����
V�/���Y%�	��^��_R�$"M �=%��>����e�e��������op��bU�6+���!j�����CAaIV�������6����dd��qyPVr��2bB��үN�<lK�p�Z!�!?��v�����X��ѓ��v�oOR�o��}��-]0����2/yRe��x�����8��\����ɸ���(x���3)!B)���S�:6恎-0j���1���)ŵ�Q*tJ�n�Ỹ��T1�ݸ-x�!KM�LM�13Xݰ��^ S�wȒeeB��n$���b�GM�8������W]�_A�V��t�pʛ��;�����ĵ��ӷ�K9�Yl!�0����3�n	�a��^�͸����A�?�smвY�A	"�y @�]��?f��W���	t�B�Th�s7�u�FQ������Fn�'����A\�IƈJD���d�1%l,�������w�˃�!4���O2^x����\��"?�*��j*\�)Q6�3�Z&��4$�2�������!C~z�ng�YC�X��v��k������~ H��� �z/��I��$���&�x��bkc�qO� =8�LPrE��yS'�<��xB��d�m.��㷪�!M���hs�="�<� /z�9p:��`�Z�d��%�ےN��g�O8[�;�����������d`D����b!�H���7�OF�k���=x=6],�:h.�x�|B��X��`�h���$e퇧�@�X�����H%����WXAM^����G3}s(勌A`���7����f�|����n��R������{Z��i햩jjr��׎�=�:E�P.����d��;2vaz��Ɨ�b�����<�&o�����3��:։ue8�t���È3��ª^�®,ID��tv��#�#�#SO��dw�,���S��.�������x�Eg�޶�Y��3��Ro�C��)�%�B m�4b۾^�ry�~�{�6ny�J~u�M*#�3�&a�zb�m�n���T q���� �7[��]CƔ�@��,~�ʥJSN���%t�!S/�O��nb^n~���&�`N{y3�D��w�,u8���˄� ؚ8\{����N�~,�	�����WaD�XT�:z^�3����V+W�f���4���J�?��:y
��)ఙ�c`�X�� z~���V*�����Z�δ�+�[;"��T�m���Y��bhf[�o����]�c���c9t�C[�9����	_5�g�y�UZ���s�qLΟ�*s&�w�*�䆞��U'.!�}M!��v�������ө��c?�v.+�-I��'�6򧜡��b�!�Q���2M�<�����)Wv#���R&8Yfb ;�R���b44˥	h�,�r$-�(��@��m���a����[���az���`z|I���~� |k����_j���
u�Ѥ�z��j�R1ͿI,0o}��Ń��?i����8���]����r�o1Y½?X��������iq�����9��\vH�7�3E�jB��Q/��g��*$¬�\^��d�1ܥp �ID6LL5��\��ZNθ��?�WV�i���H�}/T�B�\-z������P�T♻��4"@[T,xoО�3�QISd���lv�_�v",#�@�fx��,4F�b*1�G�$ S�D���U���{
[�s�K-����u�ZL�[� ���㼏_	���ԃ��k��Ɲ�z���>�Y��H��wv#�ٶΔ>7��H,�(�X$�ˍ|-R��m�	K�`�����O�d��{Fmd�
�]�y1�=>T�!e��Ϟ\[�� ��]�T=�s������d�2lf1���)�]y����u !)���wV��:٣�y�(,������e)Ў�c�R�_-J:MաT�Χ��
��x���Jx6.�̃�rhi��L&�If�Nn>,��f��]��.�d	mI�+�"�!�R� |و��=-����~�a���8K�E�x�u;T���7q;"�]����m�O3��Mg&d}5�-`ޡ���D�bPZ��wJ_���eh�%o�0o��1�CWh��;
Ѹ)S�X�c'V��e��K ��>�(��.�}�WP�q���#"��\%�(�����L�rIϴب�@�����E�D�{���t��e]�ѫ�yĝ,�xA�I��> r�#����=��w\���H�v�Z�q�����ѱ�J� �X��pi,���	�t��%�nq�<b����Ƴ�A��	����s����]��|�si:5��DﱊC^��I0����͋�T�4-�#��� �i�_uLG��H�0���"��F�0g�ϰL���r�?��>Ƕ"D+�*d�]!�ԙ�#;n�Be���Aw��`��$�dsۯ���i�Z:l ��O)ы��`�Ӭ��Q�}J5l(���bȱ��� Z�P�6���zÅ��j�m% ��q�{(~s��Ւ�x]���ƑZ�Oc-A��s'N2>�>r_in���4�v�����%�2���>��s��:bX����,'�� ���C\���p�L���!�=�1k��+��Ó��M�Z�X%��N3�A�lF�����J1���tFp%;���f=��G��w��9u���b5t6s��{����J��Qm\lu-ݍ҈QQ�3
��e�:�r���~�%LX��ƙs�D�k+�<6�	���N�8�$E���#��kp��"#�V ���,O�)[!�2e��6J1 �I�M�xb9�2e21�b������G�qxX�ATV���|��c����Ϥ��Z���j����'1����h�.c������fI<({�&��cS$B����̂��e� Ib1�N�F�Æ��> ��r�=.-��M�I�O��(��;�;mf{J0F��Lla�p����:���Gt�m�u�����hA�J��E�a�C`�����>:��-���\y#Q&נ1�����
�IP%@��b�L#Uj\gP\��ǉ�YN�^���P����p^�D��}�'�ֆDC%4��E�Q��r~E��tɕ��x^�؀��JV�gO�9
\ҁ�R�HB@��h4P8�>(Kq��a��J.{,���M�4i��pQӕ0�V�w~��fn� �~I���x9LaB���3�)�Y�b^��C�M�w)�,�V>�D�Bo�z���������1�]��a�u@8���h1��.�4ZQu��l�n��cOև~�!M�d%H���Z��?�AH/����bm������iAl���f\�Q��?��긖@6ZE���[� ��yA\�<?������ ���%!���(�,�7���ͪ��跎d�U��Jv�*b�~����D��c8%�����N��v���R�y��a�澣�P���M�t�w��`�Nu�C��3F;������{���d��������KR�En�F9��Z����<a��k���-s�{�M��k�C���pjOa��$�$��<��@�š4'+9��;B"�y���&4"���n��k!��n�$�V��[Y	×Kۂ�.n+������>U0�I$�; K��$鉧�r�)\�1�@�hB�D����DYs�y�w��r`{�S��)�'=� ti7���>���o�����r7�
%P-��w�<�a�B�t�\?[��n�>���$%���!f�����U�o�i�u��('C�� T��	N�����Z�&<�L������_#Bd�F���}��>�R8r�E�v����ӟ_��V�0_�CoC4��Y�g�>fE��I�o~Mry��?��<�B�Ld��α�L*2�o~/�2�+mhs>m���3����F�57 6֠�}� �������~�o�lkVK������͒���r�/��.��ƭ�~"�,֪����N�Ԛ*�:C�rؔ"��At��K��DPJ�jSj\=_o�eUK���J��~�� 'D^���(�o��'Bw,��i��c�#�<V�q pzG	ÚA�m��1���6];l��L���&!ǫ%e$����8��DL=�Lv��kD�ZD�4��>�5���g���^fˮr�'z���u�+	
2�ٹ
]	�����ݮ�l�ԅ�wn���n�/.D8�����C�_fC:F����M����tO= ��
>���`������Q�{*x����s���(��E75�;�g�l�X������S-f�'4~�*45�:�3=����t���=3��?�u{l6J͚����lĽ?�a I�ᛘU��#!��	�G���(f�2R�t��wD�-�ź(��Ją���/���>@��%;ئ�S��N�|j���O�ćs�&��s<������I+g�Ď ���ߋ��W��w����iNu�o��)M񎺜���}K�|�$s���kr+L2��)���������;��5@d���`0}���#D+�'ѫEC�%4X��4⃾�F�g�[�b��KS��8x��Y���9i�����y���o��x��	����KS]��il�$;'3=r#I0��p	���馝6k���`'�y��@�)wO�*�n~}F������;ǪC�sP�� /#ce�'��i6"�Th)��R����a�pˠ�^���w�W��|�ܢԠ7�M-��ت���v�A�r�(�&�G�{��}�0+�{�ʱi�R1�m���)�=~�ՄT�CXS��}�5�3VA�!��U���'O3~=Ȓ� Ҫ��aI�a�-��H���Cs�t��W��C�&�	�t���R���s吠�umg�,mŗ�v����$��eY��dEc:p�ώjzs�0m�n�,�"�Kb�=�x{VJjN�VP�(A���;79���#�<�m$�y����Z�YH�Gl�O-a�x0N�8�{�����l2�Lj[���V�[cG)�7M�É߁�W�?�8(6I��B)��yQ�Q��W�4UWγ���'�C)���uV�L�Xm[��ͩe�!(�!Eʄ7y���؜�����<�M�� ��X����aԣ7����*[�,#��LA���Ո�6Z�a���V0sW��|�k��� s~�Ak3H=`���3��A��W�ԮL0ڦ���f��b��VU�����8���b�a��(��\��ht�<J�Sr�h�����AMd��T��I������e�h(�~~�����9�Ͽ0<q}�N�
���з��q��"��s?��z����R?�UZ�(��w�b���~m:^~����:��\e��a�lh��L7Χ�&�	ٺ�-'�{��L_E�$==�=��6���6��Q��z�9�Y��G�M�K��QA�!�sdf�����.�p�~�ם�7��S3�t �t>Cw�=Ɖg��z�� ��(�eiz�b@1��x��� �"G�5�n�F�Hw��/��zC�ޥm�,�+���k��+mb�cv�-NBY,8W+�aЫw�.v�^wDP��X|\	s~�������&pt0=H�Z|f9oj���cz���tݭ@+��\�
�Ј�W5N*w*e�Jf=�-���p8q.t�O�����	,mO�JB%�G�͸���[�~�WA��s��f��~o���o(϶��P�E�_��������:�o���z-�Z����9 �QT��P#�����n$?���W��:��e��1f}�=�7f�6��d�Za���.ډT=U85�Ȳ�a��t2�4��i>z<[�Y$c���/�iR�P����WӃGB��U��]yb��i�Tf���(k}��d�a/�� =�^��hg���bdds�8�|�A_#5p�'<�-A�� g}.Ϩ�dC��8H+�9U��a�l2q�z⾶�گ�t�F��J��_%V�~i���9D��NBЕD\x���M`e�����uڟi���O��Y��h������;�$ �s��x�J�{:�M��V��;���k[�ӏ'��f�E��8�9���D|!
��������a��_����4W��!g�X��ܞ�5"q��uJA^��>�6avd�?{(/����a�F5�v�u��Ƭ�e�2��c��zu�8������(���}�U�<���t�0*�*�¨���f����	-�~�rx��o��!�eh���\�{=��T�܈߱|�����Ƭ�5��j`M|CL�)'z/��3Q�������4�_>�`�@��x�>�{9�~�R���H2���o�	!Ɣ�z�NjQ�(BR��~���c�n�d�9�9�ϩ�s��{��_���t����q6�1R2��Ϡ��0='��YD���<��q�_�@�����(?�o�[��&�SV��<H�+�$9
�]�(R��t����YF�5�#0h�䏐;�#eMQIOC�kf/�#:^O�[F�儷�ճ@"�g���^Y���Z|�o����cx):�
e��P�a�j
�M)�C���,a�kzO90�E�Z�8�вv�)�-��<,��Q�^���{s��`��1u�X��n�����OW	�S����
���cP	V���ᅕ��jd�s�6l?ybZ��B�@x�DX�tY��$��{@�\!F����~������c
�H��rJ��x_�
����b�a�i�s�X69(D���@��Y&�b���U�~ �h�x7��,s�W�cB�LH
�d�\��,<���_�`�2�{DA���������ʵm���F��FD�e�°\i�h��d�H��Z�cD��l�Ӝ�Ua(�`B#6YF��l����$ņ3n�v�?����l���皺Y�&:�|�����Q��@��ߦ�����K[�����7:w�FʠD�:�XM��1�q��ʠg��_"r��A��c� 6���Ѐ4��{q;�`Ao ��zwf�懿��}�*���BB�0K�����;�� ��ʸ�&'Cd���M!/��E�y���T��i��|����X@�硄����tWlB��
�a�t�׷����$zJ�+r'eDho7�fJ��% �V�`Òwn�=R�2ͣɬ;�(+dg��ۭN�P�Up~ֈ�{��gK���.�X�	$Eق�$Q�FQ��g�&d	�GP�z�Z;V�jS7 Ch�|R�����h�"���n�.��	88k.�ۇ���Ƹ��i�����tWm�@ZNv��5���db,B��1��INH_�a5���k^r;���l�!@���Eꨄ������-/;K�o"[oG�\U�"����Wj;/�sr���ع>7��s�����P�h2��uU��ez�l��Pj�/��->��ZE�-?C�~�U��E�������������hY:\������]�����z`C	�����L��Y�᭨葁A�	�E��6�Y�N$Q,v\����$(��C�Y���H3(��v>�2y�<,�a������^���p��3���u^��1��Ҏ��Σk��:u� �v;��H3�FW#N�4P�Bk�3���UDo�}匐J��!��f��˪��ň�.�DkR�G�a�����
�]�uܞ��_.��<�d��L�I�Iyr����h�"�E�[�*��x�oAZ􋂾W	7I 9I8rD"�ߙ<N�S�&�U�B����-VJ]>_G��s��B��.`���R!�G�-��M��	���� �:�nґ�� ޥ��#��)�zAW��/�}�5����tX�� �ⱼMnU@�Ѧ&Օ ��J��6���KR�<nx�qV�wJ�X����G�,��e�֡_��)~I~wdC��H�̈́��~����G2�ޥ�r�����O�f)��"���}��{�7�:�� �7���%(���1��wm�����:�G7T�U�Iԟ�矼�Y�<m������~�ҟ�*<�;j.CP��c���ɕ�0:ޛ�bh �H�C�҈�� 'T2��dFo-�	�����*��l��co��Z�¤m���T�y"���>o�r�9D��u�RA�,Ɵ�ۂڥ�hL )6s��3/Y���>T���3��єD^���aS�Ft��Ng��T�����vVُ��Z�N��#-��@M*��T�%�%!�E���i�7�CoXy~}$$����M�O��U\s�֠w���[���-	I���G�Q�6�g���$l�AL� �[�tp��G���!�*f��3��5˱t"8�r����H"���P�&HV�;�d?�m3hb_����)����8� S�Y�a,�؀�5�|�0������5"��o�ZmIxB�[�l���b	������=b�ܓ�0W��q��pWqW�c�b���ٵKՄ�{���-;؆�^&�������՟�3���3�cS����X�NW
ۊMH�ۭ͖�*5�j@��Ȇ5��,=�� J?-V�b�i˟���E@��*�*�t;=�VƟF��Ͱ�K��"&gx�r|M��&Ђ9m4\K܎T(��h�\~�ܯ>|���ނ	�5�5���fy)x0��a5Ϊ�Vnq��]�E�)��}�ѠwB<��A@{�l{�R	O����1͡VPʀ�Pr��2�+A5�r�q�E��q��������G,�^T����J-����/�,E9|��: �z@j�<l{L��IkzE��u����<���=l��I�K�
N������^��g�'�
���e�>�m�xF>w�T)�j��]�;� �$��1�4܌[�~��}�Z�=꘥��Z��cl�i�{z�[Ħ�����3G�[G��K��b=���;��r�O�W��L�h�,���M�&�I��Z���"��iZ�ӧz�^^�E�K��k��`�amQ�w��D�zwx>����:yU�[PKu ���x!C��mC'�Qb����I�1GC���Q�����kUV�B�)� ����w��)T|��HMȴ��Q�˞D8�H%��0ߠ��;�|\�::�8���u[DN��uc((�qz~0w�5�:���D�d�ֲ��B�-���v�[�r�"��Y��"S��{�mW���iM������zm�����>-Q��zͿϛ��1�e�p��n�f�$��ͫ���e
�ڊ!��K{���jX?ǕņF��WN�.�D����-O�J���#��G�*|�b���<�Q�˙��7�kq���~_� HG�Ba�O�Mnd�*l�^�Q��j��m~�����]Fnan��+��P������+���_�����z(^�,Q�]
p�q��f�x��Ӏ�
�L}���
��`)�'�t��G	q��w�o�i����F�/�d�e�d�����c�T���)����\O�ꌓ�u,Tɕ aS�����vWrC��E��\M^��	u&Q�n�,;�7\)����<�O�N.�k����P񁋤�;� ׿�#A��擮LUЁ׆j���d���k���tZ�qP��W����<�a��a��Y�8�m�$�sH�B��WY���[�������u>��jN�����+nZ�ȍ�6?O�7MW�4�<咱^�$?�}��y6�@vB�L���lZ��`
�1'X�(-���_@�[���������yV��!�=XRvzY^-�{�Sa*`�g�sk��D#$iq0^F�a�q ��I� ���h�i¾n0���/
�J���V���=r�E�{Si�ɲ�ն��D�ԡ�\(-�8��TiԂ7v�o44S�Oh��~�#;�'�h�4"!M���| !&"�۳��|���/�G1ө	��4���ym�R4��R��S#02D-�U�V��
,��K�DA���Gp�G��Y�\��? e���UW⃘�X]�5$��2c����p���[�-@�orU,��������B����D��;ǟ|��.�u,H�jv�U�Nw6!�1��{.�m�� �D��B��#�=�A�!&�I�A�Y<�ms�K�=ҍ-�m%U?&=Z�9�0d��m�Ã$������>����@R���.��2��a�����^�֣�s��;e=�k�n�dӓ~�M��-p'�Dn"��x���cGY�����/ӯ��D4gb3,��<��t6�]qf,������O������8q%@ͅ�"֚@o�p�X�U[h�����FM�{/���H�/�����e�
ϖ�I��!;m5�X�`2@wfh�}��
MF�H3��^��6�e�4*�/���G6�)���u�y7��w��^J���0RR���Ev���4�)Aݠ|���R|�
>P��! X;�ǒ"�jN�Z�zLy}�BM��l/8������S��&w7Oke�R�<y�+��G<&��߽E��u���AM�qrg��(k�&���.H
2�%�q�;�@���٭ݲs.O��B�Z�O��gsi�ȂΥ����g$��q��+�C�\*FO*sz�ϲmw���k�������]_�5�q�v��U6�F��2�*���<^��Njw����p��4 ����F��jj�X�"���!�5���˕���̈i��)�s'@ۀĕ�~ �����4���������T��L��G�U4�|�A2�_���8�Z�.+3O�F��e��u����hR��^��y��zlP� �9�xiwZ:Ԋh�&����c�����=[W���n�hI�[}m��O�D�T���F`3�T� ���������x8u%�Fd�Ғ�,�`��Ė[��7PV��?��S�����I����t�J��_ꚃ�#F�T[*���
{�ShW�ꎹ�3G.���|���/�����i�MDmҗ!�Bx�aW�mhJ���:��p�J��ilѲ�<@(^;2��)I�`����6A��2�&	�[�C�G� ����&O��$�˻��G]7����:}�"Z�v}����":���y0��\/ָ�����q��<pPwQUa�&���/*	�Ř���J
fTBպ��t�&l1�/߯�'䞳,\���v"�L���jݪ����q,('�i�Y.��xbK�1p|�J�����H��T�����vx	x�j kU��m�{E?�I�%~��#gU{���k�2����m���J=����%]�>�N�W��J�{b`>�ZE'׊��<b�GN.'��n�"���o�,�M5�&��^π��M��\�^�q�V�
]�����n�I�|
">	VQ;��J��y���d X��A�k�D��N-`k���9�J�F��^�,ZG$���^+�eo�gmٗ
JՌ�|�9QB9H˒*��bح�١�LR��d��v͔�m����d�8��E��� �Od���Z���c�iϸ�ᅮ�u�ӂ�&a:����\-�a�0� x��]t!_�}Pg�:���Qvg����8��ßv�h9Ɖц����H?�fi�x��X#���������E4��a'vYʠ�!Auk�0�}���ϸ��1{f���2�=�칄\nĔ+�Ae��ZQ͋$]z�����E������ʔ�h��}��|�
t�g`c�`݋E"3��I1z����9���v��@X�H���,I��A��V��/��X*X������X}�L/j*F��x-��t�8y�>��=u�q����`���ː�n��E����U왁23��I[�*b��2��.J�q������.�@�$�l�J�=�?o`�7����"	�������qߥP8HTٶg����h0�t�x0��\���p������,M��������mJ}��I|X�m;�L+6�Ҩ��ə��F1W��d8�u�Ik��R<-l��Q-�z��� �1-����hh�7����Տ�bS�:y]��_g���#������J�io��V�T܆w����Z��fpz����"��4��	��sH:��?�lX&�ՕqT��ss����vqb�P
�z�_��hiZK5!p]���.g[��!�1S����y�Iq4˗���DF~��'a80�|�!����)I*w/�[��9w�/�șR޼K��i+�=� 0L|Ei��v���(�9e�s����܊+��t�$<"�Yyh���Ko��P�8S���1i��r� �,Dmc*[����r�9���"ͺ�h?�H���F��������oV�����"mw#dsE[E�A�S��P�wIl�*˒��)"�O���U�$��+V/�JC�Y/lO�b1\Ό���L	�����o�4M28�8���I*Y���֦x�
`�4a<�4Y��3�;\R\jW������Y_G�h�x�� ���`t.�BFmH�규U�_�_����C�h��<%
%�!���'�ڛے$+vHS<���^K � ��f��㖣!���'D��n�vxtl*��nx1��'c��xV	�C3�r�%��ro��:v}���� Q���ػqڠX����gz��Z��G��z[�kqDU� �	[�KqK��K�B8�^HG�F< c�V�n�:s��)�H��XE~k��1��<:O�׸2H5�+wӖ����	rVK�P	���[�����՛i.#Q�,�~���Ӎ�-�^sy��Jd!02���g�����m��x���@C���0H�;�o�?������yp�
�3X�_���ca��7��c�i,Æ8�}�8�oϞ�M@�"�B��a �<Z��H8q����B�
p}�Nv�2l���j�StD^w⮬s���O:�2��o,p��&��3#g9�Ƹ���F�<%�Ez0�zN�6�U����7�M�C�W�B8� GM��nyTlL��e刋)Q@��{�ݩ�쾊e��Vj���0�� ���1N�]� c.t�1��_E��ĳn�PG�j�l-{9�A�DS�NJCܺ�=�ȟ��� �}lK?�;~f�?�ή�6��K�����*-�QV�X�;F��a��6�K�hĦ>lh^	Rr�ש��5��B����Ue�=�y�00ua��U�ճ�C�̚=�fG�~�u�ͣ�m� ǀm��"�����iȚw *�H�`.	<�2�l����i�c�R%x���7�\l�?R��l,r̕L�CpN��0,�C0D&�a�eq��{��<:�؀j�}�a��9�;�+��i�ZC��aPfL���ʫ(�%��1X�׭5��}�s���͢(�e{�S��U��"�ΜcB��Z���(��m�ͩM�r������q�QZ.����ɒTB�]M�e�NG/c�_T�߳���DU<gd��Z/8_!����{iο͝�Y�8{{��NوJ�Z䯽����h_]U�K�ĉ�c�x�V�*oyTxl���*��~߇�u��������r�N:P�NaJ\E!��P���MSC��1������"l�ߙ� ���Ǥg����3N~�}"N��I�R����7��w���Ż���Xss��!J^x��\G�.�\hs\fB:{�A�e̪�xwzJ�oM�Z{H���R*����r���Z�݀���(���Ev�)����uX����m�NX��`$���=y���m�{+b7F�H,�cH"ä*$-/�G7?Bf>=� בo���Ip`+������W9�~uA�4��Z��:#$"�����2V��8`j�)h���7ZLr(�H��rQiL�k98]Bu�1�k����į��m���J�U�mU��ؾ���j(`ɏ�4����2��t;�������VNV-B�2@����z���X�@�|q��̐+O�W5o�Y8}��B-�;�c�����e���-�M���쐚xl�"G�W���-�Z:�8�қu,��*"	=�n}M��:��q�]}me�H�����º���0���БԖє"�-��WU�v�ٖ����`d�(*����q�	�KƖͶc�6�i����E'�c�Y��P<앝ϮE�����t7l{J(<�\�������[�%��8�h�����/��d	N2���cN�$p�����쁶�9�8Ś�t�����A��V?�(�@fP`�;����&���FH"�O���n;
�͞��M}��+�{G_|�Ws�}~�H���1̰,p�.�.3*�
*Q���$��Ru�8̱r�*g�S�H$��m
:xk�8��9K�~fE���V�̝A�Q��R�.����@o�6��8;����Z�3�<�-�zV�?���)[�b�s��e7�ڰ5�TlC�ߣ%p�s܌�޺�{�i���L�c�D�<�	W\�=g�QP�^�&W��źJ�\�(�px=�,��v%�U�-�����a�K1D��J��M���Z�y�$M2�l]�E�[GIh���D���ݰ�1�>ߥ	��3��̰sJl���}���Ϣ��N�$�Q�A��_��Y�zHc�~+b�C�8�1᪊�بE1)ʦ]z*1��Ce��QN_�K?!F��ǨBK�� ��gʿ����!:����-���A� 'zCƱ>`��_Txw�oǞV��E���~}%�֥�mE�}$�7���j���Kk��g�p����>̯����4{Ǳ��^��S��L�b/ق�(,����b�W���x8���Z����HC�m�~�H[Ί�;����gL��w�^��
ׂmn��H_���lW�%����.('m.� =�_E�|4Rgȹ��R9��Ezӎ4��	-�vI	�N�p��Y4��qK���--����X���?�]�u�$��e�fX�E�YJl���B�5�wpjZ����%;�i�ꩃ%6~6��B�t/4W�LN�@�������/}���P]m���#3n��g���Vy����On�7�c� ׮ǋ�ƫ8��F`&.�s�Y\�B�j6�W�;�S&��l:b۶my��_:��,~;��$����{�it�Q��UV���wR����u����O��y�G�����g��^��s���/�C]��5T��i bE㒀;��`x�m�^���iv$I\��W	g�|���-��.8�-�J��9?_p�FTpw&[ޯ�b�����h�f��c�G���.���*� �����N�F
����M���e ����B�lZC�%_9*z�o�(�b��+���Q*�q�֯���o�5Ȑ_&>Iq�:��%��0���T�i�x���D��e��Ozh(���m�d�GN�W���	����jWu��A��e�������  dH<mA�����Tg����5�0�0���O|ԨH��P�5����K�?�H��\��������;���U*����!xRR�K�]�5)k*��Lh���d���`,=�6J, �L�U�����z�G[ٿ��VW7��ik��E��>0�����q7���n�"@�|�{����T%%l���4'�X~�lئ��f;��
��J,�	q��l��V�(�P�:����|׸��NP�t)��T�n�4K}�r����=��b��.~�嫘p��絆�x�A�q���n�ւ�u���X�s�5��I�ϋy�V�U/�( K$�Xxn|(�p� �v\�Y[�V��p��n�6�b��f7P�������X��t�/:шA�'[>�)O��{p��?�W���I�0����'�G?q�A�*[B�)/���=Y�R��U~Rz|����@Ѕe7��;� ������.RX>�RoX
]�����:���&�R�'ԡN%�M��W��ki�D���ȟ5Ւ�\�(����<���H��*`gB2����e���Ln	�������D���0�_'u�n������i�@4�6\[�~bpÎ0[at��$�؇�x�/%wR#��������%t�?^����@l�_��^��)o �Y.��y��ʊ{>����~`�a��;T�:�='Z�~-Wм�t���*�>�>:�;������.\�W;_�M��&��s^�� ���O��I��,ӱ��0Z��7��c�$y�����'��q��A\�aXcK�.I���Ӻ��Dq8֟7!)�,����B��bWb����j
�0'���E꾏l'�(�GT}��킭�C��^��6����*��L��Y%����/�Xe��ֈ9�x�:
�yvw����k��#3~#-�֮���RP���6��}���� {����E�)hµJ�p^Ȏ�)/�����)'ʙ`e���5�f�p'��d��h\n�9��Ľ�: ��١��"��y�Zjb7�u��T���� ]U�+�T�*M %rF�s�Gge60}+qA
9�}�^��{dΈ�iԣd����W�M�>�w�Z1���_�}�\6ž��ʻ2�z,0�� Bc4'���]t:$Od���V��_�W�6A���g�)╿p,J�/`��k�x�<���j=�	����.�xM��)�r��V��c��S�s��V8gn4�o�KϮ���jd�[�	���ːp����Ft
e�el�����S�DV`�ՠ��3Y� ?���
��'�*��4c�~C���6Z�� %h��X�x?�1M�'�nƜ
h��GԌ�Q�Cvv"��0��6dK�B95g�H��5SC�C1Ub�hZ�^�N=%�@��0�K�!�'C\������4��ӭW�+����Snl�����%I���4��C�o	���+v=)_GO	̄6̗tǖ�_�����y����t�&��K?�E^��<,.�
��kB,�)wF��98]@� a�&qx:,����1��m*'��Vr��{l���0��~-Wo�;D-"�4������ڜ��x���]q�{�+�u�y"vQn���-���M�曈��K���?��
���T	�-����fY�J�_����J\��JvՃ6�0��mP�n������>{����Y1�'�`�H�3�����(�Tg�]6f�Q�o�N�babMwݎ�.�\.q��Pȧ�w��$~�(�i�N�E,�'�B,�.�otHO���u�*���^���LP�= �D�w��Il�*�[(�A\�^���Vg���7��3��% ;(�]J|� 
\�����"aO�R�k(�Ծ�7�����z�l4^��}��]!�ISI�^�J[8�x2���O��(T��I�t�������?�;^,.� ����TW��7�D��+A�S��D|�r��28��߲X��7i��F��X�[5DD�����uS�]V͵��(M��H[���8$�X$j����G[C�ːY�T�8
��F����{����C`�k����A������HM�{$�yz���w[�5�ӻW8�(�X8LɁ����|ԡ�fr����h�pXϚ#h%�Azth����Jy��L'kC��sѐ�cٿ��}hܗ
G��nd�������ء��>8��������;d�B� ��L � k�*��+ix��?w���?֢�F���j���.T<��Z~A�����K]���	�/l»wpl��Sq��J��K��0*�@8���N_��X6]���gKJ���+qHT*ꦒA�Ywp�Ho	���eoz��x��,���A��%{
�@�����k�~���5{=�6��T�@�� ��v���\1��n�sF(&l}G�^X�C	ӣ@*���n0K�f4�H.�W�y)b��.шX��ű���#k��U�<_Qq�X!_=�"��@�_����HkK]��7��9]�[$�
O8qX����gd4�}�*ݣ�al|�>��a���3�%^+��_·���̎ouJQ��í��=l�r�����O��cڸ��mt���2/m��kjc�Z=�ǜ�3b�d�Z��kaez2~��'}��aS��:Z�.�$��e�C/mЗ�~{�=�OP'_��M���u��,��h�h2[6�����E !��ஏ���:|�F��k���Zږ��Q�3��i��'f@A8\�`��)+���z�/�R�T��Ԑ�3c�҆�����5(���H����C�Q����4앲������"�f��z(���rY���q2�|�D�cD oPa0y�H���g#�����B�Y�=���D3Ng]�fk��B�FB�PY&8�cWn2�Ii�WYv��[f[R����5���������z.hh(׮*����صp��~�Hee�V5�p_?���]���oEq���8����b'�Rš �U�p�k=��*40�txiB4�vK�1.��}!z�V5c�O�Q���d�����:�;�.����Ty�X@�v�_�8�_�!s<W�d3��b��7��\��S�Ũ�}+��ܠ�I�V.:"��e�ƫ{��Xv���>dI�s+t�[__ �מ���5�	i�I��y���>�&7�0�>uīkBښV��鄍U�X@���Za�S�Q`<��M�J���h�臘�d��B�����}��{�8O�4a*B�P�KK�n*~���O���/@�м�Q�2�z�rMF^���,$�X�i��UNG���@�T���Ň�c�Ɇ��eR�?����UTJ�H?�Q$&C@s�\��-���*�g���
��_S`{P$�ɶ�ӚQd���~X5�r�O��?@��ұN�~+z����8b���5^����)P�?B� "�1鐷���X��UՂ�1�j��&lX���2�P�f Sd�����:�?GQ��Ge2��t12u�� ��^$}�8{y$<�����Γ
��1�b�������	��n��]�Z���YK	�q�[^įmض�﹦���Vc_FЎqc�!�^��� O�=�C��֙�#���W��:����ӛ�)	T8�F><D�����;w8W��4(PnF���*̀�Ӯf �l*��S|ʋ����;�آ��z����t�@����l���C��-^��{nnF�lA�`1�O4S��+��qK��Vu�G�Z���2��$6���4�r��Rް�U����=T1z&M����Yt<9���l�_���4��[�&:`r[���_�=W�G+�ƀ���t��	��WA�&��l8m���� �j{��ǆ��FzkR�01i�:�h�*�TP"8�n�(��#�Wjl͸���9�sd�tB���4h����w��_�o�d:Y�!��A��f۵�eB[wZ*1�g-"<�,|[i~V�:˪�hz�����[|T�ֺ@x�7{��2��ĕ�D�H��h;��z��%�Qg�^E�7H�"���.�[&v�"�����"'ȏ	b���ž����{���9�<�Ѱ�<�)U���c��`�L�C���g��1L��"x�-)�15���N̅�uɨ��[�E+�F�ĝ�U�������đ�w~w��W��z˟Vd�j;�BI�S�IEwP�EP�ۑ�V������L�.���x�W~�v���� �+�8��R̓��n"A��	Y�+ (�/wV0��s�Wb�ͬ����"��pN*������YݘIl,>#�)b>��K����*�S�KXo����� ����TlKM����C&
��:f��3W���K^*+��&��K|D�	^�kڌfg`�K��I� ���O��D�����~�^|(H۫��
xQԒ`Uy���#̓еEw'nM�k��#Z'�DroY�[+vρ=hW߆3L"�0��|��[X w��cX:O}��첽��>5�o3+�(����Q��
ñ�<^�r n�	S���&��j��,�b�4V�����s�8#�\����-���-Y��]O�^\�튌�!x�4�G���3���`HLD�{�ŝ�H-�<�V~&N��=��)�5B0�ҟ�����݌v���JH�T��s�Q�Q����HN��Oa�8H:JWmϿ��b#����1sr���[��������̕ކ���1f���'*�C��@ot���^Tm�G�8�G�"�a�-��;�>��H&o#F@���K��c9��}e��%v�JHg�̼7j��sȽb�"��2�xS	s�V�@K��8�����
x �U��c	G?�2Qb�������i0<�GH��~�E�í�G�����������[q�cҼxG=��_�0&3�=��6r�Fާ w�
�$��E��۲��V����q�X���I�#+U`v�V��`x\O�γ�_����?�kZx��y�f�� D����,�7f=��Jk�nD�r�/��`�FA`���ج�����o+��wTn���o}��)򍮽EkQ�c���
;oo�r"�����L<8+�7͡��E�#BY"ُrD6������ɨq��"w��2E�SZ��22�;�N{n|Zx���~S����Y�)��N�H����]]o1kG�XG��8��Μ��:r�n� �|E�f��g�C��mV1��'��:�p1�2���hָW��o��F%��K��<�w��AI�?�α�\{�ס��߹H�ϱ��2�β�ӽ���	��I�5r�Ҁ��߆/iR]��,�YFr�����D,�y�~Eh��
��ԇ�碘]DN=�'m�eGj���%61�e��܄a���Lv�&֘�%���X=�C�5y"o������Qz�L�<7�|���t��j���l�7�J� ֤�:��x���O�R�t��|$�
��H�=:�"I؆���|��B��ȣ�jn���eZ�Eќ׹Rusu�f����d��&Ь���@�7��`�. Z.�����Atx8Q1��/&��w����2�:_����<^��&Əib�
���I$給�=ʎ�(q���}?=;��p�+�5I�{&s�?(��<��g�,PZڗmv1��^���!M�8��������������$q163��岾�����/�����ǃ.a�03������ӓ4F�Rv%V8
0�/���H�	���.�`��<�i�2�Pa�$���lB|a��j)o�?���2-�I��\,B'��WoI�捿�s�����������hHӄ~�[Ρ6O��ӽxgUm�)7�ӗ��oL�]��H�B��xj�O˿y�[1��q�H"�;0���{�y���uC�Xَ;�-AM�xZ��|]�A�Gz_s�Ԅz0g��2I#qeِ!���\SJ���0'R��O�anO��԰�����	��Ǒ�'`W4�G���_Td�Ȳ�&H�9z`˧�����ʁ5o_'�J�|�s�s,�R2��o����< 딉/ d�~;�����!�u��R}R�0�9+H�	m&C������4w�Ú{"1g�u=)�P��m����7�(�����.�6$��$�a�+��$�2������V����^Kf�Zmx� ���9�ս�Jɩ��.V|N�:�%=�pq�e�d�� ��G��9(J@dN� �|E��O������UD�<�!�������o��V����f�I�U�,�" ��R슴�M��?H u��Z��#�V*�gd����y0�v�����
<I�a�S�R�����
>s^�����H�?��O{י74D��l�U<��[�ƝܛQd�╶*�p H8<�t�*�ܰK���-�X�	E�íE�@�c�oz�ᣢ�����'��!�o?u�˵"�9�鴫쐔��W�F�Ξ��3u����.��V��4.ȟ��	��8��[����H&�R5�1V,x�gK�VlUH��C\㧵�6�2e���.��s�hܱ�w�%�.��I�i��F�)�i�e7�z�ƛ�>f�_�ExDl�-�UEC7��`Mx		�z��'�mDJ����6�ke�F�]�o��.ە�%��W&B���G�qcZ�f��C(Cl����Jl���s�Gc��\�=�ϯ5
�D�0-G$Ss���Wj�DGu
3�V�#�3�!��{7�g�QQ���i���0=2�)���9l*��X�Q^e���!L��8
�s�v<�axTί�ۻy>;D ���]I���|3 �G|u)�/�#�������L��$��@.�Ig�;��y\f����2���@�Q�@7ڈw���/���=��LEY�?%�VF:�4�cLs�%)��X�@̩R1i����p�{�Be�k<~y�9RQ!g���U?Z�ʲ����jed��q\Sz��G@��"~J0@D=�sD_V��A�rmǝ�����k�����Y�A�k�6�xK�\�PL��
c�ŋ	=�ւ[�����@ �b�?1�B�h��w7�����j�Z�xQ�bC��63 ΢|kw���:�E�AR��3w�ե%��bLDg=��*�����=d�
�GiZ��B� ۅӏ$�F:�,��S8�����L���Q�=!#W{���)Qq�_��0���qw���/!BYN��J��.*YT�����8��p����Q��'��[��D.ִ�\�7�B�m}�<�s��2�dS���uH�}��q��g0ɦ�����9�[('e��@'�U�[3u�3K	k�f7&���N]ŷ�m���9�'�t�W��I�Xҹ�e;M��5��t�P������U�S,N*�,����a��$h�����8XV���?����v�e0����"��$���]���LLꃟ����"p�G\��ڨ�-�F���Z�S��B]�@S�+��
I�y+�YLD�#^k�dc!+m������N.R�N���p�[����ܕ.D�|m�S��@�
��SN�Z@��Z�+*�Ƣ�]z(]Gx1�
ec��29�Z�Ѣ��vI �Q��rV�!om���6\���*�g0���_[���0������pdD�X�WV�% ����ٗ�R�4wӵ�������mo�� :�V�����k�?�������y�б��0ݢ��#<����]ib���r:@�"�Y���>������_��p�o��zg�����+��4~��tx�	S�rCr}a�ӹS�f��O|�<"�X<��<��)#�'�KX��f����;WE�i��͆K)�#k|}u��E��G�;|x�l��6���k_4�a�S��o4�J��QW{1;�썔82NfCZ��ր�N��\��/�U��j�s$��v�tֿ7c5�Yz�x�s�8^lCT�5v�9#'[���.F���I}���Y3��<��Z`V� f3��b����
��H���c��ri.`�}��>u�Z�l�N�(=���T�~U�A8J_mGY����/��eFYZJB��-Y��q�"{�U�H�őoL)�?��/�d�]�q2���r~\��P�x�	�	V�O�����)�$��S�o�l�@���8���,��T������r����G��?�k�=�QaM�V\��5����ё���e)t����2F�k#��E�G���)�����@"櫌�s����r�T�\��e:q<��`��&@����zph�
�J��T�1�]el��}j����F~�#eR�Lm���{��(��+��E68��Jfq�[�]2s�)3�fʕL�Y3�xvt�k���%�`��#7��BMZ}gK
ş�Կ׬���C��NI1�ubuOhDH-�(�:��b�<�gzߔ��Zby����8M��_ ��[p0� ����7��uB�"�)���s��+*�e�����2(;� ��w51FO���`F���u�"��e<t5����ֹ苢����}��8��SUU)��̵N)�Q��knץ�}���]�f�R��Ԝ�����김�<u�.֙�����=_^��0ԥ��o��6�W&�IRp2��b��!��޳w6�����
w3����������,�^�O��,���vɺ3wf&�ձ�<�V�[{6%OK�cF����v���m�Yu�_R&p�w�,�DW�4��#b�S,y��ђ�q�h�+��|$p,63 E��T0�:��J?�}�:t���4ø�����?�Y����g�@�pz�:إ�Ɏ�
+e�/�� I��A�s�F�V(�&;����>��	"eѯ7(�����2a�M.�փ�.6:��QJ���:���.�6)Zyd
�j������)��&"C$��u(��ԩ[�����M�E��;(�����=_���%1���}�G
��wԤ~A�l� �gc�[rV��<���{Sa�M^_�B�0��?�C�7�z )X�.�.Ժc;<�f��g�X6�uf���.Y�!� ,�3���`ǇxİW��[��)A1~�kl��9ޟ����![6듙4Dӎ�hB����3��3CL=�������:����Y���h��I	�J�?$$Ŧ,Z�H��]x�#$|<�v6旧 eR����QHϨ���XJ�qC� ��y��d
h-���L.�Gg�|�k��Wx!s�:�ݭ	�tN<����p�*������P>�vj	�2m�<�Qf�ک�W@�g��A�� s� |Tb�H�J�NZo<��� ��P��4-�|�/�W(���f��Ӽj̧= 6�����0�_D��kǵ����{��h�U�!�޽��:���6�{8�_�X��=&\�i��u�*��#���1cAc(ڹq�5����h�	�ޞ�}
�a���1{��O���Ֆ|���'1G��2.t̋7BG��s���}((<�H��
p����\x��P�љ� ��Ŝ�����o��!��i����j��iî[%�2Ew/�����\f(��
M���֛5 ��2���N'���6�N9�[:���
U�X~X���L��?}x�E2a�WbB��pZ�Tj����C�$����Y�~[W�#£��#�&t�����[�B�w\�#�U;E�ui�Ň�|��X0��?�%�_�P|%a����0�e>��9'�ܑ�W����ff�,�w.�
g �u���ƙ��W��5�+��
8��dZ�O�^�ԷΉ=�>�@�4r�c��Q�b5n�H1(��̫�r<�;ZoO/?'��0ǡ��R��pM�dф��iX+�b�itc���f��52���P��G'�M�v���ܝ��q�>8W � ��#�\ |x�����4qRK��
K�L������׫�����m@����D_��sV��U\��EF��ف����:d��O	��l�:�o�F�L2�#���|Ì<�zKr1g�]�:�B�Gu��|�u�����`��܊x��cڋbo�.}���k�F���e��:C��9J�?��d��IبE5�v�����Ct�2��At�7�l;ʍ���B-�r1��y�C�8Tj�¾�H�$+��5�2(�^��a��p%Rj����}�-�7�bb�P��'b٨�,�0���g��#��Z0����S-	
��(`Ч��%l�����F7��]����Dr
���'����E>�q̣�b{Q�}DGA5��VF��qf�#Д�
�?�l���(��+"������?���y���=Ĳ?�*���D�2@YV�Ö_q/2������zk�ˇn��˛�7]�0�}:�ua�ާyj���֯���Oە��w$ ��z�d.U��p�;�3�:6�|�����K^#V�뫟��{;��^�۪X���{�^x~I�g�A�[�:&檱�훽���� �q�"�o�.U��~���a�A�c� Z��R��^R/�����,����ǞN[�e�K�U�k�(�%�����#�q
4�*�;j��{�4N��]_<������Ϝ+9��)�3�"~���׺��$�U������5b2�c~:ӟω�R��ľ�C��hK�B ��:�����Q2�^� X8܇�g8)����<Ko�%���6~\�Xq�9)�J/Ŗ�$Uv�`���Bɛ�ED�ᱜ�&}?g¢�������;!��%�U�Puט�Z(�z,`�B�C�l��`	�������Nz�"�[&�
>�]n�
>
F;�Ӽ��g��.�LbuH0(�[G��˖��c{�$˛Y����ÿ-t!31w��wI�l�OL���AD��nm�8��|>c�EB�� �04�b*g����3DAO�d����1��ʉ�?($SN����ܛ�G,�U�?T��3��FV�U i+�7�Ʌ�+�����r��{Q��T�N!��G�������zܣ�����h�ɥ�<���!7E�B�����o|l��u�C���MQ��X��'�����pX�3�޲W?A��⺬1������範?�p�.*����}8���5��$z���^9[N��(EIy�}������'Q�f���q�kZ�ǒ�[����G#d�Y�x�o3�, Ǿb�'5k����OX~Q͉3<�������_9�bd�Y��	*����\�����l�}��C�Wl����^�4g x�g��/�Ϲ��)ڭi"e�s�)�S�#�k����s�.�u�é�-zz��x�����N�{�ph��f�~W�LJC:���4tNb!��
�N�	��\�Y�X�7����|��F� ��`�`��W�mx�rL�</����	�3���[��k�T��ӊ�����i��%����58)�s�w�(N�+ �\!T횛)9�ҮO��Z��,^�%ڐ����6<����o8�m����<��o�.���i����kY�Z������{~u��YG&ԯ'7_>�3/>>8u�J�%���"N�'��k�L  �w1 w�r��ʡ+�m�L��ۼ�.��![I囘x7C���U�W��e�P%Î��A�8�	&���k�d�Sfu<S��-�0a��ќ�y���8hI
����΋���T��/X��^��ҸB�X�Օ�X]�UG�����"��-���<S�Ѳnks�fo3?l���3jg� %��;%�)��g���E�e~�˙樮�����Mp�q�EWǴf�����7�f+9ط=�L�aLnK:��6|��u&i�xg�%��-z�F��|9^2�N�`Ge&
Z'C��ѹ{q����&}�Myn��~pj,M+@�4�˥���A
`O�&��%䰚�E��,{��&u}���;?w𲿥�?c|�g@�Y++��zO�*�,����Ϳ91�o���?��p�s5^����F�I�x�F���5����){�9'[���;%o�	!y�Kh�T�x;���8���u�kU]_�Es��R`��>C:���7>	V�M�.mW�%�4���|�@"�s�&�Js_GV��� `:cB\k���d���۪����ʂ�NyɲᡎAv�#wWN���(��li٭���N�Ub&
\��z���҈�ǰ�;I�� ��۫�ӫ7.[�������<�.�����3-J���5܇]�'�����j��X�	��dS4@�J΋[�B�t�xLjmE,�}�E���<?���+�?	ja�l��o��sd?<���hBQ�.3ٯzE��'!j�`��
��˴��e*XD�9�+�&�r�����}b�u��*���t��7�Ki��'����>v�LGx�$���N�f�W:�|�x�D�Ռ�1����1UL ]��n��Ls#�Y��T����A�.�T����6� ���a�jmPRg����P�K��V�4a�Y�"k�bw[�G�EY�&46�4�.Ji9�7������p͑ڤp�)�.�#�� a �A�"�Fk<�5�Ջ��_�-�o��/�/\Mo���������e���)��Aߑ���F�,͗wT|�S��č��^ =�G(�u�HL�+��Xl�&30��'5�f:�A�=�G_I�\������+�,3ez�#KW|��a���h��klܙ8�JH��\�k����t/�� G�>Q���XA����J�.��2IRL0��,���5SD1�� rܛ���vQ���Dc^���ܺ��)��ri��%�C�C�h�k�z!X2�b�FC�l�C��D��CU����0u[#Ӱ�����iDtÔ��l���D�ڊ/�"�"	L��D^���#ӏD�c�.mChխy�����k8���n���d�șf�b�!�n��')cP�!�]����E���Y�HuZ
3�Dpy�&�Ou�A�5s�����HV���8�8���T�8�LN9�o�O^�яڒ$��EXD\0=Q`���\y�	1�����1W��Um0DEH��V�T���%	���]�ᔧ�o�>̷aZ)�hH�A8X�#��/�5��$QdN>
�I��x=��Sy,JC;��c��]���N�P�-lҪ�5��8/���k �ͭ�&�Κk�F1l��(�Y�/o��K��v�C��Ū��6n_�Ѿl��lB4���o��S������|J�>��G7O�Q�!B�\��M_Y��l邫�(;���a��F*��YywL�����g�2�s�^�3�Ɔ�ovse�r�1�s|7�f<x	�&ࡰ��;G�\ w� v��L�k��3	�:����ڞ������RsJ<��6�D6���7��s�B��:o8�$j2l�sp�ӽ�)X��Q�������GW�\&@{��^{���v��]�Q�	�N/�e�2��ٳM��T��geDm�"P��V��tI�v����.
zB�G�3��-����)ҡ�7��������Z��$�R��#�������<�,��r�k9 
����.�O��BD4!/a~�8zC�H9����8"X&�%E��@��l� %M����*}:��q��	3�5�F�p�	�-�X��ǽ��_m��a���gP��P/z�<���=vF��d�s�3h����7�fCw���~P(�1|sr���ر�O���'���s�����%�!�+����r����i"Zۥ�ؐc�f/�I�`�ŕ9,�z�a�JW���ZK�<���Z�9j%���	���_��u�KN z�J�7�f�#n嶤�qs���~�TQ�v��.�F��:	�0�0N.<�[�e(��3��S��\���s���}�`eSI��``�,��<I�G�xɸ����Ũ��&�4����f&5��,9�F���#����Ii�^����T�,�]4�+�9�f#�r��;�#�i*����5̩q��P)Q^�?�wc��#�h7���Rt��p�oY���b�1��W� �(Y���m��&�Z���O&�����Wq�[���DR`���v�GX�B��_���3��
�W�r)Z�7��F&�,'�tDaO{b�#��]Cs������
��Ȗ���Y*惝�J҈L��}M�R���J�}�?%���ٷ� �����*tk=�WY8
�B��+T��KF�*�t���v@}>(���~�,'���A/���(��[CP�Ҁ	>�hܖ�8~�ƌn�X��|~�д��a┇EcO�2� �xl[�C�ռ�F�;X�@5���A��'���F�v6��'+��r�����=Hک">G�eĸ`�W���2#��3��ﰠ�6U^E����g�"5X2��#��{��S� ��=��zn?#�+��Bϰ�*��}?�h.��j�ډjj$���>#Ah8 �����Wm����Z6��yA)�E�d��C��<�d�`m/�ru�"�X8u�LѣB��e#���ǳ��*��	�T���3�7�����	1~*uc.F�Th�p5�Dc�~/�}���H���`���#"�-��N��l�ʤ���i���=>��'�X�I�K�Z��(�R�7
����ՉW��o&W�a�7��@'�N1�؄������"��:ךֿ�>�|��������Pd�k��c������@���+���@��C6�UK����ON�9хڐ�m��-���{9���ȉ�aEJF�jɄ�s)eWo\EzQ��"���ї�>��'W3I�ӌ�)����^��:v�9'��l:v�*P��o�<c8#����`5&�0Y,�	1]m^��	����+�e�KQf��n�W~zB/��ϮFny�>Z��m��E�Q�E����e�x��ncJ��m'wG=�KEȄ�>׋8�慣<���GC�$7��C��7k�r�� $�i�*���lҵ���<�GH��u�V�!�<� E��8^��"�� m�}�g�L,�,z�K��Mg�؎~��E���
����ᤆX�x�����)p�v<80�H�s�ɐ���ǂ�A�u7!CO[�P��n����GW(���H�sk	f�¨����*��<��G�S��-�v�aLG��������F�B^J<�M��d�����>����S�x�jH΋tQL�ˇ����X�.Px�ǖ�$�߲��1y �Xu!B7p�O�5]�l��Y��5��.{�.Ҋ�x���u��d�BE	7<T�\w�b���]Χ�Ė��%�BJk�����S��%8��n'+5O��/���^��;���X�H;F6�$-�2O�_`��<�� ���-��)�:�A����0ؖ�}��=����Pٵ��}=2�)ĕ�}��~6�4�g�خ����x���<N���l�S�v���";��T\W��47�pF���g�:u�d�r:� 0��l�Gja钅7y�W �������7�Ɛ�����S}hg�%k��Q�!�M�t�1��i�:#���B����W�(ђ��{XE6=��W~G�t�#��/i���8!�-:O|�ˣ��6L��@��f��*�����vӳ���x��}�j�0��t�[ԅ�rs��Zn%�gd����>��L��"��1�#Y����i��DV	Y!��f�,
z�*�.����g�r�1�ۡ���ү�͎��3�l�2��p�4,	���Ve(��ed���O��'��uN�B���x�{'B%���>���Y�8\
��ٮ@/K�O���4�6J����|RNԟi����D��,�q����K4CH;�� ��On<F=LE����fm�yxeܹ��
�]�l>l��sG�If�+	�Tf~��H�%�� �x�c�@B����� ��6U<��� ���	p|%H������~ �?�����:u\�!j�����g�);n�������\�����}�"�Nz*_9��_<�����9�F�ɵ�h|����'����~<�c���,a��,��e�I���KkJu��֔�zSqC���QE�T�p�{�1��`��Y�9�DW;ޣ��;�E�&Fg(W�:[f�Wn��eM�k���vN�8��+H���ya	̀��BB5\]u�MB�/^F��R���tCyƳu���V�h�Mk�N�,}�{?��bl����|x�B|�-��b~<�C��3=������ׯV�h(�~�~dç#9�f���?#��|JE�xi�ҍ������/��+�_LwJ�A�2���jHw��,.��uz��M�����OPIVf���2�B�&�e#�������R��E#�R b�]�s%t_1�y�Ԉ���~]��pijم����3]3噴���Ʈt�B�X��B��L}�]�����K�|36�#�� wU�gN��>��'N���Mބ%rç�{B�d�U}=nH�Ԙx��x�?��GI�Gc�xGtit�b��zW<R%0yH�z��X��j�`}J$[=��|c�j�)�S�	����
_�eHE;l�o\ԍ�`.��+iϪ��6�]�ZΗ���U'������I�9/!c�N xUz�ZK��.ܒ�����J���"]@�4Y��1�xE�y�ulg�w1R�X���?'������H���E��j��TA��zB2�j��Ӱ5E�5���K�Ba�d�A���
l6o��,�Q��7�r{dc��T�AL<h�V���"�`^5���!#QTt���Ԩ�m��ϕW]�����k���q�/l�����ߏ������7��9�����8��A`�F�²��^UiS𣆞mV�Cs�ҩ6B� e�ޅ�-��Z�U�'����%�?���vUq����� ��D���g<���ZO�
�-W��8��_8D���A�j@ϗn��y������c���zY5�׍�Yb=C��࢓^��5�2�'����
׺��E"� �=q�8���H�~��'��i��:^ȝv˪w�|g�<���U��(2�_�@���b$z�0�аޞ���vy8���)_�|6D(ݧ
������^Uj�̷gI�|��!��`�(�k���C��b9��-�p��s��x�3�1�2��F��Z�4�ƞ� ���Fv���u�j5��=LZ���L� ����1劖�Q��m�}���>f@3�o�P���J����v5���&0m�O)�NT�[	*C `v6���A�ST����Z��k��u;!*����L
A���F�U!z���'��u��N��6�aS���M��C0����K��$}���f� �3�)F�~
�@3~I��Q��񫝱�I$¾u���'~@Y��!�P�RpbI<9<�&l����|�.���?��G"�d�l���&�)i��.,X��-:�MvN��"G�*0���Ф�P;%߁5�K�������jD\�{����]�N�T�e����ɗ���c��2ϛy��{@n���{yu2�D����&yѥ���@+o�pA���w]S_�֎U�
�3�[!ϥ+��2	\�3?�/�h=W��f�v6@�^�R�F�Q^.��{;���y�c�/9���0�w9ڕ�"�l>�ߏo�����hD�@hB�a�B$�w���6*P�Hm\F$d�MxB�w��]�w��������wtA���`�־5G�0�Pr���r�����$Ǟ��xɂf�_��sE���;�vg?�y�j�%(5����|lE!���H*%D�wz9m.s�Ư6�е�t���h��q���p��dd̟���q��b'�%�.�X���u��74]ӹb��d:.�[��)^��|�z�Bm�O$����6qb49W�l�G�����5�6�>��i�����V� �{H38�E��{�[lQ�Z����qi�wTژ�U���R�E�.�{�ɚH��>K��\A.0�p���Rp����KjǗ���TA�tZ�*3��|�f'�Ovc��#�[N�N(u�jfp�Zl)����v��/Q���塠I\���\{��}���eCX�`u�d���m�b�r���T?������T�PO��g@z�v�U�v��'��)�]�'9���ڞ��u���/��^7��N�6�|>�9�;K�������Z��.F �-�Χ��6�*=�B����d:/�>���5��������+tV��~o艆�C&�d�[�yA�|#����bJI�����J���)%{��勘_պ$�@Epn�^��m�r<jb�)XP
Fɔ�^��m���_̠go�k)���y
W	�A��(ꚼ���~ R��R+��.�t�S��S[4���p��(}�ĳn7�1Nɺ�ir�:أ=;��MBG��Z��-����?�G4}��Nǋ�0��������4��xU���~���|/��Nm�����`�*�3AZ�ic�,}&������\MT��AK�ͭ��6�5ѕ��~K��X��@��r�+��R�"p��r�h��L{[;��
�8N9΁"���>3�������*z�ok�y֏Uƞ��q��3X����*���Ȥ���^��i&�4^6�m�\�0Lן.�u���Cj0���dn��E\�z�X��L&azDI���
	!r�V�A%���Ԁ6_ �Vh������'K�?E��k�}z��(֓Q����u��g��ۂD�-��?�4�TN[�!_���y��X�&�O���oR+c�#���U�%�;�����\�>�=�N�yE�[���*�������+	V��)�q��{�Z,d�X+oR<|�i椣�Ρ�4/��l����w�c=R~��	�%O B��aA��#�7.�Z�n_`ǜ��ш����-�w}���Ap�6�?�J �M�	a�Dc��We)������Z�;׌�l�fU�%/4G�����t$��>7\�Bˠ45�垦��={�?�e�T������i0&h��?��g��͇j�{��:�N#(I��G��o����Z�׺��h✯��MQ�I���Ջ����~�;F��y��_ͺ�P��U�Z����5�ˢ��/e��MU�X�����7����; �!��`U�5	e����hϘ#���7a���
c�"M��?��h*{�&��(X�u�>�����j�J#��t!��U� Vm�*yH�$�k�*;�l,t�ۅ����ܫ�H��i��;S5�>(h�����&o��AۘX�6��H�n�h�M�H��������?1����ɜ: (m�y�}H����_��^N(U���s�����_쭆V��Qd�T�����U��L`3`���3μ.y�<��x���}�͉^�0G�����
�C{E�ԎB�2W&�}����Σ�KNL�R26������ל<��= TF~����Yk!����_��HƵK�%�vYH�o�O0 �^�m��w��*�g3��)���M�I�M�"�? g�zjxmadk(��*�36�{d�9�Lt�Zm
�3�❨���ᵂ�@A��΢=�TN��x98f�&t��u��	2�$g)YR-�k���Z�̂P�B�f��
Ñp������kZP�b8����.6K+��8���)$s	���Lo�:q�Wӣ4��k28�����
F6�#e�
�C�7���Q��E�g�qr��[��m���͞L8G��v�(�s#E1@��s��҄���ג�}�����Z�7]y�'����7MIA�E�p�a���Q֑��VQwS����Y�g�% Ϣ��D)c�n-)�����{rV�� T	����S�M�������L�A8��Al�O1�0C�r!>�h��Z���O��]���I��`0a����m]Z9�S��&�X�Z��+� �����,��3�e��tw�o ,aa�c�Q�˶�����~9��q.^0�`4/�@�p�� �!�L��ˊ^��)��eH����.�l�b�k�ޥ��f��^aog
�f�3E]iV����,cVh;��}�iy��8����=��&�`@�P���{Fu��
�bu\D�Gcl~��lJ�U*�^~/E>Q���̚���O������TƟ�B�&�'�6�ʢV� (�H{{���m}�gW`q:=�1�6w?-_����,�A���ln�w������\�I�N:�[7�&��:/�Z���������;�JS��C���SB���ȼfP���e =�VV�0M)�Ũ����cݍ��l�O~z9��z�?D�6��uA��U,4g�gD7{(Uރ&����H���^%���#�K�Y6�B[:��2Vv����/t�����l�V�ܷ�V�W��Q�ā����[��DAPw�5(��&�hF�ե����B�-��SI��� �����R�]rN�P��ky�?�uݳ{�_�$*�C!�!q2�7������a��S�����^?��zvo�'F~l��h�٥�P��E�^�����1��`y=U�:?ڃ�]��r*/-h��J�nR���/�s"���'mO�<w�.�,���Q\M��|�	��,���q�鍲уT�f���>cBtRV����y4c���&�H�`�ai�[R�a`#c��&���k�֗��-�/q�����"^3��D�X�|{��]�C#��NF	�����n���4G�'Ie<�E(z����ϕ<�����>9"������i�0K�S5t���E?Sg���_���N����R��&�짳b� O�Y��j�\ӳv�3��-*�X���G�����׶�-"w;�6ϳ�MH:�0�݆�����C��e�d5�6Ck�/�#����Z�ۻ���&[A����O�rSì���+�Y,T�W$*��y8���5T�����鵄8�:�M
*h9 δ(� �Ti�G��~�u�v��	�Z��vN��G�L��u!f\���e|�՜�����8�>�Z�=��*�a�
�{ʎ�5���3��w9�Yt�&���v�~9
&�H3!�O�P��־�l<�Mr�S��}�َQ><6��\#f�d$O��;/cd�_1�A,.8Y?Ӡ�N3�8�?�] }S�^G��7�m��5���D�d2���t-��#Ȋ#����;�u!!ս�! �!����ŨX���)@�[� ��46��h�`l��P���`�����<��=��:���Ba\�-��HF�g{�~��-a��4o��հ�B�S��Y=wF��񳉺�x�'�/�"(*H�A�Iw׶�
��N�`�IJK�~])�9!_Ͷ��ZZ�4H�Bd����Z�4��4*3�Y���J���dחh�Y�v��"r��>K��>.1���Y������n�|����A�xx�Y=V�ȳj��L`|g!���c�j׿�Կ���'����).�M��i�l������zZ�YI��%6�R5$�I�گ�@�d
�*�θ�݃.���z/q+������YK��&�F�5?.Nt�A��/ϟp\�0k����V<�	Ƙ���}�<	����DJ@��4��=z��8#jt���6q���1fB�Bk�_0�|0�F����'��x�m�Z�b� �:(�u[.o7���ɞ@��/�]���4��H�ih-͓kRK
��gA�_U�4�{���f�����uf� �&:�
,��a����N���Rn���4Y6�댯��k���Ѥ��������֡�;��7���!h'��_�Jn,Kڧ��V��c|���s�E?���c7���)p�  |X�P��}J>\a}|I�X�y�m!���E+�N5\�@Af��R�̈́��@�c��*O�����An&�/F�����r�:	,x'�I���5NH��6U�X|�r����P�~3�R@dϹ���1��w�ܽ �+t�֖n�	`��;Г�9b[�����@y-�j#%���{�-�
6~��j���B�N9���I�d�fZWr��{G.��E�wa���k�5\O��9>�ǈ�V;�&!y��U��w/<a�=$�l���ϯ�StJF��d��n�1<�xi�y���c�ӫ��Q,s.7+��Q�P˫�[��*�"C�_X%Q�����.|�m�Q��O����$`2�_�P�6듌i��}�C]ل���&;Ƨ�^/i�����l��z� KT5��B����#��e}z�{�$� _1�r�[t�R���'~(X7���b���.9Z�}%T0Aڄ_ӃM�_3���L���^���HTu)uDT�g��V߻˅���-<z.{�F�l�o��Byd��0E�k'!�*|O����V���`�(X!���e�]۽`�Y��^ �2�V?j�����c��n��&�7����׎��-K�R������&�&�����t�����'�Tݾh���3!�����ń�!P�L����pL�hi������M��KF���U�E	N�F5v�Y?�璂��=T�u�������O��g�������H��܇���������a\{��@�DP�)sQm�OQn����75=������k"�����߅�"-vڔs���dr�HT��LIo�Jtv�����<k�G���OD��Æ�@L)�,e��lQ��U�
*����V��w�	�k���Q�Ǻ�8��w6��ʣ����ʷa��0�pJ��	�&���WZ�]�
:\�	�ί�BW�(���J����^#���$� ��Š(����qp�ȳ��3�I#/2�,�Zi�[�O,���3^��h�47	v�n���[u�3'/���]S�Sx�����R.d��6:+����ָ 4�uN�� ���*F$�L����/��:��|y`$wF�!��Eg�P?�	��n�n��.4�"�Ӓ���>�čc�t	�餫p�^1�S*�)�g�g}�Tm5�ĸ��my#厂l�]I��zj�n�+����3���I��r��E�xn�.2�L;�6�!�I�δ �Fx�?YN���|�1p��J����K�0���p�e#�����= 诉��L�S��tZ�$bxÔ���7b
ͥ�?��U�Ds�5	������U)����4o���7�ᴽ���F��,��s����Ԣ;����9�"a���^��Q)��D]xf�V�4�n-J2�39�ɝL���gMUsY���,ͥ>���+F��d�;��)O�4rv�vd�!X�=�D	PTy��.<w���:Qs޹~�ns�4����`k����|�����)m�k�rR=s��P�N���5��v�]w�[�~p�%�D��V�'���`��ćsj)����5�)
���F�b2o
ob1R_{��s=��v88��)37��:T�rb���b6�����on���s�7�V��8�F���u)�e�v�=xkt��o��� �EƑ�(]���V���Ko*����e?���^dQ.����P��@N��ށ��A��HH��v%�6�A`��{��U��nv���3v�.��ǯ=�~`��ĳȘ�b�^g�F���������o���nw"s9%�Urrb���q������_�o�ƘV�mc��4�6k��wX��Η	�׳Q}l�	�=�&����1��XӇY�j��1vu[����h�l����aoArB���1L3�ZE�.��V�'- }�� ����/��,3���پ�n�:�o��3�ᗵ0�y�����L�����ú�T#�U,�*7pQ�Ba��=�'Q��.ߕܜ��j�@)�vS���"T��~��pS�*h�B���*�������ߙ��;��d㩀+���l�.7�ݸ	�k��
�#_��$|
��N��S����/�JD�}e�ܱ���,�����_^p϶��O����L6����!)��dM�N�؀�U��q��W)I2V��r�f�[�~eK����:��8;`�G��T��K���ؿ�n���A����~��A����QPߊ݇�)�O��ki]����ez�H��w<=�W]GGA1DgB?���V�;L!w�<�}`�䈅m�¥���<Pf��8�C��$g�	䴷K�	A.]��5���J��[.]�Ú4Jl�9d��TZ�䠓&�;�C�����#E���:�S��K^��V��zQ�ls���
lEz���M���N��Ov�#)\^��!=j���H��7d�(<#$��%�Z�����K��i�X�a� �ϊG�m��l��K���
�`�gEv�Ћ���t��+ǌ�_���2ә	n�n�&N��&k=p9-����$� ������t��	����J!��Զ9��A��.3�`�x�4K��:�2_f����+a���1�=T¾y)u��9j@<���*��=m����EL.j�<��sA���������:ⓔ.��Xi'��n�m�Fa@l����(}�ˤ-��OX���h���vε%Klk��{��C�<�t[|��'�����\_����1�N�ˍ�ަ��OS��C�q[l��B�O���G�r16�g��_v�+�0zbߩ�@|#Kfnl&61׀`��PE��ҙ˚�E��,~*��j��J�&W�@��s��xD8��e�kk&�ʼ2�u�5�:�i�Z[�i����ed\�LU�T�V���Q��;o��I4u��p ��uF�{��1֋��Ŋ���p�k)��X���X �B8/���̳�����_W�R���{��Z��b�x��Bh :T؟��h fr�fC�^К}c	N��}�Q���
��pp�L�,�ħI���I�|ٺ8�v��w��-��UjH�1&��Ý*���/�L���,��#��{]:o���mcu̠���G)?�&=�M,��p��Tq!������,�.�F���Hi?���/�9��pk$��
���J_�/�[��˗���#��	���]Cc^��EX��He���C2����5=�s+o
��{��\��urz3>w|��)�!�@,+xخ���M�h�Vi�{�y���*��좻�12��H�|�B�,wq:l�X���Q��:�YB�>�=�S�Pp��Zo
���B���Δ:��,��F^P_5Ҭ�&@,���q�
/�S��2?�K���-�ߎE��n�΃��I7ZTw�"��>�{��M������t�M����z���0E��>�wnos ��GN��oWˊ�k�~vU�"vtM<"�mI�~w��d�@a�X.�"��} ��h� ��w(��nc��tΝ1p�R�G;�q������2�.�'m�r�	)6â��8B�e7U������;.�yH���x@���\�9�X�X�d�U�f�$�e��y�V5"��V]o���F7���7���C�&�q�?N�6"Vb�Q���Q���b�j� O�2��ƅ[auL女a.s�ï@�&,�4��"dES��K�\A�����'�U�M�UU̟H��H*Y�Y�4T�/(�*�������O��B41QLk�+�2�*ˉ�ˋe��A�dz:�����??W�(�F6��y����p����'7p�<��֍�֪e	m�7�5�r�l��0C�dO�&Z^��O��~����ۊr1��ؽz-�UT����&z�����ň�Мo��g��G�ktVj,4�?��V΅AU;՘��M<�֗X�~��{��'�ۿ]:ch�A���_
���E�[@�Ssɻ�qtj�d�[�%0�,��@��I�{��ôÜ֤��a䝕����}����ز�Pk�C�-'x���)� ��Ju;D w����9���C�v���Yz�p�&-�yL�T��uȟ&|ϴ�7�Sm�a�~�Nf�[�o�T����57����,���j
u-�.�����A����
���ul^�n�R�e`��+6T�6:�����"���P&T��MҘb�F􅡕�^�&�q�
�/L��E)��YB�-R[��M�V���0��v�^4J�=26b�^ ��I��8�*՛ȥ+��U����(52=�m0Y�$����(;�K�?ϩF���!'�lt�k���~���ŭ�
�B���nI�u��2�V��Օ�r�h]����6��>T���������'<�l�õ��3G.����	L+�"�2����L���[���S�s���3O9��x}�@���0IDF�B��7��_A��4�PFu&뫯_�p��8�#�Ak����]�E�\b� cmtܠ���0+R''�/�&�������WZ$��G�A����/�F^�	��K��#0�h)�G���+0_.����az��L:@�xe�LG@���Pq����9��&6�_T�K���4�K��*@��fkԈ2���nW�����TA��w-CW.�qO��'�
��FO����]�9� [^-M�DE�{��-��ƻ9�W�d�C �l�Ek'����������8�,<���l?`#Mp2�;��bZ%�[B���r�2��u.�2��AQw:h����<B�H�����u9=�[��Q8%ө�w���r��t ?}�G�ak, ��DXa]t\�r�LE�����:�w�� D����4DS�;����Y&��6V���J�a�	g�;#n>����E�@����\3'[DO݉^�n�@� �b�M0|���/L0+~���P'���\-�d7��I��\�5M����XS� �SO���Yu]�Z�ټ%��%Y�l?Mw���<�dif��_�}N�҃�`{s�4�m�ݔ9"�5	�yt�Wշ�d����M�@	��J���ޣ���.C{['�')��Վ�^��Dת�eGK�vs5�����B�7���Bƚ�ī�D�V��#��ֈ����`���%�2��e�e���H;&�;q̽�)n�Ԛ�f�m��{8?9=����Cgk��S��D�:6�Gg���/%b<���RN0�l]�Ո�V{��j�-%z��YZV� �����ï�E���s�n&9�}�ib++%��$��R�̙�M:%J�����A�O  �ޞ��cH����-=z>a.�T�$$I*�̈��}�����͔&]�knar���k�>f�T�]��7V��n��
����s�%�߬�p/Y>=�[ͽ鎻�I�3kTt`�J.�܏����Ш���W F{q+)��?��i�Bm�m��F6�iIP��Y�E�t�������4[�v���M;��<BW~��7�Y�ҴvH���y$36Y�+s�?�.pG����+��ەBA? �jxO�4�f�<�q@ ��@�E�˵�T	�Q�"��\���dI��Om�1��Sm����͍I���Whѱ՝�]Ͱ��I��e������Fk��>O����w��g"̰�C�)�(R�ſ������V���|XS��3�pJ��Y�/2r��e���RF{L��(��n��5G8Ѕ�Õx����dM����Ҁ;&�N�	����k�`��Pp�h)�s�M�����:�V=5���0Ur��dh��*'�{���1�4z^'aeF��Ç�>s̃, 〿��&���4*��k~��3�ȫ�޹�^6W��f���.��U�P�{眘/�������8�/yj,#� ��#�\iF":]bP`-g3Q�o�LSV�� 6����S��F�����t"�t����cUf�WU�S�0����"ˑ��%Q���\ͣDII���_Z��F�ZF��K�����S>o
C���&�����73^���jl���LHG!j�Hm�]����W*�ᛴ9��Y>՗e=�drJ��o�P��辄'��Q��v�
t���G&��I�Pf�b�5�W���5τ�z���Av�X���n��2��lq���VS�g�-�q��FA,��e� #���_5�$�':��dVMB<hۮ��rӗg2f��]��[#�TD��;�ʤj����:�������aE,_q�L}��b�[n5���%��;�R�
g3�H'WE�B\ki��*�t¶;F>��*�puD;C�%ς���=�c��,��ɽ��;98��s3�TQ����f�C����\�Z�A�Gc�~b�A�l�jV9\�/_��d\�����`�(c_���{�1O�wa6|o ��U�k��$���