��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�J��"4�=�7(�T�JѺ�ő��,\��s���ӣ�F�؏�ho�i�@�CL������xТv��m\$�-e�����q��0��������y�ߗJ�J�a�HB@�¢�3�-s��F˫�R�V>�M�e���-ѡZ`�>S��d�Y�sMA�e���~����)���S���祌�����Hc�����>�������ݶ>���R|,�TC�Ԍ��B@�-�G<��3P��B���(��Cf�Ht����_�yܺ�2���P�Z��\O�(l�HW<#�`rd�O��!R��؋�)y�x��}���k蝽��B&���/��	c�2�C�yW� x��GL�u5L�.:�LJ�()bX��\h�VW��}�3�ݡ"7{���7}ۍ�h_T�*;�~�ҡ�mWsZ�8�`���Ă�m;�w[m-)�b�S.����;|�]�h ����?�������r�Kf��[f���	��B�g{O��ӥ/V�  :ʐ�o�� ?��npr���:B�u��r��՜ߺ_ׅ�>~�27nE�k�e�ܚ�&h�8ǈf;�Z�I�7��pK�l����,V�>~��1��Vަi�)"��(#Z�,��-^vѯ�����.�����gy�0c�t��=h��S�0�9|��<�|B)��p|Ah����P�
wa�%�Pc���4α��� ��Gd�M��9�~�[6�h/��,��I��y�jĝ�W]�H��>���Q�����%�#t�nɩ`Pi<r�c@���\�8�~�l�V_5p�>��>����s�s՜�]a�{X�՞�,[�r��������=\���ә^��
\��S�t>/�^ñ���8�V�?�����OnGD�((�A\$ܝ���&�㰂�UA���(��
�+�l*K�_�S��V��H��ZfF�n��y_KX)c�[�oy��<�1��@���&��r���:��@eX��&m�6�vٜ۲� E��Y��=T&����wj�d�g��T���OL�v8�%A��#��^�_�Fa�3l��m:�U#c�G���u��7}cD��������Qt;��R��Y� q׋B�O����uq=�ͩ�ǘ%��,�ЬbmW�w�Q��x1pX#t��T�ipB5�	����
3��y�K���/KFy��,�����^�o����k�>����ro����$:��;JXV#�P�M<�e�/ \N��J��>S�n�;d�_ab�hA���0����U��%��gww��7F�M�����w?7�r�r��	¨���F�����vɵЅ`�ꗂx��y$Yf���3A�=r�~X���$��Ylݠ���aA��L)W�)!�Bچ~���a�dbU���Ͳyhf����`���2��6�f��f��I�Z�K�A�J�جd�u{���歄8�r��B�j��Vmϗy�.�U0�%a֏V�m��(B;m����S!�����ᕲ�6��.��
TT��Z��i|q�(�����y���Kj(v��K�s�1��ƶ�\��u�����H�Q~~�]��d�h�nG��3�s��1M�T�:G�89Iȍ�9C��z��#>3(:9�:h=ūcDEm��M�TΘM�p�g��n�<H�~��� M����A�b�<BJ��jWs�R��#@�_L�^��G�G7fvͭ1�PS���M&Cׂ(=(��ahv�#�4p銵�2��,6��v�@�}�5*Ѓ�}�L:��P���iB���W"�&��G��k�h�)OaA�RR��S.��O�Z�Ȗ�2{e,M����wJ>����+	�v���u���	��^pL��B0��|��?<H���p����U{�U��]K��v���Ӵt"�)`�x.���d>u�\� ��!��L$(wae>���-���D0i��6�y��eP_H�fj3����"�����g���-�|JTA�N,SR�t���R\����}����bxiz(D?�G��3Hu���-�G���S���LX��>��s���#�H܀�0�q���)�mA1�q�n��T5�0?�� �g�c(���mr��%���������4��Bp|������f	>5`g�4��*�t9�� V�.e=�i���E/¸�<�5�:��"e�X,�=a����w�9�P�9�a�w�q�C���7�/�Sę�1-�/A��Z,y2�#%�)wP8�Iz'X��\E����1�Ȟ���K�t���w%�&29rz%�<͖*���41i&#;�~y,���`l�6	{n���*7���4���@��*�#{�bEK����|�k�]{I�.�щ9h����{� ��<B:1kc�i0F��2!��Cy- �U��/�}v1��8ah�v��'K����������=2���~�����m2���2�W�D����;����~=�#���RdDn:��Q=�F����i�iX�
���/�@!>MiHU��V���!���m����_;;D��~`�:�׍]��+�~�*���<���w��.�)�'�_e��s�5�@B;�W���9)��I�1�+�y����V2>˻?F��8�l�EKؠ�9l{�Q _��{RFy�7��C�s��Yd3�;��\���N�&L�d�� �D �=�H,ڙr�%�=�7q譔�D�����c���'��_���y��jХ�������MFR�ń��þ�60�Q�S�S�C $dGq0&[���RA&���8������O��
��5e�U��c`�f���<D%QR�\Տ���i�����ݴ��*#HrF���Ա��U����<�������=`��߁:w*w �	q���ξ�e�]bF��*?��}f�������S�x���c<�Ǝ�"����%�<l �R ʄb���s�ǳ֮m�!��y��������9D��*�";jdi���B�tzj��i�6���2�唑{�Y��?L�M�WTFD�M��:�e�Ry�	���T*ђ���2ցM��: !HR�
k63�O8KR#�JP�9X�Y !	R�WC���l�!����p�7�tr��ʉ5��'�D�>����Ikܓ�u���W�����y��мv)?��D��1��>54���ޖ�B�#�)Y��`{4��	F���`S
QP��6��&�e��XC~貿�.��F>�� �}��>���%*3_a{��6�l��`��B4qx4��5�$����wd0��q�K���{`_{�)��N"����\I��@{Ƞ��ڦ�sB�-2��m[N_]�066�뻛CЇ����`~+]J���k-.5�� _2>� , �yD۪)�:E�CSb�Z�,5�<fx4��)��oc!�-�cM��O �d֑�q���D�5�R���
+�l,c�Ԡ��l��K�8��y�Wh���o�2TRnS����R��2��	��N��H��Ϊ��2�+�9�Q���3�
Z�j%/����7�����QR�yh�RԀj�U���q���`|Yj��=)�N�C��Y�!�{r���A-,�3�P�E��?>�4��кW�1� �&v��槴����Ø> ��>jn�1�BGٖ뎧HATEV� ��\K�������r�>bM9���[�3�껫y�?L��N��K�N$�W�������l�����������˪?��7}u�Of�s�e8����k�0�@�����FK�j��ݗ2'1"m�J��Z��%�Z�N �@V�z��3b�H����c�n1��4b�E�hh}4-��g���3'X0�_f�];o�� %oy����la�l�D�o�0�J�Mlݰ_n�I���H���(q'l�;?�[!k�� �[y��t:�:q6�Y!L��W��R�9�1�u�����7����=!��d)�4��s"?�^�C@e|M\����X�d�U�8'v(�g����X!��O���6��k)���Ka��4*�k�w���z�q��� ��(LI0^F+�E�AA��;ax-�Li�v<e��|t �7���;r�Wd  l�V�N�Si�˯L��X������@�r�uK���m���&?s���GV�M�R��z�Ȕ"mS�6 m{J5���"�&j�zp!�Tɉw|4\V@����O�w���n�ٷ�Ȫ��?b�1�R�N��IG��ԧ�?�x��rf��_w�������>���ɓtW��Mʉ�)�c��� ����!Ѐ\׷s7u� -J�zH�d��IP;�W��ո˖1��?�����k��՛�B�;IK�t6��e�����9P�i��c\�� �!�x�?cZ�\��v��B@i�lEV���0{�����H�J*d�}`�DO�+��B�L'5�i�x����n�� �h
*��܆M�X(;8�y Y������ai&�f1��_�
I�f��3�AO3Ӈs��m�j;V]-���}�-0���|�%���?����OG�~-���y���1���T�
k�t2���+����3b/����e�{�K��\����X�e��!�(Z���=p�ڲ���;^�X����\��ʪY�I̾�y���}N{�f9QX.E#���Nς��&;��Ve��w�����������1�`�����̄Ce� '�1�)��v�>N&�5��0u������2T��^�G-Q��pT��A���NǛ�e�(���y;b�[K]B��r4GK�~X��\߰Ӡ�ī���zC�%D�`ىD79` �I4:�{ɁZ���V��~:�y}�H�O�򸪭�'��ˡ�T�,&k;����b�R�o��+-7G����h'E1��O6�1��)�fj��ǩ���Z��, �C��k���
���a�g?��=�`0�oB۶EA���⦜���1����@���ؔ|��Ѫ�����8K�)eܿ��5�b�*�]Z�1~�73� ;$*r�������:ʯR	��h�tn�I� -#�%���"�3	M�MM�#�^�JAu����u�c��E�7�$���8C�j	l�=�rs�K��g9%��'k>F���_�|�|:�?��riC�$f��ꊮ`6�kS�H����n۟��A�0�Ո�q�ص"{fY)Q&V��ދ�����&#q]ㄦe�۠=��و��+`8����	�yuV���8�bI[/_�-�*o��G��1*	ā�&�$�_=���{k���-�&�D�h��Mg�* �w�MZz�'X{�[꿬:�n��)s�N&����iE�*d�W��<~��B"bDA��	.T�vY�8��;Pi�*0A��8�H����a����z+77rG �e	h�~
k�	0]��f&���Kf�u�e�&��c'��c��z�0������	����z�M���34��^� ��%�Lg��������$��mD<6�����0(N��ހH&8m%��� ۆ�yM��_*AI�N��8��0�G������j��S_'Vi@�)���&<�YY�[��"�;���ּ��	��(iq��i�զ�l�Y��/	�%+����l�v��nS�����T��D1%����{�"��a��
��&�^:�E�W�G|���@��[��W|@��h��s�D���$44�O;��COng�b��\噥��3���nU��0���6��t�F�N���b�� 
���SF�)G�y�M1m�p5�*ME��+S/9a �H�#K���eU �(,�c�_I����,X���Q��~���Nr@�?#�#��$PV^H�U78�����0g�(GszJa3C�O=x/W��@@��{e�G%�=9G�]l/�5���}�}�nLr;�\�Q»E*Д�7�)��^�5�����a���I��P��Mؗ;9���O!��q"ݕJ[�"�{����lY/��xc ��xz��BSR?�P���8tƪ殼ȡ'�4}�"�q�-K�ot�vO��S��e#9n�Ѱ�(���xR9ⵏ&-�Cٛ�Ј"R93�s�l�f2�ŷ�=�m�E�dP����M�:����'�)����)��Y�J�<CN4����C�Q$_4��d#G��)�rO���+	~�>�����T�#[L�bW�gj��#���`me�6؎;^����Π�tH����	��_M�^�[&�1$�d�ڥө)q��-}���Iߞ�-�F��%g�s�.)_���6�+-J�K�~*M���j����'�.����Q��nHٽ�d��w���c�����{��<@�n,]T/��bP��x�����X���لN8�"�VLS)պ�v��㽘W�~Æ2�mS e6�`�H�sr������/�P�4n�����V�~��!�&o��k�/�e��������:�2�.�e�����LrVr�51��09�a�Qm��2|�N��m�S�ccU|��- 4�5Qr2X��"���<G�lM�R���$N�gK�Pv>[�������R�����h)s^$EP��G�*��&q�6��5�N���YҏAFT�>g�խvZ؜_J���5���橖�Ha����:"�DD�5����s�$���wh�F�PĿ�-����=�vhn`\�	,�%��>����}��g^�v�j�b h�^/z5�)o�׼�р�@6�tu�7m�τ��3
���������y
�����@z�n�,��<[=�7յ���SNц'!�Jl2��R�1�6�[�.6�J��ij�%����ٵ���^=�kE��b]��o�Nz�0�X�|J�NIʃ��;��<b�D֚��9_�!]�ߤ{�^�chB����\_�qnWT��볮BDjVv�������1M�j��_�$�����*J�y���� �2��97#E:��D�j�i��[7�+�,��5i{��6E�tM\j��*.A��R^f�^!�a�s���t�P����6-����p�U#�k��5��DbO��Q����K'Ґ�2�z��/��{܇G�v= rɌ
���#
^����x�}Bl��@�iB���|������mM ��K�2�S��E�r�;CM�WH��VK�Cg&��H�mEſ��]s�#�N�[b����� �=^P� l�fR342��z�0vS�_�EV� u�סڲO�l.� IP���9#B�-�t��%:CUZ� �aQݏ������o�@h{�%V�ֽ$)�$�qqEn�Ԟ~�� �wz|���iZF��"X��9�Rd�����e� ��$���y�[���&����{pVfz~��>��
IÒ�P�¼�l������M9�]�V�>�H���}���R7�b�@+�^9��U��� �����C�+xVu�zS��n��q{O�f�(��u��+�[ �*��g��u�â0��%)�41��ugЌ8�E֜hM2O��K���`��b���9j^�y��X0��#� \�\c�ev�F"7;��v�pA_�w^�of-�+'��Ʌ�=w����8�>"��W|��CK!��1��<lJȵ����8j��á�dE�^`'�7>`�9�a�,�,e��=�I�=�������L��{�����T�ݻ/�1�,��|�2n�8�d��Y��Z������8Q�4jJ�R��Ȋ|3�V
(�)�)�a��Z��1��h�Bxp��C��?p�>ߎ"G�A�ಐ�Ƅ'Źe
��~(阕m�Dǌi ۤӯ��0%ŝ��W�@�j)���
G9dLBK@������C���L�ڪu~���9_j�Gw�R�6�s'��ḧ^,���9��S{�R�����~K���i�޴e�lX8d2�@��s+�kh�����$P�Rc��̭R�	q���1� vK�eu���ZA�C�}�"䃧�Tx����(�D��3���(�h��v�����e�H��8�P�1����A&�����5�Z4�����"����C%�q%HP
k�G�zq�"�{�	њ����o?4�@�z��S���hK*ԫ��>.���"���a�h��a����í׊��W0���8D�������K�[� ��C��E1��yZ<�k���P$�E��5�l���?�v��d��"үwT��OO�N��`:f������1(R�R⫘,/51�[����qΔ�Q0�ԂA��8�o�����Q�di#���x�{TK�F9o����yz!���2�E8�]}�-�[�e�Q���f�?	D��+��[��zq�>�Hq��/}��� >w�T�*��uÍ��N��蹐���p\����H=ؙD�)��-�p�w��4b�Ϟ��UĉzZEk�;�\�RM�>Nc�f:�9St�-���� ���p27��!Ðl���m9�J8���}�r6�M����(��[���#x����[%���砒���վ�
�j�v�'%���_)3���I�\��h]��,?��z�1Or?{��֭v���PO���v��S����'ޡ�w�����|#��$�l�>,�W�ٟխ��)`K"#��1��D٠�\�vǎ �=e�d�S!wp�X���6eu!R���_�	z��M�;�K)��/��%���J	�,L�eA�b`���
Xd)	����/*5��(����-E��!�`��J�8�#d����Q��#Um�Z�:+��� �=~e$A	F��6]��*�	�!J# ��\aj�?ҷ��dݍ�<Av�Z��h>�y�����^���	���ڜ*V&�!����|�<:oxy�6���m���I��q�"�H$k]�HP$�&D��Ic������\�|�=��Y#�Q�r��Eu�C�v c����
9/~�J�����s��c0sJ�͙��9�b��H��	�H��M	�k���>���kqɽ�S����Ԁ"#�,�a�ba�N|�I�w�,v�ڪ�qb�u��	+���83�����r:�Ӝn��.h`S�tJր���Q�*4�{{�1��Yb��|���f�_	�t�Fl�G/�qnz�Z�:�b�7i�^Ds�`���3�6�4�l��d�ez�8BP~��}�Pe���4T���u]r:��`�y~N8�vG���okYS�yaԡL�c���g����3K��M5�����1�pN���c�-�A��N8#:����Bb��tHcG2��)���nB������P"F�(� p�z|���+�I����/�#&XRTq�j,7���7!��\�ء����M���_YrN��K��1i.� �í>�Jr��0��-cQE���<���9`z?�;�LrM��|��k�i(�a��u�uN	�9F�BL�z����p��^�q�pkI')�O�K����9L���Zbm1�,��1_�K+z �gf],(��w�廫�n1�	:�H�ǏMV��O$��=���A{;/�@�z�u2��Z���|�;^�vY鑁�r߭Y��Kk`e��e�t�C�k���4� V�l�^��>{�t_^�x��D��_A�hHo�dn[j��� � �B;cӈH�"ĩ}�5�5�ZƥLɵ���������"��o��\mu��1E0ӧ���{�B�^�<֟�q�]�_>U$��%
��Ծ�lw����C��~��3J�������m/��`PָӀ�<l�9��'�$��{�S���Rll�k��$����Υ�s���f����((�&?;ݎ�%t��o��%�?�RƳ��{���#�Y��O��e��f�k�@O%��<��*R�{�U�q5�w�WA�S�}��ܷ�2�m����@A_M١���"l��+Qm����fi�p��ƞ�Z=�9BV�]Ŕ�E`�WF{,)H<ce�k�vd�|�9yo�U�Nk�5y@�IY�R8;�I���e��\;;���|&j�"�'���mU�x�Y����u��K<��ؼ�1����KU��b�����=y�C%K����(�Mg-�1�y�mP�'=a�!Y�?����4@�?�6y;	ٺ:gޯ"�L:��lC as""n�o|����δ�,��� ���ўb
��f�����l���5�l�1�o��b:d��iU�O�g�дp�����XZ7�W�#��f ,�����Oفԩ�E�oUD���!VluX�d�Wp]���}{/7�K�#|Lۋ��=�G��T\���=��:�{�؞�8�gP�7lR�Һ�z����	�M��Pܓ�>��q�����%���)0����($�O2)��~�dǣ��Y06�ǩ�F䋌u�:���)'�������X`N1���4��	Y�T�Zr�CuP;2k�]�k�t���������� 8�xp�^�٘�x����3
�!\�f!T��Л�S%���\\�'O�M(_P�:�F���00Ӱ@�Hc�z�ˤ�$���<J���P"��U5\saۗ��Pg#Jd�"�nEN����.22Zů�!�F�EF�r�ID&,Lx}��&�>�]�\r����,�����N*��e�)���0�`�ؐK� {
k�b��U�&��4�z�]�DO%G���
t���37��8��4 yTZ�0z�JfyIZ��9��63 �a)�Wp�p@���1��D��dr$wʀe�Q�ܥ���y�I1%�p�U�D�4���7�D7�os�B��͘��\�Pw(�{Xp�cΑ!?+r����R����>"�˩�J�ˤ�Ϛ��lὪEM��`�3e���%A�Gг�Օ0ࡶy}
����@��L����u��ɞU���ȥSn�tV�t�B�1�cV�� a`�'�/JM�Օ��S�`|[��9�2@Zf?��%'��� �&Mٸ�/���T�*ɾ��M^�P�4@v���ax������c�̏{�w��>�X��N�ܺ�'�{�Ur��bv>BJ�Ճ1^��ٛ�8x��P�8(�y��	9]��a����5�y�FT[h��G�6��%}*��N��}�A��:''���-R򀘧��P�� �� /-��];j�/�|�Z�{�>���Q�!o�A`eԦ��V�Fo/k�ũ�S��d[�+v�����M)�7[���S�A2�� iMqd�qzlU�J8�nV� n��"�����V�I)2e�v~����*zQV���&[X Q���m�]�ct��1��U�W�I[Y+��S��b3����o(�� �DA�q'mY�7s]�9����O�����м�j�X���������-5F�z�����z('��M'�	�K*�J�+�������;4޲����#�g��z3q!�hN�F�D��,�È��P�M�� ٪�yإ�S3MP�Q\Ĕ��f�����hK�ᑑ�#t�WU��fC�Ho�	+0�Z�����|�`��"��x�?�`��vx;�e ��?;�B&�O��VB+;����4Rn+���Ԭؖih�<�����]�0h��$4��1����T+Ol&xh�.��<��T�0!����|�^Ap��@ڭ���ۃ�	�P
�WM�s4Ao�~2�׽8��Z"Gn�>��"Pj$�W���,���L��"�I�c�.-�o�0�K#��Ro
��lGAC�Xټ�࡛l���W�
���F�g;}�� �"�b��iCb�)�[�{bf@�+��Z�[)N���Э	��-���b�FJ�ϵ����m�/Q���Fh����K¯�������&tqd�~��bE�|rE�����W�
킰
X(�0��ILN�{���Ц.�h��k�� �'x���ikz�	�'�<�`��=w��W�P���k5O�@� E?^�,/�"�4Vw�:�|�H��Io���4T���⥊��J�ܙF�b�@f��MҨ�b���AƸ�Oխ#$���A��4'F죵B�����^�Q:'X�&���z�Qߢq��ұ@���(�hd�fK��6m��q��C�-�0L(�Ay����Y?�Ȩ]�����0ڊ�4jzC,@�Sm�{����EG���!��#	�1�h�2ג�r��.6�;���8�����m!�F�bڗv�u�ta��p��n�x�i��� �?��|��`j㢾s����p�߄��o��oGG��q�B&�Q,����j\�jaOj���yo�faYӂ����9� ��P�C����YN^�j^nfɜ���Rݩ\҅4=h)q���T+�-=_Mc�a�M�>�e��0�l����Ȱi$�9�d�Yٕ���3�L�ڇsR�����[�W�h��I�rj��Fj>��mt�0��J�,a���,���Რ���$x����5R�P9��� ��!�[��Q�hz����/q���5����#�d��Э��)S&�!J�:��c܂�"Z,
.�=J�Puܧ4H��e�k�,+2��X����LOB`��5m���k���q�ս����Trxn1�`�V��'�x�f߉���F�x��X�,���fJ4pu�_[��[@6�;�m`�]L�:=W}��[�'xg+�T&%Np�,�&�K���N�D�ʪq:��a�L�	���3����15Z;�[Ɋ`���5���;�xkT��)����I�i�,����҉��$�w��fU �S��6_�M�T��#����D���H�mq���O*
�]�T�8�/-��~���l�VĐ�E>�rݳl�����jT���P_4��ki�@Nu,�:�3u'��G��tU��׽����յ;O�\�/(p�C�������\7h�;��r$ʴ�W���慿�ڐ����w!�<9ч�:%�K�)���2��c��t#�t,c(ANX��R�P.����^��DL+�l�"Ϊ!Ym�{=C��ҟt¢z	
C��|��b΍.��y,�׸�~�(���ũ���hM&��y��f|�RA)�x�4e��F��^J�iK f&C��O:���J�����e�T~��0�+�W`����j�_��u�]G+��� {7@�+Vwb�G4�� �lO�n�'N�l	_ޘ���O�����	�m��ԟl�6��CkT���7h5*+�I�t�@j��tsB���"���	�~n����>��.��y�e2Gx~�*y�m���y�+����zw)OTB)2h��퍯*��ƾ�/���S�J�i�U���aO�$7L<9&s���Τ��b�C�x#{��Kf�n�F����� :wi,��Y��7���,�IC�Xt���;���(�ہ�/�����U�|'��Of����*<s�%|ae��@ux�ܯKHq\)�h:�/�(D"���Խ򳂝�'�䤌��ObN#�F-1�2���yKkOU�:Zn�g�&�V�`mĶ���R� �������,"�<¹0����6��k���>�9�.��&��ߍ�a��0*(;`S��H��:�j��<���^)~���hK[�Y�owC-$ ���:qh�E��~��a�1s��&�7\��'�$<m1d=0�&�6�?�>�Q�I�q���\)��{ ���'��[f�{y��ċ�	��S3<\h�H�;F3���+����&<_IZHl�ڭ�*�$ 0��Y�u��G�׭�O^��z��F�O����Fۭ����"�m"I	y�Yh��[��Y���y�P~w6J67���ٳ�,ʅ٘���*ڈ]rNoy�Uls� 	��~o�^�8�{)��~Ő��GцJ����P'U[|F�)'�!�h|<|'��.Q�RE֧�F ���T�R�pQ�jNk�i�5~SD�7��M�u��T6hV�S��lW_U�X�o6fMrع������5b��9iP�H�;U��k`sh6�b.o����~yhA���T��.�������'�K|�.��@�^���֠ǫ2T�x�.�i�k�H{㭆 �n�$f��h�d~ԧ)����Gz���de�;��Eq_�W����Ma>f�A���ICV-�����C�v�]dd���ewdd�i����>ޗ�q[K���
&$��s�"��������Vܾ˛y�0�gle#K"�lx�^r�4k@l.�g�����	g6�;@�WJ���.��"�p��N���;�H��;��#HW�q��#de��c���#-�9�D3�w;�� ?�k�j G=dLQ�+ݜ�N���C�đN_�j��>�h� �4q�4^��yc`j%{�+ߒ��E������A�p
"+��`�S�G2�8½�	Ո���p��t�S��E��`r�O�)���F�(�D��� �Xo�V�;��N���ƞ*����q;D��oG<ݍ�Z[<W�F�P�X�@�f�d��:�b�����(���C����^�� U�؊�ߺ^�|��nuޘq1,H9߬�g���hEX�_���|F��)r���hT��%	&3,-zrQ$�����Y�K���Bf?�������=e�'��k�m�GK�~�*,�d�x���B%� k�^����<�}s��
���b�Fj��������S��HI?ߴ�n=<�_��F�4>��^�v�"���4+�����{�O�1�'e��.-��:8蔋�q+	�;k�fH�n}aA1|��L�b j���8Ȓ�� �>�������F=����������q@*Q7�n>�Ƚݤk� ��M^��-��W����(��"QU��핉kp��:f�f�^�/�2��+]x`z@"t�F�\�xl�<Ğ����q�Q�E�&v��ի�i�P�W���p>U���[�P�ԤW�����,���-�O����GE�m\�a���YY
F�TU$�TBZ�A#�;�?~����w�U�#�nLD~<GX�&r�U|�G��h�9
�	}k�q��V�}�f�wS�-Be^������u����7+��\ q҂�z�枢���bf�g[�'�����R5����g�8x�Fn ˖� ��`K)C ����3� !wD'�w��0�@D�!����!� ѳ�)�п\a�'��\���6�V�/� ���=�^Dd�V[��~�R�F�|x�S#��
[��_��` ��?���.��^B��6��X�5�\/Y�z�[��QJ�������l�D��sg���_���q�<p�7��"fZ�RG�@j����_��l�����^Z�6'�,����ޞ�/���Uʨ��ݏG��""��G�m�i�����ʰ���&᫙h��C �s5>=���˥��m���S����;^d��x&A��b�*,�3�K��&H�o	�����,.���F]lf�{Ay�޺�[�-Z�/ ����Au�7�ĝxdMU�~J@N�O���$n����~Ȑhv�I���&j��@�� �3�oftC�V[&�Aۭ�s���h2�Rɽq�3_+�����R��l�ePF9
���Ǉ�sO�>�8\�
�\�%�+`telq9fX��U�~��^五��}�z@H��!�M��]Ӯ�s���(���K� ށ�y^z(˫�-[�y�/���;�GCÈ�RH��rZ�� ��z`~��-�`q`e�i�����V��JXOx>�)l"�tY&�M�ђ�'��\������.wv�y��h��庌�Z�����8�8���B�+:.�z,p�$-�̭z��5L�Y���z�!�[��x?l���œ8�ݲ�X��x/6��H����x�z����Of
A�2�9��Wn�D�k��>�vl��������M5K��;$��\���g閅��� G�C���ڽ�D�p��0*Ըh�����%����P�L=��gEX�c@;*^�Q2B@�I��2abz3{�ײX��H�랏��]g�\#1���bH��f�넎���}���ל��VE/��d,��UW����͆�w6d:-t�i�^�ܓ� �<ʌ�$ۃ	x�y�ox+Wn�yz�m�����%���\��!f��?oN����(�R�Q��B����L�Dsؔ1�M!�"�1%+[��(qY���Ȯ�fxTqO����dM!{�:1|Ϝ��U&ᝢ�m.SbSS��*.�"�� ����ʧ3���i����~YWآ��z�Ň��i�a�ûP�'�
�V!ń���}k�,�X[T�k(�/؉/������L2��S�T �ὕ�^6#p�$o�U,O����YZL4c����;6��-��ü=�5�Nl!˃�޹�E��^�A���{�3���@�vø|��F�\��4oG��hEC~D�Z����)�a�/W�i[)��v�������&Z���17q5x��y	ڤ>�����Yy0�&�����J�)Ԁ��iR�S9���Mx��k���Dʽ@n(�E�c�L~��R��p.���	z��>I��z��z�h޷��\YR�,!�'��� d�����!�	��ju���� 'd�U�Gn�5��ɮ�Zd�%��B$9��Z���eq�b�s��=���|�=u��:����:����=����1��
N���t��L��k�D���m�����k"��x���}�p�1;�yM���1�/���T�9K�G=�<��4����|�!�1BF�q��#F��*C����6*h��r�P ���'۱�����@D��Y'�m�36�Q���Y��PFL�\^	п�ę	�DM����q	���L�|(ZO{�J�gc<+����< �aWz�w�N��t�nW��@	z-�� ���VC;�*<a�?�m����P��v�h�n��Y,��K����0���a�#���_���D�w4�g�K�Dy ��y��r��0% ɔ%�p��L��Ƞ��I�,#9��W]�>��ϖ�q�Y�n8Nx��@�Sg,@������a�����]���N:�*�ڌ�=���}6e#�G�z�3%�f��W����:A}�Gq�iEE��*L|�!,�Pd�\����:F"��H��|�l��ZߌDg�gɏ�I}�.d��Cr��.�<�'74���,жV���k.
���GW��^�=��݃�8M0��n�2+4���@9�󴢆��U���/$��F�CQX^�Z�Q�l=�L���J�o6�W	W~�ef�@6~eFگ���j���5��
ӏ�_(�Y�5�x���z�蟆u_��7�>M��4�#�\�T���9뗦�w����q�U��M02�Ӷ_�U�wm\��ã
7�?�2a�^B+#/���5U�bx�bT��,:n.�	1�TN�d7.�͘20W����������t9�xp��5x��K�d+�� �.Q��K|1����`��CO��¨u���ݦ���%��8�@u���٣JF�{AL���V��4�ؗY'r������[.�#c�^�'�9����Զ�KN_���w4e�*�XO�E3��#X=Y�p�e�R$ƃC�ݮX- ����w��� �
�J1����h���y�bW�m�ќʇ�u��:��m6҆lv���	a��Ql���s�g��*�S�F��up-Cli:�5�Qcz���S�afK�&�yAr���E�#����?�9�-�	���嶸����b*p`%H���\O����Ȃ�@�݄�PsH�!�)��3*>��h�A��������1α���0�vQm��k<������L5S��j�)#��hb8(��;Xp�������| $c��-�����w�h�k0�����$�`"_rr�y�@�r� F@���}i�*�>��1�-I��U�2�H���R߸ ����1q����^�H��įJ;0pD�����=�_��8�z0��K"��.�cH%al�ה�g�]�I�)�TO�W�׫H�E������
Eq%�m� ���L��;˙��H/�X��,�O�T^^sV4����ia�Dk��\̳�z��:�����ٖ�+���/hۏ�`&�(k�v�d#ĞV�yC�t��>6�,[g��$P�����Tùs�����:����#+tъ������$�|/�*�LpnT��@-�j��t��.�a��p'����3���W��=c��VW�g�}�0W~�͙%@���GU��篎�X�~A׌-w�����,s��3��w���!�Y�fvx&�]��hP�m��O�,bs���K!��d���E31��4���?=}T��4��7_7��ʘ�G��8������%d�v�<�G��ඎpqe�u�A!�#gVqn��;;�:�l뽳Z�Ov��;�3���<4�|���Ҡ�K}p�x��������,!";]<���uF����)Q�nF��j���xg]6M����V*0���������/V��k/@K���ԸSS�?���ȶ���r�%������νG�CH*B8�1#�:Z�9ټ��X��ڷ�#E''�~� ���.�7�YP�C@��ý5+	�z�y�h�LJ�w�Sم�ʛ'x�x�cj���!3Y���#�ҭ�sP�QH�g�|e֯<Z_Cț�g����F��+6"a�ߑP�Pv�㓱���*򔖺8�̃���'P_�9r�(B�x��{e3`��4���D���Yy;a�[%�B�^I��WCfB�6,Dɸ�lem��}wEr|ku;�l���௜��z��&>�v!� oI��'�����,���]�R���O�xk
���^�L��I�������h��ɝ�7^?ג�(���]�DY~6*�z�&]\Y�n�X�/��E�����7$�ԯMA였��sΪ��K�R`M6��k��^��0�ʑ��S.@�)�#i<�^���%+�D����	�)Ң�l�̅��0��t�������&�W��/��aQGO�gݖwݤ^�;0ظ��䫦#�� T;���Xt9�.N9��2r�4܌�~�F~Y�pY�Ҡ���6~4�=�~��eO�	9���i)wH%�F� �t��!A���.(�U�E҃P�����.��uРB��"�r���#/���|��>�/��M�uY_�L���!w����"qK��jvk5��F4���Eym��j2$�A��{=h��n�o)
;��<y+���,O����Q\!�2�zv��d'���p���XAaj���ݙ��w,<A��5��[��,ԵG��s��o��VO�y�%��}5��Ѵ�"����A�z��!7�ĀM_��n7{���=�=d�̟؍5�P���o�P٬�e������!����u�{�8���wQ�f��.�
I�!�>d2+!zp�v}'~R��Yn�;)}���(g�J�8�F�NBG@�<~ݬ�̡�Kc{�ʦ���o��dsձ��wq�*o��,L_(V��B�m�B��zmlb��� {l�6Bpfo���x�zC~�� B�l�~��\�	�a��Z	����:��azT}�S���ӳ�v��F��������t�>9�Z��x����0�K�7��'j�
#�"�Nƙ���Ϲ�`H*����Z8>��Z��f���S���|b8I�N�*^f���F���(n�t�!["Ypz��{+�ZO������i�{��	8���_]�Z��.��jw���-�����u�Q8���]$p��lZ2��k���� �H��H*I*�f�m;��VEd"�V�e8��ł�,oNT��td�<ͫ�
�3o��L�!���N�?��%^���气����g"��
׻�������T*S�s��5��ha���� �$(H�y@I3^�C���+nM֣��ժҳo m^�R��"�Ĩo]� Y��u��د�z[�z�����k�3`/�NV0G/QϺ�
 ��A|�D���P��������К�O��e�% J��=��dp�,�����
�ʈL{R��d˜��.�M+�39��!�V�A:r�@AB&>qQJnȣ8b���3�ޓ��(����>�]��ftDP	nv����t�&�͇�J#B~�&���5����� � ��қ�> !}L�p�vc�?U^��z����F|�"`��/�Q:�]�akp99B?�1lY$����9	�Eβ|�Wr��wz���pI�8I��-����z/2�:_�A�>t����v��{
C�Ã�	8�C`�jVV���&����)e��i��A ����3,���Ѯ�3�8 ���!�("�� �KiK*T}���LC|S��luע3�Xf�DW�O�8�������3|D܃��s|%R;DKL��*&<h�q���m>u�*l���+l����$0N�i�9cp�]0��vb�t��w���n6"I�=��$��A`�k���q��.�q�0lp��~�t
P�X�3ql��T�*f�-��7j}�l�;�H�Vxb)�ڄ]q�ꏡ��mߝ_pl(ƍR�v f�.$Z�Z"sZ�=fŲ}��A�H\M[��/��*��N����ẪMNB�����x�VS�x\KǓm�g�b��d�W�A,'�̫ '�h�6���r18�W�_zddĬ�WP����.��6�R�w"^��I�-�1�Dl���c��mk��ά3�ˮ�|V��ٗ�U!�**6#����4��H�v�rvͱ��/V���DGd%Ha .KcM�<�#���T����n"�	�y��~�������z%����~���:�j��v�L�E{Q���ܴ��94����������~���x�k	�	G�Ūb-{{�'�)�٣&sE=�fP�{��|��w6V��&�3]ydz��A쾧�QKOF&RzOH��^��tӉB�L~��F�os�3����U�H�·���7LR�`�u"��D����&lL�J	d;^$���]���g~nKk�UNR{��n��$53�
Id���$��m��f-� ��\�4�Fj�KM��(l��gز|`�B�y۽�"�p�:G�@��4��	&��6���� D�1FI}%�i�]�C��Rq�if��Nf��\]Q�}�l�� 4���d��;��/��p :�k!S�rB��B�.N�w`%R���\~/[��+�@+8����3���҂�=��Jh�
Pt�����M��ۻy��_�uu�S2�y���BG��&�l�K���N�/p�Z���'e_�F�����8����Ht�J����"�O(~�h8��4�����S	8L:��ǒ���9*&�ټ4����A����� p��f5��Lz�q��&�(����\��/��+�O�HյE�p�u\���BV�B*b�)U؜� �*�y�C�~���*���]Z��3ݽ()`62�˳�D��AI��ҹ��n�?V�M�C:���\���1VJ��0��8ͩ�(���X�Ř�%?�\�I� \�r�U�hs���+��"�.Y����e���5�wA�Y`y?=Irگ��˥��w%����V��l>��)�cW����蝍/��'Ҡt��;�y�AD�X-�}5�t[� 9H,��9�a>b5��4����ǿQ�umC�A�� �i�e�_�jƔ�o�v�A�Y"Z�..��[+Ѳ���S�Z������WC�������U� Tϭ��Mi��A��G�}"��r�
)~!���Z�Q1lvXa=�t���,��)�;N����KI�_�!S&|�G�o��E�Qq��P��Yq<d�zצS���CE���h�������t]?�ȳ��Ufk��2���J�7���c�Zxt���u��L�V���ze4U�G�Q-6�����
s�����v�>���y/au)�B�{�K���b�'���:%5qǾ�6i�pBFc�|��CM�ͥZ���HT��$�U����.��F�=
lg]m��I[iU5���<j�x+-�8܅�F�u^j���,���λ�tȱw��x	��	T��ǲ�"~�Ǐ�y)�[�$^���	���)���v�	����PY�|��3r������Ć_3�3�ck�^��[;b$'�X$�|��ޠ�1/������C�ԤY�<�T3�u��N	���:�d��0u�L��m�!��⑈]��2���w��؎��R����JU�MTОj,���~�|��u�#�Z�>]..KI�ϝ*K�r>�pZ;�����.�q�Fv!�
�ɳ�8M�g��d��]5�]AH�7 ��ݠT0�I��c�zfL�ڵNag����~�Jǈ7�U��v�Q��w��u���_��+1�r]���������ny��q��t����]�ϲ� ���o�h#��xU.�����u\��#��kυ�n�\m��&�L"��RG2��\)z ��t����r����?��&Ӛ./þ��� W���Y��:����.�?x�����$����ahD�z��9 ?8̪�w)�w��X9n��p��~��g�ݢ�TH���z�f���.&�m+)�Z���A����=l���͉��W{30Be����.��v�p��Y�������*�51�ǁ���4�\���QQ�g]�7�x!�%�:v>{�EZ�R���aB>�5ȖD��)m�`2ׁ!�9j���@����?9��rۻ_&$�O�d���+��,�a����Lp�K���!A���3�XS�co�X����`�m���濮f�R���óz��da	���4nl�h��I�NW������H��EpoF��a� �1$@8��E�e� �6���a�^:�*U\c�6v�1�W���������4Q��`v�}q~OW�Z�~M���H�eǒ?��bB�ٜE\G\=f���F��()��1��Rg?QFs�W�c�GGT��q뜭����P�o��o>�jǣ�]1B���V�� Ψ� ;Z��利>�Jfr�x!xQ�۪G���5����	�����89����3��d5q$���[���PH�	h��;���9B�J�]i67���ǻ(�,��.Ioғ#i�m���k��*T�p\ 2�T��Q �.xC-�_:.�-�q�,�z�b:u�V�I�b��+��k��C�~�q7�<H��_܆����u�;";�VQF��
�������x�"�J��׎�.b��.�D����t��
�0�k�-t,ƀ#*VhۈF��׸�Q3Q���e7*�����.y�pv5��Nj��Q�޳�V���ɤ�rمoC&�O<0�!w��:����%��G��	�������w:_�i Pt�U����}�O�E����d���P�b��t[cVR,u��tڋ�yz2��m������b3N�F��;��w�� 
�p]��yb�[��㲡��Z��4��}Z�7���c�y��DH���w��b��ρ砦L��s�GT*��DX�[+���^�׏/���B���h˾T� ����l�#  ?��.�LK��5�2[`�!�B�$��@:&���p��1%��P�X��'�~�"Č9��[�8�B�I*.�P��3� Ɵ��,o�r��3�f�܊�'9��B¼�blp�n��Q���B���xMj+^��nЩ�M�$ �`�{�������PuR�W�i�������Hm�����(�S�T�Y���S
�Cf�?�u@��� <�i�� ���7�0��xd~�"�E-OO��K{9k^����7���Z���rܟP��m筃9��n�V���FZ4>�K/��\ �z��c�DrhD�Kn��ގ��ei��r��u��`��x��W׍�@u�]O��A�(
TWR��`
	Ϫ�(xF-�E7�nU#���ϗr�����eMyu	�X�(!��_�B9���i��]��d	Z ۦ������/�}���*�G软P���2TB�fǚC��j���O�QGI��B�2�݅�U��hz~a�
8oy��ޮ^BWkn���O����z�LK�#�����pg�I�M ���y���n,[gd��<�w%?�f_�ec�JIS��*�r*`Q�4ˣ�\"�5�G�ȾS��r͍MX�Oy 4����\�ȷ��F2�������\(�'`[���8����@�/0��:�;8��6e�����A� �/��A�Pҙe�f�~
e+�B��3(���+cgr����{<�o��J�Vk y�+�S7wz�Fj<��A.}�:�5�B�V�O�9��7��K���ݵ��֌�Z������q�����UrA>�����k2M�ՠ�8�1�{.��D婊�'n��C�"��QA5�P�p\��-��p���y�q��HgP�U4��5�m�M���R�/�Q��A&n�:�Z��/t9��
k��/�n�]xnR۱},�v�I�\�G[s���8_������j �<�/"Uc�z谜5�U�t�`�w!R��k�EvsIO����jX�.8�b��K&��i�y�r�������Sm�<�,�+�����i�5���ب��H���9���q_	im�|ɝ��g#U�ڃ��^H�׻���SB�y�pVô޶�@l���7�ׂ��:�LY�0����j�,�q���ǎ�Y"��\�Q�r�`(Nx�)~�成'�@���[0�5/b�+G��de�Ί�0��',yYVn�+I� ̻��ynL"��$�l����)ШӘ����g���w�[Y�/8e�'N�W��
Д��6#}.���gW�h���D_?�9�)Gn�<:ߕk��
�p�\��<{����)Yd��ި��`G��Sŧ汛`gs���t�"_��u�Ge�����EJ ;A�
�|��'������[�b�t�)�Ϡ�a����F(��P]�7�'kI�g׏����HOL'��&�2"��T��<{�>2�>]
v���c��:�t����ǉ�)��Y����&yݬ*1e��_���.M.a���_NЖi`,00�"��卞I���N��JV b��:����_�<�ؑΑ[��ӟ*�TǠ�`\���3l3�Q��/��Enm�@��>�m'2�q[/aң��-z<������Yؔ��MD����tp#`N����ai!���0Ű����v�ժ�щ���r?���Ѻ:X��۞r���͍MAz�#��WD���ѡQ�����P��<��6rU[��:ߚ��ƞ� ���z��X����y�`�#p�'J�C.U���H�?�Y��ք�N��vnY��Kӎ18+i�r�C>09B.�'���9B��9���sڅ%F�+g�3W򚶍ȘM[�J�lE����������r�
u�������N��eesf/:���3�Z��Zώ�����>����e9R� y�j���a��p�>��#��a�]�s2U�f_�<ͱn�q���ŝ����ZAQ�^�f�-H�>��@1sRP"@�!d�h����pUzRB:�`��4� ��u/���x��5�q�X�|��d�M��t��S:�����M�7��y+���ƿ�Ȓ�TfJ��K����R���ܹ+$Nv(�&:����ss��1��'������a����Hl�+�P��Zf6p��pdj��̸��J\K����|X��W_Ns��.jj�,������o����å,]'Q@�2s7[/G�{N��#������j�'DW����3��x������LIj�W'K�"�f-�f���j&;�i��1��Q?����^��C�<%n�΋8���(V�w�|�&C#5U4&�G��Y3d��M�!���̞�l�<���u�R?��}чŲ��Q�t��Ö�~�Ri�;T�TQ�6�'u��PO(IqN��|�k�h6�ȍ�2ֈZ��"�Sj���Y ��>��s�@�ؓ�C�H����LB�?���vE�ty6L�h,{���?�J��T���� ���J�@I����ޓ�2c�f+r��M,�#��Wˣd���^�#�GV�v?H&��OH\�Y��"����c�ݼ�#�*��{U���r�,�J�%������Do�����"�^C8��de�<��k(t^j��n��b-�O�������+� Ϩ�¿��̢����
f�V��*�D�Z�k>	Hֱ�9���4�.�)�?W��|�ټx(�@@
�9e���)T�}z�;Ut��;~K��S>Ŷ�@�w�mt"��������b�U��[�A&�@T�����Y<��h���,�Z.��<D�2N�;�3}�:RY�¸�'�zO6�����ca��$�O�ɘ^JЁ2U����E�aڕ#a�t�E�I�ǂ4PW'�-�a���#X�o��)�Gi���A�ڐ���Ko�����>��)�\���hr�)�#*#��Y	��-��2]��8g�F�i0@Ve:���Ijc/>{O��|�G!`�>j`U#fOkS?�E�ʍ����]���;�*>nr��Ñ�o��@��7\�������9 Z��I��	�࡚s�)� ]�4mY�Q$&��ϟ�Tn=ᕲru�?T�����O��«�o7�����SMi�r��Z�W�ǘ�(-	Z���j���?�k~��~�1Pp��4�?��CU� EY�㥰��bRr�1��,?��ϋ�"��{��p@���Cu�hHP� ��p�)8ȃ`�%	�8m��w�;�5��۹w	���Xe�ܐ�V�K`�u9�̿�(8W���K*�+���P�؇��'1��_��B�^�����s��8��~�3*��(i�'�A��(�n����uƄ)�]~G�j�/��`�����֜]i�N� BP�Ruz�o�&+�����8�IV"z��]�a�*u�F_8�uy�M��%d5"������?�JB�a!㛵�N�ʭ-����w�!��~�B�Շ}:����/O�bx���+���o�|ٚ�x]�%����=�9iBl��x"AI�����+��gl�qq�SĴ;�Pu"��8��W����]/M�g�h&�(� ���`��5�n>W*��J�C�ݣd:#_�6H�t*��y���<M6��}s>r+E\�!������Csa����>��N�E�=�t�g+R)2y�a��7��T"�pz�+��~71����uf%hO�J�>�z25.؍�x ���������ʭFz�y��G�6�6H�X�����t�F�z�����0뀺7���r7 7�8��y��h��W�Փ�ذ�RV�\��j!��u�F�<��5om�q�d!X�Bj����p^�d�,R�0N� ߢ�}�Lk\~Č̛5emF�G�WOj��_A� ��D�zyL����g��kk���n�RJ@�ӊeς�-`��.]�9O�ty�>Z��':w��:��5
�A
�q�~�BI�L�
�Ѧ����X��>X5W٦`�^m���c�G��*t[J����b��\A�R7G'���>�e"�"7r�b�k�J�b�0��U�ADO�1퇐��, !� ��K+��}�
�&r٥����p�aj)�2�{��<��Ұ�Y�1M� $����	��2��+��go����6�䉙�M�N���f��V�*=�e��5 $1x�=5�N�b �0G&ȆC�`���80Y|d�f��������,�O ������ˉW�"���O���j���o�Qu�.tY��ZJ!�P�'r�{}ȇ�
!�RKK��)l���W����uI�������]���T��u�ll�anDB�&������c����g������C�O!�jFJ^�Q)W�Ȉ6ԚH��
�9΀��R �zH
�ϿĔ���!�\WS�ο�s��%a�;�d"��f���U�����<��`�ɱoU�e0t�#��^�;�S��4AɽƳH��(�p���8]�V`��h!+��?���،��#����8���{���cy�`�bbFg��A|V���kWȝ�y�M�*�%M��e����i��]��*?{�[�pY�� :@�<�
������Ժ�)荘�b��]gBhX�u�	W�:��']��ޒ	Irɋ}����XٍcLW��!���y1�C$	]��"G��<�l�`�K̩�-�v:T���"(kCK{.�f��S1!5gI{r3N�7v�O�f���M�6a�-�]ۮ��5�M?�`�>��"[��(��{��0@G6���r��Fp�(X�Z��u��8����X�Y����@���&�հ�� tG-�SuV�
�o�_��Q�A��?_f��%R�E��@�te	<�	3) z��{��]M&��5��J�6tg�r�e3���?+�-M^,�pZ)��WC�T���,7*X[��M�P�*�����D�F���\�jKX-�jwu텞����\��11�������5;}h�6Aژ�NFz��x�h�~��q�%����c�EkW�s��f�vB�st3��4����b_4����:lH�(e�83љ�l��/娱�K���
�L;��E��vHr���؏IC�&���tG��]��oLQY�\u`��$LU!�G<���]�e�t�nS-:�LR�}��O�j;�GTh�/1C�:w�'Q��DAK9�W>2*\:ŜS�����a� 5� �M�I�9��)JԹ�ih��.&t�0�eC��+@�B.wk���*��6�'"i��J�=g�~�y�v����=ͻ��YpX^�Iʁ>��c�IH9ۻy:#�e�e���)�W���^���k�����
SR"��+�zZ�*�7|�@3��<��$a
��i�>g�߾����ߧ��-N;��*9.U��\�VB-UH�"� �G+j�}���w]�<���>
U�{�GN��a���h����5a?름����R�c߀J��u��o�Z���R�J�+8�GB�V@�m��գ�LOz�RXʔ����/���~�of-��%�5RG`]2z?pNm��&����N�M|�t�e�m�L���'v��B�Wl��ez��5�%_�;��<���'[o�Ren���B��ŨI�~ѡ�c�y*���jԗ�>(|M��f�	[���Ddy�8q�&1\�O!��Yq��ʬz�\ĂH�5�w�<I�|�z�6����X����X�ĀI��0���K�=�Y`�Bq?᱾�KէŁ4�[v�6�x_���0���*���`�@0uy�E�Y2�6���  ������|�dnf�h'F�
����xi��W�����������󂆱���ӆq�n�Wg�uĜ,�^ҁ\�r�� ���6j�jo�<}��(�Jm��'Mş�J�8V��̂�舜C*���ZT����X�XH�.Y���R��ߜ�qY?�~���	sM:�	�c����vI>C���ēWYN�2�ho(�1ɀ�-K��ɔkq9�_oT|��Ur�֮Rg�asS+.ƒ�ٺ�(\-�!'$�*��>"��"XC�k9����c��Z}Z���-�=�>b*svʔ���
�A-�r)ig�i@��YlBM�Z�Fc';�������\��c؅��h	3�S�=l��3�eEio��_�L�"��ysz�B�t�ן��w���z��7��Z�i`��Pl�)�g�V�0s8m3bT)
׾��E3kO�o�Go����3I=TDJҿ���ҍbT�<ƻp���?���!d.>��#�M*����	}���������u|u��Yk)E�KU/x�z��� &3�Ȁ2ޏ�Ϸ���L�S �Wkey���SOf��8r�\��2>���%�*"�
=0�9]S��՘�)�'8$k�eg�;�j�ǆ�{�O۫�8�\)k&$��IQ������ �k#��[ە7�A&G�<�(�le������ʨ��ʌ�b��������#��`:�
�Q�R���i��4Q����zi�9ٓ*�4��i�Gۊ�n d7���%q�U&-ڭ?(���_8&>\XC��y�iݟT/t��?��*�s'aH�I��|:y�M�P�?� ���^�(��#�Ν<'pP{X����{��'+.�ж�k.��tS/G���t�q^�Y[��e��YѼ֑�$XN#U��G�C�
�n�dZ̮֦��k7Nn7��f�v��o���3�T���!��x��xE��gݏ<�(;Ӹ��MР���<��z�ӑ������g)�� 1���B2ڕ���]$�����Fb�ݡ�_�x�������4�|��_�4.��"b��L+���y��H���#�6jܱ�6N�"��U������^�=���������vꞸǎ�{���G��E��?gC���1C�2@��k�M�['��݄͗��9�ڏv+d�^~�^ыD��_�B�Cىr8ҹ	zH��y�%Z����9���c[��:��"�VQs�	!��s�5E�גO���}Cd���E0m/.K
6�e���5�*���-����E;vU,=hn�9����칹x�\ai �%���Q�gY�$�˰�5)8��{i撊��4.�o%�b�*�@����w?2^H��5�hYY;e�;����C���#BFaNҍ%�u����?���Cv��i�D��]�Dgw�RG��o��p�n���ng�I�|��X7lB�����(�����z�J�f��#�K��`���
��~٘���H>M��+-M�7<U��K�#�6���LF�(�d��'n��Si�m�����c
X�a,f��vf�&>4��ڰ�v=������z�py{2Q*At���l����Wo��dΐ����b�.>�d	�7�,ѐ�`Ɇ?���1��e��k�r�wl|z���o ��@X����%�a����G�4��J�:t��BT���U c<R���CdO>@�QU �n9$�g�H��*�dhl��^	��j����o�3ܐ�`A
EQ�m��k����~��(�Fq�G�ӭ	����L\�vٍ�3f0�-���h,E�j%��l��L�L��P��k���a!��k�k�>��V>ҥ��Y���F7E���k((市�j��*�@� W~�fQ���R ��@łO�fN�#�uX8�Ң~س-���N7p/I�\J�^z�#٢���L�Pw���ܭn]�=3f�ﰅ��Ԏ�(�kP&owel��9D�O����Cd�sJ����H�I� ��"����r 42ۋ���O��.���I;h����:КDA��^��t���"}�w��C\�ڰe���{H)�Ox�>�!UU%�=�5��19H�<�G�/�z[~|��|�{:�D����~��I�q�s�%�oՒ�����:Ce�.9*l1��=.�����{�ʧ� ��Z��7�O�֕�!��ł���P �[㷯�Z֛ڱ��<�p�g��a�Sb�T�zë
�Α7��x�N՟bJN��� F���	���f[��-�H	+bb�"�{ػ91W�Od�@' h�h[�#�eKS�A�ȋx'��';�ϔ��]5�hu�<t$$�;/�Rŵ�"�륢Z��\�	F�;[iZ��8�<�[q̥#�NP�\��m�kw̍�Y{�Cu6"j|���W�v WR���h �AI:�c������9N��o��1�ݼ��n[�(��m�J�(�x�j�<_���@�oK��y�2�ɼ�tO�Ų,<✟R��X_�V����e@n>�ܽ$�䮗�s���2P��,�\����h��*m\*�d�Q>�ؙwd~��i�z;d�p�8��'6&9/�P<��C#p7��>��5�k��ú.{�(��[��T2�jN2�\�,;�=�?� %FnF� ����j���B����E��ve��0��`���Be�Y��>+��f^�8�!0���c}�G��z��Q���_�!͌�#�X��Pǀ m�n�f4�T�H)�#�@~��)W�tZA��
(0`pr���*��+wz��"�Wh�x�Z���u_Ңy���~�G�:z���Z3����& $�j����7 ���M���x�^��>"�����9�h_ 2L�I,H��R%m����K!N\@Ӧt�2-1Nn^��Y�
����Ԫ��g��g�Zz?&�(o�'�1L��D�gxa������^�'[l��9h��5���m���Q}sz	�1r1wU;�=)0���?�QZ���rN ɒ����Ā�{k@���m�/�VM~��Ѕ$?3.��0��<G�)�q_0�1�Z�Rr�LyN	���k?�d�T��\���(�Aym���#����B>��[�$;a���yI���ɬ��7W��'�sB��I�6�f�2����k��B������@��cDĀ�^b	�2j�Z�X�(� �\u`�[�A�-�4H��C�to%B${��z�
�-;�ZA>��Z�z��qy�
h��)X�ҡ%�%cL��r���tC� {8�Ϯ <��	T���g��6lV��-�H���B�!`��)��M��d���䵌�Z�Ǉg#��$/YTA�b�\���L�$���4:d�T�J�,���-ڨ��BDz�=כ0��nOe�)*�"������J����_l��[a�&�1[�NMC�n���t&�*����=�\�ͷ�tNV�Mw�1�7�^�^�Gk*��!b�(L��s�68w�m�w��RaEbp�(������F>���<lL��BsS�k��GSr>�����Ԛ�R�i'�C��q�PZh`��:׳Rhc����!�Qڻ��\r!E$�#�6�e6�6�}3gf*�����ª?L��U�Ȱ��nAꌆK�e\�����̍��Ø���w���q���j-�P��y�(F��=`q���kY����:3~�18�Y�^Q;"}�SI���j��7�����󮟤�T�nFz�nN��,ǲ�4I�Q稸uūv�������!;�)6y'�#A���S=6�bM8���@�Ib�q���y��NV��Ֆ/Ĵ,���z���>���Z!�͟�0OC�����_�갗_U��ϣ�#��6E�՘R]�$�<��T�$Y���{s���Q��`*�ߚQ�oL#�
BQX��Ǝ�.�Ց݌�����a-��\I��68����}!�A��{۶���h��_��yn��-���-rB��U�$�
/|�x��#AazdHϰ�� �d�J#0
+�E�S��]O���\��֨MrT���l�������K��,����,~zq�����PK�v[C�]�El_X���஼��,p���K��|f��`��r��Њy�Eƾ�/���F`/�C����ͻrU���'Sh@����v�Mš�3l�Lb���p\���aؕ�b~/E��}3]�h�
i����|���cY�Ve�����ﱅ3��
�B�k�з<F������UI�{a�cx���Ek��ݐ�}x;j[�x/�'�3��g&�ԧ^;q����"6��v��2��d����9��t�j6{�F�/�L�y�����
���ȝnv����\{jP#@���
fpA��г�~{}P���b7C��Q%�vK�s�9j��[lOJ�@>`XUd��7�F�z�ّdûr3[�7��u0 ��-\���mΟ.��h��%�|�<�:�X"��׵c�C:'p��tc���.ҿ���:��Vv����b�R�Ȫ`��/D�+'׽a���e�!���7�dk\By����ʔ�7�<x���L�����pDm������ "]�����6�!u�SJ�ך��]jGq��ռD�t@���Xd�~������IV��@֝�N����2�ϼ?uc��Z~�u	�}���H�m=���1��Ä�pQޣ�������)����T��ʗd��dU㶼��ŀ��L���~��B;���'5�sƹc��� T����J�i��d4�ܫv�Gw��"���� �8���қ޾+��ےM��7�T� y�@�ڨe=��^y�!��`��[,K�(A�O������^��D��P�J�̴#���=7�ΰU�,s��\u��C��~ǒ�����_H���8B��O�*��
X 5�l]�]F��nk&�9r��i�ȁ����xc�#�]���	*�[u�1���fS����vn���,ym�A����_K��،R���X61#S�]��k�6e�����&��[��х�Be�����4��Y�;)=Z���ȝ�6i���\�}E�:(r����Y�'C�X�Я$(ZoZ�W&�3��%��釪�H?6���`��wqH��1��M[+����ëW���W6����}�E�C����)�0;�˓�]+�a%��T
1J�+��`��W�WjQ�\yU��Yj�6m=	�J��~��S����XP.�ck.<se6&��T���������1�)���wN�|�.>f_����4�� 6�W���`w* �䈋��7l�Yź��֎�N���V�l��X�~�͚r�]�Ú,�x��ʂ���;�F�J�����nl�T��X�z��6y�'�|V�unVN��L��Kj7���!Xu��u��jn��\=/7Cw�ZB�������tV/:���}xH�0���*��iW�f%]������5 ��Wm�;�c�����RaQ�\v �B�
CQ�k'�B�o7>h���A�,4h�{ȟ����y���Xغ�l��X�oU5̘y�c撙IX�G��x�'2�g.������ɬU#��>��=�Hy:�F2��ċ� /ÿ�ȹx�E4�l�S�F ��=�x���+Ф�=/Z�V�$��_�X㕏�o����b��=(�qԱ3첱�ۮ�5���@�W�̬^~�R�R�������j��I��AYl<� �ͩ�%��ݾ���tW�[x��"�Ǒ:�'����o�_(B�}�)8
ة��%&��	I���~���$Éo�Nm��r+ܾ�r�)Δ���(�����R�:�OA<��H}7k�r$���Oq,� �ֆ���4�A�J��2m��T3sl,Ha·���N���n<j%z\��g+{*F=ӭ�Ѯ7f�z}଼�{By�&�K�Ǝ���)+����!�Ku�����Xq6��ĔH��_4R��>���n0k���4�b:ګ��.�n)�rE�>t��kIoP�p�L��i3��%'�ΐșH��W�j*��;�}����,W׮�ө�e-b����TV�}D'l�ȋ!�m����%�B�H��'�ʋ��j%��$zxQ���� ^am o�9x6�����$(B�YPz��M/W��첳-���(ЦBQ>ځ�\��)a�: ���jSqLhH���:4�!,8�������ъ���XY�A	�8#��ڍ3&.E��԰���4�R
Sz�ϧU*�Xs����9V�||�Lj)���l�R�"@,gf��q�{�(~�?Xt�5ҕNwt�J�F���O�.'o��E��A��$��F�r�d���{Gy��.�ў3`�Ǖ�2�X1�eƪ�$�]�L�uˠj�!���Ռ_�`�s���@z�4E�E����B����7��fε���u�!V~Yc�,��/M�)T��b">=���q��A�Q=��:����?��/w*�������l"��C�C�p�
�S�w���g��bj�������@/�h�C�w|sY�y�3~��h ���K��eX��W:;֑���n��tBPPK�1�M"�Q�aI�fG?$�PU��ص?.��Y�b���6��]Z�j8^�W�U����ہ���TPP��ݖgp���)���5\p��'�/�����w�MS�N����;��6��a�I�)�(ޯ��z����_􆯟�
`h�\7�u���E� n=�Uk�&��/�KH���g�Vc��ktq�m8{
�p��P1a��"£̽�WUNI�j�r<`�C��b3D2>,6�	2� ���訂���Oɤ�l��b�۵�����ɵQN9:�ۊ�+ӫ��������&k��1j]Y榋��v�Ū�V(�țpk�'�J]zpL�	*�g1��3��P �������V�]m�$3)6�N�"�:��x ��-��c�Ø����=�DQ�kN����ˇ�����#���P�1���*�+\w^1�=S����R���-"r���tPf4���oM�<N�(u�/H7�&x)K���{�{e�?g��7��&��p�+�Y�mX*ͩ�.�z�L�����㊄Q2�(d��ǡ8o*�G�.���F��ح�XBҒ�T:шC�L՟jF�jEHb�x�㒹h,��}W�ٸ��1�A���(T)��;#���uċ���է:.CV3�)y�)s�Vb�������W@Z�-%R����F��t�!�|g����ʷrV��Ck�,k�5�Y_y4�K�8bd��Z��`�1*t��a�&_����/��$U8cq��-��\��Hb�A;?6��kK��I��oN�Zg�A�*
�P�0e��D1���A�J0� �tI�ݤR���F�b�l����d/	a꼮�������)��8�����ggWZ}�)"�n�}�SfMQ,��"b���`HP��+�!o.NG;�A636J[bbC=����
_���g	�=;��C
 �`��O��,G�U��b'�� 7i��&;"(s5z�{ �˫�]H7�h�C��.���B�r�H����M��^0�&��ś}���ovJCs`t�xM��<5��p��բ�5��R�¸���ba�\�^N���,�L��VZ��:���D|~���{��a�D�<�ͯ�%n�>"dd`d�����(�jIo)d��'Ҩ�&��]Х��æ�(ST�B��Mc��a*:rS\��c}�&YL�R傡����S��a���l	�/��dN�aoR�Wi�㰧�x���P]1{���v���������h�����Du�Ӝ�!8�%�y�i^��:�$�p0�mk���p�ע7
Q|��ɴ-WO>����������#�uϤ'��*S��9�C*��>��l)�(=�M^���˖��(ܶ�g�Xn!�ڛ4v�bq��~�4*,�ٗ�Dg-�yVd���V�f[6@���y����a|���}��G�[
|�-/�co�<\�1]��Y�l&D۲�=�yB�=���.3������VӬ�[<l���7;.�ऋ��z��=8��^>���f�4����;[H	�-_��Yy��G��'=s7�
R��2s�W�Y�KD�xl��&:�h����8A��)Y0^v �>��~�`�N`�:U�7���M�7:���ۀ��^3҄��y�Is�,{wq$@�I���m����%���ï_@	R�YA-ź_��p�sw��e#{��ia�J�j��#����+�˿�#�Ӓ��ߵ6�=�#��:���	}'��p (�9}Z���?��o�7������l�/'�^�j¸���c�fH�R`, ��ǰc���0���4-*�5�oG}2Uߟ`�獐�Y���bn�&�@j�ZSϮi~:�i����eAS�V.��;)�]����bg/��@{�Gܗ�1�`:`+�|U�l�����f�0���O���y�X��E���^Jn���1c~6'�������]�
􉳱�,�� 4���b;e�K���۲�(F[ˡ!�����I��I�4�:�����"	�*?P��{�F�C!u9�c������xR�lVG�I���r'cS~:�/��6.H�䳞`�2Y׈ '�?e":\+�WX��Z�5�_@�G�^P�����ـ`1�I�+�I����Vq[}t̓gU�tq4�Z��ES\�)o���Bf�L�|���dY��/b�#>u�h%�l��Vy�fZ�pS�E� Yu�bbO�=j�����aҠ��T���7�d���۬�O�ϛ�<F�
&�,��9Q��z�]��۩��-\��ƛp%�l_����z��F,�uh;[��7��c�4��.�ٚ���"������q���8�J�����H��v��`���Q]��ם'�0tjy�_ݞ`"���!��j���|� �*���:	cő�(�tj�m���3}ܷ�jg?s���~YZ���X^KRL����G!��7J�z��v#�s�p&il����b��рy�AԖՔ2����I�-�;���]L9���ʢÇ�J ���}��3�/��9Y-�1T_,�^���_�w�~�v�2�2ņ·�%��,H80ôU2Y%��u�~Z��>瘎y;���wO�(;��mkKJ�<A�	�T9+OO{=C&|[�|p�{B
�[�@��2Y#�
�op���q��2�Ap��Y�11�b�`����Req���j���G*IYvr��]Y8K��� �J@;���1�D����ݠi�3�9z6�2+�'U��S~���ִp۾1"M�
�.�B�b���m�f�4<�3?k%��R�ek
�$�;�ǣ� ������`@�Q��y�[�$ jN
�s��S�:�?e�����2�_h���3�)2�߹y��n�<���QI��
��j����q����uM�끱uO��˹�c�2
��@���ӂ��A�Cd��k�'��Nt�fm���B$2�%$X��T�f�yqO�ӪJ����g��^�޹`����%���vr�PI��:WW�l�0��.�l���Ռ��n�$F��ǡ\࿝>Fn�3���"M���Aao�E�v��2=�D�TuV�щ?BL!W8*������ F5���[���yT�
ƃ9{����A�=� �~9���D=�9v�F��/p��9>�L󸦎�~�^O� �	����
���쏍V|���Lyh:G.S}�⸫�"���p5�:�G��2 ���|[�E��,�Ţ���Z�:!1�Fd�(�����D�m��zG���0���s�	�p������ê��2��[�Ui�䤟��L�%Ʌ�� !�_�87�]��^�u�Z�XѬ�[�*!�Eg7f�6���f���A�Nj V:��C�-�����L̛_\s�R���(���7���o^)���z��Y3ŷ.lSq����U,5}i�0����j���&�s�rl�	G}�^?���#z!����H��B�(���^��y���57IE�.bd�@KNi�å�)�l�a��,�\�oI����̭�Y�3$XқN<Q�D�vS�ţsBf�	f����/7��{�*pO���I�U��W��♕^٘&��b�z��$�L����DJ>�K)�m��ڤ���m«��K��]Qp�8�SX'����Q���/�;�<��Q��Gt�u�n�q�K�n����s�g4��พa>F"D��&38%�ȯ���XR�sR���*�+v�Y���&rW����7��M���d�C�}���O�<��{Sv�����߲�G�E�$��̢;���B���b�,Ӄ���_���(��Y�J`�%Iڮ���2�����`$�h)�JE{b�P�hC�y/��ȯH+�apb2%K�]�h}�R��"y��L���|Ǒ-漂*8�ë��A�_��(��O�d�Փ����v:6�6�/|�-f�ӫiE�y��o -�����&P~�d�!�l�8X��V�Ї���NoP����Ο�I��D�*�x�)�!��ЋK�׽���"w�s9FK^ X})lM�s� ��Ln�UVB2YV��W/2Mz��G1���e��5,�%�����*�YQqR[FMQD�}*�ȁW|i*�b�uyP��*�BzT��R&V�`�b�8>�ҙ�t���� �Ix	o�̘cZ0x�0K{�lHb�苕Κ7+҆r�Kw
԰=_lI�$52
�l3!��6��e�bL��*�d��9LH!r�{҈�Q�#��r�Yl��$A]��b��D�@�b�����<�7D�E�Ob���"ȣFƪN���j�N�����纠3���-�m�~�g��1�_��2�O7S�^�,��딤Aw������x�A��K�����RV�P��=�,ף:�p?�rF|R�ɺ�*y[�lW.S�-H6���9W���޿�#K�\��c��s���p��I���e+w�9��:S��?�H���^[&R��Ó<��k^0��q�s�Z~|zbD'����4ČLwoN���2��q�<��8 ��Ci�(�X1w�Pr�md����dmn���x��G�%�*[@ܲ�?���Ω+:�<�]F�Q���]�ƻ]�8� ޻��Ss�Q�D�ԠBQRC�[���Hl�޲}.�N�^X�z�D�>��_���DV�?r�N��D��
gp~��TEG�^��� � #Pg&X��ɬD?J�,�P��п2@��4�ۦ�p��}���������
��_P�چ�܆9 c�Zl]��(�����n��#�H�Jv���%��;����Fq���L���U\ʹ�q�`i��v���C(���T��&��y���N8����)����t6�M�P�0+"O��[��[�R�T6��kK�s��\G�>�*&�j����Ij��>2�\�7qN�8b�[F��{,��K\��R��J)����?8"�׳��9����	��$�wI������=����>.��s��fG���������tʙz7M�8+o`tj.$E�hs�<����󕚪�A�}�u�htySf�BU�0�7�Bv���K���9��u��G��91�<G����(D>�,��~�gz�.xCU��ʽ�~F�rѐ�(|��wl�������bL�M�l�l��D����u�:s��g�~ee�~�gz6�pâE� U��!0I�����A���lc�9���ؖ-6<��S��ϰ�3�Ǫcs^���W�u�K��O};����VDm4��a�HP�wM3 F@3UAwV�%�旫t|��0)Fͪ���͎=����0�d�[,��d
p��AE�V�*�͜�$K�f�ž�@Q�Z�.�2�k
��ڭ:�\ȍ&$�y��Z/<�����$��ޗ�J���K��7��{4��Oo#%݁��m���S�W�N�Ւ��dNz�*��FW�����ǊQ'X52���Itķ��JB���H	 ���ILO�Y�=Ł�|�*�)lK9��nW}jf"�
������f��(H�?��T�wB g�f�aK�X�Pû�~���n1V&~A��BR����Kcc)�K�]i-C[n�����H{B�s�ѿV�I;�?�~ 7��W�My�
�I)6ӄ� ��tt�Wc�uĲ�@-v�`ߋg������e�醯9l�Q��\�u_{�nc �|��+����p7v��3¤��#���; �#�=9"�iq�2�n?ct
4=pFr �$���U�M� C��ɀ�!��a�ʷi�3o#�߫.�:�tph�����;PC_6�{�D�u���ý�o$A�c�}������C]�nZ�_�y����ud�&�Y4�IIq}�hR��*-�>]�[i��8;��q�z�����f~~������h�հ'���Y�Cg*��.�u!��^ ӧ�PL��������E%S��MܵN�j�`�h;%]�\�#[a�ƹb���Y`i�z0�	�Bj��plq��t�]��:Ttp&��#���lf�F0N38@.�і5$����~A}\N���m����G�9�8�����9V������a�v~8<C!�E��\~n�����<�0I���@���p}D<dA�IU��L��#q�톃���y�ԵK̤
7�c8X���G�`�J�= )�_��	-�&Ԫ��ɲ��s,��S^�LK�-� r��f:��/���4�	���:��w�7��ۙ��hE����ꦾ|	���T�Oϫ]zIZej��oY�����mL�BHJsb��P':k-���.�/����8Ŕ���:k���2=V����d{�-�����Q���* "��4����\�Y-h�ԣޖ�o��C
u��W��>:������@gPH{��#JS�5�n�KKk׎��O^�s[���%{��-jCO(3*�	?�����������v� E�#f�ów��۟�]P#N	>Q���m�f�ҟ���B�5�{�a�& X���a�{���R���R��Cv���1��(~���{��/�#ݮh�]�z�_�K#B�z��d�멨�c�#n^�R�rp3<�m���6�0���(�� ��B�߃�3g��h��8�9r�*���c��^��Ez
MYu���Ns`Xǅ�Ns3$he���qi(��y��!cd��@&1';_.WKYR�(������s���|�7������u�\�'d;q*B���1!�s��>[�i,���"ǡ�I+s%�^�8�%��8��W����h�9�'���P9t��Б>��tx�S+/At���q���0����淕��T-��E�Y܀�@�U�#Z���	y:�ճ���<�ì��%e2-�
�� �%E�p)�7����L�z����r��:�0�#��<e��>�H�we���j����x�t´@�¶���������Ĕl����܉E;q�o��?���v���p��ኄ.������IŻ��8Bh?��0g��eȾŋ��w �GgE
W{�@t4.�(!.zŐ�shP��{-*��v1; ј.��1ɥ(��� 3��H�����oU�?��Z1o\�V�:Ax��3�����Tظ�^t-����w|׻�����y��U������c�`}�]�r����^�BU6U��z�]#��?^ A�U��9?��6��]]���[��r�^���y����n�	�Gp�+��9��	���D	�,U�p�E����{"�W�u,��.oԤQ�72A�|����1⟮�k�� �|� �U<U�T�x�pzdaܵv�gCA�K�[]i!�CBy��$a�v�`F-��x�,�t��sG����5�p�o�x�#�['U&-2N৆�y����E��8o��m��f�r���_R���%�٣�z?��3�9:��E�+y���Gw����l�]sK����|�İ��������P���9�'�+�@�9��(�К�L�2Ks2Q��9!l��;�Q��w��PR.�� l�͎���i��)�jӊlal-^�l6E3�EM����S��:�ll�24��v�BQ����/m5�j��g.�U��vMv[��Ӕ^
�����1����t�ȟ���)MC��\"˥Xn�E�b�3��.��R��=Qm�R��;M=^`�s�[��h.=�[��o���5ޖ� J۵��	���
i��>h8�����N�������]r蚓������ 1|�M��u'�Ӑ��`������"c�W^�z��+'�Zl�zN��k�UN���w( ��h��d-��e�U~{��G�����D���h�^Qf�ێU����<<��ysS<�L9�W>d?TU�����(��}���z%ϑ.�>$���~�,��M�TP�Hx�W-c��r�u���;^�î��|�yk�`8�(H�5E����1�����?�G�EX6O��{����[�����T8q�/���2��w�[�X{����E-�~d��7+�c��؃ ���Y�	nͲ\Z;ָ��M3 ���r�a|��co�wٷ�F�{K����T�J��4r�#}R���0b��^.0�*-��0�X]'��\vB���z�~���dulwu��*:7��i�u(�,nG�ԧ{4ՃM�<�m�RB��Il�0Q���)�89����ݶ��"�)���7��&+16���3�~:���Enqx-�/�A���VN	���弆��c䗦Υ�d��H��5j΢V����^��8v������\;�Z�)
l*.ƻ�?ٳ���x&V�1o1���SvÖ�U������\J�������)��9v��@�n�-�b�}62�O��I��A9N�3A���'A9)�c���A�|m��l".F2:o>���ܗL��+8�Z[n�v�J�� x]$>gG�V���p�Y%�M7��1���ŃF|m���SΧ��)��������3�,����fN&W�����;A��=����0�u_E���V�F'�=� �/�l��l�Z�~{��@0��!A'��ep�7�8p �[�R<����^}}�Kl&�<�O�NlN3A�t��SjؒT@���� �G �_*���E��i�!T�W���C.���=�v�0�!�q0ҽ�!n�M�p*�� ��B�	�x��6A�f�����pRI:-�#B$nY*���E�Dr#:�w��Oޗ �%j
��賫��`�l������Lx�47��$PL��C<V
1�����~^�Mz�p��"ҧ���g��m��W���-b�����m?��c�v�Y��rKhD�ƿm��X#�E����(p�������a��i��?�G���#m�(E`����9�N��L�`���K��!��Rz[?���T ,h�U1E��WRF6�֜� 6K�_4�fl�bY����l�ܲl���6uؚ�^�"ı�piV7q-ڻ`�Ua����A��V+m�䍹�Zk����M���r�-���3UB���7�M7O����"�	£T��_Ƨlq��� ��y�w��z7Ȩc?|IT��!<�q�B'�CZ\�`�zșuO��e�{P�z"4}�6׀�G�y�(ê�>���1F�O�I� �!�}�%v~�I��ew�bA;`o*{����AJ�����{���@�\J��K�5f������K�Gqo�
[���%bF���Ma��ܳ[�ı��X`!yA|D�t$ $�+��R��,�n8q�}�j�,�*<$���W\DP48ӛ�Z����\�5���'������kj�HDJ��-�`s-�0�#�Sg z�|�#!��&�[��{���4�r��%�k'e�+�-��%�e��/�U�Z(���3���3"iG�U[�Co�s�#��>Q;A���^Y�㽨<5�#6<��r\���':�S]��8mv�Ϝ-/;ǴPe`�q􀌭f=M΅�	)��GGV��+�|�ߠ�ID��x��l��U���KpI*��{��J#�M���u���Yg�]�h� R���~*��2�z_��� ��P�2��ù�>	���hf��-P�a�]�j��~�7�O��u�^�)f�"V�(5}NXM�[��h�}��1J�
������r+׷W�
!u�쬵r%h�ȑ�@��r�U:�ޠ��Ν�]����]�s��2ۥ| �@��&���J�@��K�&�􋆜�V�7���F<���_�[�fb�	�MEثm�=W�	��$m�� H�Ч��.e�i�_��j}�)��H�`�f�3#�M8+����WI�O6#�p����vS�����x>�O��'��I,�%�0HO�cޢ6��ی�������%��&����F�6�2#��h�0B���	o�q���n[7~�ׄl��!���w��+������ς����>P�̦M��m�~\�0;�[�I�o���k�1G�*�|��4ʃ!jǬ���K�����l�A)�Iq���H���q�&?i���-*���օnem|@����1�Ep4Ldd����խ
j��r9����B��`4vX�"}>�C�!.p�<��nn��;��Ҏ8��I<*��˅-�A�J�Է�\[Ɩ�����/�⿢$�x�d��L����I�������ʳ��C��y�>1��
�Kf�+T_)b�C�>ƽ����W������&�ʤ@���3FMb�����ʊ�
/ ծ�59wi����I��p���wKc�mL��z��Y����/��U���� U{��>�]m�>S;n��l�x��޾r�$�Vm��z8k݇�9J�3΢L{\����
���]^~��H����Hč�gC��"g��r-�qn;�\g�i�f�x�1�C���j���W=(�e��!0���9eyM��t��؝S*���-<`I0�/��P,���ٿ�wfp�rd����UfB�>��ia�>-䧻.��?
Cey�J�+k�&.����J���������F��Z50�zгF����A�e�A��73A-(�<9J��A%���ڹ���R�&��k��q)�Atە������.=�D;X	P�TC�nd�3j��,"�Nb5�x{t�z��G�(>�m�����VlPT�jܼ�V��R&r���,�k���������;|��C���d,�ْ��}qO��^:I�z�Q_���U�:!մA��\>�Ҷ�-��Ox/_r��U���zJ E��V��60ɋ_�%G&�6|Hg�UW>ձdl�c�A����>�0�:˅�%'���k���q�����S�W�D_	.��U�?b��ֹ5ܧ>k{�a��2�ׁ�K���'s�HX7z��|*#䲮M�=c�qؓ	���\���N��}�y|P4�H��O8��������b� ��~y��n{���w�� ��^ �ńb:8���q�u1	�M��Ѧ|�t��̊3#o��2���@����]��u��Ȩ���X;L��Q�Q"��A��M��Z"˳2��o,�`��:/G��|pGpi$*��l�����5��Y��Q�+��I��	{��$�*�+����vꨌ"7��\�,�~]�j ����M���>���32B�iln���S[O��I'nD��KN~�ز�<S����݅����y#o~5>�O���Ow�r� Rp"��SΎ���S����hu�GF�?F>��,��g!u��W�KC/ ~�Ԗ�*A�I�r�����T�{�w���#qԡ[P�k��
�%��|5��ޤP��%0e�5"}�D���K,�9�7C����e�j��t~�\�
��l�h�ͯ,��i�.-��$�i�G�G���y,&w~H]�G����Ir�J����Z�櫗"Z�O��"��JT���}�\1M!`c��R�,�-C(�քpk��G��/+ԯH�$G�Й �BY�����U	x=��5E��a�h�o ��)R:�޾��|��̤��M�9FB�j�S`q&.,eh�����&�E���6l�4�����'���>��g�jk#	8q�)��<9/�|p��������!��n<�`�bE�(���^ ���zh������[ɻ��-��<��D�2#���@R���� R�Z�r-t��B����f6-�:�vA���<�%I@O��]ZV�����;��e�_�":�	x�W���u�G���9Oͣ���/~\~�Y�7|| �:F4q�}�+�����0
���l}�.+�\���|�a�
:��G�X1�\nw�A��e�X�j8��r�P���Ǥ�[E@���F��tf��kh��)��H?D?hD+�gbПœ�"����l4S`dXZ�q4���1]$	ڲSY���-gR.��V@��M$u��Oԕk�6JD���5�{L�+l��>�$̱��C�y5����B�Z(b���^�*Qu�L��SF��EI��j�E���o ��*�
2#"찄��^i��n�?��'�W���U(�	�_G�oo]�n�q��-�Ke�K���w���c�ZH=��!Q9ӗ'����S+���,���'�^�A��s�K<�0�3���Sα�k�#�&�A�I�b��:�$3a?����S�l�2��S�9`�/���Ki�켙���̕�oM��OY�6�an��[�a��p5b�^K*|Ḵj�|�s��b��"m�O�+�$��LF���U���x�����IH�.��6��3H����K�6��V�[�	�kG�"Яg�wZ��H�WIs�P�~�^� �V��x*]pOm����͛ƌ�hm�x�DyfG�Q1"��[��"���7!/r����z��#��6�YFC���&�A���CϾK,c��Q��~R���w���D��pQ�?`�RR����#��Ks�Y�?,7��L�ޔ���7�x�(H�s�G���~��-Ց�w�?I� �J_�li�3m���*�����-���YLz�)�y�6�'���~� �\�j�OP���euRB�b���s�|���zm�W��x�Ǐ���)���(���[*����Vb�*�M��`"M1��ch]��>����x�ąY5�`V���R �:���~O�M_��������Z� �c����C���*��*��(MI�����Mӏ̆D�<3�������]�v:��)7�6�т�	hY��u=������HTd���'S���^.V+��jL�u�