��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�P�;�{��3�OT����n/\�@���V�F�	G�V��]� z�`t���y[q����a2��;��i�t��,-��1�� pz�jI;�"<i����#{���<�G�N�3�mŬ�#�:����(U-6��K��j�'��Y�}'	T�(L��ag�=���`m%5�|Nq�Y;�:�|���Q@Y遀 ץ1X�q��j�%|�H�����la�IKA�w��H�=0z �y���Ʀ#��au��#E*��p��c��>�$0i8Y=�P���(�]hϽ�8��1���y���*��V]�t����śvrs�C��G��d@�GZXU�P)��n��>(٩�P�u�?P��xo�NmpC(\�ժ��W[�c����L��1�h�$QֻH�RgM�3-�~�U�S���m~b����/����1VQ� =���\�~����\F!I����
xjo��Ƕj8K�3��O5#�$����x�����U<#��2boc��s��J�H�Sxp����E�Ѵ��"�T��I�f�EA�Fc>�`ʡh�����>���BW撒�MlH!;q�Cf�SS������2��j�ݔ��mF��Bm�����3O#�:��|Й�l�D��|%��⾿vJ6�e|y�"����q��#b-
���BK�� �3��E����"�*E�^I,��Q�4Y�ŧ���}
lTIs$���a0ݍ�ni\|xUiKP]`����_��*Q
DW�L3,����7a˯H��eKi�_�Q _�4ND'K׽	�iR�C)f���,A�-�Y����4>5<�*�-j��tYB�T=ot*7 �pz�>�"�pv�V�¼a��@���o��}~���s'�����p��-�����F�eU�S}&�~b.(�����7`���ODp$���c�a�f| �Aqa�/�����Z�ܻ��_'G�,�YH���+C�i|B��H]ψÙ��<vӭ��$��4�q���ֽG8���? 9�!߰Z���N�;�ϖ���3� ξtS����x�r����E�!xѮ<�� ��]��s�>+À�w��=t�Aw`�$�]��h���m���=�~���'O0>���v���C��M�����󢓾h�䭡�����b�����_TK�C&-Jty;]���ش�Ū3���~���j@ Mu��X�4ۆ%]C%M�kݧv�:����?$ ��;������G����TZC��ys)6Q�I�64��?���)�t�	��i�ڊ�q��AzDB����ΣMlrf�DS-kª��ݢ" мm| �8|�Z�Qn9o��4��$:�Q7*����f� 8qqtO�y���fm?�9x��Q{���q2��W��C*IӇ���m�C@�r#��3u>�;)������wm���g>�mzj��b���h�9�����c�fͷ�`)�����'
��Y6 ��p�;�@��k=�102^�<����z�8:��ڬ�ll�&���A\�$>fTU�nW6#���ƅ�-[M� ��o�\�Ծ�x��y8vA�c�.m}�jy�2��N��b�݆�/���Iծ��7c�h�L����Ɵ{���g+�ϕx-���Z@��3�k��ؕkG��~�i�ul0�� 6��P㊣
����V��s���3�q�y��6�C�M;�u"1� �.����J:��H�i��fq��9\�Dr'�U�ĵ!���DF
 ��N�@h%���3��D5��sr�;�,Qϲ2v�-�6���X�̲ݗ�!S)��}�cfጩ�F�(.�}�,Ҩk_��=���\$��d�x�
��oq��{��K���6;}����h���L�PdJHH��*m��9��:`�4v�7�r�W�� �Z��޷�4� \��gLk>y����L֊��z\�Ȼࠑ��9�ޫ������/��ˈ��z�a0b�O!+"��g��2eQ22���w�Uᮾ��#���W}��-zpQ�6�ݳhT!*a ���@���750��ԭ�5]��� !&M*,���n
RK���n��G�冮�VƓ����������Yn�&��oZz^�Rzvi����hw�������5�3?tEe޿}�!���u�Y�*Cv�+�OL�Qnќc�0�X�*�N��l^G��ȑl� �_�#W��@�K�1���Vx�A�wl�E��*\@�
g�<��&'��E< \�*"��F̊$߀L��>k�1M�o��N$`�_B��=�<��RS�11��2/Iu	���p��� ���\��Ȝ25+e�/���������B�gq�����г\��I���1�/��8�:�F�p�৽��!��؞�����fGq���~y[�V�?n����|*R��;&`!Qk�V��hs� �T��k	j����A	�|��?�| ^�ӷ��LA?�uN2/T��N$�'m�{�ׅ:. ��ܕ%�y�����z)����.Ub0�XO�9�Ȉ���`�@sv��G��gFr:6�W��L�|��멥�d12�湙-%�ViŐ8�Ps�7�TF�����>{kU~c�(Qx��N�<�S(�^p��ua��M4�K�*�j+�1�	`Y	����[cQ���,��G��dv2�%ZG
Y�k1��IZ+P�LU��J����H|2�o漂������LOt;�(2"Ȥk�c���|�RsaLAv�tQyV7�ŭՃ�^����b��#�rR`�n/q�q�F5��������>_��6�(~D.7�|��
J8LB��rvcJ�1|��h�:�l��I�y��r�d��c1����=C�a���U)����n��P�H69Q��=�.$616�	�Ґ�Z]wNl���,➨�2�N������]��i�^	�QU�kD}�����59(��ں)���X�=�_��M��r���I�ָY��m[�q�<�lS�P�S12{�Ҿ gBE��u��aԐ��/7<�0��qf`p��x�!`�������spI��t�R�^L�|��ه�6c�jJ�(.�X@esx{�dڵn��l Xx���2���ZF&�\�C�.�.�P� ���A� �C�LÅڨvYy��<���&C���>�1��"�����w�b�L�f�h��1R��dC)��>#�^E�o��#uꍎݏ�=�P�|�Y9��qһ�p�]i�@�[	�n�\[..I�.4�S؜x)��X8\6�9L)����YGAwC����O�q��R���nM~^�(���Yw���n��g�#�A��T���dZ��T��U���O)b| 	�]���.K������	��F�w�n�%�	\@|;�8���U'Q�v�Z����P�����R@��%����Zi~�@��ȡP@��=��ַn�U�풕��?����ח��j' ��p���N�6PG����/�Ë�x�A�J[ 1��lV*\W%� ԙ�?l�e��e��4o�Q���T���C!}��9-�\}�#(q�/�����dθ'��?�]����W#����Ǚ+���/�uss�o���I-�Ui�N��^����Ѡ��Mu-FR�\k�(���F�_ z�����5ʲ�����}�Q�<w�BY�`���������Vs4�j��"�����L�`��2�L�۞t���\
�.�A��{�Lc�&�0�l�&u��ݾ����򮿃�_�`3c�]��x�[H=�L�����w���9e0w�Ǵ����ꯣ
��?q�]7a%��8"���:�vO�����B8�t7�r�H����?�i���!l�(���mqT/�D�%/v�����y��ʦք����L2o����Al�Q8�0�-��<1�UmB����a�w]jA�d�;�:�l�����'�,a�^ib�Q�\1���� ay���	dUZ:f���a��D�BWrP�<����������֭�y��c��G�ˣ��J[��T�r�ʗN�/�Q|;˽I��E�ly���B��|����� �A�6�Z�>��Y�0�k�<�'��p�1�\�:�3-���˰A������$Mh�ɨ�7�c�:�Nw����PA�ꁁރ�S��X =z'|3C��3�0�K��&8�V')½ Y(֏���1���E�\�I,%�}7@�����JpB�'K����ΖYL^��k٩#�^�NhI ]�v=��5������d41�u��2Cbrd/�d��@��si1yN�O(���&�UO�$F^�r�r7��~vݍ^GА:6��oW�Q�K��)�1Tݕ���.a���)�dy��k��-�8�`G�V�v����qN�$�Ĕ!<a��Q#��kO%���2ּ��"��_F��T�Ae^-7 �Ma.�8J�p~-�q���gVYaD8l��}��C)�5u�����v�Rc�o��gc���k�єm%43�T�쎺���Ix��`�ϪJ�U���m#hc��������o��4O j���u�5a�����E��o[4!�X*��>�,_�V�&Q�,=*\����_�4r�_�g�U�V��"�+�c�Gݍ����Dlf�}����J4f��� o���p}�!ӧ��-K�d���f�4gӜq���Ǽ��s�Pꭤ8ϣ6ewi2�ʺ�_�۽���u,x&�}�ӈ�XEC^�qu90ʤ��|V��B0 _w�t�7� ;�@j������ˀ��?�C���Xݢv�v�9��i��[�}+'Dj4���UȒ�9Z���r�Keb�9(5�:����\:w�NU>�1|C�D\~��50>>t��D`)~d6���T�#�!%���Ős-Շ��MAs�����w��hs���_�6�\�.��ʣ��p �b��Q�׊TX�~{V���y��l9E֒"��9���d�UoOޔ�<I����vF�߽�2?*_�R5�M�P�.C��SfΒ��;�%�g��7��"�,,u[0��{��e9T��d�)=rs�"P�OJD��e������H_�| f��"-5VT�4f~���z�\���]A�!߉k'R�N��������e(�V��c	z
�+dS�s��M�q/�7V�Noy��_��"u����:�m�@���E�F�nR��J�5R J��S�9w�X��G��Q7��o��7�0~ ����k=�0v�����������UF�~�[��n< F;�sz���ʼ��	����Y���~7v�ټ��+���<(�z�&�1���tn���JFoi�{�lb��N Þ`&T��[�� ��Тc�k(
(�U����*������r��r�/g	��ܰV�e�Zٷ���`�~���M�����M����z��w�JE�G�*�b�~9��Q6#n�
�Ѓ��&����	,�FN�L(еHe�2���f�Y��N�*e�Їǟ�b	A{ݣ���k����F�M�Ε�`�и9M��V�x�"���:��3>��F�Y����8�6(�Pj�F��B�Y�I�Q>ך���ۭ�C���Kj�h�uWŹ����rO8�W#t�l>�e|���\�ZG���<hXGP��%��D����I-j)��vԶ:��(|����,pO��M����e�����f�F#�P���w3�h7�\�a�
��S����i��P`ZD�e��"?�X	��>�,�\���{z�H�#��H񾦀)S�B��A�TH<��e+Z	je���t��|qA�37�O�YЗ9��W��F�:�I�>�9P�����[rM�𝁇���5�XĽgR�+q®S����FŃ���]IA$�Z�az�*�
sz�ک�/�ݱ�����ا���G�D���=_O��x����g	���Qe�Y��Y���hU��ai��k������/��Dj떒1=��{��*�x���沋����$�K��I�$�I/�ۏ�@w0%�<\�)O����`�T]]�T�v��m�|QY5ٺ� iy�9�Lu������!�+�ܹ�'w����{-�: ,k��4K�xT���|+⍭ޠg%��K���B&�h�S�*q�W\Wd�fZ�OQ�HD��)�=���p��Ri=<��La�I�+|3/�mW��pj\鯓5 S.F<k���JJT@(e�?��j�í�C<��fi�>鉽�� zE�iJ����
�y��qJ��1r��|.���w�����ϳ����g$��|A�V��� ���,TO'����_�Y}�	C��ro����΀��6��?��+�Խ�I%�V�m~?4[��bw�{Δ�Zsw��!N�7Yi����L8�d�ӗ����OA�~$U��X��L�O�V�W��sd5txX�8�4yso���}�,��:�DN3L���U�c����Ѧ�	�������;ș>�pZ��y�B �Qb��������n��lq7V���Sl�p��|k/�>�;�:ߎN�� l<��Dُ���s��s�A\Q$�]w)�
yg1kj��|�&
W�A�4�!�%�H�,# k�)�ى3 P���a�O�ϾM3z���-��y����;t�;�I�9�.4t�s�e�A���7��� ���"��26s^�ʆ*�u��i]��U��uQ�g�l���v�*al�ZO�,4l����(V�u��0��ut)-#�&��������tD:{c���&�Yj2�WF᫙� �^`i"0�B�2�+g�'G	M���2�cO�)�82�>.�W�fz&�q�.��a� ���P�EC���WQ,�J�i�_(��1��R
#X'�T&����AK����/���h�+�[��F̞%vc� �n��y��f�^�q���ޒ-z�l]�B�oo
Վ�\}���.�c>���㡈p�Tӯ���㱷eP=Q������]�>6��&Aue��s��?��EG+�c�����D���bG
,����ܩ�p^W�F�m�����\�7=��X.L���V/mj���c�*���r�Nrz'"�>��q��@��LU	��d���<��Z:y���
��kݒ�B��W+&Gއ�,"�$oN�\{�X.��Y �]4*��p� fK�' �%]U8+,����)2�� "�UY�=��Ub���Z�	�1�̴�I�1{���w�ai�o?O��Or$n������T ��>8|.( �y�5�BQ��8tDR'�մ���?���%�Z�3h��#�����McHj�G��w�8� X�]���X��㋮Y�;G�`{�_�z���A�^�׵r��u�T�M�9b��Z�O��L�������vP���-�q8���S�(��p�/�����BC����A�Ѕ�o� ���{�~��ș��Η�9��˘e_��������Z�v��mӝ�Ȼ�����5�ωA���PT�.��S�0�gY��9�t0|I1�vTTJ��B��y�����ʀu��%YLek�>�UA]F�[2�F*�m���.���E*r�$q�v�C�N_���R� ?������R���x�D� �8{C��������~w�>�C��
���y�(���Ʋ�\�z��� X�g���{W�\c%lI s��]�Dq ��]ϵٺ1;�x��_��UR�R�x��v���l�K~c���#Js[��h=��w'l��>�j�m�m\e~�/�d��о!�۱	e��m�?����Lj�_�X*�ED�2DHI_�������NV*���8����+D۱}Ǳ�|�Vx�i:�:�}�{Q
�K�v}\.��DK���`��Q����.�d8���~��Ê^Z��}������0�7agC,�<u������ݬ$�Gk�Z1��0"���c�!.�ZRW{��1P�.��̉���v��4�x��g�.&�5~��_�C��H� �r��'��̰�Be���D����-D.����9���΃�����K�2��� /��ϫ�V������ZH�d��ɢ�ϪnC4�9�q#�J���AU�4&,O�'5���Y�,��]�3���~�����Q4��eB� )P͡�P��w���`zg�_�?���.�,-�����Uʯ�ך�y#A�x�g
��]�X����={pY��1g�@Y�c8�~� :���x�ދ�:W6&�N�h��E�#
�E"P����+�����`��WN6e���߽�hڎ����� �8@����?躒|�bִ����6�2@���I���n**�I�ZGns��3�z���<�B�}�%�DJ�Y�99�3����1��R� �*Z�67n#�e}����Q�ܚ���N�,1�&�#���;�
��2���<ػo�EB�e��\DA��/�WO�P�E��:��=n�i����^�H�B�s6
���Q����z[AO��Z6�0���1f�|��|?�ᠯa�D)
6�`���X}+���o�A�3���>���ѲV��g�;rj�i$<b�cN ��Sn+���	4I�}�Ww�^GVNQ�B�!Ļ:r-�4#�K��JF=�	�����1=�s�S�~V�� qZu:-ٵ �!��i�Ez��;<%V'ǹ�m���08�7o�T1����c��J?�4��0Kt0��[�_S�^�H�ҷ��[`ۈ�c��[����[=���-B��wSz.�#�+=�w�Z��mی0��G�heǯ� ���\�2	q�(f`��:����ؑ���5C$���n�h���-	\{7��V%��x�*�k��;D[A?�i	9hi��+�����O�2��~�^3���IL
P͠X��,e�<�O�B�!uv
]�_?��J>���Z�q��`�y��*�
ݹ�Yw�}6q��HpR
ݢ?��AEm�'�',��rB_��I�@3lO׍���N�*�gM�G���N`J3H5�׈�g��G�N��K8U& ��f��� �޴YG��@Hs��X3!#�ٰ�� 	�����oFJq��p��vu���(��^��R������wAF����m�<W��KcS`�ZLw)7���B���ݒ��Z�v�x�5 ���X�db��:QXo����f2��Z������W�(���u���(���)�fH����Lz|7#@)L����xa�|��`IN#���vn�ָ���g���*)�նn���P��<�k��}�}�s��e%(~��r���8	���6�=਄?<���I�ުOD	�g/&͟R�p�0�7i��7���?��A�}Vc�3�����0"@V�@�o4��"Y�Xwj꒽�"BK��Ka����( ��v��V�[�a}��]�.�y�!��3�<J����כ�KX����T�g�y�-��q�q��'��:�/��_�0��Ŭ:4\�Ř�
/�a�ݮ����^��H��ʌ��_�V�tL��p�����aP���U����_������O����M�����!��F�U���N�v1�j�N�f��
���5�P0p�홺%�ڣ�]>�JK����.����&K��:�,]q���AF��h,�vM�tC2��D%�žy��nQ��x֮��a�������cR��͒�M�D��; ;�rGZ��ݏ�N��l�?|f�_�쓐�fyC4%�{KFC��S���������,L���1(�h��}EĲ��rtP(�|U8.�{��u�����1s�K��p-AaK�Q���G�ꎷ����MS@xX���*q'��I������uP>J;�
���y��=/��	�f��x�|x��.^̇���8g��3�i���z��<х���C�ݓso������ ��3��q`����Ɇf+�`�5�R{�5%�C�n��|LP���|�̄,$��+fa����sf=�%� Q"�����8��3S�ɍ4���v�ؔ�F��X��i�t��7]fN�Y2 �6��B]x  ���;�.O9���m��=�q�=�f-�]O��f���E�6q�E>���@p@ۺ짎���qFCH�dS�����Y��lf(��$/���h�!�8e͙�Q;��kgmq�=��lj���w�/���Apw�%�(�6�b<K,8�(Vz�^�8�[B9=3�BB�T�}�����_�9�LD���ݽ�4%JJU��M�������FK�%X/E�l$�J��f��e��hڦ�XJ\�_��ɝR�ka˭k���Y�j�0�oHvt�28�.��6��,�Rej����ã�/_�,�<���g�j�x���Q��W���圪mI�+U�g9���`4=�Lq��/��
jjև�pLAQj1���i+��J���^�{�@��F��
���¬监uyo�mI���NӖW��ӧVi�K2�B��bO,P;����u��gy���H�q��L�o&�� %�#]ln����WY�7.Q&����w� ��u�o�I����ɒ�	�X� ���ŀ�D_3�<;�z��Bݱ�(�#J�f�̙�ǹ��ƚ	��d΁`����m�c��3�m��FrfF��={c�L���}�S֚���0]��h:�ޥ�fD�+veg_:E_$�e��kJ�b���v�+ܨ!�0�P�*����*�"���}K�"L֡�Xx���:�4�P]w;�� �Y�L��|�J�⺽�s�ϳ���߅���K�dr�*��Rx�Ih]�B����ڔ j�;q.�����hvO���h}�� �v|~S���h>7�P�x�l���N�r>���lcH��J`>^�0�1�Z����"|�VIeR6��2#��5���7�L�C��<'���!	Jݻ/��"�$�]г�Zo�:�ǖ��1����4��1��=9�Oޔ>����Є�<0����N�����Iu��M��T8�S���>�g�����m]��3m� *��YsC�S�4����<
�������1�Z��n�El2��M��*(�/_ BE���m��9�,����]�����0;��2�g������[e���O�DA|l>Aa"浺~ǵԃ��k�u���V��5�
N�<$2Lx{�����{�O�^v�=��;��>�����Tq
�&�/�����\U*���|�"�|$��EU����Xx�
��2U�ն��I-F=�<�W� ��	�UGR��,�_��@���]�TKm�5��Sfz����-����E\�> x��Q�OD�\7l�n�_b�-Hw
�mt���,�a�׻����*2����'Z�w���P�|4��#�^�R����d��{Q�R!@��{��@X}��0'�7tY��彯=�ދ���>��X�g���1F�}FV��t��Y�m��wV���X�r$cK��
/@ 0\ܰ��Ә�$[`TJ�@�_�p��=�b��PA��#��R
d.�N~��:�F����I�R�F�q��5a�����S� �j�V$ �J�%��sv�1qt�ߖ� V�+f�Ix��=�W��~ѐ|yk���m��f�LVQ�H��V�U��3.�o�0g��8�՛ν���ݾNz3���(���ymx_F�����\K�PrY ����b% ஡�M�=Фu`BӳC���HAR>�6sHe��ɋ?;�eb9N[���1�-�I���,4w�6�l���lA����^�Fr*���Ы���1��
����[?���BE�'���������M��]}�)�5�9��Od�M���7"y�9�\aɵ`Z]��L�o���x���^X�re��O�cふv���G3�x�G�M� z�#
&\|���ӦXX�Jl�
5e�q/ڄ�SЄ���@��ŰG֚["7<��H7O���j���M�mi�9wS=�h����p�u� PY{�n�t������ a<-�1��_�3;�p����\�T��+s�G���t�-����O��|	W�����E���Tߩ���Y=x���	e3^�hГw� G�cr+����Y@�B}�#����J�V�4�S�h�֓���5&�m`�e�',m�R~!όcr&}�e��>\j'�ݦE��ѮL�(���ԛ=K���L-f���o��#,�ƏV*��hf�o�a%��p�H�Z�D�u�������ǡ�)��x��EKvU�xy�������c�o�j�H^�-!̽�j�3ʗ�� F�6���,t��
��C>Zh�m��;&�p3��9VyJ��-���k��A!^�k�эժ��lAo�e�+I��N�J%{��"�����%�+٦lR�����{���T��T(.[�����棬���F ФO����j���+ٯ�"��'KVwJ�)Y��G�*�Wϒ%�%}uw�l�� A�CP��4���5��8�֍E�# ��9E�sX�p|����U�4k�ԯ�YN�Dd �L�c����<�#��٦�y+Ѕ��4cZ ��Q�~�I�NJ�RB*�p��Ƒ甍������a�Nk��[�*O�
~��#��6�?�C���v"�AXk�*0�Q��^&�����{�l�pQ���y��O0�8��Wݜ��R�K�mK�x\�� M�̓��������'kط�A���z�+�9��B\`�"9��^(�#���!�/���H���K̓w8ψ�@�Д���N-ɉ	�+��^�0"���1)z�(N�MN5�s>����(V~��$UK��`���ѭ}J8�^�-��Y��e���nxk%�����YJ{@un�rW>�d�P����ŝ���ku�+��g&�	��|+7Z���A��x��ϙӇ�O��z�a�ƯrD��f�a������$�R$��j�����^l�Gd�&�}W�ՍJ ��߫7�j!ԥ"��<�OV,<��˾�(�!�n��fM ��	��psEOq���ED@��Ӄa��҆��)�T/���j�>�X
��Z��p��w�����{k�o�����tn8!���G��L�i��*_�ί�w,R��G�8�����CJA�fd��crA	-�7�2�߁¹�>V ������q�B
p����ص�U� c�����%h )���G��0�A**���w͍�m3s	~����2�O�DAq��a*�!��q� �l�.e+�p�ֆ�P�(Ɓd�хY��<�b�)��d���5M�^��r���A����$���-�,!&���Z6��*	���i_�*�qX| �Y��,�SrׂM�֮�>��S�����X��-+���&Z�Y���qj^h������_:R%0���X�Ί�X�~�Y�F��zO=�3܍A�wW��C�d��Cy��dh8��o��{a
��g��I�[Z]�5h���
�M�����at���#����HC���U���(�{�)%��$QO����R+�Y����2L��qU�Uf���8�7�I�G)?JO��c�����b%/�?:ш�6e�Dė9a�I�bK��9���mͺ�JS��S������0#`EZ�պ�>�0����N���_+����Wv���r����wH��.��� ���I������3��W�gE��lh"�����w��U��P]Y��Jɶ�/��t2�̞��8�-�!wI��U����m��L��M�5d"[s8:����@HS��hX�(^�ʗ���f3�MnR���E��dp
����\Lh�I��������
�)T�k�x!��m�Di�ץ�F�r��~5_�Z�t���C�cg���e��/Q��d����7�r����*���@w�� V۾��ϒ1J�Q$/�x����oekF��jr妈��E]i����6s��o��pW�c���$����c��w������[�c)B���5������FlG�=?���RWK�/V�rX9�.��N�I}_ڎ�6���ε��POđo�{���9Z'��,�̖��龥h���jR���ßqJ�rBl��6��Gu?icYk������Ms�f�߭�G�H'��Ym&#s[
���9c�i�ež�b<ڍ(\�k�Ѳ nX��&c}*��>���6��j56�f�R���<�@�KC��'ZJ����0op�%@�y75���\9�6z��l��K����	��
�9���jF���Z�G�bێV���K��|ci���)6��c���mkr�|��2���?�t�:e�=���s�@��C�P�L���m�"m�.t06͞����6�>MF��1~Ub6Z�MpE_7P9��h��ɢ;��������Y�Q��
�d��h��;���-[�9�3� %B��A��i���� X�"�,�ڝujo����77_��KB3Kmؘ0��*ܷ�H�P��d�L��ܒP�r�C�r���s��� ���}DX�V�l�̔.��y�*�y.t �zw!�!�co���:�L�玗��I����J��|%'S�BN&������4|�tR��-'����>�
��ˁ�w�� ��ދd_�6o��Y�1Dz-.%t����͵�o�w7G-5^���}C�lH>:��;l�"��'��TDT̋|d_�G�B�tN��;Q����}*f��g��qe�K@\�枹��jP�R�V��kX�g���
u�y|W��C������tu�-:=ZC&kT*%�D𺝬�1l���S�*�Ks>�����A�c����@�䏁(��I�������x% ��f���N��i��L;�"O0V�d��Q7���-Z7�Lp�g�=(:�>��4"S��׿ �D<� �sIB.,�}��S�W�4��\���$_T���/Ǌ�՚ID�\�k�I�Z�h�]E�q<��Ȕ�>�T�K�K@����S%'���ҕ��n6��,��وox�ٚ/�ĝL�ev�iuJBE��L��nI��0Fo��ZU�l�KbU�8[FC�o�ɋ�G�-�-�f�L5P֙��Ʀ"��v'6��*�S���TSMC�aHօ��{���P�����q��A1�$S�3,��
��5�_=>��yd��1�N:+bP�r��L̆T�X��������W�J���PU���������Ȱ]7�\���a/r�j���q���ʺ�!8ɝ����Q;��4���1D�CP�^�f�������-�ũ%��f ybrF����Wm�o2�cr��퐺�6C]�ؐ�4]%��\��?E��������%�餹M�#D߷(�h!v?�z���[���d��ٰrh�����R dhnܠ��H�za��+>o�w+ڤ���VQ�iH+�ltn�&�<-d%�ާ;~d�F��K�� X N�Er�m�ېQ6��*m�����|��:����!��Kw	R� ̺�fzG���r��Vh���KS�xI<�7Ôs�b�%�\;Q��pa�џ������Id/oз[ �78���1F����,�[��tc3���lp�")���C�����m�[�ۉ�⁀sX���t&������@�TI�q�R�x��fr�5*�EƼz�^2"��"�I����>� x�c`�%��C��ȚT����GQ5���N,����E�<kx4&B��D�|�!!��%��8U����衉�|�cyN��`1nH�;2o�A5#�Of�Fid*چ"P�R�_�j$�kz����������̒����#f!�ҏ�k�-�q!�.$���[�DZ���s!k��H�Ŝ�-fR�5�\g;*��>9�pU���'���JvX��w� /g1��Sy�rkLK����QٵNqF���t֑I��V�շ`�c)�X�h>d�S�l�L�2s��y1J�k�~�۲S����� �2��Oq=>"f�o,�&���@��P�K����LQ���(,��"	�v�/��DL�#���MZ��o] ��D�%=@�Q�_�/����L.f
��G�\d��������NK/Đ���#x@̖ݤݬ �8k)b0�r
,�)4qБ%H��H�΢Dl
��GuXʟxٵ�*�H�ٴϨյ��_6ӊV�[�j����C�v�R\�Wׁ���ND���C8O�T��R'�Ǉv�S&��p����w�^�Ќ���dÉ���D�n9$8FA�Y{HV�[a0Zx�6�]fis�R)�jg���|�� j{�st�3�(�G�pOf�'�y�"?����>Q!��pW���@B����c�HښygI�nM5�����r����eb� [�!e�C���W�j�lk����}vJwP{���;9����:��X[���8��?��A�Ɖ �B��+H�0S �C����jM���PR��X��lL��v?^yS=v��S�U��z��(��TD�I��8i�\�/YH۔�m;��&�<��㺨��r������G�0���]r^��Z�ަ,�Z�2I~��`�x�VR�@+>�G���T���=3񑢯��9��8����u���%	_�J*R:%B �4j���W���R���*��U�49 uIRE�Z���c�?�WyƦ?Y��
Я+f�I�1j(T�y�y�ta�TÚw�)d��O�f}0ٱ�8F@�
X�����t��4@�vX��6d!��_5G�0�='��1��o��4�g�GN�.=��L�y\	y��4�z���
G�YtF�^p\U)}��`����RP��#���� \���ݿ&�x�zJ��ME�+Pˠ�F����sd6;��z<�j�'R�������[�Y�:�"��� �F_c��7ʂ�x���!��haO��e�PW��Y�	�pT�Ǹ�3��K�}c><����28�J2J�@�?�?5Z�`�e�h�j�?G�p�]8}�s��OA�?Y)2�7���~��wt[������]�]k&����l�L+��`d2�@\�==9�m@�/�1��8�{��;]�,��@��4"x��̀�,�\��]�ϻ8��J����[������,w�*M��b��S�$�0|�<I݁l�G!�ۼ��J9��%��[�����|>RG.o���w��[К��H/`Y��F��G<j��*�X��{����f@�d�Q1�f��:%�n�(4�>�2<&�tS��=b�a����b t�9�� 9�����m�
�Jk<�����rr�/�U��]��S4��i��������!:��Y� ��h2.���"��������tp1�s<�X7���@!йTgZ�'n�,��� ���or���k���y'Yc
�⍫��<7�U���/�w=l6�1����<�A������P�?����ek��^�p� ��E���O�
��r�x�Sa��E��I���b��0��J���e��nn���y�s����f7��4�`a�疉o3���s/�ʁ'�O�DB�V��3gg���R~��R*�ۯZ�
�v�ԇF�Ҧ�����~Y��M+ɞ՝���̒Љ���tP�<��_�e���I ����l��N�5�%_tiDo���&F�tɇ��<R��RoAZ ʘ�G�'��n�V��&!�Y粏nb�t�x*,���C�[�l�s���Я_jK�y!�V;���$�����5�}�Sdt}K�ŭ�mc���h��v:���|������mdmj���?}2A1��V�p��F�9���V�!�~Ğ0�K+!F].�)��;������Q��~d;�c��5F��L{$c��ȍ�J�u-Er�I�����;�W�F2��T�J��L���M���(�0g *�T��_p �ˁ�t�������<>��֐.q����ںn`<3��Q����#�K�y���
2خ5u��"Ue�"�߼-Aތ$�I5�|�i BpD�d��&�cy-?6n9^�"u��g�UX;���p����߈���e���S�QڿUynȝ�f۲�\�A$e�h X�)~����|��=|��R�1OVn�N��@�0b������
�X�z�� k� h�ƿ���	�,ySy���ut챯���\���K�<�kG��ΏCj!-2LG����</�i�Ŵ=� ?��&���i��*o0��v.s�~o����� tgw��fr*��i+9e�j�oB���\�!� Q�� �N��p��'3�i~ıq�n,���^*�?��󊙽�-����%��1^��=`��I�wF2k���z0�L(~Wm*Hg>���ýI�f�6C�"�M��X���IG��Kӊ%��3	J�1*�^�Wi�cK�n��(�A\+���8<��U�\ Uӽ��8�#�J8���,�d����\w��B �]�m%�B#49�S{%��}�Kp�Z��~�S-zP����>6��TRˈ�x1l*��"W�z:�:�u�p�zy�ڦF�|��s�EZ�^�9���O@�L��j�]�Ÿ��Y*�Q��GSu���m��h4R���i��3H���"�J��i�HRx�����vs��$��2s"�%<稉�u��}|�����x
�'�d�U���h�=�[�\�)-̼	��j��f�v��y���N�ٸ��p�Wyvb��E�I��;���٘}b�>�6gyB�B�d�p��t^N?�����ѩ��+��NVP%�~�E�o��J�}�e�89-�$�����E�
bШ~��Y"�.~9���ә];�7�%_8`Cnɰ�6�DncP;Ѳ��,c�ͩ>��0��؇P"��>�}�^��;��� #}���0����J�V9���|��R�<�a�	�S\'4~2�vm���>�w4���?d�T���Sjs����n�O/�@_�\L8q����u|��1^<���F�b�0�����$k؂�P���A�w��&Ux����<�Jj7K�����]��A.�yg�u�Q���O����&�����t��-6���e'h#?L&�Q�l� 2�ۧ&�/�޺����쨞�ߖB�[��� V��d��`��_��?��vL�v*0\��@¯#�p�1~ks9L��ϔ��J�7��c�}6
��e/DK�*��Ÿr����I��f@�sQ�|���a)0ڹ��ޔ�|Z��h��FH�/%��K1��
N��X�z��1ׇ�>�ٽp��ۢ�k���޽.�)KI呴f��{[�;l\�V ���֩�@}h}&P���/���}���������nw����#VZ
)�f�W��zd����{[��5 Umzx��7W�hL�?A��p8��TZN�{3%�c�s��{���#����k��BW'�k���aE��U�&����weJ.I�d���~-+���@S��{<>��B����x%ǖhE-&��	e�PH?y<"A�Y�"�X:�&g=�g�#}��e<#��ʠ��
r�ث����y�Ɇ	[�JL��@oy�x�n���\��\�h��bY�����rP��ʞT>a���V�gw�-�`�T�7l��}���h/���`�W�f5յC���TAYN�fKU�UY�{�VѬm�",Rjkpy���ȵ
�펯)�����<V�O�@��?�e^�D|��;EKs��F�puk����Ϙj������s==���R)�%P�a��X>(�Ԓ�O����cB-�,�m�I|�?w^��v���7�E�!��y��9�9Qx(�C�x���Ȇ���x�P� tc���~k��ݿ����Zf�>����_Q�r�Y�BɤYbd/��4����?����(ZX��E����������m�)	��vq�6�@�'�"��N��][��V 0{.⁇�O��B�Q	��S���c�"H>������h;� pӸz0�
ⴧ�3酛�Ր��Yp��x:r�3y e��MT�������Hց��;�_\�5���"��������fQ����x���\�l4$0�g�s,���H��G�z���n\���\iC�1n��]�?�"s�}�t�_�Z�j�Ԝ��.XN�\�d����Hz-K{�ݫ�@}�z�f���㎌�?�|���$�[HN��0de�/���F�B:ڙ}Y�����9x�:��\�\�S�B_�HM9��g(B���
�6/zVUmx�|	r�Ĉ�b6���l"R2"�G�"zx�vf�"G��:ٲ�_]�E���T\�x<n��3W(f�R�§� ao�>bs�x�@ �k�d��O7��dL�/�}�ӳ�9�e����Z�Uy$p�3�0[�Ў(��}������a����QT��;���Z`�Kf|�#/Ah'�� ��T���[.��K����Ѹé�x}<o�i�q�Cμ�攂�0�A��&�11�(-洲���[v��/�K�g�j�����)���wǟI���j�~�,�X�:��p.UWD��ù�C�I�l���N:��h���̩�/��;ŭD�!&6�IQL�*�)|�j��T��)"O��k�tl'��J�>��@�JN��JL.Nt��F į��-��j�m{v�5�X����S5�B������_Y<���&��(;�͜��r���X:P6�!=
;�%Fl�X����O���4=1�O��G�������l5�O��z�z��=��a��+3t`�[\�L��"y��'-Y���gDoM/&*_~L�dײ��3F�����)˯�$W+�8np�-}��r;3�}qs]|�����ズ�~�E�j�-���cuL1
��Q ᠅A*�1�r�B2G{��p���*�Qp��V�j��*� �a�����`�O����>�d����!��c�
�����Jkv_4�iͲ��"����nͪi#�QSv��d�x'���54C�Q��@�#H`� ��-���$ `��ʓf�O,�}��v�iZ����\&/���G��܈Z�_oU�%�4�%�|=����4�@�7U�:�R��r����eM'��0L��1>t����e1�I4�M�N��8����Y�Q}Y��PYOR(`��>�
Q�v[����y��B ��z\㬮&�����e��d�����B�!\:��]�o@�1xw�e�	%�BhB\/�����J [�Q��N$����;�s*��	`?<�QA���?���n)u�u��3�t�W����M����H�� �����J�BV�	E��a'{X��n1� �Չ��������h̔?���UpI��S[��UDY�T�p�#��L�ubD��[��ʹ(E�p�֚K��C(�B#4׈ N��C@@s�V��+{����9���a��H|�$Iޥd;������m^o�R$�`qy{��л+���8����u���z\��Sga�Pw{G�.f�-��k�Qx��t׼@�+E�_�_�M�+t���1"Ǥ$�+��<���,�=��ǖ�� �]"��{`3�,��b$}�״���T�JY�ɦD�³�/?���X2a��[�|y�3���r�J��vd1�Sf�>$�4�)4��HV�EW����>B�v�B��>s)")W}�-�����FRXܯG~�3�=���{E�j���W�1��#��.��-�����ag��|,�vg�ϼ]I���,�i�_���0R�|�� ~(�)���M!TQU^yk:��҉@���ƚ����[&�#.�RE��+,�Gۀ/V�8W#c��c���[|�'�"�1�
�>Vp]��x_��~Td�q�?C���N��O�de !ç����Sa��7��yA��u�d�Y>o�o���4D=��Y,�����~ӿ��O���ayR, ]��R���z��{�e/,�~ql���ZG����� ���H]'z�A��}�����0e�E@hk���?�t���%+o�
������caI/dmn�S�q�鿅ЫW?ߵ'�]�ʶv�7���HE{���R�D���&@߅O��'�0�(�Kqyo��{�q.��HR�*��̮�i=�QST�^(��D���l��3�b����bP�%g^T����AO�}�Xts֍F�B͖��(c����N�-H�6��''U~���S0h�[`�j��?Ƨ��`�c0�貘a��T�O�����A��*�:`�;�q�i0��f4���訕H˼ԅD�{u��&���i������>J3�ښ��.�kKx/5ӹ�m���h.�8� �k����X/5}�=U"�-����"1��ҙ�Ma�6�%�(���Y~B$�{�X�2t������lc��=������NX�F᠖ﴚ��;,/>Ŀ�r`/atϥ��6[*Po-.�$�2��0�;�!�[6�J�h:H����� y+H���>�#8���Û�+S2��Z��Q���ۼ,[�rwV����N�E

m�����"�<����6�l�����6��	�*�e:�RYmx7у�U����ޅy���ë�0�$u�t��� ��9ｵ�>��<��*9�����*=yw��7����1������N^D�bj?����@*�U�<R ��Uz��MN��F����I-NQWwh��D��F,����Z��)�x��|�q�o$�$�)A�{oF_�]��m�C�f|$�e��<ʇ\hH��\#��>��l��
��˕�׿GE+Lw�Y|��Rj7�����0��w���*�z�:�xV�y��<Г��E�����pQm�u��,j�am!�QCrq���W@�ʮ�	O��?��_g|�fS(�6�&޹��K�7n�?�m��}/�<�Гn�)¤g<�*��p���/L�
A������f�0���������8Ũ#���|}�r���m�lB�h�)�.��TrO�1[L�^��ש�����/ل?�"2֨1�苠-�<���C
��ig�p�۪�Z�c��*C�=C���s���F.]��#O���s�"�o����J���ˎ*qIF&�&`=8$��Z�����f��9ă����fk|R�1�P�����
���Տ��='�`p��w����ަ�ɣ����:��� d��!9^'����b��m��Ft�(������3�hm�B^�S.����
�������2>�WCN�<:�{�v��@���]4������V�q	����ƂQ�t�U��)����y��ze�5:���/Z�����l��մ��a�K�[�&~,��Y��w�flӻLZ\`yW��1����
��BKL��.�/&7!γ��8ģ��RP���d��/�D]������3H�G��P}��s��b�2\:A�[�6�F?l]���^I�}te������)cՃ�GG}K���I�����c�㙗*R��jy���4�W
R�n����m�h���إ���x���5��|s��I9��|�ԛ��KC�����TD��ӄHp4Y��1��sVԑ�ǹ�ʊ��T�x%��jn�e	v�<�}��*���ݥ�{���A�I�0�1r7�ZAyQ�.�mk(�:Wu�Qe~k�Rj4�	>:�+���;~�K>�O�W�2�!�K����}��	a�|ҩ|4QK�R�*�r���������"xt�$�.;}��Ӯ{�{/]A�����cE���V��� �"�Zq6*0�7�͇#�Z~c�����1���Xy��Jb��H���;0�?JIW	Qr�x�+�m�/���QA_��iϗ�=3[���= N%k�ԥ�[zH�_s�LO���Pp�G�*��Ge��7y�=�w`��	��~���d�.0@_�z!&���<����u��!CF��+�Q������<��^购8�bl���sд6��fB^�I���86��'�{*��zq
�����U��GQ�>sz5��CFg,ه�̀�@U��60N�wzA������t���r�n�� G��!�^��k"�(�8�ٽ�/�M��J�L�K���E]�8�����=O��x�.��:�U�p_`8���c=nQ^Řw-�	��J�%ܡ���5L�_�~��h��8�Mݯ���"�+	��s�[sNu��[8:��i'<u/�K�a[�3/��w�ݜ���J�"^'?��UY�����h�Y{W��H-��Y�	o?X�a��PM090΀Jbi3^	r:<U���9T"���Up;}����c*�Ĭ�CG7��O��[�P���ΰ�;o ���e��l��r�����a���V�(u��i�mz[�@��P�`��Lg��a���@�F��"���#����!�4#,���lɊ��V�)O������d�L�]~	?�֢���/Q��h�"�6���!}��{��X���j��%>�_ª�=��7-��r'L�@��H�Y@N>��sH��,C�=v!J��؁�kK�Hd����1Z���~f�-������{��>��u�Á^,�,Z���}�]$�g�J�Z��:�A\�E���+��=�[�F�ԟR� �8Y t���@y�������Ӯ�h��`|;-`�����_�(�B>-��O/>�^�fgk@c�%��?
bgF��<��!gL��]�ة���Z����>�J|�����o�'1���+&D�ȿ��&5H�b��0�F�#�	��<�@��M��SH���l���B��+��:t��8P��d���pv
\���{�m@���69���k�d���S��9	���=��U�t�tI��_�vX�K�_s��ٝ(B����ޤ����s�)~}Ŵ�!�=���.�5��9w�UO�E�|�f��r�*ĩ�=�a\����qn"y9£U8Z�D��Dvm��L6x�|��7���)j]�R�[�օ�@�#cEg=�JU��B��& �ɕ�5S��!�ɶ�TBh�����O���;��$-5��"��u�P�<��2�Հn�M(��f��sۧ(,��%��-6Q�Ϧ��bY��~}K���3���9����s�2,�`�)��� l�CJ�a����@�Ybߊ[��#s��'t t����Ļ�����مo����C>�	&u��r�w�KlG�|�}%�T�G�_Yd�h�p�f^Q]+�,)f��R0��z����-Ȁ1�{|�<�m{��a;�Y�LU�=.��e]�]Kh�&O�a°���7�������t���zFL,���� M)���-Q�5�wΜ��ڷ�ؗ��=^�׹	���\�:�	�^9i��k����BO��O5���-�IgE�G�ʐ�]�{6;�>����s�r����iP�j!%�ߺ�
�|��I�����1�$�#�����nOo��J�(����)�U��.@GZr+{�_ʎ���_���a���K������d�������p��҆� �<n5^�~������(2�����k��gt�eQP�Ls���f��Do�8!#W\���,�	a���`0�)՜L�j˭�-�)զ~?G�Y>�<_yjI�(�k�T��_sVȀ��4���F�t1�hޑY���y�q�1Uv����tL�dpK��o���v�<�t��[���	�JͲt��Rr����ɀY|>���������Y	������?I�;�5�}��
`0�a�"���keu)���Z��� �*%�+$���dr�7���x��m����G��[/�5a�,�r��ή��
�+���S���J�u��?��!���t����8N��G�DV��'=L �KO�����h�<�,l��Z6��pS���!�IG�������ɤ��ra�$��rLϐ�e^�-^3��y�'h��~��8F��hK��*z�W2��&-6�ϳ���0m��Z�!y9(*��y�)l�Q�]� 	�j�wß&��A�'���@
T�P֌t5;�)�K�K��sU���8N��Fڒ��?j���ڿ���~c4%�m7!��H�r�h�1��}�ơ��1�ba���cvs�g|a�i��Q��?�tHS��5?�_��B��)�ų�q�®ȉ���A,�UJ��(��9������!C��b�~}w�v�HHګQ-���7�ɬ��gkc������L҃qD�h�u!��a�ː�\:�Y�Ŗ�o1)�D�D&�Gf�#9QE�
�.n�zƥ���TEnD�� �����XL���u���ޚ�������zAg��=�#�Ө`���L�[���n�U�0��G�5�]��p?��cZjf=dPz�қY\��d�4�Ҟ�����D��1�[F,�����!~DON@�_:zݶ�h�p�<�����^%���X0�����-_YC`��]ѭg[d��W�9��t�D������� oC��7��
�1th�S����5���}z����!�#eZ����g�0<L��.؇}�,���\e�a�_"���~�|�/���۷5w��>���M�e�:�Ж~��|��%P��Y���{�-5k5K�E�}y[1[�����5e��[�$���_�|�7T����JfW���I�����ې�s�q���� �ȱ6�F��/�uV:��adͼH�m�NUï��FK1y�/"��#%�������Qx�0U"��б�a3�"c[&��%���k�򯍂�qE���΀����%�1��la_&+�������&�@��� ���3�k`���C��R��C�v�yΒ
�E�%���$�|�J�k�W�M"�ݠ .��f��T^���A�U"�~HȌ5-��Q�3%nx�-��wխ�xc����w����¶�w�����X/e��G��ߐ!��˜~p�3����T���]'�������3[�S��ȓ�!��W氚�(;���b'8')���/�7Ś6Ó���D�gCS�p��XF=e<�$��.��۲fY�Wy{��m�fҊ���Nes����oK+������'Set�L�	l�ݤ�֧�84��)�[Y�l!���)i����$~�KlX9��?f��|�^���T���o�jX�Y�p�ʥ\岥3q�EDh�Q�b8�D<Z7��9�N��2d�@[���^xm(z����U�l���P]���.҃�Z�ⶥ�)���Ș��7v]=H�F��"*�?#Gf�M�� [d�d.����oP&\L��
b��V�9\�}��AF;w�ĭB�ף���>B�x���5�L�����?^>�'����\���'���8W��3�{
+ڬ7Rg_6�s�:zBǮ^)�%�>�Zam	��j�T`?��$����C7�C����&OB�*��ܓAB��s���H��AS���_0r�}��)l���5�,]����=u��j�����Ꙣ���n5�- ��)����7��w�0F�Ʊ�i���0/�������osSُ<9�&�������t����5u䥶]t��F���Y�߀2�T�3���M��2&�y:#ZǙ"s�D����֐��Dt"<��Y˒e�^7�ê\�Q��nޯ�T����YJ��������U�V���AӢO�5�.���l􋆣�}g��5�����]#�|�	B��-�[[���G"4�'aj�C��HL����X�?�N���ʑ��6F�;���E�	�e�9;!FG��K(f��K�L-�ٟ\x�o��)l�y5� ZVQ�-\��/q�ާ��1! �}�id6�OX�����M��SM�W騦�|���r���͐��e��3oD��h2��vwG~ňj��8p�ǬOvgw�Ni[q�*�t6�R�E�bUF|P�j�g���x��hJ��MVN�v�����%��I1X�v�xH�!�G�n.P��AvY+
1ss/��Z��(�ftJÙ��}��8�6�<wR�o#�No����a�h��nl;unRB�k�+��#L@��|Ŭ��#`��4IaK8viR�ΕYo�^zc�x&��Ӝ�m1����&�`�$f�mD��?DY���熪��l%˖\�`Hϐqk�,60���e�:4ro�5/߆/q�i�>�]v&wT:�v�[O.$��J��T�[?'�-�^�U������B�&i=�����rˋ��%�:�!���=H!���AV�q��C�㳝u����^�;���i #����+Cj���3
�ʅ���=�}sd�̃���Fz"<H�$���_�� ��nf_� ;]O���1����Hm�����
=Vƹ'�'�|O�3�\�D�T
�B��O,��F�
�䊶�P6�b[����7R¾�>z ���K }��.���������ά{�V�_�>�u�o��d7�uG� �n����^΄b	W�@i�ûf�=��
L��V��A�*�n���.s�⨀��߰T8�%Af��-�����BSad[�5��� /B]eK�>�3����7}}�U�%�M���K	j�OD�7�c3�bb*�_*�(�Z�T�m����Ï1X< mP̠Ȁ4���K�T�mN�-�JK��X��\��G{(�~)Sp���س]�b�bO�\�����i+:�"T{$���[�&n� @M�A6T[��sP�`4�Jl��# �v/���T�0�u�Mv���������L�X)|/h��08`9��c5pw#H���o(�����Ƭ����л{3_X�[n�H]�6ϮT�j��Z�4��<M�d���vt�c��V���z�Q2�z�('�,���M�
>��}uo�	��x+��|:q�kL�����Y2���m�</z��4�%���#�����D�D�^/�07�$�Oz�ڝMm�~+#3���((��@������qM��7�.]�0ّ�I��#m�ϋ�wc0�\6
�CT��0��+��w�wN,d�����7�:�ᯎ$��k�z�"�(�VuF����X��Ǥ��"jd<`�MO�Lh,�L�A����o�*�oϲi�Pr������%d���8hP{_����|��"kϢ'{J6�MWf��(��\�r�G�6�v��nq�&��� gR S�8��LR�4��(��s�'��Wu�[�_2lt��B��$$h�S_�SOtt+�^$���(X��B4:A��(7���S2K�RoJ��"�Uk��Nί̽<l�`���#zxu�P=F�_��C�7��� ��`�MEי���CN�~e%�7'r��X��9�Ru8Sծ'm˼�7�so?���cl��MW�|NЀ��[�����pa9B��t�����ɜ���j�����ќn�Ժ����絇�E�"9�Ii�,��ǚnϮ��r,�6�]�h�)���3?aw,��U����w'�ӫ6l�i�7u7�����0�Tn��� l�>���|ړ�t�uO^�k�	r\�W��P��Ų�DN�#[���Ǹ� �%�ʆ�v{�B:<}'"�S�!���6�b���?���%�2)����}�X�>./��G�؃de�@6�2D.�)~�cwa�!ϊ�$.�K�%��WZ�&��3k�ra�����`v�zX�� F v�IܧG�,T)S7㮑o�-B"^��3p|~j�Di�h^�o��[8EO,µ���M ��ʋ!;3��c�_�=�Aq�H�ũ�����U5n�3[@�:v:�8=�[%���|�ǚ�(�>o�S?�K1"����K����.�c熄s�T"h�W�e����%�e͋�e�m˩@I'������'��6?�~iNR��iO�x�����Ao�&��˦�=�ea����ǖ�
�����!f�I���0��=�=�c	8�sCt�?��{���`#KH���	��}G�c�&�m9>EwX2�������nӯ��T��������V#p���*��EP��<۠5�}}7̴�đ}T���f��#�XucQ�8�ս��B��/D ���X&�(�: �}����[R �7Y������ś��~� �Zy3�$���yYj�G����&�֌������q�^I
s0��3b_ä| ���X�6�}"q��f9��H�Dm(�qٖ°�.�QEa�N��$������Y�ۖ��A1���9wˮtu�k.��O�<'@�OH/�YS�#�h��B��[g�x�%˓�d��0ځGJ�����xnX'	T�?�z���B! ���E
vߨ	ȓ4ߨ.�Ʀ��޻(b�v��v�V��eK;}�x.�>/�Ww���h�F�N�BP��ܤ���j�$%p�{���^O���d��`Yo�)Ut賅H��!|���Q|:�J��O�3t=3#�,�ψ�11B&��;�>�	+�-Tw.O�bG���F;��|��l�S�Z��(�3�&��Y��b��[��;��k���Wu��y4+�O�?��7��>�F�����)����}~�0?�j	Z���#.6�"��� WU�ڭe���9`k�ud�D���8�*_h<(����j�a��7G��������Xs�l��$�C%����阐wd|�5\e���M��t��/NS�S��9ā�w���܀`�V�%��T7�J�����$Ya�+jv2&��xj��ᬯI�����(N��]�pk�T(6kf�c:��Rs��:IS^��Q�R���XE���ބ8i;J�/��<�NbN
��D)Z���I?�3���F�]��^�ʳ�N�	`�Ip�]�\�%�b���~�-*�١ �Uװ�k�Y����!����񈖫i�p�l� �>�C�@a%�u�(=���v�Uw�M�;A7f9�H9x_(o�Zt�~�mv�um�i����dH���S/��!�.�C�ܐ�"(s$ny%�S��N���,{�H��6�ǚif�?��!^ଁ����pc,!V'�����l�ܟ�oe�����/�xWi�^�U#4d�S�u ��S����ER�*�D�Y�B�¢I G�sJP¨�w��s\l�bz�K[2#k�0yK_^&fΝčn�Q~	>��h�%�jQI�8�����>���X�<@�q]!����Q�|���*�c�T�����8+���������#�X��6�|ډo3����+�Jx��ټ�=
����H��谮(~¹�ñlj@Ð@y�*�o�?�䘼��o�v�vꁦ���>�e�*B�=�I�j)�zfB��Š91͡�\���xlI��&�|U�����ڑ[�ܮv�PG�TȽi�Ȍ�!w��H���&��eU���tt��{�ب:#+8�+ا U��G�;�
Ş�p-^{T/��Y��4G�a���#�b�Oh��{{�B�*Bm_u6$�Z*����tl�􆮦�}CTh=���ޒ ����K�;���<)u	Y`�y7e>��L<���2Ft���i�m�"SéyE�KR�}~i���P��'HPo�����9��.�X�6���.��52M2�}�����F�����)8��;ro��s�>ݕ��ñ:�}\@l�&ߝ'�C�P򁼦�\����>���卄R*�խa۱$����GGL�;�e��!�n�g�8M�W8�|/���Z�*�9��b���8w>�Ǟ��� �r}��U�Hh�G$h�ԞF��6UEeG)�+�J؃�)_�Ƨ-��դ��gS|e�K�}�ͅXfx��D�;8頱���9h�|VD�X�<y�k)L�/�����b^�Ңx�=Þ�n��*�v�U8���s^��`��>PZ�g�� �p�3�Cz	��~l%
Ga����Ƹ$N 9ج��)T��JǬ�bK��5�5�E�$ T��{�A�<͵Y�&a���B����7��2%�����N�9��H��%�V]GA�����_�z'���4��!}я\g���T��R����,����d�n�f�G��Sܢ�Kǐ�*�����/�ǳB����l�#����L8o���A	��h6.�:�t�Ћ�İM_`�ߧ�Oږ\˕Σ� ���$۝�\_��##�ǰ/�vQdаXM��ZU�f'5���_/ �BL�0/3�Wbݚ�9P�+m{�n��Uh�@:$:
��}�U����K(��VMhQ�ws�Ȏ?����t�"qp�!�L�0����S 6g��x�%�������^��ßSχ!�-�V��@�.�D�,�`�j`o�Y�_˳�j���9Oi �ynأ=�U��k��1
0���i���������o�.陈̖uj �`�=4E,'f�`�E��e+WCf\����]��K�J�j9�?����2�'��FZ��o���R��;�C��Li�����Ж�ɛ3�a=w���7��<����N� ��}:�8xly�Jp1�K���6�m���MyJ�Mly�M74����y�nX�[���>FyC13�bW:�q����~��Vv��.��*�4��Q?��y����� �V�|����	e��짥�y??�z��͊j]z���h��@�,���A|�z�[D��͗���n|�JTq<�Z�l���'���`��S��p��V*%O�w/��2]$�ѵ��Z9����;=�p_�awv'v�Zm�c���d���s��h�l|q��ɩ:L�LN�E6�Y��UNO����+?9	����@<�RҔw�k���3: ��&�z?�o,��3�CS]�S����� ��2a{q&
�����V(�ֺ��5��g��|$���I:�� 5��?�����?����ro�ZK�_p�x�3�Yѕ@	���jU������Y��~�_U�]�y1�%���D�̜\���?�ܠ�Cw�e�->���E��A:�+�j�F�P\�2]ϋ#��ɻ�*�g��r��3ޤ��ɫ�'0�u�
����>��+nَ��>10���tcD\=:��
����^��%h@|���$X�{!j�Ay���7�f���ޏ_Kr�7�ӧ����o
u-�jmiԶ-�;!�\ɫ���(`��`�7�S��TD�~�G�J�ˊV��|�6{�0�
����~-UM��
A ���9�Xz5����R۝�����0MBr��U�t���Q'L�Ǖ�N)�簔��?-tԥ��H��!Vx�������<^��T_�,�~��*�����֭�p9S�a�o0(�_�j���(NA�F�[}�y���ڞ�T%rG���bd��	���A!g�6tQ���� &^�|���G��F�s�8��&��P�Z�U�yqb�?��F�i}k�!Ml�ЮX��_Rf���[�Y6Z�v�^7���Yʚ����4�f�4`�ٮ��y���_�#0י4.�_u�8קݿF���h ���`#3���h�<l0��t羬��IªBSdCyI�V�d;���>��]b0:�P�!T�ks�JU�rQ�jT��;NYAeU�,j�[�y��h��Q��9@�>�����
n��ܐ���j���ݜW�.�����HZZ�E�! ����T�8(a�Y��ZӅ|��z$�L�7Ԍ�\h�-{�6����k�ao�<���;�z(Iŉ�6�1�9/��]|<.�z���4'�5�WQ!m��m%A���(fl��eJ
�r��.��;XY�l�P?���?c�P�W��B;�D�:2X��BRr�cS�2�jT9�T�c��U%�w���m}��Ϣp�b�3A$ǫ�J��	Ώ�!<���0|�(�����y��I�o"��EU̴+��eft"�] ����@B ��ٷo���y����o����\������v�מQs��n���l�[L3`�g�w�ftr��^���M������Zn���کN7���ܬ:�-��|H� �e�me��2K������S�Fm%��Ea#��6W�o�P,t_����Y��,_���V�!�X߀�bއ��0������3�t�a2ܚ�s����Ч�����]0���_+%���\���3�.x���݆�����<��>nR�|�DV�Z�}����� �(̞�kE]X���z8���W�k��i"��I�r<[�H=[������y�QRZ	c�6�lʝ/O��~Vq�ȏO�M�h��[>��-�����Ӵ�4���x�/$\�zX|uq�oɳ^q�\��].8�KJ=|�Ŏ4&T�Y���b��W��d�V���t��D��lW{��Hq������hb����T���r�у;��5�f�f��I_5w�A�	)�Ćv�+��ֲ��P~%���~ƏWI��^}�Ő�S��5��f'��4��pc���du0ς{�6�MŻݖ�{���9K-�b�oM�Ta��]��W��J�Nr}cZo�O��Ǣ=�,ᡪx�T��Hq%�����jd�~l2�I����MPF��Q�i��b�E�"7�x�Q�f�L\�Z��DcR�����C�ȈFУ*_5������m�w��@� ��W�b�Q+�jF�-Wi6r����g:�#��-d�jʓN� E�.d�{Oz��U�Huj)w͊<<6���+oOD����z���5O�K v��Ȃ���L.5���y(�^[9?y��wH�j��6G|?��Y�IJE�~���!z����u�4�8�#X*��6}"�o�{�]+U�Z-���m�ǡ,�����D�Qep �Y���Y缏$K��*� ]J�*��.�\�u��5p�6z��1�z��� ]���@�\`�p��P^���ۗ`-t;t����U1�$�;�J.ٷ_���N�����K9gӲ5q�IS�]��=ۂ{�+�vTh�4INg�뻹ۍ�*�������[ؗ�'�%_c ���z��Ã@<���Z�x?�:N�M=r\�TV���+�4Q�9ַ�=�c>��2��u;�朒��Rs�Ќ�[,+2l��ۚEy]��>���5t�(G��HxJ6_���*�����|'b�v.E2hE��������~9r�|���]�����U��<FZ�k-�b�׊��Ζ��l�B�b�(e���.lN��3aV�x���}}]!	�E��W�l�թM�y9��ls�a��w3�S�@�GE%᠌s��?� ��v������P4T��q2��v�.��S���ܦ��� ;s����j�&�p��s�g����aUM�;#f�2�={�Yޔ���
Q��!��e_����\b;����������LO0o+8Raի�}O!��W�;4s�$�t-L)�L��Ezg����p��[�1�ְ��3I��m5�#�����;��K0�0]O K�Vw:Τ������,�<9�`W���G^�37��4x��,�T%ēi�l ��{�&��a���I�G,�#��P�R�~Ԧ������4�$w�
��q�9�_�B�̋E �,���@�)����	��rua�%a.��g_jx2�+̯��\���~\p%Ţ���Z��9O�.���_�M�s�]5d�8q��kM`U]�9ƑS8�b��];uM�ikLc����	�zHe�E��iQ�T;�@!�Z��Ѵ_=57QE�'rAP0�FRnEKF�[��kE���	�k�Ͷ6_J���E�D@/����{�e��MLn��_$3����n8G�[�?ٙ�i%q3�FGd���.	@!0��=-��w�b�AA��Y��C�̭�}�3ŉ�а���\��B\B�5��ʾq1�k��|H��� ��N@(fK���\(?�j_ƣW||�	s1[4�;��YG�̛C�7��L��i�,Xc����x����M��]�%M�Tm؝�~�h�徂׵Ox�e��-մ������V�K�jsn�yYk���z�T!:����;.��?oJ��~�	b 6t�$�i������3��,R�Qv+_JY��c��ؔ�k�絕Y!�����Zx�gJ���� (��C@�5ڡ+Bs2l �|�鴴�L7,�6���>�d;�)2g���NM�H�d�&ҫRP�#[�G��;�2M�B�{�T� �s��×j1v^]u���u�.�=$��E|�����h�N���3O0�kN$Q]�}^�=�������G�^r4D��_h�H���m+ً�3�7�\���`Kx,����g��v<F�E�I`u������L��`�' cSer�5���m
�fTV2u9��h�+���U*��=<���p;���J� qm��qg�U@��m��S������pk�5ߍ&��EO�^=�HEQ�����������0�xzS�I���u����:M�K<C���ݎ(�z����e�NO�98��Ƒ�g��[< �{5j�ݾ�܍��V�(�)��ٳ�)Ff� �aE�ǲ*�jd��H$ء��VJm�a�l�?�"~��s���pO�Q�m���)3xC����m_
�����5��?D�/��6҃��
���q�e���P���m션�� -�t�� b��;�:��`���`4A_#��*�J�dP������pM\�/M���~�/�zӲ:�^���n�%Aen����Ii����Y+GO��	��Կ]��f��c����MG�z$�AR�V�D�g��7S�s�E2�T�Y���nWI�??�L͝C:�n�y��P���\O����~8�S\�N�-�	��W�b{�p)�8��J�w
�ue�P�#w�����g�!ӭ�`ͪ��fw7���^�R�k�QD]T%7;q*M$nm��X6�D<]^�=�qxU�t4����p�`b�t��9�du�R�p��(.2��8&�8=��K��vn]QJ]���U�@tă��--5�B�F6�z��a���Am�Hޜ;b���1�;N#I�ڒ�w�Z�C&�c�.<�J˅h��<�mt=�ǻA�$�o��9b��ԉSο�Sx��D L4Y�K��c� ���P���O�*�"G�wĭ�?}}�h�i$�>�P��ӗ<�H���;��@��Q�������Wt	=yhw5Q��D�ߌ���Þr1��u��^8#XX�l�P�ѻu�u��������C	����'��6���4��h�מ�2�sj�u$�5v�wX�@8�S�~2��H�_Օ�u��o=�RҀ!%�7�LKmΡcrZ�Pk-��6_w��DX^��`�F�σxL!��1���h�oV��0oM��Z�������2A�N��3�-�^����/45�(�>:y�7Nv"��=�5�@ـ������7��p���$5J1����h��B�y)Es�MHGP�ƄD��.t�bD���$�ޢ{���z~�z��ރp�Ь�4��)[���KyT������9m��N-T�Eg���i�b` ��`(ڿ��,��=T}�ob�r�3	5cҾZt�m�n')4P<��K��O�Y�A#��#� �|�r��3�9�g蚀�����p;UNY�p��gp��7c������H�������D��금j�����+#�O̹�A��LJG�^�ɽ�vB��&XR�������4�c��d�7���� ���a"4���J��#�C2��aqU�=�o�i,f=bL�8�?�Q�&�M��)����&�ͩ�U@���.T	8���E����@��Fk��3�]쪞RqF*5��~Lk�ܴ^ �]�'����|��
�/1A����Z�S�����
����CV���!� �"��V�=���C�v��������� qÞ��+y������[�Ջ�h��<�̀�Zr��E�/�zF���?*e�e��3c�b��2�p],����Qc��p3�x�]�OF�/t����Op��l�6�I����E�ǚ����	Y��aƜp��j��������d�W�
��z�b����N���k���</z\!�I��N�|90]��Z�»��O�(dcQ��&�LeRv��=��Zn���J<悃�?ϵ�'R�?6�f�w�Ԏ���[��q�ącR7���O��uM�m{FfW>���vF1Z�)��O���9mD�;�<0	��oXz�yb�T�}��[=;�nK�N5��9z
��T�ҚQ�U����Ӵq%����!xĜ!^�AYuehs7>��^���~��f��v��ŀ���;wZ��۶��AK7(��y�	\sWoIq�_�K�ۘ���)��7�Hª�ݻ Xl�;$�Lj%s��(N�8��e�e+��L�d_��)x]b�r��tseϳ7��]#����ޏ9<��?|$����ɼ<�K�٧@�e2F�L��������mXR�Vk1]'���e�����*az��z#��:"����S�r�8?�F-B����DT+�ɋ;�7�M2���o*��{ [Q9�u���U5��ښI����8�E����[K;�G�����S��4xv�1R�g"��ڔ��b+�w|Ğ�L�����K��׀g����n	3߇8�����r�Tw���n#�o�GM�{n�p��X�`�G;��	`8AX�؄��b!Q<)��]-��}��v���̖;�s�i��B�?����M86ȏ����լΚ|�K�4E~�����$�`Y�'�^��w�dIf���l\�+9�S�[�ەW��n�zS�n���L��;�Zň]%�Of��e[�p��%Y��gϖǰ3UA��v��N�t �_��5��5b�c�D��|�m�����n^Ъ���P'�#�\���.�q;�:�eG7�1��4W������v� �F=^e`"fe���oӜ�H��������k׬�3����~U����@��{��}J-��Wk�I-O?��p�$���!�N-���c�i�-��dQ�d��N����h���v�."EF�I��#�����9w�׫��cνs��&�&�֟��:l?Q�>/Gk�7zN�O�4��1���p�P��l�3�ϊ�[��_陃.*i�\쳆9AhG�Z���-&~��B�QH�f=��{ʈz�i�W�f9��i髿��	J������^=����?������
�_��8�N"C��<r	.����q֫�	�d��{LO��=B���@�}���i��*�<^ytpG�7|�`��K���M�P4_�ㄷ�2�����ߗ�txT"���0��u��UOg"�{�0�̏����dx�O}E���IP����nz��LŽ5X�N����+uD�0�M��N@D�NR(�/�Z����Dp�����f#N
`�����X�`��}t}��D0d�zsJ,��ŷ�?��3�ې��x�P"M]��U�<�j��PX{��ˋ�r~�?��O�;+�w�2�{����Ɣ�J�x%�z����F!��\���B�<\��e`��ёѽb����ư��3�=d��5C�2=[io��E8>4�絘z�Xl��tZ��l|�g����l��~1��Z���/��%��$�B}������E��b$�#E+��7���8C�A��rlm��%Jb���#N#����N���e=4��ѬV)��'����jx��&y�o�D���6��B�n����A��F�V�0�Ǥ�Sb!w� W�;, ��h�6.�7i	��ƥ�ӾM��R���y&����l#�Ƃ��^� ���+�LN�M.Nv���U��r�r�9m E� k�L)��ʳXl�aYj�����J<M�5D�������"��H�q�qO�0{,$؍�F�p�Th�fZn���#nû��������7����M�r���1Go-�TE.v�d��蟌q���f�8�Ь�/@
��"P�Z����+�O��rM��u.ie���Q�ӕ#�>�K��w���q�*o*s\_C���\&�4�1W�5�/<NqԹ��Qpy�zI�}we�YP9�.�{���6|�k�'��c���Π,���k?�.Md;����Aa�R\�������R�L7r���;@G-�&s�28{�yn�����h��o߃A�����$�bf���$�wQiN�h�G�$:��y>�ۃ:�����i����b��\��:/� (����pB��KT��֍��/KN�!���C0 g��0�x^]x�H�E�_]�:	�:^���Ɍ�+yOBO�`޵��a^���0�&:�9iӻy6�b�F|�W��;<��UҨ'�B�w+ ��a�&aN��z��F��L�Q����XM\����U��	ǥcK�����4��G�TC�j�͒�U�m�g!�mU��!�^��zq��];޵��7��-�ӰU�(�r���/ C��Cd!~�@9��6yA�Lx~���'�ɀ���U�\�0Jv���m5���O����!���J���JJ��.�]&��Sb�!��>@>��V-�H�"�?"O,�#���`�it~����5�À���R�t9�b�aٚ0�7^;�V�%�����Ai�t��:ͲD�v���i�����	�uK)\&�e���A��G���r'&�Nq��T�1�&��TrҾ�m�����)Z-�X��H#K�	ؿ��{ �ˮW0��j;R43u�
�"��>��s������"����Tx3w�(^�fq�>Ǉ���J��C��k0E�I�!�M�(Q�"<�e]Dga���̀�~Ѳ����k��- �\�A�SW\����ዸˋ�E[P<j}���dME:{���N5��X��9� ����d���[QR)]Ҕ�u|?�hM��<R ���͝zr��(�$��DY�Ĩݬ�������A�ATl�&)`���" z9�f!���k����e��
A�j�b�>m�?-�Z9��U�o#HČ�g?�=S��J����ҷ\K`�6��阁�DN�{�.��0���m�~@�~}�կ��J��B�"��Ն�q�9[�%�,N�T<[����󝧠�I��q��N� �8�n([�U��\�����Š��;��4<����Y��j�����k}����ũ�Sgg&���pf��/2.E:�U�6v���cT���6|�==j�