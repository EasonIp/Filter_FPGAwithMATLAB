��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M��*����g#φ'����T��6%.^f��8{�^v�wK�T��fAN(.�oC�Yt���Ao�>���� �h�*��9礩[s�Tj˧��Y���oG� �'!�D!�#S��E3@b����}��doB۳��P����F�.r�Z8Bg��������K~�g\�l1�i����r`0���Sw����X՛m�ɒ��Fq{�GT���܉Ub��o#���;��V���
��ħ�u#ĳY���Ei�Տ�#4�P!���	j�c0G�'�(t�g�5g�O�U���H�x�{ؽ%�qT�ˡ���٫^�)�׶�rn�.c����Z] p�ֆ����s��b'��qw�3�Շ�O��)b��тI����\ia(���J��z�	�#��S�2%lĩ���l|�Z�V���p��M� ��2Y&ݖ�~�~h�ě+]�H%���/����!��s��I���ր{<�a�{qb���?^������Z������s!z(�Z�ɗ����(��W؁g�u���M)#@�E�	Z��M���/X�6,׽�"�Q�Dm08V����0�_�feJ�O񠞤��X�&\ݺ�Th�+����u���&M���{^�1
�_���������������+d4��(�=}@�<�_`�L���ގ���o��o���߄�7c��*�b�<�C�l`[K�ܪ�j8�R��{� ��|n�}F�X�<�n9�;�V�b;���:�U>��$�>�wr�'�FTm��9�����Ř�L�ɋ��>��4�!��lT�XҾ8[�׆f:@�G(���ߖYiH��mq������f=�R���<�f�xpla�u<Ū����Pxv*I��Y�Gy9�4XM@�v�4��݇�Uɛ.7�g�<��	��+��r��^a��s���̥N����U(FD7���Ԕ��j3,�9�/d�4{��"�s�"E�-.x����4�eƕ�ءVv�	ф�s|� ��m��)?�&787���0Ű.�nf�Ԝ�XlW��7�'���*��-�H��$3��I�HH�}x���|c�ˇY�+;�:{�� m7��mA�ˀy�!�3j��>Y���|�qn�~[��Ւn��V��p��8��k���.KZV����j����Q.8�Z��2�TB}�v5a��`�D���iO+�27�䂲i^?�,x'<���� kp����%y���V8��wQ�)�Y�LܶL��Z�������L��U��(4󲛃��IߥѴ��}�@'x��Ks3V�A�'.ߞYA9�ta M�%��ϩ��d�<%2&r@4ҋ6g2Y���=k��=�T�M�i�U7T���z���i|~Z5`�b�f��=�H�{�3��p�LA	�ʁ}����đ{�t�o#8ňejh}U���=ge�-���qy�TwW��4��Ja�ߛ�4��4e����C�>n��Tqպ�殺�bk_�_�$����~�o�G�~�s�á�70��y��Y�5��V8���Р���UTYKB��Py�BJ�TS+0͑���<kf*׷7���c�q��L�K�!�6#�f�gCO�2��JG-�_�&�x�1��*����@O��g�������6�xH�z�8UM��A���]�t	{�a�n��;,�$Q-�'�Av��*�`�ӛ�H�8���!e�=
��k�b�V�1<�0�+,�9�wZ�<ۡ��Ww6��:��`�	az��uYH
�ټ���s+�%(�u������u����I��L�B��1ݶ�zǃ��<�z�fJ|�e��yQR�{�r1����J�.�a��,Zag��I7�d>`�Q�����oI�S���Gmd��=�ڊ�f����wtK���XYթpa��C��������P|?�r�*f�Za!$L������+t�e�����[ή�N��ڑy���yMKr�%�i�\Wj	�{�`^%�2u�x
��/Z�΋���QRlе@��6 �x�"~�a���*����,�b�"���0�:H;R8r������k��7���T�ؙ��Sӕ
��~?�F��Vu?�w����F��2eC�8t�u���*sN}����
�N�<k*���S�&Ls��{>j��X�ǈԵB)£��I��T:�`��C�"?�x �9Z`��$������G����]X	��_�	�Ϡ�����ĕ�H]Z8Rd9v�ǙO �}���c�R}}e�q��(���җȞ|�лPB+����깈,�6a	x�X�%V�
,6�i�`��i�1;W}L�r�gdV簘yb� 0v�ֱ���3�j�����Q:��&Z�xT)�o'�͐"8�c��}{r_]�_ހ' �ߩ���T�����ӵ��R2l���k[�㈵��:��l+��^���pBۍ2)��j':U��gm٭{3
��=v\�Y��*Y��&�.d6�����R���q҉7'o�$����gɗU�=��U����ʷne���x�o�dj�/�\r�DO��X!�hLNz���MVE$��M��6s�K�CB�.����G���}&�'��y;3m�*�TR��9�^���D9?��G՜*��tLIDo%-�H#�M9E��:�\��'��6��5�W�6#�瑩͛O��j,AR��G7���u+�.��5ND�̌�0�i�G"WNl�Yǫ~W�I-��s�`�-t�������� ����.���)}��M%_[J)U{E�sxx�rʟa��9�!H���W<<O���_@UI>�M�RF菟�|�:γ�a⇑���_3>@O���Z�&QB� a�>�� W��>c��@�◀֑|�b�[]�/X�8t��*���m�rm���:�BdR���?�j{�O|���][M��0�%i;��y�i5����f �o�ZYC��'5�za;$�z<�W�\A��j%���4��Ջ��
 w`��Y�`p��3u�$8zV!
����#JA~5aI�Rؠ2�xKId��}S�вĻ<C�l�Cr_>u�6"��� ś�X���}d��tu�V
 ����5�/�F��u�j줢���=�d&�72M@D��K�]��l���0>H��W*�9%�G��k���9�7[S������DwF�=��$Q'H���g4��h�=��#�����m&?�[ L]�Ѝ�:F�T�E��9�u��/��p�<{s+g�a�:����D�]��"VU�BѪ��Zϵ�`.y8�Z� �y<��9-��g�۷�O��u 90.�?���9�|Ӎ@��\*Oo�^sUcC^�O�|��`[�����  �0��<�?����(M���=�Ȍ�8
��%�ub�3|V��l���ȵ�iI,��y�l��^?���-t?�Ҏv�
�����{�	Q��?z3:fu_�5�c�@��Rޚ��s��(:���v�S�g׽;���� �&k�L%b��$�/�gf!
����g[����Lǆ���Ɣ{���n;�n�\O6���Tx��՟[/�Z�jf�f�觨\b�q��~oܿC��(T N��j��P"蛇Q�U ��U��������k�O�*+@"|�d������^M}i����u���I	w�Ҷ#���FmRd��Ȧi�#�w���{���"J�����)��4xK�l��d�}�!��KGX[�=����T���˴۲��7��a蕊����'*Ym�?$,:�'c�/a�{���%�X�3��<��(����Ò�`r��b񥡩�_i����N�\�D��ˉs�?��N=JIFO 	ʦY�Z&W�I�nD�z_0��.P|*��V�����_�[��c/<5V)
��}u�ڧo�s��bP�	 �̲�??�E;v�0�X�N�@����/מY}�ӓ�f�*��a
`6\��>so���
e�:�}pj��K�'ޟ�`�C(Y�Zd���OV

y�Yv��`�
�.�.�;K� nضӭ�9Jw��t��W���G+���[:��ħ~�}&�*�%[���T��� �F9��Q��@�-P�����b�.jm ���3�~�Aק
+���ȥ����Dw��,�FP�S4�.B�5LNk��|�t��$�9���T��;�9��1>�X]�^}U�n�����Si#��\SR�Kfk�=Pm���}��'�Q8��R(BZY(1���bK=Kj��ܴ�����-�u6�Bof5�!�Q_S�\B����:��j]Ƞ��T�G�ˆN�����~
�������M�k��>[f6"�3ܙtp��-��c�G��c!��� �����+�y�n
W�Q���;,v��G���"��7z��/�R7]j�uD�Ѕ�#����	�dz��ئ×��]��V��h,k��o������3��~kɜ[�aC��N�GA��6���(3ɵ�>�F�v����S�VL��O\!�"6imtI�`����u�{{���y�*}2)���}� ��0ПZ�~�ĥ����VTU��#i{B���28���/��Z�u�l^�������� 4kM�����E[�-���^���3��h�j��p:2K�ٖ�F�/��_&)��RkW a��t�������re�m.R������x�ge���f�f�z�t�=�r�ؗߤ���q-v�1 �g�b|B��t.�=Ä#p�@jX6��b!��ms��tO%��Mx�D��&�����*��`:�?�P�[�Yй��Y[̈�v��E�z6<�qՏ=༴}���G�s�^o�����f�i���,R� Kb�����O�1�AF�� ���l��pI�
��dA�0�҂�sk�V���s_����}O@{�ʸ�d�	C��'}�o�/
W��P�BU��i�s�13BLB�1��ݸ̡�޵Q\�8�b�5�1��@C�Co�4[!���%��[���o���یJ��(��s�a�m%��֢^k���l�Txl>�Z��]��,G���A9h���kF6v���j�s�ǯ�PL� ��2��m3�Qڞ���4x����g���"boV�,R�x+�ڃ�c)�q�@����63�#�?d@+z`S���S�O�f��~�E���J�����>����B ��sNZȒ	᭙~�q/���oI�GRq��T'R�z���AxU����M��m ���e�g��D��47��V�d�RK���w�協��w�O>5��p�>�6%��.5�ЛĜ+�r�X� ��� ��l>�T�FL���Nm���������"(*�|�_EC����_ʮZ����1=v5�:��)�Ӏ�Z�,��r{���HF �3Ƴ���Ѩ�|:����4�.��(�ՀwpCG�~i�wg	��66����;$4{F�M���w��h\�
I���g����]7����H�*�:�$����F�?F�,�f!h|d~V�$�j�������+j&�& �d�M��; ���������U��H{8����Q�y9⵿)Y*J䍎y4����}n���c����ak�)[��'�y�T�߁��:�\�a���/	��	r�:r��Ԃ�̏�#\=e�t�m�ʶ�/rz&�P�Xpt|m,�>=VK8p^M�o�����`�8�[�Q��/#����v�X���e�;���q�-�N��m}&e��$c0�U�c�p��/�Y�g:���'�,D�[�P�D�(�m���b^%SC�R?]�ugf�<t	�#��̓��뛂�36T�3�;��h$a�[��������#D���*C'~��9�93�e�,���uJ������R���4���ƶ��J�_���͐\�p��rY�h������i� q�읿����f��J�4��dJ�mW.����S���h�������9oj����*}1���CpQ_MF±X�ݦH�|����q��u�F3�X���! �Teb�i���/\���M
�[�Θ���f��\�R+�d���w(�|#�3�M��n�#�3���4eIAx�U^Y���r/�B�ކ�ܒ,~�l%�*\��%���51�J�^�ya�S����L�zfN./�\��gwK�rŌ�16E���y�R��0F�>ߞ"��9��*z���(�0G��l[��B��rY��/>�6�i�Y/ھ+?[d��5��f��@
4�	����w��Y����
)���,=�v>KB�� ˂�ݭQSY�?�:���3���2��:�y��������1+�Sqy%kw�$u?��.�R���2�7�RS�O0/x�a��G_���0�Y��Ae;i6�ҠQ���ʺ-�s��oa��H�1_�(���Dn#�µ��)&�L�z���t͐�u��>�]����L������WO�]`#;BLh��z���[�ٔ���V??H��=Z�R��oM�E��=m9���r듰�o4�Sh����EWR{�072�p�~��<7K �T.�h�6�7F$N/r.HE���<���M�"�?׌4�|� ����4��-�)8o���	�&��o���b(�(�֯L|��Q��o�>��uG��wU�@OXp���`���M�/�:���˱%2[��r)�ͼ�Oj���]��J�2S�p���V�
Y���U�k�+r�]�L&f�;��ܞ~�w*�PA,@"���z[�٣;�d��G��e	E�����.�����[�c��b������2t���g-r�|n��k�J�{�Kn��z�V������[����p���W�mF2������� gR�M�$��O�>F��U�)���y4.�;� �OA�(��l=)�f`���.���6�O��kD�P^@����0�{x^�^�PU��u�ʛdJw�_��s>����E.ڦ�9Y�4�Ll�<�x�ǽ��zA���\3��A��^��#��(g	|h���zI�*�KlV�{�.:G���B�z����5��0�.�tNK��󕒸߃��I�J�p�
�kj$��B!�m�g�d�2%�#�jMC;�5Vؼ����D�[�J��h^�M��
OKo����?�$s��1!3�:�A2��A~?�}B�����L@n��k=����¹�p|buIx��e�ޥm�$Z��8P�c�B;�k�q�o�h�L�8���S+���������-�`4B�7�AƷh+r�(L+"[V����i�@u������j��om�����	���s.�m��,u%�������{&.S/)��<G���i�m���Y[?0�8�2{O�f�N>J��=��.�O��;ؒ9������f_4 II̬d T�?��ȑ��PL=2�%�rU4�W��(U\��/=(k�X8�0�����D,��� ��xԊW{�$��@�2�8��x��n	٧W��X�NV#���>�y>Wp��>�~���������]~I<(oO�`P�HN�;+5�`��@EŅm�Z	%�\]	4)�����d�L��d���M�ȭ�RR��Cb5ݭ��!%�R( �^TZ�p��.D��@!�v��`����V�Dg*�3y�\���1ո�Ip� P\��Q]��! �c�2O�ε��U�)�}���p����C��r��{�r�jbP
1��`)�do����@e{���c���c���0ED��B���2jjq��V�U<�\DI*�z-��Mۢ�@8��f���y�k��4*y{8�GI�a��qUY�uR�Xf�LC>�a���,�:��n�(�#�$��@�.����ο����0����S��Q����o�j��;l	��a�M`EZ�O�&��
�S�S:�qXU�Ư�I��-ǽ�����!>��$�d2H7E0`~�p@�)�&��p������v¢{��!�q�>3[�L��V�6F�:��~�lN�eپ�^��3����@�X�Oo �A����JF}�攽l5!@�,$�ִ�,un8u���e2���Gw���L��<�Z
���L�<)Ϋ�!�m�v�]V��xt�~~���@�w�N,E�5�~?~i����ܭ7���4ƙ�_���Mz_�s���~�������#Ϲ�H���)�g��o��F��E�;�ySv������i�A��Ry0"rQH�b��-��Ë�-�N����ZsҼٹ�<�w�6���n��p�y���}g����s�,}�}2��E������(�b��fbvE�$ǠR�U�Ҝ3������8X^B;�iA��t�h����^�vF�����>Q��;Ypi�v��A�'$�[B��%�ċ�Ab��z�3�=2��c����1bM(�_���f٬d� �Ҕ[�W8�"���Q����Zȓ٘i�u�M��|�؀pL<'6c�	G��!lq��;�L�Q�u��N���?}D��x8� ��^�j�V�\F��A��bRjV��-鱦�(��.T� 3�_{��>�9sُǿ����-'� ���+�������L>�OY�廙]�
ԑ���@��n�����K	��N�f��L=
�E ��V
�Zt���V�i�+@˒�<8��H������./���>�����6
X"^>�}�?<���&Ʉ')����r�I�v3s�4-L"�I����E1����>��o�T%(EO&�4�eȦo;�b���+�U�R�jžd�$2��vJ6��<u,XiȲM��N�<7���A�n�jxZ���_Y� ��ΔBd�o c܉����QG9�=���F2�I03�H"��R���_\Ms�a�&�yB?�c�Ű$Agэ��)��1^*���v
h#4k�H}�W�M�팝a��ٷF� �" ���-����8�"�[E�ϱ6r,�e�� f><���]X��TJ ���9߃�(1����E���1���(n~�`�[A9�s��Z��xG@K�x�}U��0�A.��P���0ސ/�0���,�Nʄ�Τ
�lف{>،��t+�<�d_ss�<��Q��0�u�`e�8x��Cb����'H�k/ �<l�\�
���*���N8��-���0,k`�oL��'�C������L��Z��=�@���}��l����z��Ϗ,S@휌��'|��+jL�j�De���ٔ%sZ������^�uQ)��^��Y3P�

����ʇN�jP��ƱO�Q6ȼ�Țjg�4��l=Dh_�E����0�r���[:�]} 7+�������(�cj�1�sC��(�c̽[�ֽ�2_ζ-��z(���B�r]�Mʺ'��5[��h��k��{�q�~`����/�c�f���O����7��ܜ����j���AI�QO�vZ�,�(q��Y�Yt�K8+���6�5��{���Vw!�9rQH\�S6MS;9e#&��vNt��@�F�,��{[����{��zYYt�b<�J=0�;�خwJ�)��ph�B��u�9�(���=���"�?/^N�H0�a����\n��49IA���a1C��/ݩd[�Y/��v'�cb�`�>����wc��&;�y�_�t�?�~���;�MQ�{b�Xl#�L���:#���k��nd���)/6e�S�R
�M�?���E'u�w�]C�q��Cw#i�l������i�����R�΄]Gvz��a�1ʐ� ]�H�{i� �7�I�qR��im2�c~7eQ����mѷK{8�����,�.m�g�l�;.�^%��ӨZ�#�.TG�pd��?'"�5��.n���Yf)�������T��ظC�==0��%}A��,f>��ۿ��A9�b�ɐڹ�ä�,��C�=�û�&~L��(s7����H,�ן��v0��� ��u	,a�|5��E�W�pT����$,�
�pa��&w����_%�hfB|���"ή���zK`�ԉ˜�i�E?_2b���ײ�Lr.�o�ʭ�/��G���O
�r؃|��S�����=�j�Oc�qP�PgWf-=��&�b�̮�A�9x|����x��T��W�d���K��SE�c|_��O�J��@���@���i$��+��Q���1Z�֨R�=ȩYS�����]?�U����T:���}[ByeI����6*hf��B��]hP �ju=�1�$daՂ�B9kw߻[YQ�"���;<�%ǔ���o�1�io��8X��a*X�gMXI�i��p��Fd��K�&��^g�0ÓE=F�!\�����"�4Ք���#����./�1���*���ͨm�f���t�=����&��r`����(6/2(�rI����h?ħ��=[���m�ju�X�MiU�e�ډL��c���A0{=�cw^����F�p�*���]�)�6co���/���	�>��7� ���3�je7K��ޛDHaU�qwƱ��*h^�W$�����!,����d��F��WzNE�";�iU�j@��
k
��0]�q��y�:�@���'���Y^S���|�z�����1�;W)�`ޗ�?�Iq��0Ƙ&��Qˬ�i��V�2���\��=�!���N�	�#�wv�d���^����3LSـ)��2��(N���KGߩ�RkU��M\n{�UC�g�G���yz�Op���&�V��M�!t�N\zG�3�1��ċ�"�tײ�U��U���H�A�L%]R��%���$ku����i0�|W8Rt� ����d����.bNY���o�Й��n��1� Q���VL�s��'��NX�ң\<�c�K�؜4�tM@�s'�-S��V�3lz��[$��j���_��7��u�����X	 �\|���2	�@�w�}��f�P��P�$��>nx��O��-�:��)���B
`���,g�tw�4�>n��cR����RdA��Xk����I0ƣY�e�PBY��SKd��4�(*��.�	�q|9Da�����k�&S�����mW��UI(w��rq|�� 7��u�F�QT9�^�taR~X����&���c����7������е�t�����4|�Q��U��E�E��-�	y��E���5>��6\���Pr���R�bR�if��F"�5G�-6^l��?*-�%QȂ��1C;V������V������8V��mD��u�<�)ݴd�D��Bm��$�4U�EY�>�wޣ`�2 ��Paռ�dv��H��岸���mFvZg����c��4�
����6M��ȷ����'0K��a�|3�a�����׹��V�;|�Gm����9���6 ��B��5Z�6�g��}�5���F���|OƲ|�*��0rY�">�2�����>��1P�;�x	h`KE>݊]~�v��Y|�]�(�R�*u�r��^�6�L���Io����y�K=_2�H�RpF N�$]I���?AR�{p9�d}������V���2�C(�@x�# �D�0X���还�T/�����˲��ffd࡞s���iE>^�t ��3��뻑�g��x�G�Ljn25�-!�Ξ=ٷ]S�����R�g\�3h���i� g:t	h�v�F1� ��*��c�@T�|�T�aX�Rn���¼RU�=+,&jE)� d��v>�`��d\�����^�ʙ ��KX룳2���E�v�� όMI�"�dFC`�j�"J��?_�:S�>����sυ�o�eɎb��J�0���8\�-�8��n	
,���_[_:J��&���K5��>qw?d@�j��-pU�����L����H�/����Qv0�kN�"hz�	0�ZAO��K�ȅQPp0�#u�����z�]����Ζ9�&v��ܐ�
[���0;P]�l�{��ػ��=b�&Ϲ������{@��mL��5�H�RxA$��6J�c+�қ�.@G��옧��T6���X:�O7KG�
��M�`��dDu �����z*�Ț�gE˙_�ou�ց�,�Jْ{�h�e�F>��%��	;�RER���B�8�Y㑊ge�D�oRk="~Rc����C��^�����J�O�B9C�����L>�v�� �Sg��+Pnq�X�5)���w`�g��.F��2��hW����e ����E�:Gc;�?�".`ō3��.�-��j�_���b�0��LO����ڴ����b��dx_:Oa��l+��7��G�
cC�*�o�3��˼�lx)>cT�Ci�z��u��|n͖��=i�ئ�Uf�o���*���@�ù����#u��s���4jH�����{�\�%�_�	��'Q���{�9 ��Њ堊Gf�����ۆ�9�z�QGs��i�@R�ba�!�8�M�|#�F��KcϠ�hkW<:>��60�R��s_�D�"V̯`u-�v'��U'�L{b���xN����%%�P*����Z�lcɻp�������R�e�k
�^�(5ƘP��ǐ��~W�o����ͭ��T� ��a� Z���Mз��0x�)q�`v!���y�|��5��r��!.���|7�e�M�sf%Q=bU�f�?���7">�1��ϰ%�\U��#G��C�e��)S?�aJx?c��5h��Σ=�v���'0���/&e3��ǌ��^�����QBbW����ʈ]���HۜXi���QVd9؀Qw�p*c���6Z�:�{L���J�����w��2v��:焊je��
(a�by�������m������(��'�9��_=u�!�`�o�U�c��Χ[>%��#�#Xm+Hm��	��A7|�J7���U���d1��gOB��,���S��I =&�X��]�������ץC�]�K�;(��W�g^�X�-p����$�d���y��$�u�ġ%̱/qn���!��1���z;�F�m��b�"� z��wId����	IP��{�+`�n�Xg��Q)k�	���2�O�@%z��
NL`6�h��nK���j����K�b��ס�вA�w|��^c�血��� ����zr����Ŝ�54�?e�+����a��E��M3��*PD/t�hC�{e
Z��F��4`qmZ�C�+��o$ͣz�puה���,mَ����&��y�U�Eu�d���t�L�3s�(�e~
�0�F=o�&��� ��t�.7z�m����o�g�@��C�!�����d��f].\�e���Пͦ�&�w]����~0n��jOY��$��Ʉh̓�N�v��"��hu���L��ҝ��PH<��-F�P�o���z�DCx���o�}�<&�Q��A<�q�s�o��*�6��N�1zg�_�����l5nJ���6�\`�
��-f�5(9����5\��,�t�^�x�dF��TXRx��qt�"Bۭ
_�Q��w�Z��<y�& bR���(�7T���2�H���d�� Z��=f~��m�%(-
:i�C~t_��k/I��첢���i?zR�%�JO]2��yP��ߣb���{�-�|�
������T��T�(�'���/��f�ST��F�w`3Ps����m�B�j??g�X�R���t�F^�&���k�d���1�s��`S���+�N��J����?��~�9_gL��!^_��vywA*�g@�QS��0��A@r��p��K�rىOǌ�+�aY�G�=*]g`�I�����z�QO��鿵����ϰ/l���L�y�2���~�$�	�u� <iDg[z��`(&&	���iLT�v�z�������S
~b}~*��釅l�d���޼9�萯�j��DP���jYf~#/�C�$��V�,P���ݸ�U��������>�*U�rZ�ǛEJ�N�}���p-ǥ	�>��},�5��,���JJ���mA��]'	GgY@�'���`E���#s�7�c���! �a�f���h�]ch�w�D�t�"�	Cܫ��N�n�ia?����N��<�O^���<Ҵ���eb�ġXKZ�#N-���>- �B����b�<��X)Z;�>S�B�K��	�*��Q.z0�G9�e%z�h֢�P�4=�B/b�
u�x��ZM�}�D�L��2����ʚ�98���{[G�r]*46����t�.1��e<��k���b�w��#���l���yLЖ"�wX�	M?S8~����u��×��)@��F��*0���:�/��/?$�ܬ�ډ�;��GG��a�8��mF,�Y�ۉAb��g�˭�\�N�C7��l�&����Sn��˲�o�Ԭ'�9ԧ+3�'�a�W2������ӡ�m��}a
ط�$V:���1�;��w`9�S�׮�w�Q��9�����
���>s�֊dﭫ�t�Q��'���$�J�a�@}������WЅ8 j���<��_o� ��g���7Y۱�F�" �H��5@��-CڏLu������-g����z����ȸ�)f�ع/������Z�6��-��ze	&Z����b�iק��i�nOi�Z��@�JZZ�1le�u'>ᮅ�d���z�m�pg#K�����9��8cJ����;�r�q�S���S<G�Ѥ�pژ�8J�!��/X�0lX�����+F��O�?�)V/<������J�q#�{�x�^�8���8��TfH����(f�D�ԙ���kD��+R]2�p�=�7T'�X�@F��]orc��s-.�r"ÆN�T]]���n:�O&O�=��@�l���5�j6DGi�myJ�{��xYM�_	'���_R<�A�����
��'��j�Hc��|��Y��X�`ƟVeU|�)���dJ��/?��In�!�(�7�������>����C��G���3��>f��m�}��kc576w���.*��l��C�e:Q���2��T�{G��&4�X��؈��+}*-�A�����h0*�6Q�����|ۡ���D@��� ��H��CX�p���`2�ͤɨ����6�#-YD~ا���ÏE?��R��`���ۺJ٥�%��ܢ}����3�;.  >�2F�Q�~��,����_J��Ps��f���)4�gs��f�.�RgEE��}�3e�g xgV��n<hf�1�����c���'�v9t��RG�=c"���n�O6��4����Fv@���Ͻ��i�f8+�Ɂ�vF"�f�8Թcqڃ~2��T�!��©u}Z��U����
�Q�l����%׍��4Q��W�*Rç*مx	B�ܭ#�E�@�.�F́�\�ܬ��1���ͣ�}B�{�L�Kv\�P�̇�^}�
w>��Z���&��;��k�Ƨ�Q^�xs���np��@w ,��-���*?P6���Ŷ!^��E�����2
����Ճv��y!�̷�|u΅)Yn��-J���NⱩ�}�+⦎:�ezO�\�l��V�%b��!�_�|��r!S���|,�\H �����fhy�A*"�?�=�j�v�]z2�~�8���x68��qj����4q��.ȈIF@��N1Bu�wp�L�_�ڔLoR�J'	A����7(�@CȵJ�E$�/5�Ϩn,������:'��7��n���,�,�ջ?�V*�n�"F�Q!V��>����6����i�@W��GB]B��Ir�Yv�F,�����CȳE7��R��8�|?)E|F��|k'�R� |?���-��������O�����&Sƨ$�&'g2\k,ڀ����p3��@�+�-}�a��Q�욼��u)<�	WB�":1~��W���DS��?�ꎨ���� 
8	}*=�ݾiC���a�!{���7?3�~�8R��@Qo�?������ mĻ �h��xhխV»gI���&>�V`Kc���u��R�C3l�ר{�A����x X6�B��c}ژh�s�Hw#|d&���WGҴI�E^E����R��xPwh'KO�bMF����'me,���3�H������%��7˯�K!ۊ�S���F��y9�jVȚjs<�,�H�+�?@��L�jԌ��GU���]65W�eb�����кg�Ϙ�RW��H$�RCB(Ǭ��C�nVek�����ؽƀA�tQ�;K�M��;�z���
6�(��ۤ���lt�i�b�6Zm��b�JA��p3o��/^��	�ԙI�T���ǭ��Mo��;��ұ>LJ��xmZn��^���a!���צ1.r֍����2q�Ue�rR��ꁾҸ�Ԥy�|�W��3�y���2V�����PV}�>��.�K���ݤ���{w�\�"�Pr��� ���)/�r�"�1�I��c%:퓕�;�����)ču�U�iWp�);3fKB��(�%�j@��np���̅\����A�^U|�0���:)�L�+�{�C��Q���g
ڵ�e����kF3�X�o���
\���O^�|pL�)HX9��?���j�P��[�g	Ո�Sj�� K=`,�n¬� ��r6X��������l�p'�I�
�2�۩`Y|+J����ÎU���O�%��UtW��&���^����F7sB�M��lb=r��ۻ���kI��o���"���S��� ���b�@�}G��Ii�6����_\@� �D'�F0��R%'�k�GS$˔$�ܟ/�O�|�=���#�ѓ9RX�N��a^�U:h�Z#�){��X�0 �Xp}��Y��>s�;�l����(���#q{�^	-��\�zb[��Y���_Hn!S�cz�U��XC���V�w�ɤ�>F�p=O1�:�jW�
/��3WFF1R$=�
ɮ�O{C��{Z%ȭ�����gB���T�7\��IT�F���t_�fy~��CKŋķ`�h�AՁ�'���EO稸3)'��ѯ�謏�&�_�����X�k�������Z��|�Fh�B�3���Bz��B�	I���3&ܮ���J���0�G���(tU6Q�l�75����_f���$��ׂ~���M�*�����p�$�l�~y���]��eK��:Xd��߮3*��d;8�{�`3^��kʐ36.B�ͤ��q�<���v��;�����/"���yA�v�b�:0CS��:���H��vu{�j����kIN)"���5�V)�����v>�Ue\d?���D`Ge���Q\��h��ʷ1�%^굍����[�)G'zLu7�Ŷ�8�A#=��T	�x��ɞ g���*�^��V�����x�U'�@b5��Z�9�e�%N���]K@G�]7z,��.���L�f!XƊ�N�0���(SA��G�<mF�>�V>A���4~a�?%+����@�\��y��v��� ,�I��`����4"���O��O��_�.=��t�P���q/�4��l[�� ���ت$t�	{ؑ>'E<��?���>���q��y[,�b���ǡF�r`�2h�q�!ݽ ˴�m���h�:+.��He�ҍ!m�ٟ��P����}��QP�Jp`:�֧��2W͝�l���8=?km␑���Z�b|��d�#���J����J(�TK��l�,����IbV��~�� bxA�\�W�3�&7�����9mvU��*
��*�]��齣?�vb�K#�l��,��7��TTX41!惄h\�������*\��Z��V�1�t�<���jl՟��j���h��_�T���1�^�-7k�*J)8�Zb{=jB]��o�cm����[j�'z@Ti���wh4��h�[��s�y�|W��r�-T��-"t���<�!H( �Klj�eXLK±��2��ld���@�G�FL������T�z��v�����X�,�x��G�vP��	����3�4H���ut0�,|�G�x�����DQH���][��V�',�M��bd��r8�Op�/
W��L�7�a�$�h��#��%>�V����t?��AWЌ���y�)º��]���>M	M�N�m�6��1վ�Zh�3C6��T�Αp���b��o{���1k4r&������(�͙�*bM�|/-�3ōMhA��(+UE%��'m�;�;#T�?X�c9�*��S A��S���4�B�%h���c�;{�n��g�[��H��|u��h~t��<��Z$:����W ��d��	�M��\0�1��s�eW�����~����pa[�C�����>�,Q�Z�i|���[�q]d�N	�[�b��^g�����zχq�����Ǆ:��3ht_�$3�B�djً�r�(?�ݿ�)3!�z��|=��d`?�����GX���iaPE;�t�����8�����_W�Oc�~9-5~�fV�\w�_�1m�<�C"�	6�����H0 ���M����l�<�*�dx'mVܠ�t>W�dBE��?���Tf33��!��,�8���ߧ| �݉��E�&��يCg����Ɠ�/��j��Xn>F�uv�]]�	oW����E�ZR]�â�.�bv�wյ�� %QDT��6�;(~ǋw��k���m���u>v�+��7��j�?C�`/�-��.�n���<�[�Jl���N�ɤ~\��1#MtA}հޓ�?��	����颟��s�zU{�.�!��D���`ʣ���NW��yߍL��/��W9�ω�uwn�?������f���L��?�<�*aS+k&,8/-�B=�x�2���FM1Li<����/�8#BnM�n��?�ܮU�ȍi���<�N�C�a��������^�EumB���
�0�=Ǘ/3�q��������.��F��Z����&ϥ#W��i�g�92.�?����F>���H��l��Q����=�&eI	lP�a��G��Aw���o.{�%pp�L!n�����}bA9��j�lwrrU-u<+�A�=�9��fl��.j�3��N���Z�jC'Ө�%8��&2�{�ǙZ@�lHX���X�$ ���`7aIȂ�:�U�Fs���T����]��m[�RR����W|?h��XU���d��w ����n헚�
0��T��ᗴ�L�S��ݼ<�M����w�@,�O~˃y���IڂJ�g���ˡ�/4��v�V�-ڐ�EI�LcB�T��J�/$ю��w��~X��F��g�l��Y_��R%	��=�9~�2�L��漾�D}���Ba~�1k5�U�V�Я��Ӱ���/����a�E���b@7c�-���u���%m�p�vƃהB��[b�5A0���A��ɡG.�_J���r17?K����`�WXs>(ڳ/���b��Z#��%h+�U�L\]ܔ�s���xhu�Ě�\�w����g|;u]Of��ۧ~?���LmhLK
Qj����LK�6��9]"���"�^Xn:}YG9v't6�o#��ׇ=��lL�|�[O������N��D�,��Z�
�_��<za�|�g˲Hh�%���s]P6,1�JA�i�q�������QMk<ow��h��d8�	���yPQ<Q"�^�F�[d����<\��H�l{���	L`6�N��P(o�]d�[��.Ho6|� qA���M#w�ni��H�^�{�8=J��/���#'�F
�R�������|o)�\F��f����^a��M�6�-sf:�pM+���+T�s����X�;ڥ)��{ޗ�?"R4%�"�e�i?  l�"�M����� :[dn�0���'���m/4��x��e7�WI�Ca ��J���3B���ѡ��G/����HWB&�ܨ����][,�'��P�Yj7$���G���>���>nb����I��**�Nf�PV5���_�G���z��-r���6,2���s����֜2�)2w�ݮn2E$N��v�+b��5Ͽ�
��zg��1�+��x�����L� (�����XE{¿\��K�I�·XQ�NJ�S{�9���a��?����l�י�|�$L�D�5�Jt�=[�f%��3V> \ը8e���i�;߬�*~#/��
����):�h�9�jY݊ւ �	�R�K]������Uz�c>]rԼ^�<��Ub�ҍ�RAE�������(S ��r|��cUm��;q��⛻V(��y+�FX L�)n�W�w�^�=�-�0|/�v\���"G��Z�>i�΀њ�s�P�����Zk���0��6 ܪ(�@ CI��{KT,�"؋���|DE��Lh`�һ,t�H�D��?�S1^�@�e�J��0�s(N�C1��a)��,="G��0�0�D�(�Ґ�\��%�cB�Bȍ�<_��?����d9ϔp�k�S�T)�� ��0��:�2А���?��{j��:��^G#	�y��9�v�FN�q�0��s�?�A�Sp V$T���������D�����A�7sN�����I)�c���)�)�a<m�8Q?���[�W���W��?�P��qn���>���:������4�'T�E[�o���C�֫g���O�T��v�g5}jL���w�ă5/bZA(�B�"i���Z���P�S>�l7��͒���_rP�4'��T�Ҏջ���81T��E�s�/d�:���5L�rC(�i]�a���p�tŹw� �2���&r~�򦸰P
��+��ʺ��X]�����'B�̚��Pķu,�C��떊����Os,}o}ьh��nh<E���-��$ـv��<�(���mQ9�p���Z�oHwd�o�6׳2`S���E�O�����K,�7�鮮=�y�L�тj| �S,�~���3[M�����>�7�R;`;1���nsN:���SE�������p���ƫ�0F�{������c�EX��I��h�6����0������X����B��m�i.ܺ!���� �X֌�+@�Q��jΪ t�<8�\���,�E�s#K�YcқcyXS��%G�;��k�\|�zSF�O�+�u_�rL�O��R)-���C�U�H��}>a�Q��{q��)�edb����*�`����KAC	���Q�X�*ھ��ҭ��a�k�2�F#�������/�^bO�),�f{Z���g�wB����^Ԕ�V>�E�fk�/��;tO�jD��O�0�)y(�"@Y�%�\wS���h7D��検�;E}k+�A��9���J���~�=�4eN��7��E�Lt�V{�aO����4�������K ��;�[���O�3?�I���=�aJ�S� �މ�1ڑTB�)i+��_2b�*۾;�冨(2�6�о���=o9�-���p3[ʒ�1U�M����CEB�v����
6�Z�v��k�sY�"���}�Ce��.���m?o�G
;Ј�m�w�؅��/v�>@/5fv�8����� 0Ǒ�I-Y ����%v&tGR���xL��|h�"�u��e�[��G}OC��o�E܀ �`1=z,t����M�i���U��ymJܦ|@ɤ��i)1rܷ�IK-2�h�@?�撣�#�i��p�ێ��ϣ���j�� OXg�ņ�[H ��`���TU!؞�yj�:�M�izک��.���~�� �5��Me�S9G��k�؇�}+��MS�.�d(sC˧�`<8U���t%�)��n�$8�3X��A���x��b�5�]�M��%\����?�~'���[ M�aф"x/����W�e�ؚ���6Ot�?<.1�����vX/|�ouz��aQ����m6�=@�y�3�a$l,����!�`z9\��J��D�.�R#5%����&�B��t��z��9j�3b���i����CLĄ���f��J���֥�AQ/�?�O��h%q�ڝ&�n�D'�lͮ�&1�gz (����c1�͓�?NP�v���?Ǭ���kL���_w�4���u���1����\���{�H3'���<�Ń���x��7ۊ��{�L �]tvզ��Y��OQUp�V�ٯ�|5��+3�ci���8��Z��~W�� i�<�獤�����`�	�7XYX��3�[8e��cg2e��k�rR��.)�d��E:X���d��,j�w`��t�<�g�D[����Q��#`�V�՟4%�E4��8,�Q�S�����R����A=��Oɺ�R9<ɚі��P]]-�&c-f\��8��&�ay^YR�,���K�.�N�0>K�b76�?��9�pvF'?�&���SW�,�>�q������졌*�A=�b�g� ɾO?��E
��c��0��₫�14@��c�w�y&_:�R/�� ??��tl��ޚɌb[�q���
\/H��ul?���rnIڱ�q/�L[�~R[��A��t���߁�&.�w�J�#*�"]�O�M��Ұ�pz�w>���]:�蔁���^���Q UT�]_��6W����/�+��aBoA�m�Ȳ���#Q��S`n��*����_h@_�4&���Rl>�wk�G���P��R�t���}s8��U�Qݫ���b��!���d��%-�����lt���C'�Lu_6[a,�oZoW�K`��1�Is�g �|uj��k�F�J�hw�ө'8�Q���turW��^����oN���K�~�s���8۟��DOGC4��-�(O�'�r�[��	��d5!�5�%X>C��?��1��'F�@��������7t��I����>�V-��fC� �k��3w���'(Sj�;�>UK5(�EC��s�JrN����5*��MdX�˜��!�	��QC�u�����1-Nۿ|���)��7��a@	I���}�M�mu���G���a�Zݍ�����c�)�;)ۺF��N|[����5�S�"�YW�>Eo�.�1�y���}k�+tT7�P�B)�������5�ho�+����5���ֱU��{1V�?T�Mm' j��4����+Fmṕܮ)ŕ��i4H!�av\�pzٛ�����TF��Ze�54�4	�I�$�%eq0�3`%e��o�3���%�?��#��[AӶ�Vl�y�xPo��OGyz�����l��y^®Z�^tnm;-C��_��o�}�(�S���6o�VJ�s��CX��F0��JKpn�����l!���_�i���o�|֖��k���bG����`��FV�'������!Uݰ�n����ƾ��	벾��G�Am1�H:$�o(�]�jg=�/P��;Sp�aҀ������R�
|ե�
���L�	jjU9%����ʞ��$d���m"m7�-�v27��6*b�]���Ỵ*A��t�4�Qs4��1g�ź+ܷ��dR|�ɵ<^��5��;� ��x�#�m	( e-�W2�v���&���HRe�:a3l�`l�(Z��s�)���U�h0���k�|t�)G��₋'l���\��CL�YT��Lf���ʱ���l�ͪBzB���&-;�[x�dm�?��}��I���j$����=�oC�=��-�p�#2֤";���)=��Ȝ߆t����g�S�i,�"@�LA��
xM�b�gs�w B�ƤDM�u h>���x2�E}��AOs�e����?g�4��9�#/���ك�3�Wd�C�����%n�O&�0u�a����K����x�t<9_ɳs��C*��tӠ���|3�,fv�|�|�`���G��fT�[/����YXV�����@!�:�&�f��ee�{"�{�4�W�L[��^XR�
��Yb��5����./��#Jw'Cq��~�tˮ{�t %���&e�w]�7c���G�`��X�A}�י��˥��)q+T�#��z�y��`=�8$]�g5�+]��&\}�����?��tpS�2�E�,����FC��_�x���ֵjf��H�3Z��}���H�H��"(v��P�*&^<�z���o ��
Nl[�L0����vB��>�e�q[��'��EBy�BE%��i��_��u���-=:*,��Gۈ^�jM9�\�O_�*��&�]�9�����Ͽ�Xҩ*�=�:��]1o}�K���~��Gǁ#=��	�y��%d>k�A�?ތ��q�Z;Hԋ��QR�d��?O�c�����[BJH���L�|#.�)�'�Ac	Dÿ����ϡ��F�`?U?�y=��s��uLVE�{�pڲ#%��
_Q%nؙ$��B����1�:	o�Z	��x�b�6˰���	o��͏�}�_umM|���? ���I2�h��������ā�[rf52�f;�4�ε�~G����h-hu�UJ�x\�^ʤ���.&l��s�<�`��Sq��k
5M��4Z!�����}�r����'&���V��Vv�ѿ�%�!��z��h����*;��T=X��K�/9�/�� ���>�W����BD�B%2~-�v���º26���l�����͙�C�������9Ș�[f!���+ZC��ԁ�)�tM�܀[�����jr�,o���+z�i]�@���|핪��c�}�~#��d�:R5������l����
��Q��rѾ7	o4���y��j���V$��� ��<���NDLW��S��	��<�	U���!r�G��n)��Ip)�d����v�{��<�a8�9]���h*��+ �V/�{�4L�+��(����jaNf�ZX3>&l_�Yz��fg�"/���	���D���-�O��mb/N�����pB���Z�'��;w�j!�s�k�T�:�P�m^?n�o]�����'����>�W�G�W9�?ho�秺Z���Ӊ����,3
�)M\x�9B~I@��VZ��9JY������K�w�ڽzPM�� ���qS=����⯥��)�Oǆ^8��&�Tx�9n8��@�����/"&]iVl�R&\�+ԡ���3��H;8H�W.��E��zyBiZ��Qk.�sHL���t���Y��n&�����eg�.Q���Z~J��B�^
�>}0���~�
ڶm`��ڜ��_� �\H���Gbߴ�ێ#jY��ݱ������\���F��D�-�S�g��R)mSX����[򛝾�k�t�X��<=�{k���_Dn����b_L�E�=��8%ⶍ �]�ӫ�ʸ+�k�f	A���o�|�,����d�Z� �x��
(x:@C�6�}:DRӿ�(�5Û@��l%���Ml)�01Gч@��J����Z�<6r�FC�E:&땔�x@��ȃ��3A�Ňn���tCM����$i��ms���H���6�3ge�}�ܦ�R��3赏�N�b,�b�����p.B��W-�̰N�-7E\|X>�|4�+H�a��r��Qp,�Ht�o��٧2I�O��Ki��k�f�y�����Ōw�w����Ц��m���ճ�H�\b{/X.��ޚ����`��p.��@-}���"u̵c�R�b��(���i���"K5$.����T4�!�����ǎj:P�~<i4ѱ.���p���=�U\s�6(�?�*]�0uk���$a�E��)��Ko��R�{0�g�}��I�����E��]��Gąt!g�۲��3�W���i���԰��p��I�XY�(���|ܙ��V�M��N�S߽H���k�ځ[?}
�,Rʧ�Qˊ��RBܞ�|�R��d+%�W��t����x�Q�±}	�Ͳ~��V1Yn:��)��c��v���o����;L^V 2��	a��43d�-��&OE@�S�G
&�1�q�:�V)u:�<�5�1�/��D��������Iʁ���sJ�]R�8�D1���
���d��h��8��`��b2����/aR10j�S���n\��haT7J�B��`e@��Hέ�0y�m��}~0-�3�������I�g�RȗoN�����8��,�d
gZ�),Q��!;��я!���u��ү�ǳ��_�b��تk�����	Y����:�%Z�k+s���b�f<�����+l���_�����7u�S����*���m�7�#��A	�b�4��f�3YP�_��t�?������8��G#�it��>eK���]x �#�#�a��J�M�|#A$na�]�+'�m1����N��e��_M��z�y�|���O�%*ȫ(5v�Թ����W�+�O���9UG 8����ޏ��692�V��|�3`%	�	\f 
7'���@�5��ڊT)Q�6>�c,����-�(b��fBb.]�#d��`��O����{��?�#v����<�e�l�*KG)��q�"2R��lI[}���c������[y���m=�%�]޷(�T+כ��g��t,
'\8�4Q׿��X#�F��Н��r�`d�W���Ö��FPH_g�_����K�.6�|�1�쉿��	�pC�zN���ʮ?���a�?`���}���d@���a��O��tY`����:������zC*7�0+MQ�$�TFX��WӮ�u�>kR�j�����ʞB�刱X��l�j��=�G��ã�s����N_��P�r4E��$���2k1B��(l�v�[J�"�=��ZTB�$�f�T��ˎ}'�F�����ı��g�ѫX͠-b7�H���~����$�d�,��3�<�tz�j�[A�C���E�Ž�y/�}��j$�3g1�L�8v$i
���m����g�Ul�	�a�=|�xܐ�S~q�޲[�+����
��Yw���Ӂp�{Jr5`�M��H��P��Msf�h˨���o �hE@����=X����U������{ �i�1Z6�^�;JU�#��
ڵ͗è���C��X)��hYb���z*�v+��}�� 9���>�[E�y=���
B��cjӖ)�����W�x�̝[J���U��l�<$�J[��Q�uf?[槖qcz����h�_'����`2�+k՛����E䌡M7���}ځɠ@�J�|��"fv��<��+�s�.�T����D%�;я&�����-��������PP�
�ܹl��ߠRXy�Q�-�5�H��P�v0���W��~���vjN\�O��������֒������	[�CR������E�]#$soSA � )�`QtW9c�'�4���+���n�=��Z'?���UJ�V��d�K����`*}v|e��Hf�3�_ZPi롮/�S�i����w�<����#��?���A.~W�:�D=}��)	L)aE�ԇX��.i}�pзǟ�ub�h��I�0�ʵD�m�`��ji(��8.z�}o�q&�O�qL��rs�b�P���B�o�ϸD�V���:�.X{]۫k	)�x��hj�;w���t�g�+�T�;Ϩp��*̂+Z�P�\T��-�,�Y>�|��_�:�D]��Tm;���&0�"K��cȰ��P�O����ri�1��ޕ�bz��ww���6��&߳r�ȟ�Ƭ��vN�a3uz�Jq����}8�.ɣ0��1�7�
�M�"Mr<@7ҏ��e��p� l��J5� 4.-0������������]�D�q{�6��d�錝�U��ύ��i�U��F1���-��-��Tg͠ni����s*P{�V��J~m);`�D%rƣE�~����0\>V��R�U�VH&�2������g���T�T�b����G-Ů��e���1�Wз�>�9y�.���`�!es�s��8=z�$N:�TRKiO�,�Ac�>mM3�=U4U��TE{�ޮ�+Z�1K�����RvaPF.�L�m���y���d�C��U2��+Z����>G�HL1�j��0ncw��y�-��,2�\�X��{���! �uM�sm��N}^◤	t��tiq��3��7����� ���fƃ�U5��w�R�ֳ��G8�{�_�{�+X��I���,��,Xcݮ��j��؎�;�����/'pkQ��!��>��,� B�*��2X&�F�{�B;.�t~H2؄X^��PU���������5�S5����J� �7��`�4<_+cp�@�|����s�-M2 @_���n����� µ5 %d�}��MP����W�M�����ǏO���
��������»��!�ߓ+-��ю,�؍�	���)�~�*�e�9�:^�/�3�������/�W.�����v=43&?�E5;�fOD�K��G'ޑ9�D��0G���^t��T���J��N�I�鏪o�p�)�A�"���V�w���"i�o�7���~ճ
<v���f9�\O~�.��'Mˍ`D%�\�3-�b9?�!1�]o��$�����0j����lK��J�A��� (�_���k3��j췼(U=�	#q�����jI�j�ޘ=��⍳惷ן��v��f��?5�L����FG�Ld�S;�������)��)��#�T\�	�U�Ez<U�J����bu�j�J+�f$0y��R��Ƽ�j�+�'7$k��tb���C}�\�, 툑3X�"�^���|7ѱ����
�g��@���*_
��9��@��l0w1�ظ��9���KO!�a`nvN ~W~��MP��6N;J�-n7�5$
��	a�R�^�	�}�I���"r"LO�G��FϜ$x4��}NAV�H��y���:�d3����=5�n�y+ʬ�����4����7���Q�U�"��\������y��A��2!��2�R�C�&��Q�#s���'�����GĶ�@�t�6�#�f�F�G�V�NFsf31��%q���0�1wi�G��L\-����N���&Hp�m���ʅ�Z�1�㵝�g�MS��݃]A�Z����I��GK����k�y}6�F��)���EN�A�*��'*����M���n��	�F��ۃr�[��d�!v�tM 56��|óz��$�	
`�*�2����'Df�,�[�g�'1Y|<�kQ�S�����Ia;"Ax���ɼe(�7�ͥ[�Я��iyq�qR�#��!b�2���f�W� �}�1�� �4�z�{]��-����~Lq+�o�A,���_�	
��0�x7*�R#�����ɤ���d�:3\�?�jwNR���hu��+�/���]��w�do/��s�C��6v^�\	'����v�����e�|$#��}�12�+���c3�w�1�z���C���d��܏�5H@��.Hm)�ۺΰm�����_��z��R��G�S��r���rL������7>�U��/��0G\O(7br!4���<�L)(�F�������tv�u�F��y�tܡ�\�bDJ������ċ��K��s:uo �����Nv�Wi+q��n'?'L,�Ht�����^��Q`-_ L.]�R��ʝ]
Ɛ1W��KC/�#Z!K�<����P��R�4{�gg����ӌ���څ"�/o�8�J�f
r�IY���v��x���H��g��9����4�Ĳ��e������� ��ӹ��
���F�����cѰ�k{Gs���@*�RB���UEhM0p���z��x_��錸���@eD���(_�o�~���J_���
���-�'⣓�	$�:Ӊt����JN��Wi1
�����11w���_���Sհvu��Nل�='�@W���#]��ؐL1]A����^�8�.ޢ�&�v^������)ꜳ�A�3��MW8ըY��6K1�aM'拤n�$ZW�zy��ի��	VR�]��)@A}����qU%
�Pk�H���W�\�D|[�=�n�.z����{�:�	�'5�n?1�^��cW����0�t��z8�$���I�����'���TSO�5��p&*;�?�-�k��A��3��c@�SJ���;����b80V�^B��T(��c�<�#T��Û$��;FO����&}�o:e	�,���ˁ���ҳߕPY�J�����%��c���G������d�V�B���h��`,B�a���$̴���s!��Z��+�-}V��b���d,K�� W7�8����[�� �zm�e��xE,��?x��ߗ�	��{
�Բ���B4-�V9~��� ̡��qC�ǔo�f�#�rC��q|�Er]�?�4����l�s�(�.F]�<�ƽh���W?F�� ǌ��n�b]�'�慠{ȶŗ�'������ME�-L� #*���0}�`�[�#g�e��p3=�#��5����$�!Q����0��^�D��>�zd�uF*���p`Oxz���Ւ���2�'k���C=�]�c�*V�����[ᇪ�iXV��x���K�_p� u)ل��s�AP\�zОF�`���{����7�k\���%��@ȿ�:ΠJ?�,�)��C
V���И�)���ۿ;�p�7���)�9�0�s-j��X�V���L.r�)�{f*�L��gb愒x s�1>���r��1�!�*�ͪ�2VU�cq��C�U�B�� ��	Q+@Gp?'�x�,x2w�=�6�Mg� t��/���ﮮͪꋹ���c,��<�9�?߸2|�I�0h|H�<�J�Z8 ��Z2��	S�W���S�����|<����(<�ӫ��o�Z��N0�8w�#�V���Ym�]��p&�d͈�z��Kf�D���3�a�]�A`��Q��k7M�K{�FmT8�X��}뎅�V�Tm���x{���.�1��3q�&�-Zkw�����H�^ �U���_�1��e8GF�	��uf�4� ���T���%|R���~�?P���.�ʹ���4�w]�1��N:�Tצ&MD`�}g����3���]���m�;#tO"���{��|u	�+;�`�k��B-�tKt9�I�\��_~nԽ �o�Q�Iz#����q?�_� ��-t/dUc���������I(SA1n�f_SGx��a�Y&宂a��P֩be�0��fj�I���sʛԇ���4��F��:�[��^66�����j:���pr?�g	*�x�����;��Ux�ɷ���ܜ�	�}�)�XY4m��Wz���B���U��$h�jRbfϵ�(����7I�����k���7�� �$k ��sJ�u-��7�<�cS&������k�wUp�b�*���n5��yύ�_��!�,;DLƨ6����"��>r�R�<��Y%7��-im�+��z��f@�_H y��%�`
|�\���s}j[p��jEvt� �'��&�A=�y��>�Y��%������Oe�4&w��)|����h[+�Wq-�T���tq}D�e��W~���Jf[	Ҧ���N���40(�	hBN ip��<�=UVp�y�-ڿp�J�飲��[l��a���up_�q�?p�u�����9lu`�/�w��J'��=A|
�x����D_��� � T��%o�Ū����@~ϓ^����W��˛Ť�w�L�kh����{J�WE���vO�1����m��h�$/'(����! �ܼѭ}!~�od�U�2��\7j(�p̒`\�̀�x���/�F�]��U��bFõ���B.-n`jG�2B���I]�����֩y��ג�
y(`>+��;G�+=��B����%n�"꩚/Е:}K�BY�ABF���_(�J�2����σ���|A��L��Z�f��J�	jy��{#��⽿Da��F�>�����y��ye�"F�ڈAZ�G���~�EҪ����|�]VR���<��92��Z_z5M�؎eFu��7�)LOp�X*�n*KVY�1Q,b& /	\�D��F<���+۝XG��O�o�_Y�?J����#��6:{��u�wn�NP�)� ���1v����Bo�����8a��V�	z�����R��_�z�"ƈ���YK�}>�vb��	ݥA���Z�a�8	�n�r`��p[e�o�)�YJgw� '�|�J�*��69�
��"�������\�!�j�~�vR����V��Z��郤Y�m@�m�W�]݃�p%\BV�=�}��39{
� ��F�����@��8ҙ2��}Y]o��:��n��-P����bba$�~�~6]��&9���ɠ�ڞ�v�q$ݮ�N�]�Ti+���r�*G����X8/����ob����x�)���S2-�ϵ
ݺ�=��M0'������r��H�v [����Zێ)�A�����(����>y���VnÍ��]�u����`�se�qNpaȓQh2ʔ�RvZ賬r���U���=�_�l䐴Z
��s��]����3k�B"n��0bR!�.���sCW�p����&�hQ�t��B$~��[�uJg��}g�2�-A����INJ��Ǿ/\�/���O�A�^ᘨPG	��C<�w�������j_X=3Iy�9�}�)����2b�5�_0�#�=���͉~dH����9Ю!B��u=`�OW TgP�E��r��(ֿ�!�$�M�qCr1' ʈ�˭���M�B)�5�<0%�0F���2���T�����u��Ы9[��u�*��I��u8,���٩�����������,�	���I�m�0�E]~�
���CD�6*y�����A&%�⋻ȕ�Z(�9ɶ%!�tĒu����W�e��!�x�!"�qA<���N�Ԛ�=[����ɩ�C��z~��Cc�jη��ǭ�=��Z��`� W��2֥��eq.S�I�D+�� d�
}�����`�į
��^�#I�+������Y��؉@G�7>Ä?���نkn�T削��/RE���k�:+�ѱ�-�}j=��&!�<����:�SJ��4�wWاy����j��Y��CK�H]?%�OW��:�_>����HE���,��7�aPG���| �E%)����g��8�Z� G�8۪��4�R3!"���Hu�`a;�T.�����J<XBt���bYQ
���4Ydҫ	�s�pa���$���C�Њ��O�=mXu��_h94��~6r4����/��8H���1C�Ʀ���l6�2�^�_��P0�<r9̷�g���E}��!ڮ�V�2�����<�v:�+{�,rIԶ�����O�@�g���x6ݒ lbItͳ=%�	Y"��j�n�'���x�T�
�:@��%w�˛�&zG���vQv7���Wz�>��Ե���lP��bd��{�Q%�����aw�M�V�A�j��`�	���e[�N��ikTd���U���KxY���jw��WM�e��]~�'y�8 �*��ꝗ���iݍ�ϙ����!L�of�V���:��uW�A�xrB�p+9��`H1o��e�>�&��p;�������j�j�ل�qW<-A 2��/��l�9��~r�0��Z�U�yR!�b�(�k�E�P��.�[��3s/rGzq�	1�u�,_�{�gș������09c�@gˉ[w�ѽ�k���K���8yp���3Y��cw�oW�����K��K{}�Z{g�����e�V�_"~���Ӎ��h�4+<5�rf�y��:6��0x�7�t(¾|��VH@ʋ��;���>�K��M�IO%H��ة�?���ۼFN�(v�~�\|O��9��������/WA1H�}մ�0	�B�	�9�	�8�$#�g�kR�>kYE<��XާM��Qb���93�).f��7z���4�5r7�VnL5
��}{��?ڀo*x,�W�A���p���t\������35�\ �r�����%����a�hI�}����% ��� �*��X����js=3�2��p��Ʌ��O�T��a�&/K�n�Y]�.A��zA����BOߠT�f�~�Q��,�R������A7��S��bGfeO �59�=_��<{�| ����0��R�@ƍ%��x�8���Ś�Q
2�V]^I���A6�A!�f�p���g[��1f�%(ҍT�^`V":Cu_��|�K������C��r;�o��<�NY`�4(4����tܮ�I�֪�	�m�<�y�UCs��^���?�H/����ٹ��zN��c�.Y�Z8��n��z�-��fC�f^��^�#�S�P`����B���SU�Z��l����>�#4�\���_�[�ڡ�jy�V.{�?H�Fӛ?�|�z�)/4��G�6HrE�z�(br�ǧ9�`����X	�[��$�� ���e-8G�G�����I�GkS�j�2O��1���s����t���(��A���oX)KQ��x�6�2EɈ��3b��{��URΝ����5ɕ݉��q����2\3���'2��gIF�ãT���	4�3y�h�qP���a����x�QQ)�j�Nq�.IZ(䱖�~q0���M��>�dQ!R���+�g�"6�X���bIF�
�,g[�H��l֙`����Ĺ�e9��1�+{�u���R����lS˥��O��(��  ,�h���2�+h�.�(ɥ%@�"�ȩg�k�ѕi6�����ŔM�b&�PIJW��C��E�aD���D#'�F"�ݗ=�=�)���2W��7����XRnuh�O����O��g�,��..F�~I�I6�I�#`DvJ�΍I�]C���M����{4^��X�ØlH���>�N���S�  ����a�z(���޳�G�Vm��e7�R���X��b�/�\,���&]Rp_�P�|~�,GkD�X^�[��@��g%�E�O˴ԁ0�UV�r�  rD�W�.}y	�|)��ʜ5Bu�C��+�Ѧ̪$�Na��V�����z�^�p7�n�Vh����D��Yk,%SRÑH��UA�ᾌ�*:�K�7E��=��e�U�6�Wv�b���u"��v-�\�W9�^w!�2xYX��.��&��y����oW��g�	*6m&j.�]�=��m��d�p�al�O�a�&�K��v��
*�:M��
l�0>�r�o��>��8Hn#��*)��k��^��C����RI��.�GޥZa���q��o����U��=Tמ��q��Pi�ϗ���[�,f�L��t����Cg����0�(�D���`��@;��}2X��P�U��Ē�}I�@��2aE@wZ�zП�](�� �]��.�-8���&b� u�A���n=Y8DP<e2l�*�8�8����p�����'�oϖ�u9�6�W9�ؚ�%r�q�!ѝ�3l/q�����E��<���i�[�K�� :X��`b�d��7'W�}�C���"�
���)`�T�wW�+7�Q�����k@�|@�'��t�w���A�kj��e� ˋ3B�}Bִ�(�����m���CB�O��ls_ ���M�O�r'����۸�_Y�Cч��(��4�O`�M��e�|����E�194i�����t�N'�s0X���rZi�g��5��3U"��p0��gs*�DQ�gU��/$���y�~���N�Ll�5�
6,FW=(h������s�Ob��d/�K��4YZl_{���,�՘�ǩ�`ᗻ�3�X<�1��|ݏabR�c�-�*��r?�wv�]ن{����&T�3��}	��N3T,�V1�>�珀�\UDX'��o��6� 3+�.f��b����7�/1z׳�^_o��*�ٯ<z����zSC�CJ���9|���&q�c�����h�����]>�k�C$�<�,�0�r�+8J^Cb��%�]�r����V�<�������X�Dg�P�x���S�{ z���ʴ�L�D��#d�0�p���Z'�<6ܻ�c�0ϕ��6zk����foQ� �J�$:eљ�}f�~�*�u����-A�K�CK���c8����~a�j�0����NLd� �Ci�ٙ����g���������k�._6�Tyb9hl���7�/'l�[d��6��&�R��M.\4#����[ců�P�qڨ�R�Χ.�G�+����Ѷ�e�`[pP=h�����2�G�.{ҕ�u���cֆw�:	T{��z�~L�lP�r�)^���~0Z禼�1��M��>Ѡ���"�FѶk/�B�꘼
�~��<�pZ'BZz	$� ��e�A��;���R���*3k���np��T9P�<P����o���3,�
4���T~=k���qԭnx�|4�p�,i�V�0�3
�ԏ��
n5t���S�/ν���-�����)yx�Mh����$R��S3���<;ƙ��x�(c�����qd$�����������ý�k-YY��L:�,s��=vQ+��x�
;gY��W���k�a��&UC3� i�5	��H�Ƴp�:٩���a!� ���u��t)����$�E2�j?�?t�V�*'崞�9ѣ4Έ\T��h��#�蝧M�M%���X���!B�;/���J�a��$�;�%��U_��*nA��Df!R1�>�xj�J�)D��!�9G��Ium����Z�o��bD#���z��k/W�[�X:��kmԹ�i$$���
���!��EOj�O̳��lg��miP�(i*����<QJ`�3O��W�T�X��ׯ��v�JB2d;7jו�.*#��|�ȥH6�)�y#��A&��b�ʔ�J�n��D]��f�x��g6�Y�\��X�� :O�W���BĲ���\8\�D�L�@E�L+cZ���
���(m�s�♤�/�'3�o��:�[~i��y�@���CKG��ϱ���/7�0R��EE��<�^��R��u�h+�e��♊�j���XR8�f�ݤ���(� �s�H^�j,m���Nmw'{=��<�23%�J[vD�^S<�+d��������$s��m�l|u�m		�/m:��@�~�v�8MsM�y�������6��{>�_z E�u��oAzm�4�"�@X��C��
�`����{@���a����0-�m7�Y�,p9.`(�z��6�?�Zn���z�l�%���ۄ�@:�qj�m�=�f�P�G���vK��	�S��aA�$^���<�L<���l��v��t��
R���x4,�ViS��e���@�x���?�m�:�#��9���PY���[���pEod�7�T��E�\fz-��̫B��=����{�?S�H�%k�� ���.k�BJӶp-�<-�T����R]����v��=�������?��'�s.�A��@JEJ��,@�;N��JG�)*�4�N�)�ܷPc)�R���[r�Y6÷�dm� �q�Y @�����F���`���yHR�L7�5�S�Q����V��#��/���(k�G����W޳L��~�Z�B٢ӗ��k=\�b�lc��Ԡ��$"�J�������i�G��������4���0��w����"5�A�Y;��,��8Պ�n���?��!��Ƭ��\�~�����9�
P��?�&~訇,�f^a7(Y�!�`]�V�%=&�/�t��o����ŭ)��?G��a��4T|�xA�@��@�K'5���A�y$����z�+Q�s&	�C��~+����%>_j�ˋ����`r-N�VΗ���J
���� �
��E%�m��uRjL��n~�LHOIx�D�|F�{�qEZ�a&�ݱ����e�(���.�YS )���c�z��FX����9pi�l���q�2���md����LU�N"!)bE�{�7���α*sGzbG�6��V�� aKy���_��dL5G�&p�<���l>��������"�k��Z,�g*�3�F�-�� xy�s%�p�c7��e㭣Y��rl�x*�4�@H�U0�3����5���y�i�B�,v�n���5dh.;�G"���N�9m�N�����J�͛H��@㢋��X�E�_�����m��0���� �f���\�5&�s3�@]=��b����X6��@"�;&�$��m�A��_���!�վa��h��c�+\�<�\֐e�O�eİ\>��ij�][,?R/��?�ZF��������,FCr��?c,%��g�:��w��\)�>4�x/��e o��W��}���3�	;	�h
�����)���{����-�� ���Iw;M��.)�l�d+�g��^H7�_�u�a��O!e�+#��.���
�u���{Ӽ��P�_H(�Asյm�R�+٩G��m� �`N���PK�O��i2TYd��v��K�ĹȐ=�u`1kC%�,pRe�t��M��}ɨ$��h���޶��۽z���d1p��7!�[�'u�4���rN�n���$�,��u�i�}���������J����!d��P�oM�E�k<�i@b�lأ|!FR=#d��m�7���A�~F�q��s���(?�����c�h�*_@�&�:
�^�Vo�.��]��'�4h8��(�q�U<�QMB�*k�[�;�uDB�R/�hhx��v�YϘqy>~��Kû�=좓Ɂ���r�g3���D�p�MDȥ�.k�ԩ��ew�7~'(��Y�t�X�N�4E<K��<_��� �D��+�^+��_��]�"b�f�[���Ŝ��lԩ�n��|ɍG�}W��Hò�hL�v���F|��JT��Y\�.t}��"���������'s��Zc6i,
<�W�=�Y�p����M֠́#.#���}[,9������>/���W�3��@L����
��Q[18����>w#�HoΨ&�q!A���l��3��T�B���?��u���^9l��>E�O�+K�����>'e3�ݗe�>��e��b��������aN�}5�h����;<�ĲPU�F�o iLS�Qy&���K���I{?i�Z��;RCp'�B���vZ�h����j1m�lf�h����a����0�|)w���j$�=��)Į�w�e�_�&�� �T�C"A�T��b�Z����:5�}�N�S�oS��	�ҡbC��f�d���\��]���~Ո�n6T�/}����A�_rI�v���
rU ��@Ҟ����Z�ڐ�5�WvY���瞌*��6&��+��,����E�;��Z��X�A�;�+y�7=�C�j��ۿb�	|���I6��O�AjL����-��2�R*�3����tԅ����++�3<pZ��⦭`D~CɘU;o!�l..?�V��[
j����L�iwxcw|��8�xr9����0�LBYֵ&����b̈;ڰ�}f�0��Y��q�G� 8��ef$�.�����2V�����I/Y��Pit�F"������,c2 �O��������:���H��Ǆ݌���ÃTEI��?&,�+L��I�`'B���J=q��e������ÄC�;"�u\�n���z�L9��� �$}\"���폿�z��G�)QSb�$������p��q����^2�j��]j-�lJFG�r{#8�N��o�*�8�f��H<�1�ێ��ܙ��������D!��JeƁ~0o��ZJ3H�<ŧH�F��F��� -
����U;c2�7H�Jrﰥ>F3�L?�D�����C"Mz�0�Z�
�&P�  6l��.�qN��T���]���Ӵ�9C�\���g�>��8�A��W�ߍ�nճ(�L��L�.\#+�24(�=C]� �q��!��y��'���U�'j__�vϱo�66N�W_$8�u�z�!ɟ�݂L�o�h4�C����8Q��5��S9y\7o������z�Y�{��"��c�ﺛ��0d�q�rWQ��	OD�Yu��{��.V+֣��s��W�����8#���+/��t)|��N{b=@W�Q�����X����/;��i�f6L��%�Zq^� �I/�l
�%bkΔ�lH]�_CiY���)Pi��E��Δ<�[�:�`l���4>)95�lh�(�+f�W�Vr�.c�����d��<��Ȯ*��,Xw�\�L��<�Wt�8A$��Ձ:�߈,S�&Y=��e�V�+�}��o��6�º�	���T�Y ?��wp�͚mh�~%�l�O5h�T�^~���`
�^�ķE��J�νu<�&�&�b�SWn�����SF�o����1�W*z&��7W�~�;J �'Sh����w�L]��n�@�Q3�;�"r����<��_�Ks8������M:���^K���;�|\x�9��m���ڌv�����&�p���8c�Γ�K�����š]��S�����;�uX�n��W�A��#��
z�U.�䄾^���4e�d�&4���:ʱ���� l��#)�tV��l���2�~�����kN��5:�k����Js��.e��^.�_�2��9wW���Ek����t>���܈��~JQ�:B�;PAD�st��JnP�Ũ_��FPzN�&��S��F0� 94���SW��ݠ1��������绵σ�&i c
��M�� �.�j���u3�1H�Tc�"�R��A�cU�}:z���d���P�
����PN�kY��S�����gijo���H֯�19k��I��C�K]�GҶ'AX�ᇭʶ6D���`Cy�+���@�4��6�I�"@�w���?L��2�i�W%΂�e��(��{:FX#�Y��J���z5Ծ�39L�E�˩�х�#;������/+��YL�/�JJY���5��=	$�I�t�Ϫ�[ږ�X��k�T�#kA���s<�1}��<:������r�mӷ�ih0S�K.\aѺ�GE�b-Q��$t\R���G�ȱM��6�U����4<v{Pd��BM�	�����|*���4J�W�	A�ҵȬ$VA��X�Lo��ۙ�%�Re�	�{�����l�R����q~Ъ#ݯ�֟��Cq
�~��l��t��M�\(.^_d�e*�^��ٕ[O
��
�aA���2��13�eO\���(� �#�����=F@���n��q_�5�{���t�P:'M^Z��Ͻ�(/5��:qS���8�˳L~T���-��;d�>����1Uu�ɹ��	��5� �M�|���E��q�m�4+׽c��1�8�G���?��zx�6k���4,OQ�!\;��ll���Q��-���tԎ���1�heG�5b�#��A�<��&�_6O+8�Gg�3�_5[��`���X}��ڜ{�:?�P����m�pɬ�p��{ټF��8ƻA/�.Y*O3@�꜍#�(�_�KD����7�w��M�V�bf�A_�,����yk�xcT��.�}�~�)vŻ� ������� ��h�u���@� �ι��@����,Y_w�&B��(@�m�<6<k8i�SE�{�C�'C�'�;�my����r�26(�
��<p�k��L�U�h�D4�9��S��_Դ<�u�E���-\��T���ob(�O�v����C8W
}��>KW��"#���D��B\��-�X��k����{9`��J_o�k+nf�u�Q�D�?J
�'��m��gM,�aHҫ}��PR(V;��B��#`�y>J}��&���M&ph7K�Z~6�����ݮ>�2�p�뗊��Q�����Ӎ<&A����ӵ}���l΄)a�A�����?�W�]C��*�^���8���!�`C�y�&?XD���GI-��V�ȣ����>j�m�@�`h�7�?�.x�p���ޗ���$���=�CZ�[�Ԫ�]fd݌e��F�߅j�
<��1�#��C��]@y�