��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv t1������O٘?�)/;���;�+	��۳�c.�Tw�R�.���js�w W_�k����|���vY>j<R��ZL�����X�T��ã2�ސ��]4x�{
r:����_z��F��Qq��uZb�sG�rv�Q2����=�Ђ��&�=�J��0����'r��@r� �Ӥ�ujM2ER��� ���C8ʠD�'v�3c�c��^��\J�1���_Q-����`J]7�Ƞ�y^�T�T�}��2�Y�f����ǰ�G!��,Nn�	'j�$�� �(ɤĩ01�l��\�wU�v�q�YHF��l�F�$T��'�����\�`h��e�>\�iwzG�Y��/[m��'zG↤w ��I�w���kyfkg3��y�x��T�j��ke�V��~y�e�G�\�ֺ�RdP��?Q��]��m�Ž�Mc���6�����X�Z�^�
Z�
x8����_)�h_X4 �g��t&���4���tc��fpfG�E�]�C����ͼ������*���&|��Єe�F�S
Z�1��E~Vs�x?
�u�t�rg�!�^2ײi���B�a�:�F���6|T7�y!��y�҃Z�t�=������%�ߺ5^XHp�?z2� HƋܵ
�q[�I��_R#��pږ}�`�sW�H�=l��7�h�!��%��"����*$�nT���Y7��Q�ԩ_��>�_P{�w�$~�m�gM��l��oww�,�Q�?Z��VJ�]6��i�z�ӗ]��T���Ov��P��rr�5�_���$E�Tr~y�S�=v����`�rߒ�^����0QfK����8 ��c����Е���Y
�g��i�ߎ0-���I��R�"���X��/3�!��c%����[���<�C �W�_����/%f_�T�����nd���j��1���{�s�:�,���k*T�NY�v��v�CBQ4�2��ʲo��TI�Az�[R?����{����0�%��a�5�b��.�l�ʸ�j�S�~��c-�T^���Y��D蝢�)���jJO+��؎Rr�&���\(+�l�Z���67��S0ߵ��@���w���2�02���K�p��8��.<&3ZBn.���L�!����B���|���Ѽ��vM�f�Tl^��O��Dj��UDb�9����ߢ�:�ǯaP�l}'컉R��?c�ESZ�w�p�J���p�d8��]4�iV=�J�p<�e�ǙeX�;z}��2� ҕ�Ig�AV�N�t�!.\�+���J |��Q�_ �4��J�`\�I��A�j���I�4(j��ז��LԱ]�7؋�!n�M�"6���:2��8�n���\�*%�o���:����ax�|7Έ���k&o*��}cȾ��%�g:��s���Oo^�m{u���Ԣ�e,grV/Be�0��%����h�W������y0������	i�4�'�}
L���Tx>]��$+Q��m��.Z���6jra{���}�_*�b��cU�Z`ig`�r<!~�"6pN$�lEe���1u�	S!w�87d'��^~��9��a���*. ��Ԑ+�y��,�H�FfCt.aOzɡ�^����r�	&C�׉d���:��Qm���ڑh��>��Mj���*�vDjN�������*1��w頑�yN�Z��v7R���5.R��.XZa���k?��Ke������t���yl���t�[�]�U��A�]�%ވ!_G_�[����-)ߎ@|�{Y~Ƴ�OP��9H,��m��B�'@є�K;-��8�|��#
X�#7BU���c��1��� R�(*_�
R����_�������n��G���B	����o�����貞h�mEۖ�z�����r�x�TPt r��e�����s#+��j6=����	?��6b�8�؉s�
�����N�P��	�TZ{"���%�a*�2b�T&�$�@y�Ԯm+La�eҺH뮉�3/C�����P��F�iuw��S`^ϒ���6Z�f]`q��l����b;�y(���/��B�#�(��$�l����C,�L��x+��%��"��pȈJ��8AD�U_��.kк���#���Nj{¿�F�޶rJ��.�"�K�ڥ���k�����I�����k�SY۷�(�҆���Up�pz���C��L� ��:�%HF'��GɄ��{��!z�	w�h���F�Y���"�F�p����]L�7/���c4j��#D���� L�wh��u�,9B�Ԓ���ÒA��֫����Z�ƃ[*�
�@j8C?R��~�y�E�ӅBlmr]��I4�K�������d�knFv�)�%�-!�֒�_��cµ/�NN�C�0�k�"RL�'3�6i���h!�&�c��',��5	.d𵅹7=��&hor��c�����BZ�
��Gx�s�r���:�����kC����i�8�Y:h>2�\��'E��s�ǡ���S�I��};�`9@�>	D�$�=7��$���J�:���P7�[��3�Z��P��q��M��2D�ؚD�N�2�a�������kt
1"������ۻ�h�����q�������I+��>	i�Z�:�����'�bya�\o��n#��(<&�l ��X02���IT,�`�b�1��NZ�&:�E������E��i���㠫�1��t�WǄܛ���|��}��^�v�"T����pJ#k0��<�Ll����դ71�4F����4�/xw�b�b�(�>�k	vf����B�g�nsם�t�zP�Y/o2Y�z�B(�upҖ�.�X���ܿ�a��T`��P�Sg��9ZO�]e��"��=���:���~Sэ��я�s�^���(��Ӓǵ*�	B{�Q�mE�cw���;Px?Y�\�!p���6�njuJ�.��XE��v��ˑ��n����a&8��R�H�#���y��4+k�T�9�̯<�^⊚z�Y2�Gy��#�T9�ۥ	��U;�����N�e�&�\2��>x��BO��(K	�}~EYn~׽_�i�+W}Ҽ���Ӧڏ�[�R���RY#�B.�[���D0mk<�+�@c2�YM("��ǳ��j3c�ǑM�6k.|+���%)�v��꘎�t;v2E��$�R��\�Ҋ��RN�y�D0F�GvRzVqP�����v}9B���a�<ۀC��>:Nfݘ,�g����^����z�4\d2�-�Q�.�0-E��]���; c� ���R�]�_��\p��	ns>[@��S��h��
���s�+�Y�l�n�K��;s��2Ę�N�4�a���Ӱ9�C���?���Iv�������#6	U'�}F�2�ݻV�B%��-/;�|�f5N��
��(6j���-��ޢ(�.F�<o񓆋��07��L�-pϏ,Q�U��{�R(N��Mj�I �]u��y:�T��TiF�
�=�>z @�'n9���t�'�H�ۥo�����(� %�.a�sNT��3�"�>?�ޫ�q�����[��<���ɐԤ�-�R'�꒴lQIz�/��/�jȸo����LD���"�Һ��.(2]��Y����tU�VZ�쩯�ZzF�[�b��6�i��P�MަIO@�\O	��Kv����<��\nL?Eq�������v7uipi?$^�t*<�{�{��ބ��@���˶����%m��͸f���$��D`'
���@LT�:�$*w;ב�o����&51E�t4�5Su ȁ-���8�,����|Ng4C�]�Y?�I�tj��PYap0�h��W�z�oC�Np�3fD)�|�����f�[�g�i�8Y�!�X�4���Y}�A�*�}�$��a�^�w�{'�n�?�2Z$e,�[ڀ���>�7���#�wJ�z���a�\I��f���f�ل��СN0�D��$�<z�7������h��y�_��=��T�L��A�3�>'A�C��w'P$��*K�`!�L]��"@Ȯ�?��� �M�����z�d���4Ŷ�丷�a�!�T��|0}k�ƅ5X���2�paP�z�}��xjy��J<��ogV��D�tOݴf�ם���d�B��pZ���q��Zb�����:i5��5e�Ox��N�S�A����~]�jR#��!�{$h,��K�sZ4A�jM�,`p����]�,Q[ A7.�z��?	���5�fKǃ<�YFI�V��M�#��ٙ`�Q~$��U�
�cf��x���q���ǧ��_	D��v��\�zY@e�V]� �[��f����\�mA��!�X�)�!� {I�p�D�a�+�T\����*�d�q8�7�zW��c�N��
�jQ����H�xKO�J���P>*�����D�\6�VF8�.*�W��6���+}S��߆�Yѯ�X�u�R��P7d�W�ķ�P�U��X��Z�)��Py��_Zn�PQ�Wڊ�gsm�v��?�v�v��'�d���%*ְ�_�xv����8�+F3�F�:����9���sYd�Z���1�]�7�PË��f6�fk��p@w�^R��A�R�� U�x��W�;���5�f�ﬕA��?fn�ȬP՝���+�����sT�vJ��<���WQ��\���Q�9Ӗ��z�r+H;���',g@��,i���Aߧ�W���1Q5��uO��F��sb�A�و:�q�{����I`�oŧ�ՙ�vxe>�܆2� UC�I�"	�m�ծ�P�l��h�c�F��N���� I��\#��M7!h�SҜ�:��.�˚��CY���� �v�� c�\�a�ͷ��yI��w�zԣ��?%���L�����Q�Q�ޖ��{T�-zZKܑ5�5���\趪_��n����.h��&�.�`��fN��j�:_F�~�̶s֋[.�����1b���@o�V�!��mI����?W�l�­� ����z!�j�v{����m͇1q���}~/�3r�?��>@�ߩZ ��Y��W��!��,T�jK͒�z/3�Y����}:���CB�(�5���Q��D�+s7Rވua�fx��,.��n�����SR��k�-�	|�͉��D2��Z���#0J�%�� R��?�#4��U�L�Y|B�_4��?�kK��^(����f�uQ���4��\ ���}ڿ�m��B�c/���b1�8式����U� �.ʌ�`�n�,�F�&�9�{�?V�%6���
�u��)���?�S��p!��u�l���͑�7XJQ�:EAp�=jo(�_�03�l�����oT�q�cT�6%�2�1nUi:j�kV/ެrc�0�x��k���( �0G�n�?�2d�Z��Nx��P�Z��?P9�z����Ib���&ɫAq梻�r�S���
a�Q@~� m�]%���Ws�6QB��8�%�zKD����s��5(��ފ�kӂn|�d[=����P_�ݗЬ�v���>DI�e�H%�Y6��t�E��z�%�zO&72� l},�+����ъ�?,�vA�wQU��5y���Dn�tK
�#��Iqqz{��;�U�p�`ՖQ����-vZ�ks�#$5PK��۠�u#��}eǋ�tN�~�/S�� ��r���3Z�V=q5c%�p��m�;��%Zf���wR��.s=B���J֭Ȩ;6��)*-"����m�SS��Sѕ|���Z��M��4���$^+��j�ݷ�@n`A�Z��}��o('Ϋ	��'zV�IMu 9����>���t��F`��� �l]�T3�X���R�b�>i�1o�#�:��Tu�2MWz����z&~�u��:A^��z	�*VZ,qp�ޱ+�Z��qة�RZ/�4j>�|"���U������-!���r��`��x3{�}e	6����P���Ef�SQ�v���j.��c�5�0�;F�!!~��ic L���>r	v�Q�[o��u�dc�j��0d�G:��lXl�	SH'�H�*SlE^$�2��� \�(���u���M?�hl5�[��P��J�<iݵ��B@�ݞ=��.dKFK0��ԣs����{����br�f{F�@�Fr�d����+�})��4���{[�p	�(���¥���6Q\x1�Еt����Z�&�e@��W�����P����	�Y���[�O�eJ�\ߗ<�)�Oו��
�"�-���v�����O*��D�h"X �l�H���'���<a�7�i<k��� N��̊�=I���}
���8��zFد���}�>������JU��
��^XW7�Yf����gM��"	W����B�1��ĳ��§`kK4\F�e�m��®�aN��.�p��J�$�[�cp��	W���L������^xK�ۈ��>��HL���RSr(@NL��[&um�a?����㓳�Ċڐ��轃�V#$�Y�5���=���5\W*��F?��kО���RƯ�^�D�M1�gW�ֻ����u�.�+S�G�eVs��6~?��~�sV�k}�������HnuS����U�ݪ��$�IN��B�J*o^��P�\2�ˍ�K6wUZ9$�|�Y�<;"^�v��_[]_�Iw/B<���:8�X��5������#s��(��t�ls�luU�K#��.?@�E3���>�2�:!��ap*F�vq�8�족���Z��iy9p�^�������r�rݐٺ�;�|���'�����HѲ!d�	2��w:M��*A"C�${̜a�c���ޕ�QC[��������/��6��H/0���5u���2��4�&��M�}�S��h��8��G@^g���j+w����)�����[�V���^�%6���v�hПL��7yc���9(I�P��)�[�Q���_��Ͽ)#�<����#g��M���@���m\lL�|�&T�'|�T	�>�o�� ��L
Қuo��,� �G�Yr�6�n����e�3�U�~��	�Ґ��A~���|��$��3���Z��YP������M���EIbH/���z�]`����/�O4��o�t�̂(Y��9�ˀ���m���V5����fH���s�.�>IȂ�J`�|E�*��h��G\}�l��!l��5�}�f��Dj?%�օ�,E��׽i�tA�,��T<�叝-<������������WxR��W#f�^�����U�Ѳ�P		d�Nﻕӑ�+F�W��&A�{�.t[��҄����Wb�`p�!1�c%s�:}��(Cq�@jC/V� $H��L��'u�'� W�2_H!=���D�r�
�9��	�$<�"w%�6��W��	*L<蹴�Oe�F���@��#�} y�-8R�Ц {��J�k���R����A��t��5M[��'_��4�--�^��!��6���yA��վ�#�L�1��g6ź�l�K���D��cY��TT����%o���n�_&��j)OJR�2֪f^8]o!�G�#K2]�(�؞��8�L����'Z�"��-[�P7L���c{ns�H7�`~>�UyNV1E*İX�D%��j}JaKnY��J�Nx�bgP�S�T��!
�>����g/h��\����5a|՛'�5B%�=�%|�\�q2��=���\��0��<iNt��і'�@=�8���Q���\���;�˪�8Zj����S�JUu6Ė9�?�Ҡ�������N{M;8��-	�%e��ynލq��X�
PF�:)+o�(7m[�E�>1���mw�c(�_����{���NZ���-�'��1���3���J{�>�)�Ж�}�t$�!T5w�x=¾�:�yI��ɑ�$���ޖ�e�O����T�a�*#�����,���iZ͍�8a�08����m��m%��C�t��2Ւ�A7��_U��|t�<�j��,���#�آ���h�g��x_UEN<}e�'�B���v���Xl���#��#WC�'KT)~��Y�\;�r�{��tk=�Q��;y�{��]�q���#�-X�4,-��� �S+�N���i����P��b!AAk�ִ׿�`���֕?y��v̵w�aY5e��Z�$e�X�xg?Ð���8AB�>75�����;�Q���Lx��y|��dq����F�|�*h5�v�IK=��<}�ކ��3�+���%��+e�꿺6@u�#���w g&����x0B�y��<�׍�w
;G�)�&�ֲu_�"5�J���@B��F�e�X����jZt�}�9��Q͘�WB:�����$���F�nwa��"$r�uk�Hv!��Rd��o�{�< ��������	��jFҧ�JZ�La �2t�lp�A����NȒ� ��J.�-"���s<���܈H�Y�����o��ֆ���S(+�bV����{��8Y��Lt��<J�?s?o�4�R5t�S\�;;h��`{6]~-e�Tأʲ��е�u�KL�sD8N��<2$���k�R9�J�\�A�4�Y)�%`�Bb}R�.�V^�r�k��E���R��Kp�gsN��<����u�H�R�3v���}_g�����*�k���5�?��V�1�z�!������T�i�b���;��te��C��:�:�EPt��@s:c�D:�Yܞj�FNw�\G %4��?;	�'	6�X�@Ч��E��g �;���1��}���]⧁�����:[�Q90g��V�9IE�O�{F󍹘���˾*�Ӥ^��vp��P=;j�ߛ	��/�k5���LC����sO����1vG����X����s࣬��us���)Ս�h��X�t�j�*3�v���=�� G"*`=��`���/e���ֶ�n9'`�u-�	^�@%8�Oɀ��O�7��1���Ykqz��)�ѣ��9�,"b�<*~�LE�]����W��0����3��af{�Ѳ`��|�4��Wq���
cRj�E�(����m\Q;�^�c]��RSS��R9�y��aC ���@��C�p$�'����l@�-�����^i�/h�c*��5�-#�J�nB's��XZA?�*P��u+�(���gW��c�ѭCcX`x�9���6.��?�)e�&�� ��ߗݭ�{�L�U8 �P���4�o��fuڊ`�<m;H�k����i����g�f��O�R�L�WEٸXWv&crg8�ht�z�#�x�ҷ�Q�hT��?������F�������ƮE�K�E�.�cڣ�����4���9H\y!Q�2t���H������ȥ�sC�C��</~�z��Sf�A���X�_�ܿ��v����d�6�J��|��e�˜}*�%��B�n�?QX��M�sf�gQϖ�J���XQ�ͺ���b�>|c���~��&U��`c9�츮\�1�4�ko����J�|Y3i	s��MF����&�ش ��B�T7B�0�2¤�k)S���P68a�b�╽�i'êǢ���-[	����8G:j��r2򵡷��:|�����-{�9��q�M��{�Z���ձ�iK��4�����v��6��CIn5��e����3ٵA?y0(�q �'�ݍ�Y�#�����fS���G����8�+Qi�e9�vOܑ+�W���j��i����� y���"�̖��ph	)_6���T@?趛�>w�|�ICE�>��w6�=��}�EA�K����̄�\A8fل��^�L�0�v0������'ᴼ��0�/�L��ؗ�s��� �4W�V�rU�iH�
by��f�����.��Nr�!��P�k�H�2q߬��s��g5D��tX�r�'Lp,@ZB��!n���`^�+J5Vb�^�
~ې�'�������כ��d�`��n����di��W�&��cC"�'�8.����qÅ Q8#��l^?�c��U�����%؊X�^�^[�j�E���E��c�|�B}1%ē�}��R"%:6�� M��7�������P0e\F���;,ү�c>	>��|w*M�Ȯ	��m��������O��,e��h﷨溪`Eׁ�W�����D[f�S�)�3��:x��(]�/��&�7G�kD��a_걑A!G����NC�����|
�1C:�L�CGR�Ž�'��!��0����7.
0�
:$�h�VQ
�I<�x�i�",�{�L�uD�/m!���1R]��Nex9��bMLK��Ɵ���_���;Ё	� �a�:��_�2̖�
��I����Ě�+�������9�����v[��p]
�����u���)�iIf��f�)P�_ �Bd4K'�<����]�t7����ϭ4�M�	�JqJ�Ǭ��Y#���.�Ie�P�M���>J,|�5N%@�3������ˮ<N�Q���d �_"�?�l�s��мg�G��(O��#�R������e��/�M�~t%�UU~�JuZ)4ji�����$��Aߕo4b�[I/�F����đ����w�'?ǈG�&�
A�!q���#z%�C�ǥ�%j;*2���~�Oֵ������cD�i��cŇ�ԟ�QC�$J�@�3>���3sT�@�x��7����P�L,[qH��?��ӗȽ���#�������{)�X�&���m��:! ���=�
.,Au������m�<k!�F�'KB:e	��2U�4[�仩��/B���;��ؖTS��3;��)��i*��\��Lr��а���ّ�_(��ۇ�Z;��S�J��Z`�Q%�;
�#�FJ��e���g���ܩLs\�2��_�fs�?�'�k1е�S��e~]�&�9���T��y�:��g/�B+ ��n�����*�l���Cg��O|G^čE�_6'�:���x��N-�[D��������|�HDlV�q��=�$�� �h������e�5;k[���!�c�ޥ�!���k��|L��lH��kŜfO��-	h_�Q�gAȡ�����!���Pnԫ	)�d: ��4@���m��o��N[���l#���9�@ŸD�d�鮫aGɇ7AX?@Oa��Ƨ���f��E�5�������av��
�Wy�&K�b�L�Δ��v�<���b���击� ��s��}
�"���r\��R�,F�<��tb�:���q�$��1ڶ�d/���bδWi�*Q{x�`�Rt{���1��ߓ͖`&5%߈�=?�k�N�����e7�L�d����5P�5筡���lh���8���v���������>�R��&�XB�B�i��Eb\��J�Y�Y����i�z���ˑ��5m:�}������,�(��ζ�=�P�T��!N8��'�����0̤��-9z�hE�=v���|9��IDK�1�0�Ղ}���6�����K��O���|tX���e{2��^w[�5�}�L����ݲ�H`'[�HʰH)N4ѓM ��k_�82�Bu�����o�ױ�]�eq�Gr��yr_K�O�j\�#J��]�§m�����:L�H[h��<��'=8Op&P8<�bϰ�)�����R�*��c�[��o-C,#�|�=�_*�$�R��R75���`خ�q� ���"��bӟH�sj ����F3�����H�(iR!�*KJ[F�&�׽{����1=H�q����T�p�"H`ea�ETw�F樉L���u���om0{����S�OK�s`'*kcz-ԧ�ŧ��:��� ᘛ��$_�u7�#��=��^XbW������q?A���"�R �]h�y�nŢ)	y��&�QM�@���F�_KC�=�D�}�/Av�'���-ͧ�O�����N��s]�~3�e��⯞r�49�?xRn�x<}������S�ʘL�H��#|k��A��}|��Dy`!���CfR�|/j� ����ѱgm$��>a+ϮG��p7��9"�ُ���X����O$��{S��P~MoJ�ҷ��ƌ�W� @I?Gw�f�:y�9�֗�\� 裲��U�ø�]׏��a��'}�tK� d]��J5+��C����9KhZ�a���7���jfa�7O������)��Jb��	Ci�����ıj�p߻6J(�HN="���*t�Ck���.��(݃� +�Wz�$ᆷq�d�þ�:���T��𧙛�7x�{�C�Z��}X�1���
3k;@�v�G+)]&P-pu,���]�Ԭ�.,р9䰂UV�%��8~�C���᲼�7��J�tO8����1�3�vt�F�D����moͰ,���@�Iߌ��;����~��N��K��6F��l����+��"��'�L�z�Xх'��e�#x�	��'���Z7:��~�A\Nv�<���M^���F��w��Ǩ��k����h5� �hT5�o#���L�#dجޝ���OlƑWO	7��;��n@"��,���#��R� r�viRP5n���-��B����B{M"l�L�(޲:?ekm?.؊���=U:}�'$Z����)�#�ڟ�5w��h�pH�/w��"Й�}��D`X�Ň�Gj"~^Z�eL���v���%�%U9i��١�� @����{L���	�t�u�ɵ�&
:�𯳩AYhE�Z��4G��� #�Y{�7L�r٨r��l�{`�e�m<��ϋ��P�zC���ۇ�����&#�w>EH���T$F٠]?�;H��mc�M$��rGVG���ޭ4��I�\���?���˂����o?�Ǯ�HE��F�8���s!,qJ����ݻ�ua�3BT��H'vK�qE��7i���M�3�Lvn��NF��|�W�x���:�!�GH����-�0s��6iԬί������	���La9�J������'�O��ف��j`8��s4�{/ �B�W0��.�e�&����_��S��g����@I���bmXqj ����q	ej��6��I�!+�\E#Gn�h�O��9_��>�{�2p�MWߣE�v�O,:b���#ܫb9��,kc���5̝��)u��T5rٚ�h,M�-'�|�f�sqfz�V�iJ�������=��_�~Q�v�Ȩ�c�5b�g�_&/��8���wJk���͸����%�iq����~�ƚ���@<ߚG�u
;�0l4ZG�e��Qs#:���Sֆκ�j���m�w-=���s�|�������GcB�t=Ҏ�U�7�ӥm��4�K[W���z޲$�л�q�º�b�7�-�"���WR��Z���}��b�N�Y��}	 !/�>j/���N��щ0�̪*�FxIȷJ`�x/���<ٟ�q��z_Q�S�8�I$��1�^�E�4\��r3T�/!LD"�t��.G�ň���܁�n�q�MxV��T����]�����u� �A��3t:�CS�S����CB	��
��It��70�u�m'zDY���8�j��&}!�a��/.?[��rR/�۳�\F�P�H=����4)�Mq�Y�(w��<O�J�CnHvk.�>�@��J���MXg;��^m�:֜�ǉ��PY(DX�R���kQ/���Q���	�7�=�v+#��&���$��K)3Lw�c�r����� �+c�XR���D����1�� �dB{����x��Y�yG�՛��N[T�lg4g&(+�ǐ�4�cŌf~�w�x	�R��	+0b�>�������^��R\=��:4�}os��s��o�p4M������rn`�&��k�!!cę�@Da�����&�{�'J,I�2��
3���p�R.��~/c�Ӌ1L/⑔i��Б����>gf�8��<��0uQ��F��*ـ���J�k��� �gnX�[b��l�Zn�+�td���R�N�7yj7�Ž�vr�D��@�SX�j���R� j�6f�@�#� ��e�N��>�D��8�	��J8�F_]�^�R�p_G��N�[xT����$k��X$�!�yE}g�m��4*U ���%,ܪ�Go2u��n Jg/u4�O�Ah�f�Æ�/�k�ap�(@�� e��^�B����;�ܐ�Uu�D�lClp\ꫭ%77fES=�J���g�!��2�Au�!R�C�a�­���!5�g����(��z�{��7� %����?���,L�2���`�F?�hb�=�����&����4t#��}�Ვ�+���O�tƃ��"�A0�9ܡV-3����P�@���1zU��1k�`�^4��T>rJjx������Go�t��zcIj�s�U�DH
��5Зp8U�F���1'\�1����1������pl��܌���<���EJ���բx�2�Ps\��)�~PƢ��F��K}�%o����*a"ѷ"Ur{t���_�/�@ ��C��N?l�g���%~e?A�w�� ��Tj�!Z��=��FX���`�`a��9�ˍ�aI�v�7dOX���]�z5ȂzQ�*��KEsSm�^�.�C����8�ɊcU�F��]>��H��k���ٕY1��,��0^�NIag�q
hLK�ғ�KOVd�M�`@�km�@S��-E��a�WQ�-��j������s>߯G*(�i�=��2�dW�U��� �~ʢ��ƾ���JV��ݢycK�(��`�q��S���vy=zNL'-�?�[���I=�]m)Q*,����#�EL���#2�J���g��`�JM"�,d��W$'��j�N�ǆ�㣟�|J*���p��I�A�=�}��g'>�z��C�/&�KB$R� %��9 
(#�#���n�R�����%�j���Tv^�Ȼَ�
Z��m���=��n���x��a@���g�ODi̲���a�P�b2$Xe�l��pfA�DrUr��a�'�/�{�*��T��"n�MK	���3ĵU�x4u!e��9��#�c��J\S&�Cks�us1�A���!S�K(��ҬYo�N6�Sq�gm������&7�M%6�6�� <�x�g�#�(#vȞ��ꪒ���s�j�헟}���7/�Q׌�OD��
�'/x�[�$ ���G�_�_it���]=��Kd�e��]�'��_wL�w�d�i�]����m��@md�`�@n�[F�h����zb��6�G�ñ4͓���W� �9�5��L1�Y> !��bw�l�P��^Xq��������n���I� L#�hD^�
�Ac�B,D���TY��S%9ӡbK�os]a�IЁZ3g6ʰ�
�lF�5�(���*�8��|@��U5,�46Ʃ$��]��+a�<��ܷ�U�z��6^�h��Ĵ�A%{�.��
�25轈u��Dv���176q�H<Brة5���i�?�g#�Q�~Q�/6P�/�A��Fns��g#��+BP%���#�5�a�]�u����|j����͋%�J$���Ɩ��Ѫ5T`Gڍ�`'�*�X�S���\v�5���}���zg�`��e�}�*��'��H�� f^0I�����j7t�`M0�8g����> ���l��8|&Pt4!�"�+�	x�?��E�jq�S����������)cЭ�*5"bVB������w�k���x�NáZ�� 	6��|���r���ذPl�u���y@YT�U��bg��w0����2v�/d����I<0���~4��ذ5�߰t���LLV:�����;ra���Q!k�x�DS7�9KLA�������� �8T�Z}˴��i�ʳ�?Y�2��^U�a�8�ʣ?[���,�+NZ1�;r����cr�ls��KIsߙZMn( &��Y��)"�&�M�(<`M�
ҧ��^��1���QH�	[/8�\�K �ާ]�	>�ZQNq��e�Ӑ6 �_Zq�/�7�c���Q?|���[�4�aY��P�V�IꞶ��g�4�3>VBvv4�ZIB#/��C�$ز�=�Ʉ6͸��l4&�HsL��w�˼�M�z��Aa *L�'��3�pwu�v����B�(iP[�p�2[_J�}T��rS^Fo�9��u�0++�J�U5��?����2"=(f���~5�D�hIj�W1��?�8z#����b�:1k�pZ����6Sb����;�2�b��'~�_9�ZfCvVWG���xҩ�0K�mb�X���Y��7��G~8����b�����9d��ͽd��"[[�M�p|0��,��d�}�Eao���k1w`����РV!C���w��4�󋼹'�E4�B�}���Y{��u���id���P�%:5+�Hp)����!:B	r�Dca%B���21U�\�%��ϯ=bP���U�^�,��w����a�����M����U��Jy�)��A�^O h�L��y]oFO��Sux�c\W8r�8Bǣ>�FqZ�Ly�(\��t�Ĥ�Om�Y��]��W*����7CY����;���E0v��W-$��KR/�dG���!k0�5NS�H�nr��GH��ۘ�������y��|Up)f0!)�=�DB#]S�Cبt1D�#�y�	����Ŵ�%�y���s���m�ˣ�F�G����:Z���N��!�`�
h4H݋��A���pݵ�-�CtpQ���UF-�eBPԪ{���b_s�8�2���?����J��b8�����mb�줤yݪ��U� }ޘÈCÈ;Q�1���ԷX�\�_�M��I֘�������m㚘����M��q�+�\��BG`D$�_�FG��Cc��[�O(89��h-DT���d�"�:,Ɔ�����L�Et� A��b륂*ʊa0r������67/IZ�!�����JX����Q�Q�����o8���O��Z�[&��e�%$?Nc��I�Q�F=���ת�	�� �|$���������:0�R�^<�U4cA��w�����q��4��ͫ=�2i[􁝕�_���d�/j�M��Uslܻ�.���r�G)�x�DY���3Gl�; �8 j{�bb5��0��6#��E\�pN���bX[.����S�}��̑�w�J��z��2��tE�o��;
�k��z����ޮAixC⚰�@S!hu����s���m�`�d�)/O
V���� !qv>vn���%ΌF}���qE�.����.5߂�f��R����+�-�T?O;Ru�L,��܀�%F�d�O���"�)d�ZEa
���Z����J����b����!���U�nb���y�y(!%rmsF�:�m�O��6��e��Z49.	�{q��:M<����):f����XB�뙃	f���C@��|ܙӏuo׊-����[&��V�}�Vk���
�n� ��6��yyâYߔ2�R����P�J63)�n��$ �|!��p�]l���LaP��h�b�3�Đ�Eњ�HKw�����*���[围?��K�->u�?(��� �W	O�o�I�S8O�}����N�W|����K�e� �����_��a�V|�Y��ܬc���N_~#�y�a���h���,���F_�7+�;��D[,�E����
[��a�3oW�א�_�S��+t�T=FVO�H�;��U�L�1A�Z�9����W3�ŷ@�ߓn�8z�<�����K�p���֑�(҄�I���Z�O%	���p��[j�F��݅6�'#���f^r(A渫�����"�B�TҐ�r[�W�#<r�S���Ƣ��j����*e��0C>l��v��m�_�y^'*��p�ӽ�5x�"0���)1/ﻲcy�_��$Zr��j����	����b���nЧʏ�mG�.��/�Np�?�7����VS:AM�f��������9j �����5����U��H�:�������f�FEh�ңu
�xx���,F����Hڷ��;
.oA�(j�1��JZ)/:����ʄIDֿ�
u�u�{��b��p�6�1Z�L���P���^pIw�Y��� #�q:O��dn��g���X�Z'L`�1������b{�#5e����y���\� ny���C��-~KM
7���_Z�q��<��2���.gj6�l�v;;4�&Ώ9�jcҰno�+�8QXl�<(
�`���\'���lLtA8�b�}؁0îR}I�s���^�K��G��3s��i�0N�B������rb)De��?�%�s��}h�����Z`ǂc�	)YRDmt[H�R��Gm��:�lK���h�� E��!�n�V�")e�iA�.Ǧ�.��V���3Z<�dT����A��m��mx��l�X��> )y���<�Ji�>�vr'ՋwB�9>���?���O�H ��`>��!{�O�&��.R��O4S�q���\P⏉�{G�	���@T�7o�3�N�yy]�~F~��� ��k&軅Y���,ia�d�Mx���K��!�^��7�I��і��e#` � J8w5��,�jq �o��t�����x
����O���u�����gV��1�S�4��!u�8_d��;��2X����h|���s��x�1,�V^6c�����}��♉������|E�7�N] �(Ⱦ��3��⪨6b�e��#t����aί঻M���4�z�!�D�=����{�~�^�/��;���z�K~)"���JTx����r?���F��2n8��jUv}O7:v�!�3+e�L�B}��EA���K�w|�������y���e� =����
����/Ey�\ץ����S0�n�W�n�����ls�ܢ�C��fZ�n� 02�%�%H�S�{���.�$�������6kO>��E�O�]���q����oԅ��NL�6�M<��I��:�hb�'t	��k��M�X�]=Ѝ�����4����&�Lb6%��6T�����2|���y�V�9��:����r$Ž�y���R����{����1YH�^� ��X�e�/Ht(�G�C6w�D�ö�B'��iwpw��̙��%�~�����q�T0�%����1�s���n4=X��4mm�v]N?�<�����x���{~��-���_�aȤve)=�%��#KA�6�l���V���H�1U@jP�+S��'�~�SɁ�	� S�z�N <���("�(�Z0Kn0`^j�*��B����6!�����)����ӖZ5R
>��.��R���$�9v�g*���/��n��Gx���$��Ӛ�>���&]��o5�2}n^K ����@�x�_.d��ښ7)ø���l�ۍ���;J,����NM�V��j$�xts/�D���,q�X��PJ������M'e,ִ;�g�Ţù=Ū|CM��[�&�fDr�N��h�d�D�>����w�h6�����6��V�;��4}��*-�^F�(,�)��'��ar.7��U;G�{�m���>*G9����z\NY�o�of��D_15�Y��C���Fz���͍&Z����=�1g�j������� �*w�d���^��H�)�����}*$�k>O,�a���L,&,�z�b����v�أ�E��� HSFY�o�4���4q)+��7��������)b��Ԯ�o>D��;>p[��'�R�3�n���7e���dl��5J�vA#�$�5:�h5|b5w�m����I���jO};���Y��{h�z(x�;�Dp��@�~���aH����[�?$����T�),ıh��'A�����Q���#�.D��j9����%�+y]ګ;��='�Y�4	�(f���!�aM?)��e�0��ݣ��]�n�1�P�4�ȸ
�C=�<䮃�� �I�K���Y��XSA��){k&Ŝ?vw?
��G��<<������9�G�)��S[9�l�B�mw���3��i�A.i�Oښ��q�VW��=NF�J��RoS�L�q`�<�WP���=j}6����2-�X���-5 D��r�
dTG�����eL�FW6�OD��T��<���;H=M� #��HX��E�"OL�����{Uc{#�:��)2n��/�;��8��f���k��_��vQG��\j�<)%��0M'��_ ZS5��U��?0 ���	�l?kR�y`~ψ����Maj��:1t���7b27���ug"���u+Kg@1<�|�;0��{�Uu��#�m�$
x�曔-j�-�����M��I���<�9�rz�㈺�Pd`���� �(�T��;�=���HN���$5^�+(k�Y�!�FQ8a2�U��'T�:2�{�3U��l��HX�/M;i��[�z�J��<�
k&V� F"��]�S9wh��H��<r� ��B_�{v|�w�e��G&�&�����m2����=zk��8�5o��Z犵;�p����ԟPLUPd�"]ʴD��c!͍�Tٹ'D:x#!fp���$���G1]�T�ώ�{M�F��X�8Z+H�v�w���c�`�o� �iG���̯I�	��0ML��7�v�I�͔��L���kŬq��0SREҿ�kk�r:<ɔ�dӑ�����Ȑ��������Eb:�֣k�ug�Z�K�Ӱ*�[2��Ů�N�"aY1t��{p���*��>;)��8z(	�M�^M
���#P��贇Q��&!�1�������ڜ!�UyD]@V[�Y�JW�#@1����h�m�h�
v�Ş��Yp�SS+�n������G�D�~n$:�7�cW��b��d�qV"�w�����kf�ꧣ ��C��]�r�'���TG�3����9�Ͳ���`� I�,�2�jn�%����)ü}b�X�@�q�=��$([����
x7���'w7DA�dք`T)Vw�c� � BT��<H5�ѶF�SV�e��7�l1�4R�/�a�WzK��+�\j!�9*�}���Dkʫ��|r�VoZxp����9%�J����@�,~@���ycu^���`�q����}Hٛ��e�As��}�5�~��-V��P��%ۖ���_9oUQ0ofU6EU�l<�I`�S)�\sB	��̎<��!�\B|T�ߚ�b�+7m&�o���"��N�?��ml���:�����i�c�rjdH�|����"�ar��5�0 �ø���x6�YAg�=E.�i7<��}��jb�И��\��K	��ĻBVt!�)Æ_[����ˌByYx������|5/6A��u_�ϊ���ٚ-��by[��v�?%�z?rH� d뫑!���-��>�\.BÛ*?D=�S1t_w�l�Hj//-�
��V�@��u���+T��U�h�(>��v��a*�����R�aГ�~�U�G�.)��˶��ѶG���>�����mB������2����T<f"���m���m:J��y������DϺ��2�@8�2���s����E0n@��7���h�\Oź�5
?a�j��/u)	&�~� �NY�; � Ǻ�'W��B�׌�]�vو��_�e�Z,4D��_%NlO�*�Ӊ)�v��n�L�4>i���荺�s��꧖MB�\�ƾ~ �`6m�y���D��Hw��V*צ�����'�Y���D�C��I��i*|Pے�T@�ޔ��gj���%se)�������Gj��4�jxv7sP�i����z�ُ��Ft߅)+}E��} �D��]�cɩ��}����;�x�ISe�jG2��M�eN�74�k}c������[س��S�^��ϙ��b�����:�&3���mRX�Ʈ�T_���KJ�=���	^s�x�[��p��e��ۈ7��W-ø��u�:W�|p�7�j!k�ㄻ&�"��7���d���� ��R�2=�C�;H�TfEgx�w��04���
���D�/�R�{��q�\��-I5�kP�J"��?j�����h����=��(�>��x��G��V���H��]�g0+)��~����겭�.�|_���O�x(�y�����H0���F�z�:,n&��X(�l�=�|���u���Jj��)Nd��ϭ�,}(�S'�s�h��1����<�.ò�J��l3��T�H8�t����ʋ`�I �\�J�j���TM�2�a@��ʢML�i�Z�9?��[��#�pd��9zB�i�0�;<�xB��XF(���0]�)��c�Avo��.�vF�#��#����ff�F����H�{�`7╅��;DVe��ld�r1����D�Fo�f"��� ��[`3�zgA4<�^�e���@*��wk��C��I�v�h7����5�/�=pO�ݓ����f��$�^�R��TI0�,�;������r��X\B�u����&��IO<ϝ�be�W����5�_8��RWJlY#�
~_�eȟ�Yԓn{��#�C�y�-�8�ncN˩m�w7{[��9�r��^�"��N�"�k��w�^���V�pi3���wX�v��	��P�K��E��$X�9*4�d3��e�B[H��9����d��-g�+�.�Ġ72wz��x������2N6�[�ڞ�^��M�"������r���[��A������'Z�)1�� � ̿V���Dtt-aUXZ��d��9=�98|5H��]�6n���D��f�s�p�7�%)繦��F��wyߕ��