��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$���b�����ؑo&!�yiz�@�RF�����ǰL[�K�'e2k����m�5w��)īqQ�<�X�L]���z�浘���,U�u���G��d�K���39������U���s�A����;�j��:S߯&�q�i~:��&�r�(��*�9CP��e��-��|��mZ�?}퀚�������[�:ߙ�(L4$�Ǉ�Y9�ř1,�z �Z.�d��o2�\	f�ssbo�%w_��jڒ�L�r��]�-���F2c�⦍9$N�$��a�M1�pؚ�K!*�+��d$:Y���;��kx/�U@�E8<��w�{&��D�a�.Iba���G:�f��,��vn�@�&�IT<?f�;�@�Bfp��Q���I©��5�ӛ����.;�xO2�%5�7�=�'��R���)?�K�<�g��>�Ƭ
VR/8�S=��Djԏ��@�@�ȧ~�O�$�>Jn��B=у�����84��ʩ�fO��uuA��tl��@�e���f{�	��_i������#�I�rWߙ���xy
t������_���P���teT�Ɍ8e�R*�'���0tR*�;y3���2�<�u����3��IG�ٗÚuK��_%/��A�kh���x�����Q��o���~� (n4v&����fpe#�v	-�,��-�	������JG�͖e�(����	�+*��"�V�ލO����y�)��$PEU�����?�pYD���yQ�x��l0�}ް "��3���'?��I��;��͇�Lm�Xz�W���1�B 4�A�V�b6�ˀC����(��r��>s&�!�lr�/{��kV�����?��-<6; SG�cj�#��(p�z:l�#9.��+uϓ�uT����,����v>���`3=ǩ6��	̝�̿��н���]9�SӴ#�M<zz����S�Ň�i!�r��1ݓ��բ�zG��J�����3��C�� j�-ƻ�b�?v{��=�~>j)���~L��O0��!{0�P|��$=Lÿ�٫�ðϘ;����!`R���)	�cG���}���3�!���;Z	��޶W�N@����CWT�yע�#�wb���݁��n�?M'�;�j���}��ER\��8�i�Ȩ�YM��/뎆U�Z�ҵ�Z�k���~�B\�|�0?�����tF��ݚ����Ǌ��ْ0e��w�0("21��_L���D�瀻�VM2��H��:[+*��n�i\c�{ jT!��^�	�ai�On*eŨI���d�
����}�g��g�m���f~3m# 'O���.�b3��.3T���8��3�s���1�#C�M���|���r�V''��B7?}G�o;�B�n����6���(��Z�ЌN�$B7'9Bk)N���;��.�p���7����=f���Ĉ\0��LĢ��F"�����Nh?���p��
'5���5�߈1�S8�O��)d� �W�b�vu?�����Z�$��"!��uD)"��:7R"�����d��H�aEef���G�E0��>\H�_����/�ܼV �>661�	'-��|ƨ���v� Կ4ANN�oQ*�ޔ�1�u��΃��b>\��E󐉝��`p/$&f��R�R�XSP&�x݇E���4��ͰK*v&�4i�F�~�wh�#�k���l�_Jw������!FŅ��U����Q�D���U��{kB��~�&$f:N�t�P���I�}�>@�����]�G����|f<�]˰��ǉ��k�!)\��C�Fl�/ʳ�95��{)�#�����f핹@(�C�3V
�g��h�J�""�P�h�T܏��Ns.s>���4$��Y��s�f���l����tx��f�*�կ4,l�����6t��%�����c�y%m^�3U򸣙�&�RYEJw�r�]r_k��������*������X�b��1R��(3X����<@��o ���Q��kB^G��DÐ�y�0�����J�][ύ��[�@��Ƿ��?۟P� �h�T�Ve�cf�Y�ow�)��a��E˝��q���V <U���Z9%PRH�����{�fi��aw�5S�l3sa�N-�8G�W����!��=��C׵K��G������wt�'�f�X��Q��p]����8�Y���E�`t�C�*{o���s�G�-���&;�n��5W�~05c�^�_��J]: %�i�����y�I���F�G�9;�ݑ�ݡK�W��;z��h��K��*��}dX=G���8��U?D�E=������qҐ�R�s�����̱:<�o����T�W�ӏgT.^���N�[�n���:IB	# N��a�ASn%!-U�u2��A���"���E0�Ȩ�}%xW`��;ҳ�)Uj�U��j�������$i��g	j���#�s�_��Д\ۏ�*
�-`�;�|yz:\HJу7��TT�(YӶ�����X��\�$�A�_�H������gЏ|R0G�аd��y���ς{\B���r2�>k~ i5�Ư�4�έ�"�o�����P�����cl5����&�Ƅ�˨ *ȡ��ls;�y.œ5�[�G�6?�|�kM�,c��!bv�&.b�ͥ�9�蓏q��tY~�KF�kv��F��DV��24�I��v�c�33�v0ǝ�ˌ�t�7d��0A�����fɌUO"<RH<�@�a22	����5�ɖC��KF6�ay�'�P�_5���˿�Yk�6!	p�@��?��G��(G��ϔr/�S ����m�QOCZ���Is!?"-�m���7M⒏����ǭE�H,�թ���+**8in�"EH�Ӓ��J���1�rT �M��&�,w;�Vg�̖���`�ӭ��3�)R��܂Wf��y�7�)��2�7-J��q�L@��q�}ZB�&��S�$]H��9
~�j:[l��sa�^ޞ���ڝI^�x)�x/�.�e�Iϼ�*w�^�P��=���Օ���vN\�\`�{{d�����PI�خ���Z�e*��O
3]X��`���;�]f�U�?_4�`װP��R�9=Y	U(_���foM@����sJm��M���ډba_�Jm����f:����Y5᪠��p��Ŕv7%@� �K��jT�]�F)�����kY��?9h�����~(/��b8'�8�j�^�X�-[��J�8Z����=<��1�d�\N�/ܡ����a���7���,���v�'h��{{�Wmgj�[aCR�3���tK�j��4�� �p�v6Բ����PӋ@�{���Ӻ�<�!�1���ؽ�՜�L�M�@��np��:ʗ���q����8"�
��W6r��:V,}����R�;o��I�N� X�:U� 9N�#J  F�M+�L��$DZ�]��)�M�*�2�� �|ּY�u��b��C��,���Ǝ�CM�b> ��ںF��v�;6����~����H���[�y�;��s�J6��o��r=���M���䆀%�ZΖY	;A�o����xO<��Ʊ,��2��T��I[*q��Q��t�oR[B�UM!�D�1&d�e٥J
`���F����]��|��x[/�ߩI ��ݠ')�������I��ĸ�<���K;���<�O����5���x���1�z����J�[̛خS�k�m"��t���)��脴�b��i�gf����Ѐ44JA�S�!JWU\�e|�y:Ge����0�H�o�N��~�\�+&��[m�x�,��C�e�4OGE��c�+/�@:�P
D�-s�s�j-ɃC�,���(���;��Vl��K�������<��G3l�b�x� ��0�(n4L7_uq�2Qq� u3#�P;��F8��.�|4'�㗪�;�3��[{���7���y���u:H��uDt-�6+9&[g{+/��%R�	��y�V� ,����4&}���;T���{�r��8f�6���j
W��e[_��7��.�Ep�ާC�j�-%��J��qj��S�j�W�.e],_�p��|�Y,��=�!��i�K����n`<�cl+���x8�l5����&�H<���,=ҏ���D��m�7��_I�m0	@�Ȇ���(r��x�FL��DǷ�RΏ3���݊r�C�种;9J�	�e�sa]E���Z���,S�(����]p�;z˓�"�fg��|I�x���"9d��V2���v�y7b<�^��x�1�W�@o>d�KA��{)ʅT��#7��E��/ȁuޞ.������.?F��A��M�`�JI�����}���Zr�e�/P�!ɲ,��))�\�Q{ ג�����W����K�XI�߀�ƸMFiqg״�qC��}���99Xc�x�������	��D����mz�*�~���tL�xA�f�ƣw?C��:i�n�t_U�?GD힝M��ې|�rR
RZ��� �+=�:BF�z��Ρ�vֳ	���� 3c� �v�:���_L�k��ܝR_?}XB�v�-�L�oUŦD��[��:��:~����D�������5!�y�]�QO|��M�Y��HܔRg*-2�LImH�gُ�:>�i�V63����DR)��3Й�c!�!p�}�8| Qad�R�e �)c9/d�[��g.E�U�}Vs}��g;p�ŧ0�X\t���u�O��+��r��}��+�%Ɇ�� ���L={�ڜ�s��b�.A������W�����.l��I�l�p��Z��fQ\c&��-�^	 �`�J/!��z(����"�<U�!/b�b�f9�'���6ܥ@����/��\w�p	Y���:*�׉p��<�`��F�,�EK
;�מP�.9�,9\`Ϭ�����R]׽i�����/�]Ϥ�҆a��+UÄ�/�`x؉��UA���S����o~�Xܾ֡��J	���iG�����/G� ��F��a܈�r�8�a8������|�|T"��u�n�YJ^{��)�؈�2���U����f�6�rn3��S�Nt0�ူ�<�e�HS�/5z����<���Ü!ecS�"��d/��r�6��@����iˮҮ֫�=���~�@�K����`?7n>~�FyY�R� h�ȍF�N�s��z+�|?eƥX�J@y�#l��Ty9�4�ܒ
a^X?ڍ:)��&�2}��@�.��#�~�y�g�H�5>�)�pE��9�����ip+�K0a�?]��uV�Pu�+���{Jr�}Ʒ5\�H��m)p��Rp$�
����6h_#h�S�V�(g�l��qα�.m�b�}l		�5Fݦ���)-Y p3yI9aNӢ���z3>5����t�t��%�w�#Ƹ,JN!����4u��Py/�0N�K��{퇢���v����7O?"9�~��uڛ%}�����0�:��� K��[KA=۸>Nt�z-�ý�@���L����O��_��#�lú��uX�#���=��B���?�ڥ�ϓ�(�v
tG���M�rD��όgN�~Cb�M�<��]�絶�ujN�K日T!��AE�)��0��$��|��X�ɏA��t�o�yAO��Kg���l�������x)����\B��E/����׌��=D�<=6�P�x _I�x�Rռt_�Lg��7;d-�v[ͅ�+�暬fx�F�U)�=u4����Z�ڦ�k[��!����&@|�o�.W.�����N�h�@���n��?���@���̅�H�|K���}�!�w�&y�R�*�b�<��": �>������]uc��:�~�
<�4�] 6�����Xt]ZS�����315~��2� oIh����A�%@�e< �Sio!�74�o������HLG��M��3�3�%"��fy�SN�5J����l��&_QT*�bPC�7��ߪ'K�xQm&�����zrJ��Q���-M��^A��T�H"�:
�b����J	�I$�.BZ����
������dX�S�8w������|��=o�~X��J�_����ۥř4�B;��h]h���W�l!�?��[�wi��t��7�T7��� �c����0 ����K7���m�h��S��^Bi<)�	�n`��S���n�!\�6,�3�ڒ���aѤ����m���g�[��Wz{�d$o��83����-��4U�t�v�*�]��M����V�(!!)�亷�s��?!��������$���:���IxB��$�l������wl$���
 �8'*$5a� J����X���1,�ѽY.�/%�bUI@r*!�r�0W�#�����M��R(
`� �eN�S�SNMt��|0�ߥU�p�F���S>x'b4Y$�pʍT�!5���9r�f
ǲ�AFv� �dC�SN�]���}�i�z�K�`jr<�<�B�תq��p o	bO�����@rD�Es�w�uTfk�c)v1��V.@(O���
��I�f3�%�3b
���ۗ��4�_��c�=L��6u�A
@X qbcL���0�l�����7*�sɻ��͌^m��l9��i����J�y�)��e�� }��h7mu�;��:v<hn?ӣ&�=�������_!�3�/�3�;aߞ���
�����ܔ��Ó�kZ8j"�0WPY���T
S�;Jg�6AaQ��I0����6��D�sU"�5, RD���\�R��@5�=c�N�C���~rd�@��hp�.q��������j!�O�� '����'d�_�<Hպ�V�^,��P��'&٘�0C�z���+c����}�,����P�:C��sb�R������ٞ�(�0ݛ]^�3��N�+ڽ۵�nF��5<{�������`���$��}y���l��W�fxГT�l�w�,w�M�2Ls�X<u,�ep=���ң�"&�x����04�:�;>]��c����Ŭ��_^�����V�N��!��ѻ�+hc)�n��>l���x�I!�p����U�G��b�K[ڥ�L��?1��ީ-���n�*)Q��M/��x��/���۩`�G1g^��$[Q�U�I#"j{���S��/�{KG��d��4���f��;X��-���n&Wh�%��l�j�`��^�5����,iX��Ͻ�����<lE��ʍ���	ϰ�Ć� ,Rnܐ�:��zgv�J����S�� ���K�m6�5ה�<X���`�Cojb�@Y�P�� 㪣�lqŻջ�`&dt���
`&VU�N1�s1B����;�"�_�lpO�Hb8�DU߳/��e����
�"x[B���K��?=�Ӡ�V;�������sE+f���q�M�}��ԡ\����q؉�m��ݹ3@T��g��̘��	�L}M��h�Q�_��� @���D���,���g��� 1��hx���O��J��v�>68
�҆�(���-6R�r	T?1W����vm��j�\��BgS%u_N�I<���bt��X�����G��x*[�&}1B��Rl��RA�*L�+�=e�v��t�uL��4���渙��ЌƷ�_�����9���ߗ�hc����7��-�2�	G؋,@�+y=�󚎺+��������d.����L��Қ]5��;�h�R5�i�p8�oJ�g���p�	��t3e��&!j���d�N%]�������ޒ�Zc����.=�VUQ�/y��\X���
b/����'+`)Dt����$�Ȇ ��&ݜ��7�W!�M)�P����kD�ǲ�rت�L��b~��L.^��\*N~���w(�_Q�_��3+AG��u�����s��1��`����][6ǖ��/';��rK�b��j	;`8Se}��*�>!���Ǟ�:$>��=&j�O�;���(���8ɜ4�g�t�h*w��^�0h��N!�$� .<,9B@�D�}��Sh�2U{�l�&s���)ݏ^)8�.y���,*r�0��1�j�aU�Yg5��7zW �(�� 7�7�j����_�G�r$���܉:��Ȼ5�"��@3 Ϥ���"����X�r�z[�I�&O	�o�����c���[GO����`�LbR��]�)ļm�|;.+Vq�2VR|�s���1i�R������b�ā���]�j�>W��� ���R�WDi�,|2e=&����% �� m1T$0�L=%1�&�1�XƝ�Fr_E:�FH� `x����o����*:ш��ֿD|"#�S�0B
�g���C�;�����0��g$¡1!N���7S7�%��G$Y�Zxn��b~�3�I^*։��MHb�R	�}���%,��o|̈D�QFPٟt �'��l�<^U��=,g�ps1��F��<%R;��U�Q��n`Ѹ�	 4n�:���Y��#$v�4��K�|��1�cIˤ�6Λ.#JY�o�m���v˃cwj��.mf�;���_��싯�O��>��ׯt�a��_��i}��������FW��(�>:����}š��C�1g�k�&�c�̗	�4�Kp�|[P��T�,���%������+aE���3$�����,�e�s-
j
�(��!�{��	d1��b�-���;�B;�Z����V
X|g� &����_��S9�4�`�
����o8l� �/�ئ�50��=�A��.xacu�v�� �a"�td��Y��̉�f
-l� �'4�ػ�Ty�{-`VN�zy��wwj�����v��rd��/~9��ׇSd�
	��d�^���C2C���m$Х�%3_�c��%M�`_�E���X'ŏ\K�RQ�GJz:Mt j��B*T&��F����j5�W1+s�L���5��ݜP�
�4�$��7+�,4,N<��|�m����rCGE�K���Ө�F�W���D����^�NU��ƽ�\h�k�������8��UvЊ (�=]��m�T:\V�|��FP�i��6I#�:DG>*E����P��=�d�aaW
�i��̶���6Z�������>3�ۉ���j�����#^�h���+��
Kt��/$���Z���+V�C0(�L��9�z�  s������ v��`���X�]�xC����>�D0Q����Ë�Ā5T�Ҙ&�;��R�v�䔅5k.(�J}]��0kt��Ʌ=��;�����0fug#��׃�Z/-z�
\���C6���.����~��x싂1�mun��dJI�J�>����j�͓k6 ��6у���q;��6��c�f4����M�u�mLX7!Z��l�^�bb^q��6��Mg}`�{θ�Qˈ��_VP4��آ����أ�f�ϊ"*ٞR_�\GL���BW��=Z��G\�o�)��)D�şQy�}�K�/j�n�j0��a���v4�I��Aݪ
��|��$N�A|X��n��F��}]@����~�4S-å%�ګe�l�~
��?�,EG�Yj)$�k,����oU\^�:��-�\��[ծO���`Z���|�m3�1��,Ln�<����NR����I��oi��6�����p;z.nJA�y�є�OPlJ3�u|FA#Z�3�D�\���adZ��"��3�GV���RT�A֙= �����;���tō�Q\2=�22�o�H��ųf�J b��Q��v2���<Q����=R���漰|o�����zI� ��NZ,�`T�8 ��[��<�Ng`"g92���:��b5z���k�������̤�W+	�S��C���]v˸�:n�m�R�7��f�G�_���荵��ˢ���}.aX�Ĺ���.����fm�Ռ���z�{�8\˯�#�W�Ч��K�?�����%W� �����]�r�M������H�	��`�z����uz��SVA��(�.�k�ɵ	(6�⁐�%�'�~�x����ta"���u[%�,������F��RѸ���b�0�#j��O�����GB]��i�CJ�����!5�3V*$�@�JS��y���[����ʭ���/���>��+��H6���G�q®T+�&0����6�"強��:{���輕ʽ5�!;t^3�<�غA�j"�m�k�XbF˱�3�Fꮌ�K�k%9�Lj~�R@�~L��x���A�Z�_;!Ƴ�j�~|.�q���z�t��P��wR��ǂ��0<7[vw�<�VT��{<��!um)�R��&wJ=Db�^�UJa��'�b y� "yz��@��a���F³A�|������e��?.��P�.��7Ģ��,�'����"���� UD8�::�s����8��Y#��sbPRA�˺����\�9eٚ�rƥБu�בS︭ؖ�?�o.+�8CT����mǊU+s5�n��}�DLm/�)<v9
 �w�������4�ɾ[�����%� ���@�D�V��Ä:�bc8���e��)tPK\�5c�n��w?�U"%�-�<f��+�H�tT���J�튆������� ���V́��\���K Hފ���������8K��p��I��Lw`?	= ��Er	JY��ٍ�u��E�#M������3��1���۴��焤��@�����6wBp�OM��T�$����R����{�F�5ۻ�X�`;xv9#�{ZJ(=W��F�7�m��f tbѫ�{h�h�ٟ��`�b�*7KF���/����'wI=�,Y���8ުj�
��a��S�T_�i @�}ك�6�y���0L��,�K}G�m�N��Y����x,F�$��#<<R#�`��z�(`�'�<F�:��Wga�e����N�� Ϳ�4. �$�"�I9{�؛��1ѹ����4������<����T�w��<�"\�[d/��/|�h߻��_CZ4$�=	Ժ;1DF�߱?�����E)X����*�E��=��}p!�ѐ_�A��ȍ�(?��t��h���\�Bت/�Ss�Q�J����\� ô���`�GZU�v�%��W�!�^�m�6�I�S,�f���k�p�)�AlF,�cD�1��g} 4��ع�p7�ESrG�6E��n&	�>}nA�N�#	1΍ĥ�,�U�	�b7�^�NF
�bX��y�m�U\�p����gf�~��Ŋ�b���s�f��P�;k1ꛙȸѳ�R�]�5�����<��B���p��~�Ѽe6���5��U�e����c�dh�뵧�vL�"k4צTYs��������������o��'�CT����A��ߐ�޷v�V��f3Xd�3@!�H��7z$�Y�޸`�'9�n�ꙬL~Da��<����>�n�\�&�3꧙��5���=��,O%�c��n��!��W��hD�A�WQ�v�Q��c��yc�P##5EU�&#ݶ���$F%	��U�J���4���9���U�$,�`�W�����?C�m�3�tE�W���0�w 
���V���ë,�{��Ϫ~{�,�Т>�a�&� �'�P�����>9$�{>f.���m�Ϟ�|`�s�r����vti�%4������$%��q����Ig�פ�������sa�����zM�).�C��ķ���RL�M`�F7�b���|���h����P�Gy֣-<4�v�>�oU����W�9�q�~�DF��)���j�2�����U%�=�e��=��V9��?�ʻ��{1֢��<���@��B�yl�H������+ڎ�5�.���Vǈ3f6?�����D����� an��"�G�0����R��b�jI���q(�������*<�F��Z��>nj&I*{��7����v�����5�E9e
2����:f�e��2 ��Y[$���n赧Smc��<��4�E����K�y!"p�O���60���=c)�\tq���I��Dj�`�H�����q�)��><��D�Ҷñ��E�`>��H�7�v��"l�uSC_���L-;������%j�̎�{�D|m�v�G_aiH�^'S���T���^�_�n�"+�Y⣼#ɯ�#�8�dY��^�7�uh4��4�����|���'l���;=8A�DO�(Lpp���֘<���9c��F� k;$��\uL�Z_��Z�&����}�D�"V�B�/ʶ���7�O��J��W�O����-�#
��z���]4�ݸ�K�z .Vu<c�˵M ��B��Z� �M)�4�s}��`9Y�?:9Rgfj�w®Ť ;֐:cO�)�ǖy�U\GI{��"!yp�G�� �)+B��t�V�!�����)�f��q�SW��?׶�_ oVÓ)��q�{�A�+rr�tt����E�Z�Ƽ_�d��@�T������p�EI�8d�\���d���rm)��lQ(� T*�a�`;���ZY5O����Z�=>�@�Ȼ��$���O�3�P�K..���4E�nf*v��3�P����k�$���+-�x�Cr�t����A�g��(6h*���������C�>���m1A;i3�?ݯ��䚔�wY��⛦����%��d�'�tb�,��X}�?'�O�� a8!�Mն�%� ����C���q�i&rcv��+�Ns�up���3=�{Kϓ%I8�����\H^�H�Y�MFZaԓj�l<��z�@\a�����A��͠�By����1�� x�my7�(���"�W�Vp�8
@-�Dp<�'Ԉ��Ynj2{��n����_�k�'o�!	GL��^����B׶qL�C�F���́h�1M����j��U�������uM�g�����@"F�+h:^8bVt��w�^ҢC)�*����?����j�8�p��|�ê���s7K���W��z�����4m��Dg�X8K.��>��*g3���3��c�����h�;p���=2�K�lz_�6��� ��o�8�>��ٺ.�	wK9v�����Z��aF�,�A�ႢǶ����2y��1w�����g�X]���K�<BN�]?�`��<g��Y��*��+VG�-|�>
=Q���@�,����;���`1�$\@�L�;���l)��**�{�O�v�_J�8������i��BV��%.��A�w�+�܎g��pd̍P���)��"\{k�|��'`��^�v��R-��Np�^MK{�ʺ{%��8j��=G��B���P��,�D�I�����s�&-�.�۪���[��&�WLh0 ���%���|ILz}m�}��շ��k�'`��a�E�h_��4��NS�3����m?x�g�X\	:b`�&�Ojf���\��!N�]���z;<>N��@'�S�f5,ʵ�ct*�TMѨ~�ˋ+��+\�-���zzLG��R��,e�c�=}�8���_-�+~��� �J��7� ���%���@;��!���5�Q�b9��؄K�����8�a���ͳ�'� <c%A��+	C��S��:m�@J����u�sV�� fk�4�їb;�JB#�Pʐ�;���� ���2��/qA�w�ޱ�ܥ>��UnZ0>��p��d����Gdh���#���Z��g`g {�Ǹ��\�f�e�e[g/�,K˜�����.�Ĩ���.�OJZ�D�����	�{�U���Qz?\6ǩ��z�Ѵ~{}��N2��?��8�vvu
�$��ա%� `����rD����I��#��<)��DFѭ,� �d����tj�3!�`�=�0�p_'�1+�#Q�$u�T:4��2������i����ſ����/�0X�n��fo���!�aT��)�xp�W�m6c�.5۲H�����K�l@�̜�{��3�:7C)3�;�(3/�
��W��aG]D�鳕�u=$v�(�݅����a/2ˇ��jq�3b�+c=@�6��%$�(��?��Q a�3�1;����2h�e�c2u�0���l޸�N]���Pȹ �:+��<Nud�Y�ϔ���zRN}��SĻ�TmZ���1����C��x��*fY_�5��]v��i�q�lX�$����T=ޱ�(��-x�H h��Ǳ:o�g?������d-=��w��טY��j�xԊ�NJ/_n]Ѣ1FZ"Cn���b��6�Ԍ�����b�ǅ�=�9XQ��v1�;Ƶ��Z��qv8d��|������.)�$s�b���$@zǠΏ?�,Y]�5�f���,At���Q�-h5��¤�6����f���j�s)Io9+
c�ΙXPj�{*:�U+|)�;nKWvY_ �|q��>O����?���E|�����F�/ʏn���Wdf]��{5��fZY����lj��0HFZ��(	3��l�[�릣b��u�g�j�T�8�7i���w����z��W�L���`�"��U��Y[�2&��y4�{K4�m�
�c�:�>��o ��IF�|�����+u��Mԗ���|�Ԯ��y�)k����L�{���W"�Dmo��{�f�Y��mS�Ԍ���5�[�ǭu9��&cTs�ߢ�'O16�r1TD�����J�zUF�	�\ct?��
�k�l�0��wB��u�+J����R.��<M��&z�B��`�`��j����~��Rr��*lv���g��z2<=/zU�1D��ҕ���Xۗen�f'D-�!dm��\AP��5%��W;S	�������4Q�B�ҽG��|K��q�]��J�e�~pU�:�aݬ@���U��mĝ6ȍ�D�A�c�i ���+�D{W�"09��}v�1��R�����\e�g/�U�s.{}>��j5�s�T��9���Ɏp-F�[œ�3�`(�5�܈oU}咨;;�,�Y��z>�DOj�r�i�l�
�~ToƲ�����R�)}��yw)����o�NW�-���+H���u�hX컜�4��ؑV���Cܗg1H �+�~�h6VCE���Quۈb�Yݳ�O��.�$o�t�9�3���کQ�R���?b��b���p_
�Rg��Q�#~�y����9h�PV<�/w���q�]���X��݊�|��H�/${"��5O���B����.YՈ��"9	y`�C����k劬cq�qߺ��� �nl�)~|{�a�yo��}�Ԡ�QG�MoB����7,dN/�+!��V|Ȗ��}��5����7kp�s([e�_�:�O�x����c[U�h��n���h4O!Ix��ƅc�x�sN�0y��A{x��p_г訄�|N;9w�/N`A;��O�L'��"� Xn�Z��)�.#�J�v\@�[?�}9��_[Lج90�x�h�����3ꛀUM0?�PS�`_;����4�TK�r��`�ŻVB`��V�I���&�?�>�3�]_�k��KD�s��>�C�m�������!�^���}���WX�`��3>�R�(u��F���HU��CJ�m�A�p�~ڽl��->GpX�RPYvls�w��
H��&G���F�F(��ur�*[F7�m��m�m?�<ov-�	�x�y�\���Q��74Z{z@j�~���6g<��)P ��jJ�E�2�HW�Mui����A.�Sf�O:�=�D�P3VHR���衬3j�KEy�2����'p��6;D��y���`[!ѥ���>��p��&5Gǈ�f]���e�:J��e��L��뇕I���.���RZl֠�(�����W�QR���+z��S�.����O�FI+���$ ��39���'K���X��Ҽ��N�̉Qj�!)����?�m������;m��F�M�����.��k����^�����q
��0o�DQ���E(� l1�]ΧZ6�;�+�f�i�0�s����:�o��T0�o�����3/X��8̣W�~Xt��H{�����8���g~��Ta23���6�8�i��HJ���ni������� R<�a���<na ��.��6��R��l�֙�QxR/�7��Z�(	Ѡ+eFXITyoE�r�~�l��?�$)Eܯ�Y0��.�߻��4�u�B�J_�q�6eVw_�(�+|�fq8�=���=�+CF�E�ۜ6}�:�g��(_�	�^���q�!��侺���ju�\��`�_@�;|�cVQ6ʿ�ѿ%3A��.������?���ZC��5{3b|��o�3t�$���Og��a��(kyi��ؑ�)/-|-l�M�~)�)"�����&�@T��
��l�\�F%Y�������Fh�I?��b�r��v��L!�}�C���Jt���kQ�44(���m`�Z���4�1�2f`�tð�8\ Dd�j�V�1�~��r1���(|�@�o�#���Ҝ�6�I���y���m�o-���LeY�P��)[fS�Ж������˳�cq���[_�h��5-T���:��?u��,��Ĭ�W���� �W�-���v�6���P+ӕ��نK��O=&�<LKǇDO�� �+c�p�!�˥7���/��l<��Y�U-�!$2�r�9�8Iꏷ[_C��3V/�=�t�P�9��Cl]Q�*�f��$j�P�_�r�=Tz�Л�������s329v�n2��m=&��b&^dI�7¨w<�"��!��>�6ֵ\4N&��`�AѭȽ�EX��5-Y-6��ٟ:���ۿ���'O�21��7g8�B$S��O;REF.��[��@{�V�J���,�zZ�����_Cb���&i5y�I\����d� C�O�\�+o[�H�?�;:Ή�Z�%b����|@ҐXZ��p��ۮ�7�y�b*�,Ds恰����=�ǜ���C��G��gDЊ�X�l��m'������S�����7��Ju�{�����[�j�H�J̪�%���X���.��܀d�u�%����qeD2�܍�c织`dS�Xa�l+0���m�4HO���G��s�A�4�5w:K�e�x��������'�C�ľ1�C�]T\�A���H:�N���h��S��0����mU�����s���(1�&���7>�QY%4��$+���r��Y����c;�a�	���?�}e�N�Z��S��\{�ٹ�º0�ư������Vg����ӶS���Ƭ3}5=hq���cD4����=��C<\�[dVd���Ø�-�?�)J~�`�VA�z.S��t�e	�����S�1�-�M/M-��{�:����༬<���~<1�?Z�f9��'�]k������$7�42B��A�hH�h@�.�����P�#2��{��� �y��H��V~#�~��90�����oc�_�"�6-0�NRߑ:��*�����%QM�oуKص��u�A*�,Mzh���W��F�>�¥�c�<�f��2%vd�G�˰k�Jn0���O�^���e����Hk@f'���1"�[���W�"�7����F����7�,��wd2���hDu�J��sk"஢����E �9ϛQ�E��{�����%6���%e�loRrV��:Y��},�������v���Hg�l; ӿ��~FtV��C��_��c�f��b���6+�į�8MYPg��ⲗ�l&��i�[-k�Pkw�?��J��=��0P--8/kt��~�l"��T���7��e�T�n�cM?R�Z�ѹ�Μ�?��M��Re�:ZU}�|HS��%|���Ң�~i	O���f��.�/$�(��smJ��-`����RsTp�M�`4h|�I��,5���o����ӟp��HZg9�%Mۼ�-�:H�u��|F!��m/Mg7��3J{�����w�k��׾��4i|�ˠ��˩�t+���2��gUkGa��q�J��J��ɿ�Y�E��p����Yb��T;[���:�w�v��i���GyX�����*]����܃��Bj/�n�U�*���S�+����{A���`%��58���`esHYn+�\�\���M����6Wy�oG��-y��S�����dZ#Af=�[��5��y���*U�J/�y�6au�h5Sy��>�|&�*k.U�Oqպ���Au��e�ɨ��:�l���}��[ˬ�n0���LMӫ~D{�cץ�a�_�X�"o;��3t�ط5�ܤ��I��_{>~�Fv�Bw� #6�G
1��'?�D�I�����T���w0k/�K1n�mAq$�b)�2��#���n5���$P�\�36�`g��J䈺����H�X���������ce�bM�����3�EU�tX��C�f�U^H'�6[���nh�B���{�xZ֡�ɳI��F���ƙBޣQ�$����q�ܶRKQZ��m."�f���U�vMW~�����yy+/%�����Zؾ�:�4]����q� ������}vs���R�QJ2a�vR~u�Fn��m�ܱx^ZmY0��$N�6��	X?)���뜥$�3t�yP����KB#8SSEE���ߙ��{	͹o��]�|�/�}D>L*�y(�]�N�����a�[&!��&���j�4�ʈ����w�a����38�oO�y��ߔ��g�3���K��nt=O~�>M� tw���k�=סڤ��k��+q�U����h��
�6���uF.��@!�������;���Ewu+%�"A�Q��5k��K�'���^r�x��[�m3����T��jYO3�EŞE�A-FG��|G�_
#��g�r�<���� ���bk��y�A��H9�\V��ʻ��q�\LV��-½�����߇�Z�ui���,�O����#�-5�ͫ�,�v����][���(�>O�^�w�`�v�`-E8���^��nx���?���u�|\�=�7�[�~�خ0
��|dҡ���ۦ	��?����n�K�l[��,+nDk��9&0\�[�Q��/?�b���z�S�vu)[�X�SJ�,_R>~�%D�K�9�$2�9�w�p�nđ!{K\��_�v1y�?!��ԙ��	\k?&i.��%yHuu vpX�	��|!fΗ:X����Z��THژ�;����랟��Zl;6�G�,_��	,V����v���02�[�ݹ��Z���.�޿6]B� w��&:Y2J(A6t�iv~ΥI+�QԦi�����+��������{���p?#ٌ;�L�Ң����B��7�y�(췞Ň�7��g���/K��Վ6�6���d����-'{zq}�u� ���6�H�y-ʽ;Rᨺ*�g��?�\��� �:���ܺC�z�XD�RxS`>��=��]�\��dS<L��u��0q�|��Iy�W���-��eu�X~��`_"� ��`#aJ�nn��m�M��G �R#�5���$��[Do4e�����������~4��(�IQzT�&�)7�)�O�e�Ȼ�j�����/Y+��`��Ë�HD����J���v�ڙ�0?/����=-����X�pi$IH{)�uPx゛�2�ӷ�]L�ٗ�`h�rO1�\Z6�wԯ��Gh�⮄����kx����l�� n����<,G����ʛV�%�U���h:�rt4Y���	��}j�^�#�5��YV�{�*�"�b�=b>��E	�������M�x��?L��~U���	�d�/,ҏ;���T`l��lR��"�	ڵ�`�ʼ2[����Ӑ�s��S���W�'H�B�#Cl�v�I*�xfq}����z/�������a��u�����|����ך���)c,�����	�"L��q�M��OZ u~�[�?7���з����]U�<�� J}ݒ��@���Jfh��ߏő�s�����Nk����C9s�~�Hޠ�vn  -~v�}��2k�X��p�����]�Ub���,k0���zi�`�S�g������y��>���ـ̦�g��Gz75z,`��/��t�,�,ny��.m��1㝱����N��wog��( ��� (�4�4�t�[vm�-�%J�p8�2����T۠N�oY����K�D�ܗ��2�C��fk�o���H�Z(�>��19�����6
k��2`��Mh�ޅޅ?�����lҜ�_��������e>IΣr���CX��hh`�*�t�����1�'����E�'���x5�-�C���Wў�4��W.��V2�n�յrCn����[�z�Y��h�,b��(�s4��1�.f����:�x����yҿQGM����:�q뚷�ڳ;'R����=̞Hϛ�O���ć=Zc�AxV��ed�L�B�=(I?���v��B��]��J�lrtz����l�*���������_���	O&�Φ���dn�a�kAS�@ M|���@�u\���N<�ƚ��"����UC��p0�I������>���=u�~0
S.�Yܙ��](F��W=�dG��)u��(N�8wU���8�]̯ N��+�0ކ�v������[.����ف==��g"�5�OB�߮�r�_�T�~�/)+�+��#|& �T��ս��%>�����h�b\��e�X��?���Bk����@)�#~E�L�;ej9�������^��+Y}���>�#[bm6����TW�0����V�T�?%[�6�3~�g!�aŧ�!ܨ��4�N4�|��� J����݊:]����+y�*O�rfU�.���<�L�K�>F��{��$�3�:�����1��+"X�Šs��}e���mHm}*��BⲸ�_��s���y�kF1T�c��/��}�p�.6,�0�����9�	N���,��@��0M͆�_a��e�x���4��6]Bʾ	^B���;a�^x͉�6��EgSIC,)��o�w��ﻳ�[�껫/�#S5�х�$g�2l�|y��C���W�Sb���U���R�	����B2{�+�e)���}�V��>(S8��
q@!f�:��<�6/7J��2�#�g?�I��g��� ##z�q̊1��f����[Ԍ��%�j>�+շ�$��>�Z��Y��7��;VS�������&:کO�<�"֊�G������g�̍�H+a��l���/[s��5O��0.�G��og7��mr꽮�T��g!�:S�.�rlߗ�Q���H�wN;m�Zd�1���Ps� �HGoȪ��0X�C~��m%�gfL��a���r^��N�X�ڋ��qm{{�f�T}��Z,6�ݸ2' DՊ�g����
|���@�CG�8'=$xЦ���������/����%������Fqؘ���V�l�W�dyd>�
��j:��RG����$���P����P�Ιj��_��8��~ܔa�m�71	9f��1�A�ܑ���!��s�V]9����x�������xD��]�X�[-�=��H�k�΢�s�T̩9��0=��А��&�E�@��S�G?�&0��n<�4I��y��:�����F��,�u���$%�BL9�Aj1���=� ��a��d������fp�ٓ�*�Q��7T�컎�=���w?δ��[o���J}rb-�k��؁�3�8�p�Eq�Ч�.%g��N<m��i9g�j����B�8��t�^�p*�RJ���w���`B�N�1�`��b��Y,L;.�����;yz�2ܦ���BD�O��������}��3�w�KG�0�tMu��V=���6૕�z.�j7���;\�G�.�Fe�Wl�.5O'�ݸ'7�NL��I{~c �[���Z��t�S�Q�N]�w�Zoñ�U6P�\�W[%����bréI�4m�C	*#nW�:�Ϝ�6J�D�\� ���l�ȃc��ru�˞쯣Wo�p��)'"��i�Do��
�^� ��F~�{��u����P�
�mZ:x#o�Y�];ārR���*�J�^�O*�^�����3#��	q2��'2\+�X2�ű������w�8m!f<��q�Ձ˦�-��5:�+�����J�}�)�����o����6'#�B&�/e2g$Gx�v$L0�� ����������(Tޝ��&5�[�ba���:Ĩ�kR+VI���zD�����-���4间C������kʇxx�_�(��x̖:�V�)U�0c-y�8��b��g#J���1�	~7�|�Q�aIG�c�:4�SK��㊆�:�}{�`,����q�����WB*��F���r3i��4�M�x���n���Pfu$Yw0Ϡf��v'�!���5��o����ӻ����m?�_��'�%g��&��:7�^r]�uh ��F֤��x��*'UjV�Q�Q�Z!;��R�J�t�1Z7tcI�E�d'G�k�l[�rB]�W4WMWܲ_��8Df=3wv�5���b�����G���k���_�<��x4���ٿ��ҡ�sΔ�ӕ�B�`��� �guHF����o;��[�$�;=z7�:�'G�:�o�� {C{ܧ£��v�n�L�$c�ύP0ZOH^�9K쒷�7}�(gܩe�3`���q��x�e�s�Pz��]/���g�������Zm�#/\�^��[�2�����٢��Ҭp���w6�!�H#?ӭP
�{�|��$Q�1��Q�i���8�Ae��l���q+�p6�ƍd� O�����(u���9�5AЦN���͉��&�5��sd���Y��de�(�i��)��_$!MǲjJ��;sw�Ds���̜"	�ko� �Àr�j�]|���e�Kj-��X]��rOx6����tͽ׫_j� ��7\S�I�3��؟���i����EL>zsb���0�-(.y��"� ���,����0��)u�F=WJ"�*wS���~�[�Q�E��M�	�!<P	w,s}�#4�L�� ӆ�'�
�ļ%�c�-h	�\��S8w	��Om~6l/YE�N�Y���g��|�r��Zx�f<����b�a�����;�G3��`��]��Aq3>\dɊ�q����I�4X�_���G������ M�
����D�I��3����D�O��C*#��k�{`���� <d5*�9-�8Jɨ9�iש�a�i6��C�1�@)��/��3����냭+T]EG^�y?�+4|�Τ���&�k���\��r���#��u�x��s�/T�0S;�<��.kR��o��>z��SED'H��1��wn-��u�J�L��6�:��o��ʾ[l��7��qc�7)�/^�8��n�?a��k�M��Sy�\�Vۑ��¨Ev^�LC��"���xL
�Y[�l%�L3����i��fAn��d�k�y������y�<ɏ�S���Jq,C�8���ۮ�x������*2J��Ӌ��қ�5�� ��lW4��\��`,�+lR�N��+cm�~���/�+���UNt@���rr�-A�P�pv>1�
[�Q���yF�jJ�į��e!^�ޡ��3-��ߙ�歭��9��_C2!̻���^�����|	yl)C࿤k�E���]�~�Z6���<wUBWp��>(f�Ζ����gޱ�f�|���:���T9���:��r��E1Iu�ս�8��j1��xnv��}��ы����%���@�?���e�H;L�z�:NpgB����؞��}$j0���=:�&��JPr�F4��U8qm���p���<=7��epԱy		E�"}M��.0�og�T�g�zoQV��~�Ň�1�;i${o�!]!F�NRl<�g�T̷��*;D��)�n��٥�x�HJ�G:����%����P0��OM�'�'m�
��~�*<��i�8̼�_�s�א'p�J�����j�WIyt�M����db_w��%��k�v~&/�[��p��o��`JO�}�'�� %�B:,q\4�$v�)Hh�˓ơ^��%p��@���-L�ް�l�[��������_����ǩ��}��dɪ�@\�$������5���$�mb�v�H�(�~w6�H��0JbL�Zv�)R�<y��P����J���%�1* �~�D���Wr�b��U���8�󒨠���(_��5�V���
Dp%@4��T��Ǽ�?�(�9���� �^�$��� �%
��01'�D�E�O&=|��x�S�̆۫?�E���w5�̴��޴Q�"�1������?,�r���kF�ԡT�%�#��:\�J��~�>@ ��(R/3����H3H�)u���N���XgJH��#Up�h���4zr�&�U�w����-�A�*	������[=c�Г������˱C�ϖ�jS�4���Q�)���"��~J��)6�jI:�)�12�[� Z��7���N ,��4B�a7���9�8�v�.�n���k�~�V�k!s�����K�Z��*����CY!�&6tIM�W�*C�Ѽa4(��|d�)����v4n��km��ޭ���:�V���8�he��Cԁ؟�G��cS�Y�pN�\>&�<�<����*�(�[_��t��E���ߥ���ů�(w��%�x?Mo����,���
�t[��_RJ����t�l��� ��rOFTO���3��pdy���s�d��W�2c��i�&�fN͌"⤍XX�����5�)��a+��.��+]f����h�(o�Qo'����s��� �N����������}��n���$8^=]|�@�J��~!�aU�P&"Y.$D���)���t5$�`��i�:q@�(�Q��M-�i��(�]�<�D�l��#�*^�9ٯM���{��ʣ�vD�o������Δ��A��`�cZp7�%��y7���@�Ϋ��RAy��$0��3T7���v�pp�x�'3⒔7�m8U&�ә�A����t���aj2��]9����~&�-�����a7%k��3<�CQl[�r)@���F�'F/R����i�.T�ͥs9�GP�3���r��PF��xж	����%�A.c�ab���;�Yf�^ж��OQ��Z�0�:��FF�m$�u"=�����cd��AʏPGM>��lm����C��� �h*�!�(���fwO99��� �;!���Ǒ��M�w؄�����9hHL;K���Ƴ4���� �Q, Ch��Q�V���Y���{��M��l�����v?ѓO���+>;do=�GKhL]�m��9SX�(�@��(d|8�,�
:�M�P�2b����=��U����9�⸽)�iٛ��7����?:+�8���Ĥ{l��$�ǚi?��z�[���j)�h�SJ�͠�&9���Ŝ�Q�i� ˎ �qg�lae>�E�� �ˡGєgVI��O)�z�O;�P6�!���.��vMN�-�y{g�7�G��D[$l�z:��D�̃!��N�l� d���o	��R?|wq$�Oi>ս����������i�_���ptXy��L����X���&K�����I9W�E���%A~�KE��qb[��B�V��|jr0�ꑮ!���uK�	��1����vK�m��t���M®aL�tW%��?(BK���)�n��W�W���sM	�3����|$�"ޑ���Ybp/�«b�h�59=E������2Z���p�ь�3�ʄ�4"���
��K����`�g�Z�&]&��������d�� ��"��P^�ܗݐd�{-���d�h�k���6K*& J�3�f!�Z"q��������m��h{���KE&��0�����.�*�Ҕ��Yh&��+|�����7?�Mf/��3�����}�1uݣe���}��TΦ�Z����Қ��B��b�ܥ/0���U�3�r�_Q��y=f$ǔ:���>Ppx�[�՞Uه�f�[�<M���6�U��k�6N YW!�f2�y�Ӑ{�`�bN`��扴o��>�UPJ����]�%+A�X�,J�u^�ǎ�*Z�'����#������0�b���0,�!�:jq�ŀ;�X"�ǹ�=]����sq��n'�����p=sN��>�a�Z&Q)X��#��Zu�=1������m?�A���E�Od�ы�z�%ġmҭ`�*��&�5�Y�k��7�~$�	�n(>q���_."���z(�S3xrpw+�v�'������'�?09�	`������o�"+���@-���Ua9H�H��R��fl#&�]�B�%}��ˍ�s��M��m*�4�'��1�<g3YM$�0	���2�_��A2�x���$T/x锏�"��������/1�ʹ�b?IHfk����	��!�C%>LZ�7����=^������Ow5����Y��?�0����=�6���g�K?�a�צڞ�8��qK_�~�(}� �Ee��`y�Z#��P-��x^�0��?o\�>�����ƢHk��n�Zٮ�4�����\Q_ݐ��N��B���nϿo�[
r�I��&<,��H�@��Jf~ �z�p�V�ݒW�+[Zao���-00 l��'��c�,��ڼM�f���q�v���kr����U��38�͠�Y+T���@8p�
�8)R�D�jz܄�Ϸ�ք|�F�V�����Yg��|�	k���N��6������Ԑ�������HT{�V��۴�kn:,,e�F&J�m9���My4sp�'q��#<ZBf�[���H<�:�,����_P	�Cˊ�?����M�R��Z<��Xo8�F�U�B�Zu+��+H���o-��'z�����O�}��aĩt�ł8�.'_��z�,�j4�3�|�V�8dDb9���6P0�hl���E���yy4�;�3���7<����?Pjt��Ti�E��!u)7Ddsm��'5���趪>��R�,g��[���ݠ��HB�g�]O5�� ���37���������~��F
ɖ_�$mpS�N F,M�s��2��0 ���K*(^m��Ab
Q�:^8LH�ʄ�C���p�{����4=^_�,עy�XY���7�A|�49~wpv���f�LL�o�����WY��J"DH�b���Ӏ�kdC�7m�Fƞ�}>�;�H��SF�<Ri�9�mB^\�L��ܥU�#���[�r1ǆD̀Ӆ�:S#h
��A5C҉G��^?���c;�Iaq��-xN J�a�9��/#�k��SCm�5[c#oHD 6��k��҄��>��b�$g�?r��,_0TK�������F�J
����_U�Ξ�"�X��tu��54c�pUi���y�Z��LT�܁qd�5�{~�D����_����Ŧp �C�[���p�g�̊��x2��A�y��_�����2ނ#PF��#��+����;�w���FoyZ�a#��c��o�U�c�%�*��rv���%�)�izo�g�wg��OR���5��{���Ri�^U���E$�"��x��/Z�,�f5i?ad�m���f5�b��[�����=HYm�N���z���:VEH@���-Ab!53X	�����Ò�{\�$��Ig)�fY�$V,ǋ�_�i�T9IM��U�Z�7"�ۃ.H0yk:$�vz�/e���T���V���r���~��T�����a��4u��&���f�:.+��0��k~�(E�~17۳ߖ�S���z��.gP����\��D��?�h �0�2^ʛf�E�?��������zq�`�4��:�C�ƹG;C��eM��[��t����=Y�]Q�yT�|���|�= ���y��O)@��8�/�{Ʒq��Ӱ�i�y�>���+�y����#<3����&8�.����Aٞs-���jU{�R���[ ����0�?bߟ��.����`���T�-��tXL��	�׋55cW�&��3T'���ckp�ЇG�zn��}���fn���.Y*�ܪ9�v������/�k��c��M��q�g�opm��C^4��?7�I���;����E���r�Ȃw'�2���ѳe���ܱ�@�8žo�!�'�r���>�����vn��g�V�Z�9�6Z&��af�W���&
#J�c���\W�,����k��0�����@��1VĠ�Y-3u䞇 9��:��7�^��I�4�ϓL�.�C&x�Ņ�90A���`}ɜצ���:�^&��=�bm؆bd��	�QbXe��&�����dc�VE��l�;:��u%t�/}\O3�\�ř>>�Ў�j�k�*?�d��}dbY=5���� @,b�d2B�s��{�޶�����0�<�]�Q@�p��0�A�qv�=�y ǨLׁZ!�ګ��c�w��X2�^����>��Es�v�̶[���*�-����g�Υj���ȷ�W��
`�\���>�+��`�VSa�ݿ�F�fT���tE�a/�����A����h���u���;��QU�/�z��E9����q"��c�6H�I�#~B�Ц��Y:L7�����z#a8��4
;Ғ!fR���k/(�`��2��2�+�����L	E�K�S%
�$�X�Wd}D���!P���։d�s�6����s��2.-gY���ْN2|�&o�ׄt��ܓ~Rh�����G��؛�@B�-���
�֛Iī��_t���ά����{�L�1R٬�i���^M���a�N���[�`�l$P���9���!(;��u������d)?�_����rL8��{����P.5�rM�M�����ɚ�f�Cݠ�c߀��Q7 �褛ۧ�O�Ń��ҩ:WՅ�|�'3�����5�����CȡpZ��EF�>�Mc��*��*M0,<��25¨�$x�K�E-hm��XiK��D"��Iҽ,�𾕔:U��QR)J��ógI�E�ܠFB}9��-=b;4U��Y�9�h[�
wuD�H��<I��^KIq�ei�9���XD���?\)�}`�|
Q�9���8��4
q�g�zt������D�l��J�1��ݦ�5��U{�-*�I���&F-:aŸe�S��6�S�!a�� 9%�m-����k5e���P۔^����k Q=�A�L����@� ��k��.N��+��f����8�&?��]m��Px�\�mؾ��yAqз���R��G
�M�R%�0�[�1��ܗ�Q��d{&=��8X��%>f�O�H[K�͈�ʌ �1][B�P�j��1��9���׃��6�ݯ{B��I����o�������x6�iN���N��&f�Q�#Ϙ�~pTo���$T�Zʆ����p��*jY��W1�0�}�e)��N�e��8[�טqG��e��`a�$>�$��L&��d}�1�
�+��	odm$�'('i�֞ߏ����)4�v���!L� �9�� TI�G��a��]�8�Z������Ik�!0�����ӸI�{���
���a��V��b�>�X�ZFPW>���H	�a�!�Si��#}����<z5���Ns)A�r}^h(��MmG�0#P�i0�H���$TbD�雟�f: )B��л �Vɡ�۳�Xi#�Ȅ�Rn��Z���[d$�ǮC�`����A8�_P���V��{�	
�A�<h����o���W�	�n��ر��ie� ��s���}r����YO��C7b����Bih�]��H1K�9��T�T�b�)>�y������5�u3^��D^�>�:bR�]�����'��}�`w�4��NCL��kC8Lx�,!�QǢ�Ai�O����7>���G��-�_o=�5\#����������S�W���F��>W ��0
<Y����'V���FQ�	�l��f��VM^=O�"2����2�ޱo��&ݞ�>uG���ZL�*���nh|-�	�^�ݡi�H͋˓i�����9A����;�eBx�X ���j	3���Y�S�k�G4��~s��C4��wpb�
�����X'�K���5�p�ї�IS8�!���/���O4Z���H�U2j��v`�l��γ��i)��wJ}��e�m�\q@C܄�k{O��@n���l�)�j[�ө1����`�,���9��c���轋|tXl�H�+#����������.#�T1���p����.���]����1�v~��.�y��������eˏ���0/u��n=��[)w��EQ�SQ�D����eIh�`���(�~�oV[��s��y!�EP��MΫ�ׅ��2���w���ҥ��Ax�,�u~1Ԛ(#G��ΙX3d�A�`���9�0V��K�`�7M`�e|�g�*�dm������I}c�,�3&$�Da��[e�A!��<�	�Wf��hAo�t6(hd��9Xc�/�g�����O��r!#v�Δp���,}MII��)CD�t)��7.b�Í�ڰBW��E�>�7�ؔ*���i��>��"Z��b_�*n�p
��+h�c�"����>�`�.�l�������d��S�m���g��	��(��jq��*җ���_6�����i��k�s�^���^@q�����?U_�A������h���f�~�Dgz1n��e{���Ln�3�x��-�`Q����s�+��ucʻpm�p��M�RQ�� � &4B��P_�=b(?�eF��	&.J��D��u��)�7�\&����a�.�,�=i�t�<��cp�m��<E�{)�j��l�!��cDd���L�mz��b�E4	�$J{U�k�w[ǀQGy`��޵
�4��2{�K�[�6)V����m�Z�Ŕ��
ڛ������yHq�����w��P�ʂ����6��ZS}!�4��g�H�K���o�R^�!�л���9�aý;.�a��j���I��&h���kdՠD[:Wa�l��J���m���s7Ւ1f�@�&"Y���+�g��E'	w/i�Bjʌ{]��~
?�#�<� �B������:kǡe�O�R?���$Wa�'i��N�i����+���4GM�ֹ���UmN�����I�i��͵�-���P ����b��a����pƿ(��A�)�=̒��r1�c�������X�15�4�
��������v��F=��8/j���-Di�EͬE����;�@�#L�԰�RVw�� ��+���yqA��B���z� L
��G��G�7Xo�C���[1ܜ:4�k�Ame͜����7+p�%(���>J*���?#[�#��	�%� 9eg�r�,/�}L����)f�hGH�I�5�<g}�%x�dbw�L�o��#�북��������#�� ��W�֮��K޿�Bɺ=�P!A��檽��~&s]h�p,ʇ�; N&� ���c+�ڲ7����:te��IZW���su���������y[eQ��&V��X�k���%���~5m�ϠB<�P�N��O���Y��Q����cGG�����=�Ӓ����vNu��/[���*���U$�DU;�:� �&��w+1�h�D�f�8�x�$��ؿ���3_^�-[�Bh(�J(���	�F��ip�D��{��R_^,�"�V���ߔ�+����Vd!�R�hu�A-�&��V��4�����㩯;�.M�͡��#0_��?��PB߆������x*�W@��j-H�PdC���B�pg'���|ۭs,��So��r��Z�^�1�:O�u.Ӭ&�2,�_o��\��y�[��O쵯�,�m�'���-��m,����C�:�G>�SU0��f� 
@I)����)��8j�2M[��9'�����Z��=����U�pL�2�r#P ��X8�x��z�92ͻ�0e��&̀/��JZ�Me���U6�͜)����@P�񡛉}ƌ8�r��;��ڧ��8XL�/����
|����UF�x�n�5d��)���Բ��T%�?�0|������8o����J�赝A�_oPɝَ�2��:B���1/O y\g�Pr�f$@i��<�KJ)��e��Re+�~.�۱�(����%���b ���M��ZȪh���Jk�:��@�W�X�lݦ`B36�ȴ�P����u)1���y�) R�_KF��X�v]:�u�MF>>��J�c�omp�v6Kz���A��Q�������9�껽,Ù���c+}��M�;ʭ�/�&���uW	�9�1��Q�*�}]����F���#BJ��\@�Z嘋m���6��Z���U]�4ew�����8��)#��mYR�D)-yC��O]��P�N�Fie/5}>�M��v{���5`�]�����'Z#�L��j����o����c�w�ꛮIK2dX�� +����Ɯ�ۏ��*	3Tl��R� �E��#�Y;j�-�SL�>���"��N�!}>�*�+@�<g��v3 }�M�9���";U�{»C'3ՂrFg��P�L�Gt{�K�d�. �o��QB�O��Ȁ ����J�}p:�t�t���Y.���u�z�'}l�o�f�������W�aD�s���X�D1m���f�0�p+k�.��� �X[��`�y:J2�|��Vj��I�$`��Et��:���#�U��,�gnE"�RD�R����ث1�����Rq-�Ӭb|(��R���/�x�2�� ����s��A�4$���*��:ϏV��Nɽ'�2�H��>="�W4��"�T:�x]�z�،7�T���K��E�dV:��%!���C��C&�m
1}�r�F��<�N7C�qVFZ��R߻ a�C��K�ϱ>�scM� F5P�V���C�*��T�l��JG�-<��pRy ;N��I��^�Tf�:���Ɍ�Z���T��W�4�D�/�seX�:A�������J�,up+e�R2FOwU����.�p�nz����(�m>c�J�[n)v0�u2N�����'�%�7��z���)���1��΋D�d�d�%'��j����J\��J���U��O����=��qj��08h��y+f���;|4�0�	�ľ1�n�C�K��Yƿ��������������Fa&y��i��=�$������#���P�@^m�C�)zްS�5��r�#�!�ڧ�D�]k)�W����� �����T�DR�l�Noty���	**��0b �eq{�R�����;в��Fc��DQ$�}�<�,p{l�l����[*�6�*�J�6b�-���놬�Ĺs�ت|yQ��%Y"R��(-�f݊�<�+Y�s7@6�XM�QX&a���˅K��a�V�y�x�)�x�=�=r��H��J�e*�j{���z���8`R���JS
���}���j�e`����L�����XF	i �Iݶ�m�1`7R�Ax���6��Rޘ��G&���H��Qh��:^�(}�y�
��&'͢ �#ɳ�4<�ċ�2l�� ;Q]�6��˨�)%o�5�	���>zF� �-T��$|-�< ~�nǌ���>\_�҃{\2���
��A�b>W��f�=G�՘��)��w��ԫ��S�)4�s|*2���y��#�wT��/�0�Q���y��d҅��a�o���~����\b����2��ʴ������� ����	>�������YM���N�p<ĕq׮�,@�[�K܀��Ce��$n,����z�����*����xKVGz!]]��YL��j�KT�}�{��'�Bi%��p9S��tެ�OY��8G�����3@(m�X~uy���v�����/eia����Q���E:�?��Ic_��|T�v���@I���\�0|�&S�]B��ڥb,��G�_2��B������(��V<�t��\�+q�6�FW����B�f��QgV�|�#;�,���g:͹�T�%�|� �����Ѩu�JHF�Ĳvn�+n෎-c��*�B�����<�#� �A���q�Ǣ�ō�i���?�\�7��(ý�Ct�r�O�f�,�w�nfX� =	D�vPH���7�l�FC ��X�-+���s�{X�ܤ<�V�f���ص�?�č���
@����U��9e�e\�5�p~P����|j� BF��3A���UiJQ����~��T�&�V�ݔ��i���߂�)�,��Ԣ��6o�PK�1�\9r�
���%	��)T�V�;E��h �v:?�����S�KFh+�C����^��p�-�N�^]�ei�1;kA�N!M(��i��ov
sa�tl�n��#øg�МB�d��F4�q��J�9Q����e�6��W��.��5!��M��3��	6��7����%I'ϡ%�Ĕ�Ğ�q̵�aU���|»��Y�m+;x�#r�k�J�3�����>�	�9{g��&7;���� )�/���Ȯ���`e���P�ly�Y���5϶L{,8n���!�=����VSª��Ü��1)��Q�h��_O[s,�����GJ%�z����a5�����[�s�x*J}�W���$X�k<�d��*������aBB0�yɝ�[�ά�WA���[�6�N�
��H�<�0/'�"S����Ю���s��~[&��/`kh?{.�`8����Y�F�!<�E������lIw����sB����6���θ����U�3�X�D8��i�3�EK˽���3�����!��8�c�m�b���esp�w���q	����f�H��r�u�W<�a���P�ö�:�8H�
Nj� �@���1��+3��'J�"y�-�=G�Ṙ���<b�۰�{"����,o�k�A+!n��gM��=wZ���/uwkY�mA�N�]
�u�jJ�h=k��DOӔP� ��e]�Jv�Y��c�sT+�jY����j(@9��Ύ%����o�ϰ�� ��=i1n�x�л���W�15�|�۫#�w�Jcn�>a}NҺ.�&������|�P�I4�'��u�����.�8
qƼ�w�e<ڹNn�YwWr�p������Y�\�Ӫ�>*�e����U�b{��:Sn?	R�Cy�����@u�]Iŉ���g�H�F�Uˉ�[�c��XDÛ�դ}
��%�]��#.��O�+��ؿ- �ۓ�7������"
.��D��'Pcrq����w{����Ũ�P�'��o ���s���j~��n�L���ѿ�6~!�!�����A����a����f��o��;l�,�2w&08S��qf=�o<{����1��6���s��!�_s5a��*��d� �NN@TPu*�F� ;�˯�g�V6�������f����V��^@7Ի���V��%c��M�Lľn�����w��?U3"���UHP,����Z��i�	Ř����Ij������4g�;μ4P.�"3���~tۺ�)�qMM��N�j���w�`��C���#�em矲�����9����W �c�w0;ő�*�:��j�Cns�c���̗���H��=��Ɵvl�q#Fƫ~_u-�`��� [��`m�^����\���ri2J�|�����k/��[Jg�>ǡ�i�mN�:x���K-hK�o����E��1��M�LxG��x��9�?�G^K�nC��0.�X��5�y��I-�[�g�sj7����pK�n�F!�z���ﺡ�[��g��{=V�`���aeZ)��@+"�bu�R�����gO�������N�WR�8-����+ֱ%�r4\E�ͨ�B�a\��@��y�~�i�Tag�nsb���\�@Sb��=MN��m0�䍓�T2ZcO_�������:W�'i���D>�@h��)�|5 �α/���Y�~�S �����=m6��Vc)^p���,��6�S1��m��<���0�W��2"[K=���8���2���p!�'p�V)�ϬY�S�@:Tm�L����6cc
�LJ������=DI>ca=W2��s��w1!��1�7V��8���#拼F���=V9���:���5�ZzK�p��ȵ'0H3���ِS����HA`
'�̷{ݪ���ZIm�I��dz��ζ ��M��H���k�&����*a�����h��u���@p%2�[��.N�Iw/FB����H3��m1�&��g)Z�w�㭩�2���t�'���;vV<"]�g��w��n��8{%������w�!�w[��̖b��l���M�SK����@Q����L1��������A�4)��������"ȓ�"��*a~ɺ��0;��g��d ���VIy؟%N������1KZ�>g���v�$�NiH'N��:��9���M���?�o$�_��SF��b��n	H�"��=^�3m�	_t��D�5l`�U��+�u�v������t#��޶������14t���I�/���������ĬF�0&%���7�),�)C���j�.kOt��yT2%	��b�׿���v%����w�'�"!x��]p�O���Z�Q)�Sb����s/��d(�����N�z�U�09{�c��$YF�;���'NAbM>z�~8o�Y΋ k$rM���ˍ����/��A�Dt�dR���>s�l�ɼ5S��CЭ��1K<��������y��S$b�~�s|��Hr��)</�^?Xǉ�m��o�A�d6���ʂ��/�Cށ{�i���L圏�-��^���j�|k,|ؓ��@�`&�Mn,��ǲ1�a���j�k�/���-�a���V���b�l��_�C*R�DK$am*�m�c�AQ0�O�'��wx�ѷJ$@	�~�X[����8
z���`�u��@<��T_w�}o�ReK%S�5�JU�8p�a�?0�K�/���Q�|/K
r�F)��n�� �Z&-�+=z����r��c�ɺe��[\�*�r�Ry�|" ���Q�~���`��,
����@	}�>Tv�r�>;L�QI
�^L���`�$S�}i��7\�Z�h��J�m�������M�Ǎ�7.,l��M�"Y�r�q��5Y����\w�y�����h��ё�@�@��X#�W7M<eGR{!*4/��T����BF7oU�8�]���
�.y����0A����"v�Ϗ�����Wou��~j�R�K�ڌ��̀�/y�h�����L/y-m���cl�[���k�7	��0U����!F2-�fXuѬ)�7M*ˇ����qۀZrI�;�Z��#c����K�$ސ���ڇ� �a��3`�B[	��N��Ja�]0��x�1��U`ԭ��Q���j�{�T��(Ya���A��7[���MRr��Y��w�|K��<�k����N��m�"�Pd�*���N�1��yݏ3��N�z���������ᔬ��I���T��f�3�Ef��\�v�� 0݀�2���
n�w���상�b6�xXN,� H���R��,��+c��ڔ|̰3���pQaZ+ֈzXa�@�T�n�U��c��[7e��V�kt{W!�C�)Wm���
�Z�>x�����l�o::d��:�=#��b��ģc�SiN���:HW��v�P�^њC~�|��B�pc�F5{��� i-�<c26�g��b���.E��v!��Wm T��)�zJ���������������S�^�[&D�����ܲ�����д� � �_��7/��P�LW
@^�<�b+�i�p a-��bv�Ho���G�H�N��;̢_�_�ƭf�רAi�t<���� ��z:�i���h�{�<8Y���.R2w�ح?j�◔huf��_Q"Ci�d���w|�k���N1���-ȯ�pQ��1ӝb\s~���=aU�k��kF��A�
�.��I%���30�!�(1��"��Q��-(�0���\[�΁����8�~�M!�9y���/U��%|Yg�P_r������^F�N΁���;�I�o{rF����)��з������W䐉� E�@)WDf�82��~I��$���I���Tp�L�Yt얝�J���p6g�pCVj�9������sߢ�H�	�΅���/���zR�O��~�8�?������-i���v��mjݽ$�2&gK�~�B&0,�kuU��U2��]��h���D�U�gn�_p�����s?}���g�^�os�.��e�1?.����l�:㤺���J����Rb�ʋ)������\��R�J�Ƅ.L��?����ߧ8N��ˀm�c�V��E7��4�;#4ޅ<�g�uzT�/edb�K�-��O5�i��ɐ���r���>��P�Da��	P-�@�M�ޘ��YmÆ�Am�tC� ~�3Q��Q�sE�Ճ��� A[t(���S��'^8�����)���BN⽨{/�ͷD�ߍ�������X�d|,qH��<��@��
}?�\Ւq�B9Q����Z��>�? pT�a�;�뼿�Ί�(qg��$1O,l8V���H�sx���w�?��jg�?��N����.J��6;�*C@M2϶[YԵOJ��W���E&�~̖=���x�fG��/�&x���u���(�%� P�֢�#�'P��$�0Bk^7[&[2E���
x��������� ,���F!��=)���q�r��P��d�|D���Y!�ip�%�i�k`m�ă���%��33aTZ\åA���3?Ud�nh%��uF2�g�y'g�ڎ��VMRLx���N�uVחj�1��m���lJ��ܮ�ߕ��@PC�,�J(����P�G6+1�0��O�>�鷺!���r(�l��Y����C�}e*�ሇ͙�a&�I	���e��٢
P�wz�C8�x����� �0�V��|��� m���!��j�Q.��_I���a�CB�=���F��,�Ϻu�'��v�uH���=��00!�����X�p�P�Ϯ)��΂�*ȁ]yT3;��~�1t9����	��9&{�^�#�^��+I�/���e�"Wc�D���&U5�����_��.b��[���K�wt��u�l�U�
�.\=T69��4����y��sÁ8,^|>�P�S!���/���W�l��tU�������=#��������SjxW[9AQ�+���ɍ²�>��+x���,]�,%���_��]�,�1Yv}`cJBhJ�3F?i�����r���0��N���O44�D���2:Ro�Q�$k��1^8�-e�xBҵs�5FH�� �z���'�Vs_�)3�ᘌ�j'U�R(����ԏ=�P�V�eS��i����a;�c�%ܽD[���n�>X=����B �s��g����RC�/3ߦTJ��S�Vh4�,���<�؋E��J�=�
��D���S���Ͱq�h�t��f��|�M0�65$?t�6�3n~g�t-/dn耖,�BF^�,U���3�#�Yw�)9Yо��a�و
��V��_���~��7��Y�m?U�jr�u�nޜ�c�:2.Y�{3�.a'�L��J~'젅�zz�\��|a6�;��}}�:��%KQ����ڸ�lOjo-�!<S��-���q�*�T�8�2����Fx^#I�u�'5W�0]k����/��rg�r�I͐ڊd��z��G$S��K��l�-��LK�� ;���8����h���P/]��H�5�W�0{�Yy{�v�6RS�?��"H����Z$�	����j3�k�����")�x�y��a�v��ӭ�n]��cn�3t�$����!@g�R4K L��=�m�T'p��UZ���O]n95�Y��@X6�G���hA0#�t'�J5��[�4��`\�,O_۶S��O���~��577/���pI��ԟg���Px�NH*�R�LW��}00���BD/C÷S�a�������#Z��ZS	�A++�E�)�����2��yw),�K
t~�� HC����Sq�'�,�C;KC}�4m��AA���:*�����1
�4��l<��S���*YI\�~
�,T��Kvk�� �K�s<��u!�0��c�{4��V�g�ߒ�Ѣ^�e��̢n�+/X\��-,Cu��)�j�7���z,hW��4�%H����vDtx���;R��\��9����7����z6^�H�asAd���X|�v��\�WG�2]s���y�kvFy�_�L�X���Y>/�C"+����AV�30�TC0���j(yOn\$D̠�"���$�"4	V�#�Q��9(xO�v!#��N�����C�0y�i�9�ބht�T��R�Y����\JPx�z�ش�XNlBKV�5��1���t]��&KIE�u&#9C9�ڞJe<��1n�JB|���� Q��;HVO����P.ة� ܛzv�"a��rYi�nT��.��/)����B�82
���ωN��^�Nw��u��gv�	i�.�%�J�y��}�y��bx�}�.����&d�sf�,z�g����Ԅ�-�u�l6-(m�zi)$f;�7�o?L1�[b��W!F�$C:?�ec����Ɲ}��T9�����v�� -�Yv;
�n�Dd��e�)ۨ��ܥ��� ���҅�q����5�9�9~�ѡA���� V�"v
B��G������t҂�:g��z�=v�s�_w]��,���
�	�� j�:�,j+��E ���^�5�u������v���`�T��%��4ѿd�Sѩp�)�ë��S�N�)���"
`Z�B������<��W�%�ҥ�gQc1!�1��]�q�{K�e�Y��2�� =������9�)v����{�߼LRK�J�C<D%U�����D��[�A9� j��>�8������0�D	��ש��]h4`�k@p��3��������b��� �>*s�AX��X��J�S(}j�|�Y����+{�,�vk�����X��:�1G���0�żL!����rR|�ݵ�YW����oG�u���,Yw��F��p�G�r��>E�j����A����bۓ���E#tb��t5�x7��t"[�^R/��\S���{��:������|�4���;f#�(�]��.8�xMn洛3g�I�����7��QA�u�FP�[�-��~���{�/K�hb�.K�+�y��&�"9N����
SKSq�Kr�y�j�ת�s�K��;{��&d�3��6G�+u��Ry�[�@?o�$��;e��i�\��@37b�R�b��BӅ��4k՚������Y��.��,���[��ɀ���^��C�g��e��ʖ��/�mé�,+�CDk�d��V嘔,b�U5���/Qwzv����/,6����]2۞�c�{V��7F�os�,o,~$�"�����=O_�ff��=.��sl���k��%P��+f2�˵3���F��5b��0{�^t����{K\}k�)"S�bw'�g�$��ە�Y�9�Y�&�
�H�glI��nÄš���R(�ܼ�m'�����H�k�sP�m�J�QSí�d�h���f<C�?��g� �F�*ǂݔ��~�2� �3=kG�9���i�6�(߁mֵ��$Brh�Rd��KH���l�T��	|uז�\�ȀF��h�n�D��=q��h��q�C��:ϓZZ&c�c��]������3�=b���5'B8<yg��;�왝gI�P�G��q�Q�+�9��2�7��#f��E��*��e�MR6DOG�gma~+��?���cH�_)z��g�S��~B&��H��x�C�S����<�\�}��J�A6��Z�z�"U�؂���(ͅ����t�ڣ���S1��ӝh"3�LZ*o�l�Ġn��:���6$�Z���SE� �M�/���wt;�ć������<��E⬥w�7EJ��F3-/�����4��A��t�Կ��7\E���9�A�s(�%���n� s�"g�� ����RI�%�@	�����ߐ���k�Y�O���%
��F�����g���|��{7�6�5V42��������Qi%F�d�Hh*�O�Sֹ���ً{�s�P>)���g$��ܩ82�+����Rsw;����V�&2:*ܶ�`�chE�Q_J�����)��;\^�5�~<����Y@�2f+���b�u&#����X�?�����4Td5f���+��x#^���!Cn�&�?�cA$���q��*erf���|��71�H������ꔺ�nev���	k��[����ρ*ɮ*���eJ���b��_��3���vb�/�p��_`"�7��+���3>N7���8�b��c�Z���	U���Q0�% ����^�9��Z�\�޿� I�`�ۄ�U��ԣ/����h~T�OR��(
��d��Pݾ����V0Vk�d����b�N�~�3Xp]�8a7m?3���-d}�'?�-{�����"�/:i�R��*у�|�)��,cVY,��N����#k���h�/ՕgO���){���LXw_H�dE��90�20���5����>١ǩ�z������Н�B�糨t��˖�I�����nx��g�a�c֨� $�j�׺^l���M���ve��
��V%,�d���*�}�p�D_G����[>m�nj/� �մ]@jm ��c�љ�+�����i�Jw���V���|��xx\��b�G~U�`hr̚a��S�+I��ȀőqNΩis�H�I��&x�*�z�����=Od	��v�?'=&��¨8cM��[$�G~>�K�Aj"nS%0JL�w�@�y2���r���	Z{�a�o�W�7�Ѫ�8�|�����N�r�Z���H�ULmj�X�{�$G�:�k�E�tŅ�-�ڥc]7G� ^'� 6JB��8q&��k������w��4�l*���z�s}���O¶!��r5KP��~����?���1�-=S�u��å'	v�~��(.
1��}w����dPUاj�rR� 8#9"�x�K��0�諴_����)LMC������-);���>��e�@��3=Wkw��Ϯ��h��i%�&g6{�
���'z��g�Dg]��șᅊݻ�xێ���C����)�]�"���SߏT"i­�^L]��TK��UE�K���.�u��Z�J-55�l�Z�3���=�x��u�j~�4����i���\m�� ;>{�C�?�q���{i
-�	p����_"����S&S��v=n��Z\�Nm�MS]vﵹW��F	�>6���̈́4Y�٭K���to�O)�2�]ȡJ*��ҩU�F��綣���۾:�e���7�݁��,��I�U,�'��!?���ߔ֟��sφ��J��>��7���I+(Y�%T����x��V&�}c+�3C׉g��hy�h!��x&��a����gkB���^���,su��s~fV���!�6����h� ���U��T����ɪ�c��~�'T�:�0�o-�\!��&zk��c^�࿭;�Sm���V�A���,�(ߑ�Js֢��
���j�!���5�A�)�U���� �0r�6xփB���}~��o��7#��#Vtl���H���ڨ�T9�{�2}\�U[�}Cpu��)k���Т`�|�h��`���}ngؽ�_�2r�;n��	����/s�q�#�ޞ�oB�K��	�-�.����ֿ�8ǝ��_F�b
��[$�5.L�ǡh\Ï�mԞI�a3 ��R&�س��G�$o��U�����l��u���\�Xc;�*,��i�Ω��m� .�p;�]�y2�3��\�E�2t�m����AowG��=�6���vȝ��`T��?�Yt��"��aʃz���qI9C4�+��mX��%��D��w\�!�ѳ��bܮ�sj�5R�_l�o�G���R���!��u�lJjQx	W(�����UW���	O��Յ�G��FV�#_��_AHV�*�,�Set
`����d�̗=��';�K�K|3=��E�#�Ѫ w�b�D}�)��Y7�5Jη3#A-s�	��q��KεY	���i�߀�����)�"��^�r��c�C�~�i�=��>���w%��&n	���K��+������:�Ls���o�ʣ�P�&�a:��@�B��6�-�k1���i��/z�A�1ل���\Yq'Y�Y����xn�8H��F������\��h�c���"���E�l��CAOt;�|����h��Q-�q�'��=<I���R۔B�G��ޕ��~��S�ֳ˼���_\{����ż��Q�3�P����jΣ$�(BG
`-���T$��~CFKeR4C����gU����{� ��7beXA;���W����6�+O{q$.�-�f��!d!���ѓ-%���m-��ؔ��9��Jg٫��<�0�ʖ �_{;6����x˰�*�����UU��m�7\���Z�
2�,g
M�����%l��i�G0i����[�/�R.�*}p%�J�<���P��+��`يMֈ]�O��_�-}D��
�Z���n^�МC�|<,���~E��� ��Cr��Yo����Z�؇���k�t�Yr�=`
�x<�Q�raǞ]]n<�b��(��|���c�ͪ3��^@;]��������a��r;��A#�GF����õ	Ck�6,������
G��-s ڸ�p��`!�=J��&�sϬ<nD9�;dl��R�A=���Ļ�S>J�bH�����֕��Y�N�kg1f��U@�.t�9ךMɓ�OPR�M�|bl[���H򃭾���c�������d�ʍ��n<��菆	r�y���-	]�~Y��G,���:C��
n'�T4�JIY�\��5���N�n(�2��<�����a��z��.M	�������Adu>��ڷY�S:��V�4	��l�k����s=��_Bv��<�C��B0������5~�'���E�������N��s)��)�2㒑N�+OK��SiMX/ݭ⪅
TCTLeG�DMl$=K 4����9v�RYR�xi��\���46ӓ�m���5�~���i��_I�l7�r��<_���Ea�d7�Աb�s���W3Cu�\�>���I ����}�h
﮶$�٧��4�z�"���4E{SR�s6��}�>j1�Q&�`UsS��+���~�ޮ|�G1nƾ���+���#��S[�)���=`��=4i��æ��V%U�Bp[�-�LF��[������Ji�yƠn;�&�t��@���"����$P����M ��	��3�'�p�4P6?
�ʝi�3���B��C�l"�s7~`��;�Ko���t�O�ժ�RU �!K$N��g��c���HpL!ʦ[�J9C�ia�������!$�F�<(��^�2����T����X0n8����x�����Ǐ�_5�޸�������ͬ��N�N�gv{�=�pZA�����ʞ �u#��}}�v�g���vD�!�%����~[�2��}�X~���P7��(��+�?��J+>x�t�|�s<8���⍏W�T  ���3ˀ|^�>�|�h�D�!_�⟗�����A3z~yb1���>SI!��-"�U��)�Lݤg����س�[���U2 ��a��RJ;`3<
^(}R#F~#N�NX�&��J�.Ӆ������;���jz@��j�g�2��T��Tk�**$Nn�x�j�H��'y ��>[�mA����)�u��dm����G� F��*}���^u�-�GQn��!a=�'?���Vz�@�������̘��� L�et��{A��=	��f��U����*(}ô<0B���}���ڷ����Y�%�x	�nz�N��^��D�Npy�Y'G��:��spq��K::��v������JE�}iQ�%��\#hE	�C17����T��ϡ�@E�����R��C࿨��i����i��m��.����J��T��ԧ�I��n>��f�	�~���H2�Q�h;��nb��K�zg����;2)v�}��n���5ƷH:�l;(]_�H�u���=������qm2҅y-�]�D;�IF��{[
K�ɫb�����x��0�R�#��D��3]�W�M��O�;k���ɱ07؟v�ӺQ��Ү�6��Ba��9�*�g��B�W��i�)o�R�d5`ʀ߽0�����%���$dh<�+�R�f���Lrδ�UX�vkz��p�:0�Y�>5��'ی<S�`��H��&D���O~��,�� p���6�5�T6,R�bOQь)��Kd����7
0♡%��"�`���+�[��U�%+�\=�e�]�%������-D]�w[^��t��ѩ��ft�`gh���nL_�)��֐h+�~'�3��F�r�G
rq�{M.Yb�H��9����[C?���
a�z�����Rj��z������>6�r�f��詄C����9����Э��HqH��)(�I��=���Ьz�N�RB����_��8�=����;�������\�*�+��}GƮ��g�gMݒK�C  �o/�C��>[�j	}��k0�q�I,n��#���YӬ�dk37V����F�u����H�5�q�.g�aGk�P��-�w�hk&p#J���Rt-��? r��*�]��x'�ɨ୧�/��}0Zu��l��̪�g+CAl��	�r�a����0�\�ْ���~ڋ��WhM�}����o��߬�7z��9Y��N�&���pt��Qΐ��,�,�`�e���*E�}}���o$%h��P겎�7���t}�����9O��%���4��H��q���lG�~����{z$*��؛c�0#���/.L�V�]�dV�RN�"BVu����@���4��F���"��x��U|C�%GŪ*�@�7�jcz{C�X���Gy�&�O����{�J;
.���k�b��Jfv-�旊]��h�����%M%뒨�r��,c��.��ɬ@��;���`�6C�i�"��G����ˌ����i�2wn�7�O.��]�3XK�Z��|Esd`�V	\�h��i�w��-V7��6�#���п�
%��zǀ����y/_bȳ�nk�Y�D�����U<\;��Z;I_+������ȖՋY.��"iΤ���[5>q�˭.�k�.U�F�����$�0�I� �� t<�rM��}�A��H��o�`J�-m�B?�����W�Pajײ�G��oU3��0�����&F�,��w\�uƉ'���?UB�7�����:�(����~��_�o�t��������>�w ��8�3�_F�d^���h��:�J�x�Ly7�!���/D�}d�B��Qp�8nÂ���8�cJR���I @G
�Ƣ�j�c�2�o9�lEϜ�?��Kv ��"I�۞	�E���n���D�gc�uǤy��? %Rg-w}ʗ��*��y�l&�.��)P��Ovװ?���S
��*wc몼��lF��>ۂ�m#%#�6O�E�H���	��lײ�����ʶ<�Ղ$]Zڧ��RhL�%�"$y�T����Y��UbH��0��M�7�#���$��f;���gr��H�9���r���t��2bAE<�QW�W ��y�1�`�?�G�����:o{i{��ʾ�p`Id�����<�����F�1{[A_�d\�[(Z6�cM�@Sң�.@��x��%`b+k���Y�s�(�j�y��)۱�����a���ܾE�.�2o��\Yu7�_N	 �^IJ-��j\�aUYMh����o�:z��_�G�G�x#�ҕ�=�Jz}������>6�$x�&�2t8�XEY� ϛq^����d��.R�.23�� ���������h���/�=�+d����D�MwS����0���]�����=Ӣ�aN@���]{�	�j]��+;$K����H��e;��9E_�I��[��5r��",�YZ&퀮���޼F���x��S�_�J~X�7����Ŀ��r�S�L����jd�`S��s��[�.�G0�@��t����Xz�Zp��aV�D���� ��Q��[��-jb&[���S�}���GS�������Q>�?u�b$��*�s��b��J�S�G�m����i�^���m��s�O/������3	�dȁ�����b+>�r0��0d�Q>�KD��-WT{��DT�8(�~vu����0o���k.["0��qo�	Z����_ܟ�v��Y��G��s�۱g+��O���q[�@q�k땰 ����j���a���I�M��<5��I�q��#�h�~Xjm�Ɋ�pq��ci��l���z9lcK�c��� �J��CHv*������hh�(�v�V��i��|m�o&�` ��Cj��c��5���>�_�����dWt�:�FV��
�#8�g!cif�v�:jz0o�<��do��F" ������:;�M���{�s�Q4e��f8t'�ّm�7�V�1�P�|/��32�	����v� gR�.���Vy/�+1�d�/������=$�_���Z���7���m=��P�����Ek�5�^��9V��I���DvQi�,ֳٯ�ut�GS�mS,UD%�*9d~��� �e�| �Hj��N�o0!�o�j0��/WQ�|��GzO���L�ֺ�7��˶���S����ԙ���M��'Ԩ�Rl�w�Fˀ\*K��R]}b�wp�@&�I���>��K~j��J
���\�Ut����ů�mT�y������p��WMg�uZ�/����2�d��y�
��_DZ">��q�/����K�le��0�*܆E]��QP N��j��0��������rH:�LA�d��ҋeޜ�E�`u���aV��Ŕ�7l�����
�n�9�&rx�4_cH��=nСռ�������7��7�WiT椂�V��:��O�������� h��*��-�'���+�3��;���.9��"�6��{�==�*KD���~�U��k9��H�Rq��f��*�dIլq7�m�D2��Pܐ_P�dب�ܑ)�|QvwC���w���2b�[���Z%�(KJ.�����V1�(4�^rXu�@�W@���� NZ��Ȩ@����>v|��\T��V#�<CJ�5�sA��`G$���#�7�B�#]�e?F�hATH*x˙�1
��'�Pb�!扸!� �z�r�?�m�<<;H˯.����2�?���sύ�jH�5��-Ǧ����"�K ��\�<��ds}b�=�&t|"*h�k����+X���`��S���f\�W�@�>]�x��a��E~8P4��' X���;3v?.�[�0�����DsW�� j�sl���:4cυ=-�G��;c?)f�r:A����?jrV��$���w�����`���L=9`܄每��Yj�,�4*X5��D�	�耊��b~��r�Zf�kP�韠c�*�p0��+e��������7�9��|��6q�#ff����¶�b��U�-��YUߩY� �ׇ�´�%,&��֣uZe�? ɚ��Q���a��0�'�m,�Ă�G:��]8?1��F��"+ta2W�#�֑��+�ޏ8��6����#���'C��=��㳕Q�UoV��r^��x����(ؐ���?[0���6�}�4aw��0 ��-�O��V�i���T��sO�JL�M"�̣G����PbB�_�ĈMP�hj]4�,�}JȐ�����>AU���"���Օ�y&4��hl��r��:T.� Ÿ�e��B��}�>�w^�^�U��8J��X��nh�4�msq�G!�,�?���u"VS���OT����zF;^O�~L�}��!�Y��W��g����%%`��Ŧ=������^�0���I��zž��<V2!�\�o,P&hc�}p#��5x��A{C7��$���d"�P川�b�+��[��ή�$�ͳ&	�y.s#arհ2ͬFSꇦ�4�H�M{��u|���\�
e5G�y!{l�Oۢ��d����5
~����x���xnMj����/�W>�1/�_��%���F��OH/	�l���`A�� 9�H����z\X���u"T,
ԫp�X8Q�;��J}?Cѷ��P�}e�+-�6sA��_�C�<�J|�k�MB�py@��xԚ�f��ʮ �O
d���*�N��.��jKLf���b��G���Ayk�5O�:j�-B��8�S�udNa�b���m:,���m �v��u���G��ޕ���be4�XK�K�L7|���a�(�fDC��Taq#�R�
�mvU���}���OUK!���؍E�*�xZl� ��N�5En�����'�%�ڈ#C~sC��N�p(�{g��	{��T�D��NY���m{�2��Q��)��.�s	��=��s4���=���q�r]�)�Ar�	s� �oZ��_��@�P�,�zb$m���lSl
�aӖ��}㯸�t�E�M���ǫ����^[��F6=/V*������f0���3�N�apcA�����]~N1�ؼawDN����?֚!�kK��"�RB�����s�o��y�N(��#��0ĵ�8�bn֞�R�� I}~j���>��3L�^d]O=��
���K��p~v®�3.�ojC��	�ɧ�>�,&Z���x�>��@>՝U���=�O�a�_%g\4�������1�,��a���\���ٛ���Q$39K*������mKG����R���ik��(&�T��O�)h��EST���x�����]	���ꔫ��T��6l��P��iv� -��G�v���{w��� nƠ��>�;R)�8dv�7�½? ���/11�~����4?C�B�08iV�s�k���'�Ӄ�d�A��$ب� S�o��I��[��XW�h��Zpb.����RQj3���<�ȭ� ЍpW�v�ٲ*x��_���/��0{Yz�o<v�Oi��p�5�=�"���BI�0��Q���!�;rf�D0IE�w�Q�Ti�+��ӥ�R3#�t��I��������	h���B��Ł���_h���?*zp����rǧr����"���],�������(<�,v���|ѦB��8�]�sc��Ū���@�Կ���(eks�
wW����O�|u��N�e|o�I��|/<�J:��zJN��X��*����!Q���y�w"Ym��gH(��-�y�� OX>��^��z���c�Z:��j�)d��N�
���L�xm�%L*{"��:}CqJ��	�]P���9 /jny3K9Hʏ�%����rt��3�~ԅ�9ez��o�?�6����OOR�@DA�OŞ�BP"]�k��$~uę���"L��ܐ2���cY�y_aY.�.\=��8�1%�[�,�e�\?�r�6��I����uKn��4c�4�!M�W��_E��ǳ5^�Fᒎ���q��:�yƟ�9�aY�
���
��f����E����V<�X4�'����铟:(2u:#G�֖ʵy ��y��?%��.hpmLʼ\'\y���4j)*�r ��p�1=>��>ft�N�����'��;[�]����~����g��}���L��61��V�:{�<{>��i����]�t�0��kG�|�C�Q�v|�֔͊�U��C1(`�@/�t>\"t=�3��.���ٕ��`�#���j��G���{}��k	�Z��hFM���6���'�K��(���y^Ze��H�MEt��j�Q�C��?�L���2�.6bZG����2����pw괁�RV̘gjE��Q#϶�'?S�[M����J/w	}�J:W?M�m�t�=W�?_FMq~�&?3!�W<�*�kO��bq��A��=k�#	a����8�X���iѫ����������?�����|V]�W��Vw/�z0ߡY�����E��mh�a����|����X�Q���BK![�|�k>�lԉ{d����"�(*��3�8˾ȗ�.U�»�l������֛V&@��*t�M%o��
����i�`��7Z����I��L
��`v�ȃ,��&[u��w��l����Ϟ6$|y�v"��Z���=��	�
�]h���������o�f#��󲺕I�B$�K1��I;F['z�:r���duMZA�I�R��-����L	����!HND0�i����jИF����5�����{G]z;��7�qdڪT�4���0�Є��Uu
N4=d98�Z�� As��wc ���x��@�l�ϱ�|cA.Dx*�`�����Y��3F�7�u�`�H*���uP%�w�w^�<#��{�p�政ONQX�`���pt�u���["�h��i!�R���=xwP�ً�k=�	P���i$ϋ������#̯n*�s�+��r�ѳY?�x�h�:�:�>�]��M��3F�"$v���軚�p�+ʮX^M��A&�4*�+�)$�bV�6�u��O	��oF_P���m����,�t��R�f�q]t��"�%�0��u֢q���L,3 Q$�'�ڈ���H,�u������hv���D���^����Brٰ���O�nY��U/�1s�pZs?|�_?m��&Ѥ��K�Svsآ���n�>����+�;�[�?bt�δ��W��~��N��(R~6� �Iv%�I�!�k7�j��f���f�����n&4Sk�����q�HpC����b�p�SJ�ޣ�ɶ
j�"%l3�D|����]_L ��g��u5��)�Yd_��c�uw�C�*�vv�ǽ����I��A.�>�@�x����v��E��2z,X���~3�E�)�RkΤ�8���U���xf\/W�?��s?�=�t^����H�ϓ���R�7�o��? 1a�v�;�c��=����A~,�?�3ҡD�/�)( p>��,��GKׂ.m����3����J��F4� ��]a<�SC�`�=A]�3��B�D#�[Sߐo<;*"z;��Y�����l	�#�Ыl)ʽ�*�x�5���i��{g/
�bs[Q}����,c?'b�<}�y~��#N�o��%�/�!$�{�Uu}4�4QR���h���#hZi���4._z̦�;��'��c�J�an�J�r�yw���1���R�7�N�DS� �E�Zݙ�'4o�`�N#�%;×o]NJ��[p�/X�x߸zk�oY���PKF�Wqk�Y�Ę�97r�5 ����$��tH3X�~�P���-�D0�V�?�|No�d�n��?�s9�?�^��g"�\�YR��HyE��=Z���]�P'P���ċ��^�ҳ�r�\��{�=`?��O(`�BT ����`+���<8��š�o����"�B"�A��Y�螐�K䄀��3vZ%��̟��������Y�l�&Ӡy�(�eq�-Pbբ��íL��_�P�����l�����v�w��>v����e.U��'�����"Q��a���Z�GcP��V�*Q���6C��P�=n}���gF5ׂ�LJw]�GE(��/�<�����？����1@����:)�q�;`{2����hE>���o�bO��𡢹�'B�橋-�r�����|��_�c��h�nj8)�6�E���K��q'fP;��,I�E��n,��A�A��H��~�vv`I��2̣�D!x�]lw��ƺ��
a��}قW�Uژ����Z#u���H��~�#&�5�5�o��mϲ��;K���ܣ8��4@��m����w�����lpV�G8�"K��&���i[���B!����ӊ�Ӆ����MOz'w��7� �M��nf.������H��r\�@����+�D�Լq�#��i�;D�f�9M�u9���UD�C�'�~��)�>��d=�b
+�ƯC�B
�|«�����I.7��&\B&���9��,Ht��o�C��o���Xaf���k�N�_&�nM�i��
�/S���FxF�!'��%�o7���d`��/ 3�ګ\Lݿ�&G	��*��ߚEt݋H������K,��?�<��J\�F����Y��FEXk/k�=��$�$�o3�m�NI/�|?�-ܥ�啀�e��Sb���q����B^�I�y�p����Lt������46�k3��NU-�˕5��m1�,F��>_�N�z5kB�|mҔBb�.�d��M�@߅�p��x�����;��\�k��n��¸gh�d��TS����!��"KE	���yW����?�yi+�5JU�/��#�X�a���w�;G8+X�no����+⹷�����~t�,8�i�`%�+��^Y2��8�!��Fw��vϭ�E=4~���,�[?��X��ؤ��8W�z$N-��Tu�.��jB3��?�LV�޴$�k���N���3i�~�ܭ����ޣ�%���#oV�Mdt43E����<'��#��FU}		c_�cT�2Iyr ����|{3��X�����6o����պ|ۇ�q�a]C.Ӿ�������7q!�5��l�����4�Z�%`|���_.~.���j��ţ�g�EE�,u�'Ga�=�u�	�B����\��b��֭ɦ�αZP} ކe��]r��j���Mn����}M@���#�UhY���}:�]�k��̦�/�͡m�x�b��H�YXe��X=�--�_u���3pO��a� د������Ǜ2�_P�*�f�ϡ���s�scv,�:�T'��MkJ��Ok{ �?ȑ@��p�[�����f�v�>?5	z��i�ZV�,Y�������Өl�#$��{�;�T�p��SƻZ>����F�䧯�A�{3�>�U��������m��?������5�(E�u�CO�<���/�T0�����0��ۋ�4BW:m��GI��*Z��00(���gn����r�a ����fk��j=}���9+dd����ǴnI��zu�,�{(Ӵ�ϊW��z4;6�t,dH�.�>H�1���j:�{ �CМ�]s�e]�`�
�X�Jl]1���@0Wb�'W&ֺ����Zպ��(Hqf������ۄ���bU���ީ��)Db��C�~7u���/Mj�ì���OaDY�K�(��߅5C��,5뚾���v}��m�Z8�瞆 b�� MO�c���1������1���ǰPEV<��@�Y(ae�D�4C�aX�p�M�H�X�����\EH_�~�w�!R����^����bo��£P+�$wy��� �	��AC�]ļ�P����*)ᔴ�>0_a���`;�Cp �~�nmP%�;^�x�Y�u���{�T����]k-�8����:8G��_Z�KSҒ
!�0���v/���&�u}�X-�Z��o~��5�wn^ �3��q+mߪ!�;S��>t���%�OԪ�My:���e�(e�.L��ȸ�M�V�ɲ���M$�4��ώZN��ȓ�_|O_#q�#S,Iq�K���݉&�D��0������`iZ�!���=	�8�����r�V��d�N��Hc��B!o"=�[Hl̩��_]C�*�X0��Lh]*W�}�����p�b�Ir6z�y���wzY"��G#�$�~��B��vy#��^}��|/W	=$�5�-Uѡ�;W���������pP>�cr�.���J_aX�\�_�2��Dn��u8�m?�6i�YAU���o1K�ےK�J�h��V���_��c�7��*4���%��*�j��l���
�-�'ɼ�I��3��g���u;�=���ۑ�"���q�9xT�y�\��UIͰ>��?�D��L�P��}�Z������ҍ;�߯�ux�;�ǻ�vSc��Q���u]��32��*ס{����t��M����N�t���>���v���K��Z�$_�L���� ��l��|q'd�ԙ�{�t��'�xBx`����.W�Z��匮4���$��:����+��]�si���Iz !G�ʆ74��8��n��l_AEQ��̤�L�컣0�]z�K"(��{P�e�Ѝ��9D�J.�@q��<G�Eh�2����$o��6�|�‵����%Mh��w���Ñw/�fS!� �Cb�MN��Pf�\���c��\�������nԄ�_����I�4\q
��L
��/i�쁾 �|k��lr��O%C�x�\[lr+RvK���8�+1�^��/M�\<�$S��dڂ�G�h��8��{��O�s�����W}2�,Y���<��OB��G������h.0{����b<=t�m��M`��Ԋͥ���>a���`4Kײ^ꍤY���&N���t*�^��nWܜ+^�f
��w-�	j�
}�F"�[�j^/GBzX�M�Y}@ç�+���Y�9y�`N�iˠ�㽥ش,��8nG����6f�_��$Rbksnz_�h�(���{�l�t�<8��0��.d�>X��"�an.I��b
K���TC���Y�����D��e�?�n����੾�:z�(Ҿ�_��I�=�!�ő�5�`�1%ç�(@WيW��b�)ZX�l���c�4�M]���i���zG��E��ם5���2ƃx"��>%���Ύ�@©/|b>�E�Ũ�H��ˌ�!㒭![,]t0��CD��WhĽ�(��8�y��㊩�a��ٖ���`���Od�Ɩ�s�+T�t|� �<��.)h��l�]�jl�O��.�o����H��K�	�Y�������!q��e�����DZﮚ����7�X��|t����;���$�Ԅ/p��fo�i��/��BU�̄��0Z#mkߟ�u�6=��Iu�"�+y���X	F���rCx^����N�g�W1?����w��lL���\K�:�MU��x;�2s�<}Ų��g,����*�U�\��M�>%�ͨ�(���nFS8�/.|��T�J�7WA���{��jK/�B�x��!�~�5_�q-�4d85M9`�xN���܇Mbż��a�O���'!�M����q�;�>�+pd����P�'�0�"NЩ�Սu�L�GI����k@N�ev�ϔ.������+�F�a��4�Z�
���bq�H�2�-Z�@�F%���D"�b
�ZJ.NQ�,��$�g�b�a=� ���m�*�3kϢ���æ%�^Kw�y���.�뉶�eux�{X���Bb��|�1nkE�V��?qdE (�ި45f
o������)]���P���{/b���4'�0	b@��};|b ����@�;�ayJ"㌃�z�&��>�&<b�N˓n�)�Z���h�$"���=�3���ʑmA�}��1O_��z�"''c����XhS�W��Y����8�H����w>ICR��v� ���2�|��Bi���^����83���l`��oY<:�5�Ӧ��Ǘ!ʚ��Hu�E��	��h(=bw�Ԝ�ލ�r 0 ��;���\
mU�iO
{�@r:>���6jt�z�0�xWc<��B��"��~f�D��G�D��!Crr��+}�����[a��	�i���("��d_�b�V�w	�s��h�����0������#aa�K���c�Y%P��C����K�v���K��;6O��
����ϡy?K���5謴/l�1���h�u�/�Fhǖǝ�o�{沈g����|��[?�� ~ھ8� ���/�Tj���?[%��e��i�G,�C[�b�{��L�=j�2ߔ�pL<�!�r�ؔ;6���1�� 'xU��V/Óϗ������3��Q��l��3|�����'��ͥ.��B�D���	_�6����#@�E�}A7 ��s�٢t]��h�*���c/c�a>�<��|`n<�0���_՝3�a��J�HVB=���l��*���s�;>��!��� T{a�:���6�$X�'����V��[ } �C����|2)�#�W���b�x��A��ɩrk�B�աhn�Q��1���J�^��`�%)vR��r���E��yH붐�[~E�9����91�Z�ww�G�3����U;��	�������o��{��V늴� ��-������L�'���E�,��r�k� ���*�\'2eÝ�5��p�Yc�J�u0�	���s�u��m�5�G���B��+V��5�������v�3�M�3���j�u���
����E��/��%U�&c��ڴ�Oѓ������hf%�^	�� �3�3Aƪ�mq,��B�6�3��L�����_�����A�"ۏU�׉5G[���^O'_)Z�6�$�\�.�؇�qRC^����e�2W#�����G�aKe=3���^��ܨ����W�Ky�78Ց��{v��l�J�}+W^��������B>�Cq�soA!��֔���k�5�4	]�J���pV�=
n����s4���y�:K�]�v0�j�2�Fv%gM�z���s���-+S� uLA.�ɸ�q����c2������֤� �צ�Z����x�|rQ�%4
dI��u8����ٔ��hU�,f5��_��a=��n-OF�����y�4�p^{�;E\��i rJW5��{��l��Z�!�o�N�j���h���hö�������Umh�
�V��"��n�Vo��Z�܄��Wu}��W����$Ø�N�D�en���f8�O�"�]�Y�b��C
�|&��߇�����Z�҉UuW��>ք|��x�ݓ�,�jo�b�F�8��Q�>Se����ly�;	5�oƯ]�Eb>�xf}���k���+�����ʓ���i)�-�/���E��^«��U��7rU�9@I=�Q��v!>�U�	i��(���Y����SZ��9$��p�C� !� S�a_oC¨n���8�9�p�C�׌�F�,��#3a��{{8;��3�fe�6X`A��/���~�w|Cʹ�3f1�-~���Jp� Hjo��:�r�p�)o�u3���ܒ�el!~�}�^��������pҢ�	{@�|K(�,쏐��cj�8�����L�W���哦C�$`d���@a�T��._�1�K���>���E�uBfA��J_Dd��3 ����#��)V�[���<}� V��"x�k�=w�v�汸�*x$��YLً_��к'?�f�-3u Ñ�4�E���gE:X&S��+�i�^��*K�G��yj��Y׫\�+s����~�d��#��U���chO	ՄX���[�M�.�9��D���OM38�c9�L�vhI��LyK,�qk��
�г,��e#�q����om�ET�)J��Fjtk|����� �W��I�� ��tY�὏H�+.[:$>�>�,��TL4��7�J�?���Ԉ`�O��2 ��vm�J�u�1��9�A�X�w/��K����Z
��	[�}ή~T0ז^T��K8��g�/DeS	g�$e��K�����5���\�$ZՒ*����9v�+m��l* ��#���������'o�u(e���=�K�l�^��i��ǜ[:t�y���]~��?�Y�L���y�\���7�t�֕p􊉐{ �<0��yy�����Ra�6]������H�p;%���S����f�Ϯ�){������`�đB�I�	��u��P�Z+ �n�b�1�����?xǿ��Q\qv�d�d)O0�#8����Y�{#,�,$�����V	Y&�d��د����i�T�Tx %���@H_���[�J�u#��:&��#�a{�Ũ�;2K;��rjU��Hk/1k)I���&���u�J׊�9�M�Ѫ���6�"JZ��<}�W����O��ĩ�x�ߧQH�N�\vw�1�E(/H���lt��yʼ�����Z�)<g�r=�{/����WG씎�]���a�h	��3ayX>��4��`+���pl,twͩ� �L�?�J ��lo_$�ͪ����C���A>"O�O� �Q2DiO�S����IR1���7q���j�	_fs|�2����G��b��0����U�a !CU/+��Hu�^� �,i�bYjq;I��~��K/9�<�[�� ��3Ym[s@���Ȅ[�rn�)P�w�Z7���~|�	�������@w���zr^ ���e#�^����|��my� ^Z)#��6�]�9�itW�8ȁRt����#�Xji������Mb!{L��Wq�"��է�/-���n��,wJ�c]G���O!8�dK�,eʤ�K?��蛙Y�
��~]6f<�,x�L�	��x����-�]��c������찪g̚��v߶n�"4�F,o	��Q��P�s";��4��d�5,��]5J�]��$�������JB9��tY��Sv�mM��n�.��+���r��9��w��G{U�\�P��Cw\��$n���[����m �|��=ŉ��=��=]�	t������J��r�iD���� � ��2W�j�akEkq�B)�����LZD�rRc���3��62��Aw���(�`�#�FW��4�Ѣ�f��+O��Z΃zyP�\uą��KH����)ބ�����!�Sܬ�t�Y"�@��������K�	IX��b(oN.�v��P)��Ûd��V�P{��&)�M3��EJTf��n��>a�eͽȼr�)\��*�E�H.��IOV����uZ�%�%M�r�i}���a��'�|�>�Dy�3W����Y���h����®�C#��y�{�+�^7|�}���b����t��{�=�.3RkJ�|�:�112�D߂0��x��}b��S��'���q�*0�|[!�ƣe{@���.r�('q(8��Z���)�^B���5�yx+Qg�jU��Q���.���z>Ӛ�+��V�Ф����D��l�B+1R�[��3�vt�6�Iȕ�����&��h72�t�|���.o���Q(/�"Y0�9ntb����B�����I�Νȁˡ�was x�c�c��fx�dپ�B���͝{�rXo���_������.˒5�}�i��Ir3f����n ӈ$L��a��Q��Ӿ����^�q֍�~?@w�-3��*�hX*�	��f��mǊm�0��*���y,������>��Ac�ӂK���S�EzP��V6nmN��Z��Q6=:{�R��m��4w�O'��uH"��R��$-�=C+G���;o�����ac����ĺ�0�x8+m�����qoru�tj���)���9��}wX�`������W��L%�ks����x����-�b+�v3��+��I��k����p��+�����:' fٌ|�)G7��"�1����}Nܱqe��-?���˘���8��Lԁ�u`��r����
	 `r5 ���рɲ��<��2�Դ��֝ͦ}�"�!d����T���sP?H2/�8"�l�'d�|��-�ޯm��]�8�\�֑� %�Zx]�l^��r�r��s�J��r�U��HM�<C���6�O��~C���]���p�r_��MD�����j��j�
�����{��=j}�
 �Dd��M�����1xb�tX��q$��	�t�r�M٤j���6��Zi�.�%�S��H8s:����=T+�W�smȫ�K��'n��,z�L�(�V�s5���!L5$� V8ֱY|��X8�o
�)vX���|����ł�Eh�/?be��I��}`z�s��yk���9�%�bGת��suZ��^����e�66�%�R��f�����S��1Ʀr밓mo:wF�V����旁��b&�H>���)>��AH�H�m�:�w���̽_oA~Y/��+�S@�ȁL�R�n��kx"��iX�4����A�`n����B��~�_�v���k���Ud�� �d�lEc���xo/�C���M�X�H�Z�$2J˨���-%��h���j~d��>�9$�)�C5>"��}��o����X`�d�m+hR࿇��cF�5��/�8]D@����bD�Ѿ��I8d�는��!|��,�}� ��a�o!s!ZKC�Z�\��)��ֺ�dٺ���q��iֺ�l��&��PB�:�`��v�t��}5$V:"έP��P�e�ȴ��'���d�K���p�v��H ݘP�ް�Q3)�@Y�_�q)�����s�w�}��aƵ>���X2!I2�-~�+p��O��p�En���p�E�Zf��"b�{��+��*�#jAn�j��+E���5�P��ppJ�߈7�߄�לj��G��eB�D8���wB�D�U�߸g� �I*	D��%_�	fv9��=I�7�tJ��>c�E��nړ���f�݅�t4ܚ���>��:��E�����}������A�����P϶����m3]O�1���K��(7y�t I��Q�ҵ��= ��U�
�Qa��#ْ�	������U��Ae��!ʻ��q%�@Ŷ��N^c����8A��%J�m���ybKA�9�1�w�e���T�(�*�R�� �������#���|_IQ>nx�����8�+��ܙo�a���R��wu�>r��1����`�Ff�)4�o�w ��<��v+խ=*W~��oOZ:� ��dlK�٧8-' �Ҟi��[�ry,d�/H�ĩ�ʽ�dA�Ȳ��[2�W&eY� '�2*~do2`s2x%юk90�ή�n�n��@HE/��8�2�%��8�qW"qm�t�@��7����(�\�a�ySH�n�ً��L�����ha`zk �e�ꞡ��~6�<?YY�U*��!������+�<W�Ce,!a�٠�y��J��I����F=@Q�c;�󅸑��q�N�w���$����WJǮ�G@Ѕ����6���
��6�qD�n�K���C�2'�g�7�(TJ�:\�${I:�$cP"�������-�N�O�$�F��it}(��^��*�h��DHe�)�����(�i�@���?aKN�Q��P�t��6�i��[0�:Y��f㼫7�p�Y*�~�Q+A��f���RJDqNz�˿���G���VQ�o��KGt
v�
���T���N|O}�T{�P��9*<#@8���::��Ĭ
�P�����|�_��q9m��,���)a�ut�22B����ߧ^� ��|�&�aˌI�;���(����D��9��V���`�e�4�>���"Ϊ�4�ST�^CUZ�6L�<%lUe�b{̂Vdր4�L��Z�-Tb�:zvR�+nМOmv��ۏI�K��F<�To�O���|C���h�|�wߖ�}0it;v\J�29�)���+w���3l�11P8I��b���7��A;��)c!�ۿ�jBl�~c����ӂ�I¶"�z���4|�xD'6y~5f�iy�@����ލ��J慡Yߜ�'��	�{x �d*��
��F��� Q�.$�雏UÔQ �T�"�(����"�
�-p�dI��,(06�Pw�h��]9K��إ�$9�c ��g� ��W�ƴo Y��w�+f�o��Ic!������j��l�B ��V�����W�
��V��h�?�o�����p�� �a���(�n��]�i�1R����*伻,�Q#ej3~_H�'lP�E���$��V�]	�mWͼ����
��	�������^	-2�	���_d84kh��z����c�E-�;aa�c�[xC"hJ�$��Xq���7y���=˟ �+�d0�Ͻ�(F��2z�*a�I-`��)���n�Ð�~��� ���%��⇈Ԫw_�|���^�Wϓ^C�!�F�Gs�f	��U��@�B3��D�l)��s�dg8q=.qKZ+�T%�E�X��T�*�Hǐx�Z�fg+W��|mH�(\E��6`�����q8YV�y�t�<Ҭ��nV8�2����=�I��D"�ԫ�H�i�$���6�t���9s�u���Eu7Hub�s4(s�.!sփ���� �ŋA}��?7����裇Z&�LrU�B��|��� H�c�&lu���Oâ��Ӄ=)��,A��,md�5 ����#ci?^	��H��x�^h�=^�V�S��zD-C/�������R��/{"S�0����V��d����M���9y_Hu_��X��Z�l3H#����ڹ��jG(��6ͩ�<"#�-���>�YR]}����]Y��)t�FǓ۞�hR����$���k����ď�dx�_G�B֔	�����ދ񸚲��r
��U	Y��z��4��r�^�4��N}��Z	H_�0����qU��X����� ����b~�E�^5�ԁ�k�%]�^E�&�W;/')7\�g�1��kܒ0�@容vJ��*�l�ͱ�MpW���>�|�=T�b_����.���D<���HW�$�9#�!:�,� �z�O2,��ީͷ���O�!��;�;�����2@da�Wb!��p#(���>a���������Qa5�8��]H�W���A!���6�<��n��U�lS�UW�5���
Z�ޟ�Q�z8�
�P;���cU���X�K/�m�f<dw`4�k������T��4�E�����y+x��ٻ���6(��-���y�(���m- ,�1�ήb�ޛ��O	�VGC�U�t;���;L���v�&,�K�ա?(6����>
;
�@E���#Z{p� �թ�6�ܷ���7Ռ�e��X�G�8ܩ ��b�DD�.?��eqY�����<r�І��� ��U���zCB�x�J����G9�p0��d�;�d�
��s�V�����Z���K�D�����U�/_izsb����k��G�b�t������9Wb� aZ�,��̴ԟ�~G���Gz5�g�i�6p@���B�J�=�> %-Zm�x�z'�Ġ���<��STS�m'���z�W���{�|r�ˠ��F����~7��&�!��NGI=6/U����X�q)�n�ǚDw���M�C����FG�*FV���HY~$^b�G4����.ڜs:����O�����
���֛3��p�]�L�hz}�n�P��=j���e-Ӎ�i�*L��L2@t4�:���ǭ�wqbnh��Or�uR}�e&rԅ�>��]L��cW6�sY�����!&�[��HH��7'�8�@CIm�S��Dؼ��.MV: ��N-��-N��Q�Îzx�F�q!F-��Y~�uT��	(*W8'!q������.��!��ܐ����t(j~\����>4	Sbv���{����&��d@t%O��[�u�	��S��N`����1V���tNj�*��Y��}m�+��-@��u6B�eP̴q���=٘(2�½#�[�i��9�lx���)�!.�3v�9�{���?d%�-pvp�T*�G�S�z����&q��
��1�K���ٝC��E��� ��r��v�X�c�<�9:�f�>X��쑮6�Ո�߱�N���2�f�I[��y�W&�Q1��b+��9�rn���L�1��S�tٯ��)�"`�ZTønқ#l�;`�r���p ����t(o�f �k0�َ�|S�h��iɴ��.��1���KI٭�ad�!>+"DMWu�6X��a6ݡ�.H7�N���wo�^Ŝ�����0C`�$b�;�ܨ���$*��7w�t/V�U��<;����rX5��󪐫���
]�1-ޮ�`��.��3���ªt��\v��;;�j�Ա��h��j�
�4t�(c�����Z:��+Rc�f��\85������;��=}K�O�Zl6�I��IX�z��qІ��*��LT@�~\�s�62u�i7���� ��t}��;����K6�j}�Q_\�,@�AyGS]�ݍK乁��~؆.�5�tk�<)LCtYI�&'�^Α������>��İv@�ӯ�ҋ���\� eE vHu�Y�M�����&�F��n�4�KÖ>FL��w������Qn�s�-w��9�\hh���_5漆�Ja_3o���˅�"���M.���Ց�T��q���F�eTa�~8��*��	
<R�=�ڷ�!7N^s�����@�
W3���8�"�����.�
fQ���b3$>b�hҜ�"���:#8� S�@D�j�\;T����)[ ?�9��y�U1	�E�J/�̅N� ��du�_�
�hn�ӎM�/.��!���`������|z��V�`�ѓ�����Eҁ
ozM�@x�f	t�nO$�Ds7���~�W��������eq܈-�=�˰��M����������%�-�mu!�nRV��J-�U�Jy{a��/w��iZ�V��@�*ѳǹ��{7��`)ou��ghCC�ʿ���C�[Q�`������NUٴ����ȋE�o[��/�Io�E����&@d��Ѐ09P����ȕ�:�Z�5�s.�X<.v����u 7ۉ�5ُ5:7]=/�(�l����^miT&���\�{��t�Ar��:�}�2����=i�ӽZ���L��E�� l�%�Ah_td�N@M�~��2ƛ��NPB$[������~���'ow��A6�Ce�k����t�Km���m���Џ�X8^/�=�n"�`9��-aZ謃��b�{=E-���n�Q�[��h��5'1��1$5�\�q%|��3��>|��c��)U9+�r�D)�9��1��<����n��s�4���c�B�JC�掔x���!��Lh= 9o霴o�Ԩ��5ք�`��a(��>����/�w�ea�ps[�M�$��D�6%\Xz���J"�RK�dhţ����E(�fѴ�@2��_fÓ������b��!@ ;�ب�����n�Csk^&Uw���s�3K��U-�Lw����4���h~��1[#	|�;��L���s*��ׇ���g�ǃ<D��W���ĸ)8���eR�;��^�9�ƞ���B��]�2pvǼ?j-:@���(��#��m�Vc�W��|����1S��*�Y�<:�&�$@��m.TcP��b�u&C_�UD�~Gg���"��&�����^Av}T0������s|�Q]@תC���9(O�8z��u�����m{ص3p^��TX~ ��HI�rK���v���ȄV���i���z���G�<�}#"ZϏ���2<\"�ct��Q�I'��wc���cB�4l�p�L�`���9U.G9�yilz�7 �g�'݇�0�1F ��":���F��\1[�/��4C1x���[�?*"���/[�/�ǜ�*����jOE�&� n��}�-'fIE���ۤ��� ��q���� ����M��LNx{T�;<W{M�`T2v���E(+��hK m��V�^���R��$�-Ƿ=�tBe��	�0/ZBK��u��?��p�.c-C��"��s�t�A$2ȝ)����g��,s����6�׊/����m��T�j5�H�L�
�_q�>F7�:1�=V/�ev'��d�t��=%bT��i4�O��q�X4�h{/hI<��]��]q���ؓ�
�>"8l��!q ���K�����[�n*��y϶�ǿ��