��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$����X��2_=Q����6��R& �e޲���(b�A��x�q��z6���E��f��-����K7���΢cmY��[i�b�\�e���Ρ�A�dt���p������F'~�����FH+�V^�y��t��{)D�|p��d��|/yQ2.J�=Ea_(v��ߟ���#X�/�\XU�����2�b��m3���FC�y��u���*"��l\�!?�f�~����G�H�Ы�!r�qe4}�m¬�-����(��?���.�=�"���B�O�OW���f�o�"M�P��9�
U��"�1�(��)�ma/�/�z��,�:�<Ѿ���t�����{��Ӓ}h�;%=��qz�E�� þ=<�;����(�7{}ط��NR��ڪ&��.��=�)j�PqZ)'_��c}�?�pi�\(�m���	}��rp^q�OiSr@9�Lc�^8���U���3NMJOd삪' )l����N1s�2j�C#�)�@3�-���D�����\m�V�'S�l3܍�f,���z!trW��Fⱸ2�g�bc�;(��)�n,5������1�c��!�]�Ĭ�X���Ni� ��H����;2��cũ?���.�7��v�YZ@�d�����Oak�>=�D�bS7��7 �'P��c����U������u�@gC�a��09���֐�S�o�j�BA�id���j3��H�F��+P�}v|̘Q�t��g�:Ж�EBY|�����u�I�p+��iZz}m	��ǟ\��0�R�tU!=b@��c�"�$�����Q�H����^z���}R�ZE��qc��PV�|���[�Q��rt�!K��_pyH��i�M�T�����Ұc&k^�CjQ�t�=O��_~h_�-G��Mz� 1v=u,)���F���-�B��t�[��ob�_Fy��.bm�}#� �~`���$��]B?�d�(���b��˓�֛?��ｘHB�\�j l18���B�%.��{���%%��D�tX1���=�&���G9��":r9k�ڕ�}�3�~�"�5�ʆ���,{�z��������9�dFb��vkH�z��i Pぅ?<���ᛯ�0�l&-��=��;�kEo&b�&��U���C���k��U��XF�����;R���u�.�n����HΙ	���)��7����Hs$_Q^Fz���o}�Z�AW��!�ԝ�����lH�`Q��t��p��)��]�G�揦!�R��=�p�⽏�P5g�g�<,~�U��G�g�ob��}�O�i� ����⓿[Ғ|��=���YغR#K����k?C#s8�:yU�W��e� ���⪡����Ŧ �15�	��b,b/V+���+���-1���M��Q��4p=�m��'э�/dѹ�Q,��oX�$|�"f;�:��'s/~s�	5p&m��lD��ՈL%�ҡ��AA	�˖���T���i�z�B̌F&$��x����!;X�(׽U�fP����R�m��.��x!���*\%E2�yQ/�4?"�v��tsV[�*`4\�5��K�	H�(�x�i�����7��	�S�@��G��_s�1�M_|� �a���xp?��²"A��k̵#�dI|q�i�O3�]�j_�T܌Ԭ�IQIi{��,g�������yP�W�N�����2�\�|?�}�lx+�����)�d�'T>7H=����-x�v��s"���+���Vxq��EM2������M��>�O��83�7�z�R���U`�N+ ���0��ci��f����j4�-"<@Tgx��UYO����m=({�#���l���w��9�Yϊ��!��i�#��y��}D2���eL~�$��?���=,