��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,��.��̡�+P�FuX��d-��N��$%�I߽7>wN����u�]��j��ܹ�Ucל�|�=í[~��k�5�P�ؐ��T�5�����#�p"&�l�z�Fr&b6��,���Fԟ�Z�_�X�;���93	�����Ǘ�M�~���٘�2�c�D��������f� 3łߥ:ա�;kv��ތ(�}��r�{|�Z�LP�����!�Y{������I��܊7Է^f�L5�:�	�͎������W&��b��wD���Jݎ�IK��et��1���Lt�:��6�Ui�;F�o��!b��\#�Z��k!�Y�#Ao��U.H����Ƈ'U������0JN�]�[�萙��5��!M���@gb�t2�&J(����1<"ʧ�#�_�8��^���i���$��a��If�R�p�?"놗Ǌ>=X���mςspI��kWz��l�3C�j
��u!�#��?ۢ_4�2��>%~B�L�Y�S�I��T��E���|�RƊb+߳:�2���U{O��?�A�+���S�E�U�b��=T��v鮌2�c<J��&�su�14f�աbv
�S�8;Y3��Z�]���,!���$v�U��΃�\+�әJ��ϭ���ǉU��}w���,�ٞɂ#,������;��_|lp�BTuo^�����ԧ��3;����<��Z�ׁj%�ϣQI�0���ޞ���#(�*����Y��c��s���`th%�{n�~�x����˘���V�'k�����S�{�(�燅����:˪�\MrO��������t�K�R���Zq��Y�>�o��]��@����Y���%��m�w8�U�<��{
HK���,���T��J��*.̑=�"���� 6@�0�^�����L��M�4��+�%1s����M	��#+�0ִz��<]��̞�H�W��^����Qǻ��`��5�˾?Hs�l�-�r���}�Lt�\����p8�*�~gS��D�LI=�xw��R
U��nm��.h��h���znu������*��>�Gy�B�ߦ���Pg��D~7��0��Y�M�����zֽ��A�un�V��8��i"W���t}�ZO����͇�4/PϽ&ͥU���z�U�a�O!��m�6D"$�}$a/���x鼐�T�E��ŧ�=ϫ�$t��2.�Tfk��`2�8+T��b�4��м�4�ل���m��傪�T�>��0��zd,G3����ɿ��L0��[ 	�"~&�8�C������� �~4l�R�]��m�y-���*�E�������&�[H]�#d��5v�!8׀�#��0_w��d���UpC��n�b6���# X%�]�m�c�D��n7 1za�A!�\ik�b�-��?@m8��/�̖Dۀ7M���ʭ��uK��� -in�{(]�7���t���a%p�9g���9��a(KW���"�8S67�W7l
��H7���{���R��#n�!a���� ]��1�#Fo��*_��A���gåݏ�1H:����/�����W�P,s�q1QG.����LS��Q��;�M&Q�y(md�����nOB��5�v�"��A�gr��\���];u/����j[�M5����q%�
��Z��t6@��^��3y��%ܪ��D߾C����q�W�6>?xC�QMw�h�k8�[GAq�S�tC���n3��q��ظ,�HdN�idZ��%\��kt0l�z�hǶ�}��/&h���SV�lg��� �]2�9����<��x�J�EUBY���e�v���5bްx.01?���t�����Ӳn���8r��2	�U�n27 �Yf����h�����o��um�vT�8o:�Zw|e�f�א����|��s,c{,�#J��t��b3�����eq��ۍ���dIW�u[J#��	��J)n��6�hk
5��}�.�R�7v���o*�`*՞/;O+�t`A�����'�"j���w'���G�
�Sz��kD��C�3�JQ��0i���mQY���6X(X�"A9��O�ǽ�#8J��.��IIa��G���)���H �N3�'k�!%ڶRN��n�͑������j�m���b�'0ʾ�p>�	���쯋�Y�&v�FQ�\�n���<�z�g�E��H�y<�&�WL:�G�+W\fc;,
㿂)�4���XU�xr��c��~�=w���&d�����;��늁�YV0v��g���
�.'I��9�ʡ�M�ɉ��6MY-�eL�$_���ħ�[u�a��2��sx���dgl2?�c���nB~c�����-N��n���v�|���!�oƃu��f��bW}ç�P�P''��X���L*$����ɕc��91o��G���������D5�B�[��*C0�Яq@}������
 ���iש�7���(�M�ú�,�Ϲ���՝1���u���n�����k�x����[бS��: ��Ԧ���3�F&6��B�����!�