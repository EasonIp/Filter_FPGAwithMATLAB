��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�J��"4�=�7(�T�JѺ�ő��,\��s���ӣ�F�؏Q�j�U��uA�j}td���TF;T^���~�l%�,c,k��wG�?4�_C:��&w%�w�>Ik��c��(�J�\�<V�{Q��,��S}JUS+H�9U�M���#9�[)�7b��]i�C՚�J�e���+�K��s�]�
��w�����k�`������������/��b�p�s���Ŭ�� #Jtv��gA ��N��MHcq\d����&�w�šS����gR���mb��#Gǆ;�X�"���;�� ���t�t"�0�M�ߗ���[�*�7�\&37�MވZ�X}Sz'H�d>er��|�_=�U3OWiq��4��5�� tU�S��#�l��YV�Z�E����8�>�*�kp� ��Gw\�������Mzi��v��ox�HP�ٺ�5c}K)0��j��D���]+�J��C��;��6��z�/�]]�\�޽Q0��)ikoI[~��n]z���ϑ�i߸��Ic*7R��"�`^_g�ȱ#T�Ļ4i�[q��P��
��Kŭ�T�ݘ��=�6�#�A�b�tZG�j-�栕�� u8#Z8���\�4���>J֮@ф$���lA#��5s�3NAE]{���ਂ{�;�\!�x����"@6=�؇��q�4�L[A�����[�A��e�M��[���j���7��SR��9����H�X������!��O�>y�<C	o��%�H���U]_��ڭ�o��kF��~fX�P8��*e��1�*Ԧs���J�����������Z�!&L�%K�\�@%h�cf�''�@�O]�}�ĩ�B(�`���N�)��I|��8�b�*g��<q��T���kK�i���l�Ҁ˔|�'$�����i��Uh)Q[=�� �Q�IK��
JF��^	��)�mL���~�s�uC��Co���-<-�g�FZ���T���$���Z]��j��'�i����R���$�q�b�	A�+q���E.]~��}�����W�ۑ>��Z�ie#"܃���K@�"0�@ 0���k,j��T3��0m/
�~�}6"[��/0��+Ɠ�N���j]!Xp_����r\��,��c�{��Bl9��o'�s�
�V��.��P�GT��u��
����T���Ve�<#.�Rr8�:�*�1wo���<�ES&*����!Ы��k�Ǻ��u�'�}6������j��̧����j���ISX�
>T"�&�?�Y{A�mT(Gk��q�F��'�:���	���s��م7�.�(�M�G3�O�ȹ'>��aYV���ʭ�]X�Ȓ���oнmՏ�NH��[�������H���9��)N���4qB.�$"x`�M�P��<�Tc���V\k}��&�o�� o<vcz��k�j&�?��zih���WH_���秡L�~��=��s�飉�U�Δ�y�I&L)������K�ƻ������Y�>�h����	�RD\�y����Ռ����$�r���5(s(��li��V��n�͸2�ܩ���$��	.�a��%�l����u�{8��rⷨ���\*ȹ�"��0S�X�4��̢�Hc+�4K��T��mۘ��yE�0��8e_<�= {G+�/;z��>޻Ƥ�����X���T�w�챔�	��ו��.�+����g4��T��a�kM�M���X��}T�*.i;�ƌc���0T�}}�p�u�Y�U�0�w���O��g6�Q��9�<�q(��s�"�BF�Q��Q�?ֳ�/��5¼�o<rk��H�?t��G[� �$2ɫ���ʳN#m�֬������.��GΝh�K,l%?e[���<��[O�Xy�~�ɠ)A�6��N,�� ��9��5#\V5��Ϻ;���)����I�v���D�xwP��MeQ�TɍV�i5��8
]i�P��Saֱ�B��k��Qk���jf����f,��#Nv'R#ţ��g�9�O[�[�ڀ7�Uk �fA�E�.|�(i�K���A�̞�����z�¨�~!�$3�1y�U���NOM�<�Ľ���U�7_��+$Z�^��?�+P��vm�b�),���_�gpI����=�-��_c�0������78;/ct=?1����xB}��Z�'`����x�*�;��D�N�ŷR�rNs�^=A��t��͚�3ض,�	ل겾"�Sl���J�x
�4��G<�*���*P��^���D�sg<�7!�Pp����JbBp�Tz���V�������v��j��ɦ���%�h�
Sx�eԭ���@�
�@E!��9�������to�n��<z��^��Y����@ �O�N��~�-�w܀s���>e���O�����UK�醀�����
;����[�b&>$��@�M�����ݒִ�p��#j�oM��������������C��ЗG��g���5٩b�#�mU�f�ً�(���Mĕ��O�s`��1�x0��b��v�>[1�p�������G6[�_���$�p1L]��A�p�fc��Ԯ���aw�s�iY����*�?[�n=o�	� �f��X�ke�`.�-Ic���ڸ���u@c:�F���̗2z %z��8� �;,(�g��XET�|����^�"�g���;^�,Ա�"<P� ��d`����M�Lh��x4]Q�RT ]C$L��ٲ�H�jfm���~ �F�d/n�gX�O���G��4t�U.r�r��V��g܃~ #�>���qAY���`	܍ͨ��x2Q�9�*�Ze�}M�:E���ڙ+��*2EQ	���w�;yY9��x9����4y�U�u��.�{Z�6\��p�䅕�P��ё�CT�� ��w5�sz��~͇8m��;D�r6�ޞ��a�o�z�� K�O�,�ԯ#B���+�׺�RM�ϳ|��9M2T��[��O�Q�^�"�߿Ss�Atj'A�_l8���4P2<;���+���6Gvٛo�b�����5�:a�*d������<}����O4U�'2�����İIr��2�m$� ����fI�����~���<D!��w
4��w�p.�ӛR�["�j�g�! �**}��/��͸�4/�5����{W�O�`�^f^N�.uR���4H��~��ν~&vk/�q���dۀ���-A�/���zvz`M6�ȟ"�w�������7~�l���4S�~��t-�H�v�[u��{�49I�D�y۸Dm���ᇉ^k�v$?Ff24�	.�!��BE/"�w
�
7��"�(j{?�2���>�!O�I{�R]���a��OȆ������xEk<�$��*U����`�/r�-?]�_������{1��L����0���)��ڏŖ�����[O�H�D	�]��8��n���W��WZ|p�}��i������x�q�!�l
�tKk)Y�y�*�b"þs��Ta+:��|s���Jо\����P9�Tm	�]z��C���m�dH8X݀�+�"��]�;-X�T�h[�G��MB~i�*�7~�6뭣`��t��?�������yx�8^\��O�N�`���e.�%C;�d��t�?CD���棟��	<ҰXV`k�Qu�{F�ب�a}��-_:Q��p�	�C-�?UM�"���Өv�bs�uT�ۋl3�6�&�ez�Z
lI1���1���N����r�#��4z%� ��!���j�� ���	_A�����wg����R@K\8k�Ɉ��g�D��]K��å�n��ﱟ��{pju���]�l���h�*P��6F�&*�$�R��+��8_q��ӵ{�9���������u,�+c͖��DI�/�������ۂ��/�ĊH��O#pc@��3F�yg���C��	�,��P���Y�fQ��!=��X���L9�T��G�o���C���� o��?HO �F`1J�F+R[d�eE"���\Q"���H��)UcJNF:+C�~'M�V=�f��?A�B��[��La�&Yw8��e��Dzκ���/ް�8�Ke~�0/K4�9������S=�6	,��N�l���|���m�a`�� �g��K,e��o5����ʱE�QסIL�O�ó�I+�$/V�Z��*��G�a(j��ݩ�d=ڔ@[�+[(^bȴ���zm��h�np?%^~*z+tIS� �<%ċ�� ��\^��95�^f�� �
�I�38�lOǽXUrG���1Ր5��8�,�<�+���f���/��6\����l�A����頋�C?�2�6�Dvw�0�f��U��je���Z�R�l�LXX0��=/����Q�s�^ѕ��ӟ��9g�	�X�E�I���P �b9�0<?űAω��r�@�1~'ц���%�lb������� ��(��o<쨆���u�n�EB�]��G-��ٕ�����@�����ޠ�ᙖ�Nn�@`��ڄ�{�]`�i���˩'���NꝾKO%�N�����D�`VCj��7;(��յ`g`�����FJ��'��2J,�Ԡ���:,\��px�J�����k�;l���}������CU���ddx�ΦaJ%�*F��<�
G�IQu��B�[30�^�a�����v2�׵�zi��|{5�ꭋsd�z�!���������`����@E��{����`Gn�X^��}��c�Q­�A������t���Q~���+.��TO�R7y�2{P�$����k%�������p<;޻92��7��	�kc&�f)�T	Ӄj"C��V$�p� Fgҗ��:	X��.=EGA;N?�,�N�w�5�;#��{C��UoAd�ČU֟��0�<�4h�l&�7��r�T���`<�v��㚬��̖k]Pߙ�6�m\�5Ş���%��J�F�����Of���/)L1$E��~A�G\�V̊�q����2��*U�O��J��Ns�fw?�i1mX�Zn!b>�m�����7z3��"
7�����A�?�{�y���D`� "�Nה�i�kS�z���2=�U4��?z�0w���o��<$meV��Fn6׻B� ����)��j�)�\�qqA@�!��9U
��-Σ�#H���IH�.6>i��B�L�!�Ȯ͡|���EE��㻱ɔFK�he^�*y19_EK�g$>R�=�"��#����S�Dػ���}D��X�_�lq*,>p������?Es����?� �$��5?̡�����00¸)}�M�U�QuD�mV	����?S"��<��9Ɉ+:T����g��&U�U�M�\S�b����{1q�o�hAߒ�Kx�3����� ���]2�T�M����9�U��yj������4�fc�6�#4J	a���)~��i�T�'��1�9��%�M�ˁ��}��t�R�!]r��r}֢ɣ�u(8,��p`��`��VK�7��p�;/��(�-�n��ʆ����Zn����/�g�.�%��zs7l��R�ay��T|fX��!ݏ� ��g��"o�_r+>]h���α�	��������0g�d������ S��G�m3�f��=�[��쥣����`�wR[�*�e�<Xi΢��Xµrr캎{�V���q���dZ��>���T�^�N&J�@Ї�F����f��Q��/u	��ɓx@����T�L�p���τ�Nz�bX0C�Տ��$=�z�-Dl�t4q��A��H�p��WF=��7rZ%���&��?v��f����d�)-��_N�z9JN�=Bx��_��-���e�8<[<G�A��]�>�ُ��� ��ڏ�}��w{��E�R��`o�|�Ak�A+�I�r74I�P2
j�,����`m�c���	=Avn�^LP�Ծq)���b	g��(��a���������С0��C�',s��A�ʺ����}���0�4QX;�(pA^�01о�<�X��_8��������SjDv?!l��~�"�Ɲ�?a�qfp�{uL��d��֦���Es
�����<of<��ֽ�ell�`�4��W��4bJ�+�JƁ̸BPf�5F�2˵�l+o��/-�k]L�raD���ҕb��'^ݕ'��4T�$��ㅲ�sP9��R޹�@����J��.�-s�&���`C�K�	q���6�lM����(�V���7�4 )VL��l�oSǬ�s����6\�9'z��H�і��C��}Т�� ���]���l����+r�?��J�Ԩ�Z�uN%���)/��5�ţ,K�����8	x9�}����	;9w��<Ɋ��I���7��X����z�p�����h���wX=�F
��!�	:�d�O��1
�Q�K���ܼ��`��f�Y����a�S���{�� �i�l��@�G�}��W��]υ�:ݵ��75��z���M�[����.<�֊fH���%�C�:0?o�)#,�8����R�bq�-�#;[(�p��e\NI�ޣKj������R�&E����0"��~���@αM����t����]��Y;b���!�n�
�o���,���Ё,0�?�n�K8�[���L)�K/������m�u��f��o�0\�&ui�����������o2��� YJ��φ&%���-U��
�O����^ͨN
4+GK8ep1�o�p����t
D��� -���&ƨLM@_�03[�s��Mc,��sZ��b[�Q�~y[G��>��G�/Y>�#�d�]��(,v��rq� X:�E�����h�6�h��q�"8˾�9�pHy�F��ZC��k����#Ay)~���/���Q/�pE*,B�)���:�2�'���<i\��1�}��)�ȡ����ʳ���gn�O�2>z���\��(�X�&���`cķ�[;��v2�6\�Ka}=&�5��f#�Y�����Tp� 0�����$}��5*�3m��R�_���? �(��~v$ug�ݿ��ck j,�!�3���/G��g��h�c����D,�����'��q�Ȝ���UM�͝eѯ�̃oc��q7:����рK8�^@����*�>�*6�������&�Ȯ�;����jٯP�Ó[�[����<:4��G��VH���� �"6���=H2�e�-Be����{9 ^��Z�Ƃjj�|���yC�E5&0���F���?��1�����bМ�~�G{�̉�!�*����L��FU�Y�Z�����x��B_>sV��"o1�L�(c9�)ī��z�M����
�M��t��g�_����}�-��\��9�ʱ+#�協��}�j&-X]�^��j��9�����(Ko�����g(7Z',S�\�)]p!\b�.�&@�_6y;O����S)�m3��?�C^ӣ�,p�Y&�[i�}��l�����5�+����n+����R ��X�_��, �e�x�ǹ��}̵Qw�8H�}�j�.��7�}~Y�lp�P3S6�畭)|�J+]p�o��m`�.�v�.�s�6��Q��[=��4~�J���R�O^���d������}�G�ٴ4ᩪ�@,���=^sbĞ����F�iv���z�	�H�A��lpC��KC���L*��
 0�R(#n�(�z�y�S�swv�y�O�sRL<�@�+�[o�����Fs{�lF�=�g^pQ����(��[��*����=p-(�2�!�����bMH��vJ+�Q�����F3��d�G�(̍�%}�O�Ή>N�V\���(Y��3Wr! ��2�E��.�N�zP^ �{M���b#�X���:���^n��P.�f�#��VV*d"��Q�U�Y�/���2U�v=b�)S�DˑŬvZ_҉n�)�9v�ǵL'�Lt2��)KK%b�99��i�䝠�7�X �i��Y]-7��)��_<��/��z"�c��4��mWI\{>يX�p-u��v�_�!�K��l��GcdU6W�i�P����U��b�R�^؋��5J�Ja5�6St��JN=���d�.!��ڕ(R`c7%��'9���obc��r�O�N-��s�%}�q�E�E>m����WxGuE���e�$v:�Um� �M�p�٬)(��W�+C|�V��	!Z���'���B*�\oD�7��e��t�' ���},�Ҟ����gѧ�����v������)|��{��Jj-���=Њ��W�ӆ��val��m$+8��09"
��6	��!���5��� .�K9�u�g�(z�Rsۖ���x���ȨJM�wE��ơ%��6�OmC-g٧��� �Q�������r��6�%��F�B%H�Uw���zcjdZ�|�`6\D����E�����7?>LD*b@���j��GzĀ�t9�>q����Qv��r?�$��A�B'S�5�Xi�
Y4���-O&��{s��*i�͏_4��Y�c
�?�Z?H�!g��Xꁂ#���#r�~2����Ƅs�	s_�N��7���8�e�`�_���h8���wk*��nH_Ɩ*#��|������{VǞ�k�-��n���ըj�.��^�E��	WƊ��]�պRA�d����,��3!�֎&�uX<Ib�%��牕C��+��@1�]u��L~,(�eIX,x�� �٣,��q@�i���8�p�1!◞[RK�x�m��QuebapV
��ށ�?�}X��O^��-�/��E��#���h�U� ��c��~kCH����w���7�1��2S'��6��QN�z���	��Y�G�j����-#��S+y�(�{���e��G����Ͼ$����-�����P���rE�R��aky�@-V�xU���i'I��'OC-��TOc���1������9 ���9�+�r� �j���$ۓ'Y�Bjo�d+�)!����Y8��9���TǷ�s�[(
�jG@?�]��*�n�ܭ�����B ��7I-�'xd���"j�B�Ԋ��".K�CSFsb����%���Bj���9$���[�6f�����H?�8�6������l^�P�e<c���ˇ�:3"hRJ强`ܻ��Q2u�+��9�#�'�ri���4p�{e�g��Y�{ej�>��)'0 � ��L�I�u�؏A4�� ���b����It��w"� XxA�#��yM�*���"�>R>4a  b��af4 �#��ob��vh��b]2Di|��<����6K.c��e!�u��$7��-<��x~�T��IԘ���u�a�*|ghLmӆ��*�����[:S���;��gÕ��h/("�$
��IT��d�ྨ"sl伝�:����a�I�ߟ��~0��hC>�%8P<I$)p�EiD�#<ݥ3j�ט=�(��E��.Gj���nu����d�JV�et�7[T�b�Im�����e8��?􈧆e9������*{���+������Ck��{�B��ᶸ��0)��顚l�|�I�L�b�����u�Îk\f� kl��u�^~I�وV`a�����,]��[8|�t�6;k�萸�1�|R/�BQ�2�s���&�.p�,����.]%id��Xو�F ��R�h����(K� �Q��3y�'�]��Ȫ�.�WW䈳��7�G��}AC�e:�擥lu3D���U�C���q����.�D��qrk5����?p����[�,�=���V��z:�7-=��u��4�d�I�9YP����M��|6�ݤP�z�9���g�t�ym� �:W�B�<���Z�C0]~��E��b���`�G�	���<�m>e03���l0��i�2o�
j�1��Gh�]��Y�9�*5ǣd4ٵ�f�q=�xz����H��ׅ������h��qrD�[D�������M���2��}uzDڇc�Q"��������"�����o
�`��q]X����:Ⱦӻ0W���AW����Д���� l�0�4b�(��Q�}ۊ�d��:X�y��	#�c%��cnn�f���a�|� !	4*O a��q%�E0�aK��؝;�K7�!@Քe�yH󶤻�Y	'	.�J����6�񽫀�u��=��ʊ�x�\*zh��x�s���2�Rp;�ւ�+>�x.,5=��w�z.9�ՎK���N�|)-0���~�	��]g�^"�^s��ә�1�@�J����~T���\��1��X���H0���V~�E""ȍV�ŋ\����]Y������>N�"�wO��#�����]���A(��o8��Sl5�>�P]���R�d>��ͮ�����sj��)H��/��!�1�2��u�z����#�<3D@�q�\�����enwE7]��%��}�u��<\©�z5scg��%�i����R��w�""k�s�]�I Nǆ�&���U�,0ʙ~Q����[��AǑ{�+�w�)�%��v�|�8�В�k��v���Ԭ�(��Aɫ!&����)��߇���~)��[nf�5�����6G �q
űɇ��"��A�!��
��B2�&0e����Y�vo���.���GB4'��6�E��Ζ'i>�����E��e��������R��S1+JE��}uJa��t_BI�M�� �8����A� Ҁ�厈6H��g�^�f�CL�N��Y���3����A{��
a�/	]+�� b48���G��C�
7�L�1(��� S�
�iն��d4b�:dI^&[bvc��� ]��w�h���l��e̾��2���PP��P�-*�7xGr�) \�S�נ�p�������Aw��tqa������Z��;�G��c�3ѻ^R1�V����K"�;�5�}M/�F�h��`�+�
��jU%�A���L��ü�*�
bL8�.�w�	ZV����b��J�������F�F-��#x�?���BN�2}��\q#*�
���n=�KOɡa\��A����1f���Os�s�k)�l4f��Z�er�`��ۅ$�8�[k����jfA�]�P���1��!B^����
(��B��Z����&�O�!{���.�甾G��oކ���X���ӛsQDmB��rI�����[_[��c�z��š�y�X�+�7xev�^�Nz���!��@=ŊH&�g�dX�w��Ķۣ�"���Ͷ"�C?�d��K���q��뷆SPV�-�6w� cS����S�i\�����ƪ	r��*. ?��t���A�"��͙#�Rڎ�20 ���Qns�Em�6�?���#BhzZɾ��q����y,�Q��TTz��js�X�E5��T:d	��Vϖ��6f�B���% ���.��%nԢGuuG���{�.��z*�צ�R��K�sR3��\�%������	~���s�X��t����i�*�;���z+C��@*�������	���B�B�5S�4w�r��/)
>W{B�����[�a/14�ɦ"����^5?`fI���ʟ������I}MD���S��W�s����QQX6(f�#W�?��s6�-]m�?��F�H��Q���;��� Ԗ��6��&���/��b��S�X���`\���Q�e�맊�]��+��=��@�-[����Y����+�=Hx\Hz��3/��Fo�_�k�i�u�ͱ�>j�\fs��od03��8*��wJgp��.��O�,�J������OWP�JC&w#�!/���4uN��ݞ���w�P�/<6aP��T�d�J��(zK$�����A����F�0�U\8��~�G7����5��ؿݪZ��<��j����S��v��>ө�?3� �<[B��:�y��K	t-)���%cE[8�J�{?���� �Û^~g.��fvȡ=�CBbʁw��]E��)G��2T2��:��j�h�IyށZr� , �(DIHn�r_�n_0����3^Ύ������HU|M��,hcy��&����W�~�js�+���ܺ-V����TE���e��5�Fj�~���:t�@�.	{�W[�s�����ġ��d�ܻ�%� k>��}.�S����C}�2�\��ۨ���~�W�7{u�����|(�+!B�$;��e�W@ݨd�!���?OG��n4Q�[�y�*mccҨ��� I�׿��8�Q?;dN~���	�YIJ�C#5�E�j<�ˮSm��$4�]?��#�V�Qɩ_��=Xֳ7TSȡ��O5ZfVQkD��[/��v�� ���`;��V�ZB�64�َ¼��� s;�yn1�����_Q�O��=.�'�Z�P;�
�xκNP��{%ۋB	jF�3aV����WFE�78%���n�wFc1�'g����G�J�T����(T��3s�9�qx@9��66��g���u�����t��D����`��|vg:�q�����0"�+���!��7���JO����$Sk��s�5�DU�d4�R��ZZm*�Jr%lPb�F�`�]}v����[��^<u7��h�o��g��U,b�'�	|��.�="A�6�	������r]�ޮ��%���NM�QE�q5��l�^.�Yp<�tЃh!F���P����vqj]�],��]��B��8��B�ݩ�PK2a�f2��&F'�_��Ɛ�Gw�!i��P����E����9	9�ꇬ��3]}aF���>W��c�6i �"nxIc�W��(�%'�� <��&��P�Ɠa{�� ��P})�I�bz WӸheM>�6��5^���
���*�=8�ubU��k�����p'��y&��~�a�T�P���x[S��K���E ZG�~�!E����9�0��k����B��������59Po�@��"̭�X�Uh�d���SP���Ŏ`_+�2J�lc�
���L�����6�`o��<@8p��zom;�7�1�|�����4o#T�NV��������df��/22L�!�P�e[r�$�7��w���1�͇Ɯۻ�=!Bh��$�W�3�TG�������K�]Z8qoI���mj���GL�����hY��G�dy%�"L�%@�����l��~W��;Z3��=��4�5FĭTS�����V�5+��=i�g_[�Pw�#9n������R�>a@p��������(U�e���D�㔤��.�|�ڟIm~�����r��94�q�'r0���6�m�p�
Ȳ�{8���fcm,�����������h�w	���ĨP��#����.���v'B���R�7"��1=��x�q\8+�u��&qh�z+�f1��Hs�X��Fd��r����K�6��`����,Mu�N��0�(aL!�(�I�E�5���5�U�i2�
�G���+r�M@�k�Od���;��=?6���xN�T;P�5*
?`;ƈ�e�t�\)R?�zz��-�����_OPj��טE�R�Cj��$c�#m��Tʷ���+�����bv>��>�����gE�j��zaxc嵢@����a^S^X%)��Oأx����u3-���Y߲V�L����@K�[���Y�YA����+�������jn�(z�a'���UUH̓��~��\�� �d�
S����Oʤ[��+f���_f	�[��5����L�+j��)M�B�D��>�\�e�H�/�RljQ�jg�r,G<��;�[�Ω�����Fi��å=4uw�����q�*� �8��g*�����\w�Ĕ'Vk��u߉��z�խɜV�,�ǐ!��K���$X��s�2il��ߠ� �m(		&d�W-X����E�L�"nP#�������̹lJ�\����mCg%��F;1R��d�^��=>+��!�l���t�O�ѧ�	�kx�n�w`��;�.�j�-��E.a����:H�&v�1^%ob��>4�Q	qYG7��R6h���c�8Z�̇G��칂'G�
ԕ7���g�RޛB�kȓ��z�_��UP!nS�Z�·
��'�Ǒ�v"
��M�5rL\Kvb��n��x�ա��?�'����]S�j���Dm<����	�2�Bf�����;u�C�8YO�vK"�%8�Y�.2����k6�[_赓b[��'�^��m�O�R�5N��-gҁTX���u��Q���ƒI�)9<4�'m�K8$���	�����y�5J�&�Z�����q��*�ᕞh�<E�d㺸eU@Ֆ�}g`Lύ9�$�����5L��o���Nk���*7\,G��wt]!/2q�/�u���#p���B�R� >��Zv�O��W�->�����c��m'�E&1��C�9O�l ^�LBb_|�}\�:ǣ�y1�P���[`E
��1	�,x��Q��<I�N)�?����;�D	��דt�����Z��Mc��r����5����mN�~N�9V���4�y�ד�������6��D�pE�iś���˵vOC��H�ڔ��LE9A��~.�?e��W�-�69w7Q8;�	�}z)s���W�%�{�i�G�P�Dy�5�G5"f-�;BS�n�!mo��\>��=e���Ɲ�1��@zt\>s�/6�Y� ���AH��C��.�9�>$�n�Ul"&��N1`�ġ;�T@��F��9��ko�}�fx3��;}�$;~~I��;�����H���W���)����S�UA�{Ӟ1v6V���0��bfJ8�9�����,\�<x��L��3�$�����i�I"��#���7��8b��M�SWP���]zG�u�����OK��A�����`�@�?z ��Tx���H�B����?}�����{�n�8_�i�����qY�6�[�ŤF��7tU�nk�?���16{���e3��=�Ah򣈊AFi��g
�a�pD[��o�#�Y�^e�_�ne<|�$u�L ��ʊ�?�Gɏ��]�(��Ʃ�%f��N�n���4���$�Fz����±^��`,Z[Nd�*d�x��v���9/��M�f�%��	C�ѵ2д�1�B�_�N���EWH���#k�4#`�:��	�Ze1w���[�w��c���b�Q:�2�mmA�V�E�&�A�Р��^�KU
�/�|��R1����ʮ<-g�%���I��f~1��S��-�kH�����oQ4�Wp@�Fa.�.���l��>�݋��a�-��'�{���T����R�P�ax=�1�`�n�b#6��ߩ�v#ԯ�M��w�OR�zjne}=!��.l�ug?���R�]�#���1�a|ߤ�:A�;	�h2���Z�I�R�EV��k�#-T��ۿEﵭG����]�k -�Bb���&��Q�9�9<���?
��������$≼uhK	΍�/@+�����0�	l\ձ}���:���ೄ�y�Ok��&�D�Ŀ.2d�F�#��/�8!�*q._��z��l�KO�f9�����rp�HU�WX��,(�0�"Y	�,�Eʥڔ8�^m	ʺ8،�l#2����p͠�ҬhR�8�
A!L�?�����_����Ye�Â�0,�sX�^�ڑ'ܿ�3QUJ^`�
6
2��L
(m1�]�wO���2�������M�[}jte��7l�l����t��Σ��a��8��� �c�>��/�A����iѳv��$4;�پrw���9�&>���508��g�������k+����Z��M#2�t ۯ/V��U��*6@����0
�`�k�N ۺ�сpXX��I 8�Q'Q��\��$<G����L����Y�0�"�'�K��p՞m@���c�L�G��;M���Y����)!ײ4�>����M�@��%N����4�,1���L���3b+F��CFt>�.<wC/�j���AcY�Ny�PE� �`B�Q(��E-+�ø%Gt#%(]t�U�c]ig3T@��G�M�Jt{�l^nb�OG��T�?j�s���"s1[�e�<�?E��3Zn�i�ְ� �ߕ�'���-��	��{�hD���P�)�|9�BUy��R
�#��o��ڳ�C�D?dR�%>Y	�ZJ(·�c��ݢ\7��c��@�|j��WT���k�9��)4�;4}O�@��"����MU�A_�r�{}N8��:I��&I���	�c	p[J�*�t��B�4��vozK�9�6C�KS$m8o��B�tIoF�b]h��Te��6�P�������,4�b��]Y�)1#�g1�����x)��?��_�}�ڝ̡��!�=�8(\�Y�g�]5�>�$(�*ԁugZ�}�?�-��PѓJ�B6�X6OH�H��JU��W�M��蠁���\�vǚ����L���?�HbuQB�2n
�����"��ayCs�qW����3/ag��SR��Q�P�S�Ⲭhl5>���؜F��!]
��7ʏvP/.��)`�b^���d�$	�=X �h.�%oW���n5��A7�$d��{~��M�d{OLC?����!ƨ�Aΰ�<d{�Λ�`i?����o�E����L�y]#�}K��[���H�0�#����3�w��:��H���d%f��O��o������
5P�咃�(u�Q[��D��N������V�f+H��i��{�CiI/���ϛ�կL��<�LQJ�L�d�j�P�q��;d�9�;�!5�W8��N��ۓ=r�4���b�Mv�`�(-G����,H�/#������P�6ڄh�.x���N���������_�y��yw�3=h Gt�����H2qA���h���Bb����W��J&9�14�Y]U=2="鐷� c	DvנE0��~����h�R"���耞`��@���g���?�?:.��鸋�#��H��{z�[��Da�ÿ�8_���?����-�~Pt[��=]U-����@V6�*�q��cj[k$�.����#�IƠ�#�~�|��K�꘥��S�I�X9�jdmtx��i�}L��F�s��tt5�y`Ӵ�4�\�G���l@e�}�������m \���%���ۍ���g�|S��/5_w8SjŝR{�K��P�s�K��=:bOY�J�}Q��{���>x��A
p�+����^�i2~��d�6R��o�8c���U��K] �x�X���7�"ʦ2��9w�fp1�o�8IBYy��H�m��1��o*���k���~E���15�c�fW*1��T�9m4�
L�Rb�o����={��t,?n��'Egm��O��Dp!�ℂ���6"eU�������%���)�b�<ή��ײ��=ˋĴ.9�ɓ� �= ?���¬{89��CH���O?U�Ÿ�9R߂�6�<��ر@��f:����V�Z3���R��AF�S�U�N��S�zt�U�6������i[��;�8�7J��Ԍ�r+m���²�?�q_���톞����!���ъ5�*�@�㞨��8`����H�	l�7� t�k�GR�m�CRsܓo=��O�D��ғR�{Z���{L�ߵJ#��Ҏ�,��ʵ��^F;��,ޝ	(�R�`�_��������B5�dD��V/~Z��i$�!ƣs�N;�˃�r�a�N�km�Z ��L�� ���Z8���?"!/c��-�a�$�A�ӜJɈ$��{6<�A��Ϩ�b�a��I�*�!`�:����>���f�b9�z9Na��J�x�=�|%i<�WNs���82C�1L��Z���#�=��a�	]R�擕&<�|��0��1c,�N�nK-�!	;U�{A�z����|��KS�QB^�@S������=���V:I���$��<�4�q���*I�|J��[}�����q��(�8��`�����9�-���ԑ嵗/�CX��Ù��rw�4�|��z��X�q�'?�ο��A��Ic��"Cf,�0�w=�f3�L���T��k�[���~�"$�}�˷_��l�i�3�Md�b�,Pn�`*S �7ٚ�O��&S(��J�H����&=�v�������������q=������E�[��Z~���̎�InĂ���dFM�Xl����� �p,�m�{���+����ɱ
/�h�: ��p�M�i��9)����N�X���YH@�ϐ*�3
~�����c@A�	Rr��0yS֫V��Hā�b��,i�b�Z��nf�\N�[/-��|�Zf:���t	Ԡ
:'\G~'	oEU��l�O1�^|QP����;(�l�qdm`���c�t����@Y��70���qI4w�e&�a�T֪n�aS� � ��o��4'`�cxeW^�b;a�>EJ�0��2�IR�Jչ!Q�3��ϭN~ڔ�:|�Z�t@�3�s���$�j�A�H���q��%��7�8�
��#��%:bВ|�|'e�������e#�� �͠l{x Ԣl��܌1�#������C�vx�Ւ+3wlQ������f�Nc5����|�1|Y�-���XbbI��*�k'k6o6N�4����
W�-�Ɩ���^��`���@�����^`�*��j~���wc�F6C������k.�GFe��q��B[2bW4�~}t�����K�\�a��������ܩr���6������>V?g��pÌ�\^d]�痈�0SP)�Z!n��i ♽$����)w��$�3>�?C��Z@�Fx�LC���WbP�E�:3���������2.-�s�{$���\Pm��'�5��9G��ӃM��4�	Fs2�x��m��-�c��%q hNO��ލ}���u7��	R_�6\g�`�GR����@�Ƙ�ot����w�EY�i;�{8�&�鐻�[�B���L5cΰ:�a���Ɏ��08�	���TX��굩	� ��l2��������WJ�a>Ea�H�u��~i��q.��V�R'~�-�	$p��_"l�qL��,��L����1�2Tuуl>�x��C��̦d~��Z������q��Yj���w��M2�� ��m�ūRju�2�	�N�\E3j$����~~���xǿ˔��-�����ꎝ�= �dV��ج,�k�3����u���f&� ���!�(�nT^ʝ/��|����EKZs��=�Fcn����v�1>P99�]㳮�!�Lr��[����Re������4�3v���͐����O���ɟ!�����s]���ɻ�Ԃp>��P�F�Ɵ�ѝ��O`���54KP�퇠�xr�Y�(����:��A�����Wvf� �������*tT��,���_mFC��")�d�7w�J��!��lA�T�GԊ<��s���h�	��!ٳ�^�����+ �*3"�lk|���,9�B�%� E]�����Z��|؄11��A7+�s_&�88�Y�U�nY�t���=Z�3D�A��~T��J�Z��\��2�!��OW2��2�vu�P P6-3�U��ܸ�t�w�x�|�"^��:^qS��{�4+='
�>�8
���{�����\n��'v����p��������ў��+�߱�����v�k��dk�Gx�ttB8+r�Օ��.�3�ۑ �l��t��ڇvX`�	��1[N@�%��U��$�fn�ϑ�Ы{�����x\��B�L֋�i�H����Z���B�e܏����S�V�\������|7D��6�;�h�ٳQ�WSl�Wg�C�zX����$��GC�j�Rc��? �V�UpM�k��u�I}��p��������t>�ӱ\�G�T?�S�n���љ(u��	.]C�Ǌ(�����O���D?ֳc�r;H' ��S� SE����M�l���)���
���0���l�����á��X�Z/T��U�l�=Ҙ��z�̋.|Y��C!�]�]��D�z�Ty�2�fJ�;�o��)q���a�Bu5'-���5���{%��S��6��5��p�kX��H��R�E���[D�QB�#�xhLڙ�he�g�{2���N�4� ���f�\9޿a��֛;�;L��&�:[���ޔ�(s�7�e�h�f���gV�?��΀i�lM��7���/���A{JV�mE�>�!r�,��p
�Q1�K�W�Y�}�AVM��H�m�0����,����ݏe�ޗqrA�~��})Gܺv�p�-Q�>|�L��#Ơ��)t����ܩ�Ua�/2p>�u��{��B�3e�},�f-t�m�c�����j��Nf�TԀ��p{-KlE��~S0�O��3昦ڞJu�<���P�9�Gʤx�'�C !�E�,�y��}ɯJɟ��o26E%1dW9L���W9�}L)�I�w"}8P��<G��C8�Q���j>S1��%����o�WH���Rօh��[�y�U�vn��n=$@_S�K��������6֯u������V�=���@�덺��Q��.4v~�hr�U��$���\|E��[`٧��ֶ�CJ"���<,��m��+D5n��tJ>�5�=�׮��w���F� ��Tx��Y�v�%�;o�2�o|А>P��M� �M=w���f瞅h�R=��d7�/��A��!�x�Ѵ�-�
_��Y2����,7�R��٣u����xot�[���3�ng0G6>�m�\Q�~���c�4ސ8����o�7�@�VkT�Z r��� �D�Kgl^�|��xZ��G��4�����cYp9[z���0&��s/V�3���74s�Jr8�k5��[��(�1+��>�����)�F�L�K���Y�����\\Dt�_ͨ��ȷ��X.�%m:������J�'�]��&)m��?�p��le7B��(�7�=��I��(z���,e�=���Z0�H�BT'-�Q����G|�����2L�馁
���5��ɱ�[%{�г4�*�)���O-4Y�d��%����*n��ܷ�n`�@S�1�RV(��0xL�t�����qlu�X�Z���a�T̍%'~2�
?)�j8O��t��p�C�����"��V�4Ք��c���\�$��^��etYЧ���Qk����ۃ�x��I�d6jK�.:�T���Q�TF<ɘR���Ĭ'�����@�R훦 7�0Q#�
�xU��_��m�G�{�Hk����#F~��n�!ȶ'�B�]���#�I���VA��,T4��^)@�4?�m"�0�r�?��2�Z�/P/w������Mp�X�����
K+(F�7��̖�0���ئ���4���kCX������T����UxO\d��7[� T�G�O;�.Z�5��� ֖h���
P�q�U����+��@��U�ˇ�G0vR���}6���W@u�<�����U��q4AS˝�J�
���bs�wj��(�A�L����S��r%`h�Վ�89�F}/7Z̋?wBk_� �@$'�I����Ӵ �p2�՗C-%=�w��f�@S��/08L�n�t��Q�T�*��<^R?$�5[U)�����t�2�q��QP�ZSPws둝�2���S�M�"�nO����4 �"�
Vf;ʃ� ��k��Jab����JE��/�$�X´�ه�7��ϡ��<̠��f<oʶ�n��;��5uC_��Rxjؘ�1Mɠ��AA���H�b%����F��[���_l0�� ^�z��p�4GE�s8��N�3��o�b�|�J�y�c!��JYK� �C�95\Z�#�NJ�u�/���X�w`�~����:%*�D���,���B1+�mnѬs��Y`�����s�)��s�J��ܲ/P%���/���zb�Ȯ���*m�˵��a
����I=�ŋJ�4(
�Ӟ�!b�u4��(�K�����y�e�A���q�C�O��aqQgǲhq�M)`;���\<e��q��a����=)�잛1C�SCZ��;�c51����Z��s�@�a�=���}��y,E�0�uK�=zut\�������@���r����[�?�!<g�Tw��r�O������4szs�Ә���d������E�`ZC�q=N@��=��Y3E;4��I
z��dv�ޛ��r��!��9�w��u�Z�f��;�e�����"���p��v�c��F��e#��E� �M�T՜[�iG�Qs������bC��!��o�6֪(-k�H�)�������o����ӣ�Z�,ẽy��h�lː~7R-	@UI�с`T�C�{���SI!?р-+p&��% ��dV�k���B�5�b����kɛ���V�'�E��X� p���(Ri��;��8�e]�պ��|����N��,&a�r�u)�'�@-�Bn`/�����z2�V5��N�Ŧƕ6���b����m�_�9��#�������6��a^�{�O�x��HRh1q_��:��)��F��8;��k&Tv�ւ�W�No���*�#��;,�j�����ԕ�@A�6_��;�\1�� ��G���\u�#
�b�L�Ӻy�ױ@@�|ӀVdD�\�3"��Vsl��sc�5�v�jNډ"�����}(�s�e-;]I�i]��*�d_�)AE}�2���w�ܗÑě���o2��l��sk���|��*�]kǦ�ϠN�n�sӢ�є���Ɋ������qVstucf_ŝص�7^`CP��$������������^��.<gfhY���]�a�}���l�}E����� A��ĕ�U*D�,��_R���_�/�T��Q�KfR���@���}��It��v��>e�R~��`�(0K%����x����擋�=�����̏�ۙC?DSW 2[J-�#Bnw�N��J�$]b�PX��}_c�L��BD�B�w6��t�~�O��D"�