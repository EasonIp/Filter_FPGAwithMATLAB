��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� p�X��Y��!�����j�V^�ʳ��*
�,���I�)/��� �����{�4ePs�Ҋu�b'��j����Bw�>Uug��q39�NPU���>��Q�~�pC���ڪ�- vӏΛ�9ȁ��﨧;�2p�kq̭��cɇW �??J���=�#~�$��"k��,�Zz���h�;��89q̮�b�d*6�5����Rd���S펎�d8���)�p�qfƻ5��Nj{c�I�����eTo�5��XIID����u�<	�1 ��!g�nD�%A��
Z-Cej`�d�.��oN]&s�����d���?�L鐩��ԟA^Q�vn[T�����w���sN%�H���7Z��pz#�t4��0w߫�S�'�]KJ���
���>��u�����u��h"s[:	�G��m�k�w,����1D��i�r�b��zꃯ�, viW����]��ɢN�S��z���E��aTO���5�NZ#�2I�s�J��s(P�7w��lRy'�<�?ӵ.r�ĺ�5180�`�"`=�h�ې3�n�˶O��F'�8H�I�)��]a59��wiﾗ�F�1�ZE�c ��ӑ�ǉ?�Ҹ�3F{�M���A0���_B\jB�Ӆk�gm�?s�k�p�μ[��i�����H�M����ZH׮M�՝\gU����u9�,����q���L�Z�����;�G?",	�:��mSo~�"�<H����7�<�\��v�\�o�@�a�c��ݷ.��])�VO���\���6\�G�P�w��'�Fr��� /U��^��҃�ZP_�[)l[X3����\�+hd��N�L�C&�~�]i��(&� .$�"6ku6�`�#�ec0O���oc���|��|)�� ;+�2Kb0�!C�-C���
�4�d~�e*S*�Y6��b�h�J�������md�����-H�>�P^�����i�g�$a�Z���;�x�H[���k�c�8�S��b_���x%@���oπ�~�!�	�۫��A����P�RO�YϮ�a;�E�@��1�N/VNT?���H�)��-U��? i�/�^�UK�r�R2�3�B��d��c� U�\'�~��/�C��D�x�Kc��i(e9�Y��`N4�m����K�%����S�6Y�k
C#��E��)�L�.�f5��x�c�_�z��lr�FΧ��WE�=��?��g�4
�� ��Ĺ)�,����KI:�� z��85nŪ��v�3,�e�C�=��t(R6��C�^��U`5�9��4o��\�d�d�3�8���Y/?N�%k�,|�}�|g����+pQ��1��k��o�>Q�pF2,B�\���E����!Z �u��3�Mf�W�/�rGJ���Djd(����~�Hz�W@[��ӗk�h�i&c�O����1}賵!��Ͽ'Gc�Z�����i�l� ���ތ���[���\H������A��iZo>$.��j_��,D-Гk��6��yM@z
���]����~+$.�b[ZT�A��������'ô9V��ύ�u_J����e�:^Gp�_�a�_�9��ne¦lȄ{/���Ō�Ӌ��	�(�;(��x��xx�P�s�!PK��M��o�_�`�5�l��;L�h�Q�@���ϋq��)Vg�GN�;���4<4���W��`���J��Q��PD[�e>�&r��^I�]8x���|�<X&�[��ś��@̓J��A'���QX��4�
��t��^AP��P��W;�T�MF�;�;�w1^��do��eP�c��ㆫ�le/��c�3슲�b�U���z��m�� �P���(*� ��/PqqI� -�������@�V�L��9���"C��f�7��pmx��^�#S5#�+�ѥ���B&)|l|�G\�+�n-<�]���j����9���@!�9	�m��V.�r�����9���~esVÅ&�)q�jaB2̗���[�u3�TF�<��#P{��:����ݠ�#���S��s�@|�;.;bV��?���$J�F����Kh� M��1�)=ԑ�wip�Nl�vu}Y;K�7x쏏��L�s���ޓH�~�%�Ei4�OL��.1�*z����<_y L�b��?㌎]R���43�/X{Ŷ�	(��hr��k'��{��=k�gs2L��F�G��}J{zR"EU����������
y�t��?�k�gr=����p{����
��9n��,�d1tkL���:A��P�Ff%��ړ/y�Լ+-��T��p.�CѴQ�{��l2�D!�xu�&�����:�g�}j��\`cԜ 
�}؃)c�݁|�O	5�L��? ��lQ؎�`Й��f�o���'"�(�%�<�n�&����rw����&-�
��5t\��g2�&�k�C�@V�,�=����2^��Y^ऩ�K���R��]܂N�A�r�Ʌ&s��n�1`X���T�V���q�����P�D��}����\��1}����U'*]�)$�vQ(S����`e=I��[�agX+d��p��O�Y3�����d����Da�b��F�P��Kh�s�����71l�I��rSų<=���t����lr�q�]@�<�!���O~$X@�B,���ԝ�˽'�l��I�� �7R;9^�ܺ���K"������+��"U�yU��^L�g�������'���`aC����(&�~��Y�HZ�,n��d�;�v:�ܔd�*����~iA�c˧����إԵ5��%K'R�~x{Ϩ��<y�z���x��n)*D䄚L�	�|Xӈ�  �����Ǵ8J��N@�Cޫ`[��,�
�����٦�y�2 ~z��Z�x�I\�.�r��St7��\4���A!,2�8�ҽ��d��q��uD��������^�zG����S<#b6`D�,?��p�����8�򄩛�� �CEx�5Q�2S�R2�� D�����(�ġko�wʬ6�Oq��C���?헼,I�x��?��I�u ]�*�!�@"`˷PK[��	�Э˝���,6l��J�=⓾\��q��%?f&�����������k~ ��簙NB��]��b��@m�j��H���O�p��������ۇ��\`{��F���u�X�ښA��kEۇ��d����c)�R���&=9r�cyAE'�P/�Z р�s%\צ6�Cō�ԑD�"۔�&���BlD����'k�F���n����f3��-��8�[�u&�d�[7P(�@0n��/�FY�AF@�����_apIն��C�sp���p�����Pm�&���� 9Z�x��)�bÀȦh���~�u^q�K�5�
H����ĥu�Ĝ�
���7З<��Ps5N&x݄��ʌwb]�ِI�u�$�d�]x�̟o#�N-NE�"��A4
"��m��R`��f?"�CKt�~<�������SB/\r�:�'�ვ���g�v,�ه��~�5��bL_@ځf�tX̵��1�.zd\�|����C;q  �T����B�Vʞ\��n�G��t�)TMxg��\Uiv@����+~�8d��8��8 b����&���EnbX��W̑$B����XAΩ
*�b���0�:b:\��е+��]��)"ꗍ6q>;����t�n��떃f$�)��Y6m#�};,��$�Ν��6o��3�6v����|����Ŷ'���fP�{���p"'�8b'�=�K��
����g��>�!u�����	B�f�YX�>���O@���L>��M����������8����I/�L$E�{=���&�e��b��:�"��I�<Y��9�aСΘ6�ײ�>ُ�M<�Cu1�&�Q�.��� o_~� ]�>a�f��
"�%�f�q9{��͠�H
uBT��!�R�#;�nl��яm�F��B�j5�=�_9�w���>\�s"��[��h<�·�:U�s�wB	b�p��vEw}����6p"�*�l!�r�%	�:�nm�0��V$��P�R�9S�S�Y���yȄxF{8����2�l�N��8�߁KM��q���-J^�*{��/lf�6x�ܢd��T��J���j,]ɗ���>��Ҍ��θ�gT3��6�@g�E����~\|U��n��U]��J�[��<+�dWZ7V������Ss�1|��%2�q��l�S��ٳ\U@�@Y"�ڧc=�&�O��SF���*�!�4�3�MA����WK�P����6��B���ɺ$����7�=�)]n����n&��� ��[<���|��ҏ��tmq�PYrtB��K/{"RXH�P�.㸂ۈb6���X�� �?-D3��.��j�Ď]����*�v���*0����T�OowJY	�qw��nGW�d2��PMHa�����X�sY���)n�cg��}�h�4���D���Kf�3�7딲p^��n���o7������	W���m�������Yb#��Rst�>���1�����'6����`�ԗ�x����E ���H���0��?B;�w�0�H�@���2)υ��8gЎ���23�!c.�K�Z	)��y܋��B�C��S�>��.T�n ��,U>7�Z���s��B��;�ʔ�gC��q)]�����9s�)ؙ��)�P�0�ڭ��&�pj�Tw߆���,"J��N�L���D��S��u���bЀ74��l�+��j���u9&�,���^x�bU-�c�٢���-_O�=�~@�a	�p�m>ܸ������3h	��L쎌G��>�U�M�BY;�A�~@��6Rh�B�|p�;KS���W����f�S(n,�f�%���,j!O�B�c%��Ѐ8wg{�(�̶.U?-���f�� m��vW�@=����b�ɧ)kwQ*%C�~:P���E����%1��G�����S�B(flH�x{B꾹�B��PPI_�����p3�0����H����h�:�<�����^Vm���>���a���hDO���0���.[���#�F��PN6�t��^`�ʎc�X��;ea���2���t�X�C��L�m�I�J�����W�r@��`$���ZU�}(�&�b_Θ`^�x�}�I�땛����v6�3�}�Oj���71YY8(�B���X6uP�~���*?���㶕~�ƪ�[�5�V�%WDv�\Cu���ʗ�������6�-�{Fo~�W�˺��&"ai�ȫ�c�RX�hN}S����.D��D��j1F���zJ8�&*9<} �	�Ǖ/L#T�:]��B��� �gt����S�`�R�����pɧF2��R/'>"'$Au6�~�	h� Z�_�`�ǁp�ik�L�Ѣ���� e7��_6xIZ����\^���a�ғ�'�h�g�=����J@���JIR�kW"�2�:�u6���#��I�����%��8R³%}�Sa�!��+~4}�l���X@�Z+�O�|S�������3�ٽ�l���`B�3*
�y�)��f�5�Z`�z��I��M�\���}��!�\HF����^���D��I��gWt\6P�5+Z�:��%U��'��/yb�0��h��%�����Ԟ1itl���˰�85��Q���X% 6f�U��·r} Y�6�f��P #�_8���-"|e�y��'k8P�4q��'S�O
7����A ��7����Y�Wk%��p4cR$_�ZS��\VW��[0t��t��
���6x�kgȿXc����[ɛ<W)�Jq���6W}�2/=�-Si�n���@�pe���I'|�?�}X����g�E�W7c��4�Gq�����|���--���_�C��*n�0�g�c@���`J�-�tĉc��2�@G\ͨ�������,��O}�BaM�ֵ�Q���I�0����z63y���ۄ����<�6���&��ۢ�]0���jh�kosr\_�)�.�\䡉-�d�;'�)3xZ0�_���&��e���{ң)f�]@r+j��}7�t*��7.�8P�tl�ej����K��%K�@��n<Z��t�:�+=��u�h�X d�?��3-�8�����[EGB�o!�}�rU�~Q��k���Z�9F��1��ƕ��	��g���a[#m�`�2�hn0:�������ku�mE�kla6{\S��X�]��4�i@4B�lx�Z��+-���\+��WC���8��T��=釵Yݡb�PL����Ad�x�� �$.��	�n����V �&�|����E��k�'&���֍��ra�*�����މ"[��k��q�F#�2���s��1ȭΪ[L�`b4/t�Vն:k��&i,C�<M/Se��6fA	efV1Ӭ[�ں�װ��}��g�}��`�ƞ5�RSU qρ%��������e�g���$��t�@
��M�C�3�����,�`LȌt�J�h'S�/�I�Ti<�����g��a_�B���s.�AnP$?�wh�,o��[z'M��B�]<�0��W귢�"l	��oZ<�_�֚H��q��*v =M]U�Q/~��{Q��}������f�5C��YL�e��^@��0\"����%J�J�L�2���tL�����)d��6��y�L/�oЫ�%s��y�6�r"�QǷA��s>[Aa&!4�T�:B�F*����|�P����7�x�5���B񯉖���q��nꔞv���M~��J�Fx ���fJ]̸�w���c�A��L:����ܫR��W�P���d�8ɲ�KK��iA_�p���f������b�5�����,��Y��y慛_��gP.R6�TA���7tR�m����Q�3��+��d����{���y��VP�V�"��ꦲ�wL�� ��a��D>�����`��j�`E��^� �� i�.$�j��+蒪~Զ-��KV� �������:��I�{k������m��\��P���~.4pf�h�Uu�N������B��!�d�#��Q��TzFkH��8��@
+
B����"�-�&�=�����L���S�8�0 �Rk�� !>��p��="qy%�!�!��:ω���r�gr��axZ� Z����GY���}ڙ-���A��iP)LR��왷_~P��e�&S2òߛ�v�����	N��ڞ�T������yyN`2;3�C����V|.gj���_o-��S})�-Z�����CZ�x�/�=�X��c�v�2�-]��y�Eh�p�$��_3��z��3���2�@q������I]-���ҁ�g|�F*܇9+Y��SԊx�J����)�+W�1^^ 3��1
�k�'C�(����{��?|�nk,�%��4Rn�:{+II>j�n��ٌ�+d�3�h��&��~�wH8�r�k�? �F��ޯ�u���m�Wx\���
��#D�g.K����d��V|�b�h8X]�^�aX��=j�I� +8%�*��"����v�/$.�rԕ�/%fxK��<�!�}��R��{B/�'��F n�E���*.�}����n�54�7�4t�=�~��e�@U��^��( i+^����C���&5{usJ�8�⽎�M��8U�5 h�f���ŧ2tn���~����P"����,ek��q�ԋ<ި�Ytr%0�P8�¶�<\_�BiF{�H"_O\'�P���k/��U7�蔶� �ːq"�[W��T�0w�o��v��~A���$�����;^$�i�r�N1�'��
%�$v�0Б4���'�_ؒ�)�Yu����0�":ǔv��Ev�Ѝ�=��C?��)h�K��i4['�������2U�&�Y3��F�c%��]����"���QA���*Sa8�n�թݘ�?S� %ZݲԒ��5ݤ|<�_,VW_�?����*��Ttr�Qo#f_�}�W8�x�?�9�0qE�@y¹�C�aN6\z0�0����/۽�S��bZ�B�u
��ſ�ŊfXSk�m�v�C�V��p��	�3Ǹk�,�R��f�~d[زR�(�DS���˸;L�JP�f��j﮷7¶��=nZ#F�.��/��_���R�o'`
����!����>3�6�t��G�F�I���|6�ku��:�BƁ�4�C���6���r���W��c�H]__�V���+kk��[�~��Y=Mn*��p��+ʨ�S������:B�!��S�>o�aן��j��b�9F�sٲ�S�c��rޮ_��B"�w,_�w7��ED�z�O'��4��`�Kt�_A����ې�-a� H`�u��ɣ�Ǣç���}(�>t}9Z*���y��-+��D��(ĞvT2vL�[v��_��NZ}�&��%&�Dq�D{��T'd�;p%v��Ҫ��\XV� 4��d�#�}�P��9����k=|����D���OCR���;�IߺG�����4�
vA���>O�l,NC��o��0���ձF��^�v#�����,UY�>|(�K����t�Q���h�#��5},��t�����h�o�p��r� �1��4D����?v/�}�-�<���z�e�>qU!��w
b8�y0���dB"�liC�BH�S�gִ/�]>�e����z�ṯ\Ra���נگj=""G��Ht+�
�p�ʐq��s�^��Y�T��%ض-r��)�4p#�%�h~�:��/��֮,���7#�lkK�z.¡AOG���Iv
��`�Q����.X��T�;��h��XɳP`,u�&P3XN�{��O�I��:�=�Lو9v4�S�����d~�3;#���_\�F-��k>�t�4{��x����؁ƶp =����~��]��n ��k�p���[D3Эb��¹���)��F�����|w����ܒUH��2+���Dx(G�EL|�'��47^��%x�<�D8*�P��h��2�4��2B�
Oi
 ��LP#��#�`x �#*L��t��d}v�a勧/�H��d2v��֝��,I�ӥ�1Mhoߡ�!���m��1��%��]�_�f|	�'j�O3��ƯL��5,T��s~�������đvZlQxdQ�@>B>����@����Ai�Z.�٤�]+0/D�r��d��L�OA�iϱ�bn�3��o�f?��ۼ��t��=!��*�3b.��N�AET����R+�h/�m���1�iw\TH��GXX|5J�|"�BwBFZy������ݙ��{ �!̑������Gw�XF��S�:?'^i�{ZL+��e�I@����]� ��{�Av�A�s�c�\D���	��'X�	s�v��q�u��1� <���t�O�A� ��oS�ս?d���Ӄ��E��J=���@�	�!C�)p�����Oj�8�<��d��Ę�J ��J,_1��� ��흓]x�T�LeΤ$`�*�!V���ۙ��R�����5{�l��k��Z�k	w�?�YX�`p%�:,�=B�Wąv�]-e�i��/p1��2O5��ĵU�/ؕ�Ҽ��� 0�ª'��@
%�-�����N���%y���i���W�m���|h���	ҏL�B>y���B]�,�ݠ��x�eE�ћ�FY͂6Y�_,��hV�ə.cQ2?��JEIv8��L�"埨�?zI��ً�DM%b6�/��߁�xhUo^�9� l��S
�
���d�;�_���W5�W��M�j#�O��,��ȭtA�xp-�(V�q�i�=r:Q����o"�ݚ���h��$	��^!C#B�N�����8|!��;q?&�.��TB��(Ĳ۵7�>Sgi�f��,�@���D�?"� ������r��XHU��鬣���@��F;G�,�|짰�_W���38.M��F �0uS�l�qF>���S4�҅Wz'AU���$��LG6�����QGx�D_�:z,Q�蟆�m�
�+����rC�j^�gp���Ñ�7d�#�7�TP;��MN�Ix
3��l''$������3�x��Аgo�� X��A���/CT����]11�����л�c��i!���L�l�	r���Y�[ Y�� �jK��V��bNe�9w�Y����Z{��񚪈:�d�[���1G*��J�&�g�'�5��7�{����a4l)�&j��.~�L��=�j�*�%а�8���C\@d�Woj#tv��~�� ��>��U��b��d�f�@ޤ�'�3N�s2�W�r�������̍����b�~Bm��Q�F�T�afA�8J9�I���J�u-�����e�ha�.~qg��;\�
2���F��۽98Z�hW�o���_��Ёŷ;�-s6�*B���gz����e�@�u���|g0���7ׯkT�������D�/ek �Z�hM��|�Ġ��h�Kx,����4��p;���j$�I�l����L�l�8�u�Kj�Izc(B�I�T�K8,�Y\�=&���`�ox� �Z���������(��u���Vu��	!2�+d�GF�x·��
���IX1D�S���W7p�1��u��Z?_��2 d��e`|��4����]��Xg	�"DM���	�tל�؜��C��?�U��SI���_�|م	�4;�2轊��y�9�%�*��>��r�����[��L�����̷8�8�Ʈ�3�n�M
m���m� l���IJ	�>Տ/��:�Gά��)[,*����;&8��zu#*��)Q�����R�'�>����3{v���nx*�'��!v��t���
H٫)����<6�z��M��M�a���S^���g6L��٬�I����z�b�YW"���.$N{w�WJ��g`0�=�e6678��n��ڢM7qU��Q�uX^L9�3\hT�K�l�+�w"��>�?����A�ӛ[st�������C��P`��<�Ck-Cq���|j��d,!��S7��Ȫ!?� �EB��rT�gX�� D��Ԇ��^�k/m�*���W�u�N;}A�u$R� 8������N	`b���89BTFѱ����G�0�Ɉᢄv�[��3��z����8�"=�->k,P۹�g����j��(���}Dn��$��,et���0��G:r�w�����ԣ�W�q�"�f�vm�T���x��|ᙻ�D�خ\I�FS����+6|��@ezU�è5�j�,��53�^}��L+���P�S�U�崶b��f�7>�??��ny��p%�;i�\˳��L�������p�S茣6�=A9����w�}����^ �k����ȷ���0�#&�l���=���.a1x�uvT·jp�ׁq��V_��c^a�lyK���f����T�UՅ�b�Ua���e�^��JL��{�*��ƙ�T�
��}���qZ��l���DKð}�=����0�ّ����ֱ����NY��Ѝ��!"!��qr+IC[����\H�	�ْ���-~�L3��JcxJ�z#�N��,��/t9�I]h� )��t�(]fzՀ�b[��ݫA�B6Z�5K��N��x������9��)��d�������
��_�}�2l��IG)�g��P����)�2�#��;�`��ȳY�[�c\���`�
XD��u�u��ʞ���,����dZh�H�@��-Ӓ�\ţKu��J;tR#)S,:�$e͸?�,���ա�؝��y���҃W7�Ċ�t6Ґ���y_�~g���̽�N�S�P�R��G���+w74��v�=������T��9�<������ҵ���pFry������[A�}���nY���z�]��:i���
R��{���.j���-W��n����k]g&АC�	�0�#O�י�&M�D�X�{�׸ܟ���ď�޹"KU��.o�ڐ��gΆ���$	tag�y)��%O\�~|��M��#��y G���7�W�=ҏ�i.vſU������U~3�n��lL��d����n����1p\Մ1i��N;�*e�X���^f�T�#>��y����{�`��v6a�3�.��q�b������W09�N�DB	��-P N�X\�'�/�u��?��*���0Gr�W��O:�|��������"	��;�c��Lz;�.UH��6�S����n��Al'p<֋���]��R��U�4uLP���3.z�fM����ئ��]�sm̹��5�<�얢���i�6�*�����_�R֙��׎���7e���^Rϙ�#c�<4�h|hm�~v�	�&)v%���i��;�|�˧�@s�>� R
�*1�����/uH��GW�w������ ��~ 	yg���9>�.dD�*oR�	�Dy�Z�P�򈧧pd�(��Y�zv&��d�<��e�Q�b��U����=K%��䙸t�K���n� ���'�D;��Һ<g�me�.<�"������ר���IcY�!�����R����;�u9dE�ƙ�q��2w/�/Z�U\Qvs�J[�o��J����4�iu�b	
l�P��[&M9x���lYE*Og�І��8�Ǧ#|j磛k����m�uX[!+�*b�����M�e���S�b�W'����)�F¥�:ߨ�h�%&�Q��X� 	C&aˬB�o�������T½6F��8�O�Frz�\��`̆�{Zo�l�����R�0c�9'�I�׿�gU�����"�z��d�u'��Ҵ�l��&6��3�ӱܻ�͵/�(R�f��3x��Sݒ�s�����31�1|[�S��|'��>4�Gh�5gsO���$M������.<�>��,�Q����xt�S=�6z�qF	1� v]�S���6���C�x�}�G�%���oZ�l�t�X�;!t�4��'^�[�.��Y=!~L��Uwr�"��a����$�؎%~m�N0�KH�W�at�m��}���D���<�����9�9�(�dU/@�D6O;��Ld$|=B�o"-Y�(s�&�ǟ�������{�i7��`<rOѣ��ԅ��
�x��a]��L�Т��1�T��6������,��7���ò�;����+��$��m}��$�[��nm�c��(�w3VK@����!*��8Z2�QGl<G�E���h�S39����L����Oc�B���?�sj~��f)�ߍl�\-.��ж�^2/+?�Bo�!�RQf
3�~((��D�уmP�>��/������~��V���=aɒ	.�4��}��c��^do���	���"]���i}ъ�Ԫ3���&���3��nZ�A�Oqp��Pw���4P��r����U�q��H����Ѫ����E-"����X���g7�5Q�l.�[������)��׉�[�#ق^��~��7o�ITm�H�L"�5Q,�p�I���qx�,����Fؖ�����l'h/2�DGHJ�����=����q�C϶���c�w���_����9x6i�\ul����p5_�{c���J�x���q�q �/�hB�]n��¬�H�
����"å�>��N*#���yvS^`�,����C�`b�~1;9x ���T��}x��_۽����Cj�h#%������r�|�;?��Y��T�{}��%��Yꙁ�E�ǫ�rXN����<)��Wsln`�5�s6����1U�,Y����E`��.>Ns�0+��qZ˳�Cx��E%N�\�H�iup/�,́��e%鲳�yO$�r���N���0X}�i�]��Sw����Ray���K�5<�����EC����٘KԢn�E��,�j&a|�k990ֽ��������Y�}���կ)�|���|"j�~��⚛�$l������[��X��U:�;C�!��xR��|�ЏYrc1�v�����g����l~IM��m������]Z�P�U�� Ͼ�9A8@O�REN_3;0)#��\o�9�!��:P_VO��o����h��5�Iy��\&��k�����Bz5�7��j�"hZ$�}�N��P@�ѭOiuм=��ј�
�ͮ�ik�-�¯�,��a�*W�EA7�k�L�����;1No^� ���6Zß���\�Af=8BD��'���Y4F/f��L��~g�dFV�mi�i:.}�/Jʍ�4�s5B7�,���C���h5��_f�D ���Vo0r%?����C��P6C�݋�`��~Jt#L���ٰ��y�w����ɇ��*0&,��X�Y��'0�\x�7�2Ո�c;�%��ˣ�e63^��Ҧ��� �C�:(.@-T����.*R�ړ����Pz=Nj�B�'�(��v!�����Vոz� ����څt�p ,f����i����np�N[�b�.���n^L�	����'h�1��;58� ç��N4 ̝cXŬ��F�껡U���JQ�`�膪lrw3�����Ч���_��;�`hҺ�"�,�. ��Y���y5>��RK�)eу�W�Ķ��l��!\A0����X3�V��}78_�ȭX%,)�)����rq<�����Q~�` ��. ����X�����j����������Ե���#x�hM��P�iM��ϣ�-��H�9G=g���6+�va�'�+~�����;E(��.�$׬���M�b��*�����d�:�����P�ΦJ}J�AZ��5It��T�BC:>��k��#X@4��Ahފ�V|6&wjˍw�30����"���X}aj��y�N����C��zD�Fb���^�( �VפQ��;	���#�VK���.Ks�R) �!��DhP�B�u���HQU�<kI����FD�2�NB�	�~:m��Rg�@<u����Ρh^u�4U-͒F"E�Ew24%j�F�B���<��&sU���q��.-g��d..�9���v�2F�N�?<Z�T��E�=��W����p�-��3����\���9Ux�t����Q��hEŠ����~��9����y=3d�,��\z�}���0	�W&/$�/k�\<A�WHJ����p�~\C1�MB��%f�e�+�Q�a�n�xXj�.�@9���X���XSk~nX"�`�����e�x������t���8�_��J�	 ��NK�@�T�;�1l�Kt&�4X��2�"�>?�F��m�H,�'�-�mY�V���"�u�T%�Ǉa?_�T|Ooьh�e�]�c^�����������w�2ͥg�7�G��Y��+�t����h�Y�����Z��]��4O�"��)wE�,����n�T���AG�Is�F-�x�Nf
�l�� ���d�ރ�ڈ]���d�d����'�`�s��m����=/�[��r� ;��E����>`�#�]��
�V��˪�E]��Ј�0�Y�!��6(���F���~��+��5#��[
Oü�06+X5��ػ�"���P�ͬ^�*FܦO��������)�eR"\�C�[b�=;��oA�G�;��X`��DV��22Ovw�.:�o(~}���i���{�9h(9���Pk�N��Ӝ$z4'CkP,5������3�)ci�ŔL������``6i��C���k��Y�1��yOg�	�l��J��G�9�"V���ߎ��|�x=*�Y�@��H,8�
I�|wHF�y6QZ��ڐh�bj�jLM\�Pe�OY���0,���HPl�}4'+��4#�W�(�Ҿ��6�_q���bC;���ꂙc�=�*�`ȋG���c�S��檵䓨�K�E���Ґ