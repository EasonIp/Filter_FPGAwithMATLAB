��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$�ʰ�E���~l���>,;N����L�� ����r��E�)\.��X�hG�+bwf�!��o���r�wM�i'�����&�s=3p��^I�s�Gt�d6�|�ŉv���I�X��l����H��X��+�~Egr�c�j���\�m�{���{/�납Kwu��Z���G��V4��&���ɭU@���a�w�4:����,�y@t#��8�$���*׋�}�wS�l��(.��A7̵��OǏ_Թ�ҡ~h�"�Wnz=��hx�u�"�� �}��lÐ������N7���\VAȜC�/�x��D]�t^�To�|<}|~j�7هq��p�JPĭ����5(�J�X��� ��Ҋ���m�d�.G�!��5���3@��z�ǻ�����ߠ�o����#��3��8k�~��ec�T����hd����\l�.�y{��7P�����h���읫U�ؒ�c��rMs7�,\)�X���� ����s&}�YC�!j@���.�ب��ƶ��B��O�W᛹b�Ŭ��Ϻ7����&�Y�b�)�g�����_cmc���v����y��w��ԿR8��ҼrNҎ"�� ":�GcF*8h�	z�(�����Q@�'�U؞��%���TS�ݥ+��1�<���C�����nq��5��I�[M&�q�K�x�� �Tϼ�.O,�$ߩj�L{����ބ��!u�wnG�4eW��	�x,]�Oᤞ@��z��1�}]��`���  j/|� �p+$�����E%�-[��L�
��ˍȊ�e�8F��E+�����ʥ{����'��>sK����%��5��@o:�H�42l����i�S��QL���
x���,B������AnE�t�8�oґV���L�>r6h�����eh�nIln.�����V%�ث����J���>qS��79�9�_���x�s��������w�ί�?�M1��̳�.(.�т���g�O�X� �=�b��KGd$�(�ޢ��<�b��+4[R5�r���),Q
��fX�l��ޘ"�L"�K����PV�b�H�y�l]"�]��s�>Ev�8^�g�R�(u����V�viȊZ��)ZO�F{��D�~т�6����� uz��}�1,�uh �Q�
{�0�Eyj_��t����P�|?�,�g�ݹ��������J�t�"W�5�t.�B�pz��A
NFaD�/�PX�����&X	�'m��{"�|XɌ��7��0�T�(*1%@^��x���b�p�/<%ykѩF"��.�bۺzQS���8�]	ü%k[Y�je1^t��u��>���[�%��K�<�����tx��9�g�QDGn�v��v�^6���JD?w �g�#֮�F�=J����l�C��8ZM5�HU��?���
�I�o(������Í��[l�1�5�~م�ɛ^A�O���Jc���}��3�nDƭx����9 &5~��o��O�N�G�6 �+��*ax����`օB��^!:�I�P۳��]V*EZJ��1�.�),���/�x����'��	��K�'���]g�I��3�iV���s� [�ݰS�Z>r�Vx��!��-��X./c.X[V�&�-K&�.�=R�(@�o)�ʇ8D�f�Q�����ŝ,t����-�:����N\���M��Ij:����д��&jg�EON+��:=�v�?X1��݊����%N<������k�=�c�ٖ��3�]f�e �Ǝ�ٿY���tE[�"�:	�;ϴ�F�b�]G�b$�5)�e���v!�&��6�.�Sa���J��/������-(����l{,�гc�ۦ�b�R� 5����Z ws��g���U<���Q��!^���E�Fu�Ox}D2�l5S��KV�)W��]���x�Ýa�O|�y��P?���ܵG'�un���5x�"�ԡ`��Df:��D�=�P�)���B:u��'���z�3ྐ#���W|����}g�#�����V1R�ș�ãϮ_Hu�YC>�E͵�����]���^�q$��4�~^*lGӸM�t=�@͵0h)Ă��ߡT�'/�%��L;ج�2�'!O}.��p仁ު�g���1�AЕ��=@c�>�[�R��H����q~�з����î6p�������-vW��v�h��(ɉ��v5�2͸et�aK�������DP��̾��6shX^�7�@�L�~��SQ�HT|h���&��ޣ����)/1 �˸��	Y-�:�i܆�6a����FU�����G�u;�0g����d䖯<�]e
�*UR�,���eՑ�}�$>Me>���PiѪ�j�N�x��ߠѼ>���ح�+��������
�"��_�y<�L�*3sږ��s�K2�]i��6�(�;�K�EyÊ�(�������m���hHMA��S��؂��m�Q0b-��c��X:���1|��zL����D&�'�#�0��c޳/�N��vG<���Q��&�@�HT�%s-z���V���Jr�<p��H(e(��?e��7=Z���Ȗ��Q��ؙ9i��2/sA�;��w W[��U��K����+p�U�'�E�� \�?�;���v��(J[��a��9��<�:���8�C������g ��)�	+씧]dې[��U����=N�ԃ���ϰ�����'���+J���M64���;��ۀ<������7���T3�4�bM�Ϟx��RdlҮ\��;/�ibk�U ��X�p8s�:>���4qi�)������/&�4����L�ϥBz0�1��D��q��UQ>�cL�̯�����v+1x-[��ŅG{�{t���DځSPh��!D;���60"�١�TI�"?{u!��:,�������Ý�X�^_{�
ո�_�AH���Ӑ��*:�>g����s�����}���a&=i��')�@C�z.����}�����5\m1N��-�#�%F��g��Λ��k��������y�v~
>v�?�ɑX(�����^���M&Jd^e��(�����^�\7���~�C�Җ����������uW���,�V��V�͝'-)\�UF����Wi{}н�͓N6�7¸���Ϣ���0����k�т�*��e����@3��T�Z*B<���&�K�m*�\�ܮ���e�,����|�χ��!����?G��/(T��f�
���Z]H>���_c�WM [jy ��"� sp'��皓<;v)�`.��DV)~��fd�mԜ%jC�^�f�ʢ�p���ԓ<z.����:��R���ϖ^��[�h�Zn� ��+�7���(`��
�������עr�Q)�z"b4�S�|���lPH����7�(�3���7�n1�y�vM�B��o��m��|���By�¼�i����W�0������ĕ��!�[�����Gi�\��+K� �@]W�{�1Y'Ά�d��nmO�8��� :O1-P4��S6;�q,7"�9[\�Ma�9�o{$����#L�������^&�\Ȣ6!
�O��"M�����Y򀵄n�$/�Յ_�,rA*8�݋`E3���+!�m��1�F�/[ME�3��$RM��};
v�Ű���a�h1�$o�<���ˍj�æ�?���\!�[R��W4�ڶ���k��2�×����lm� �Te~'��? ap��tQ"0����[ E���5�\T^��>�*��:f��fV�!<3�N��ј��5�G[o�2���=�wnk�24f���q�"� e-�}�w^�V#�,��d�6H�J�����m�,`0��FZ�N�е��a)KЉ jW��;h���������*�~3�T=�Oj����Ǖ����s�~�=���)hJ��i�hh��s���z�K��(4�ʗꕶ����R4:f��"C�#KA��u���"Vb3���\��%@���w�Zga���}d3r��Ϙ�.��b/)��|�4�\�ٰgг Ͷ�"u�uR�GS����ek�����bA���H.�?C;���.BMPC��s��'��[9]Ǒ#x���ԩi�(lp����f"�C&���A��淰%��D�YrҬyS���J5nc�zZ�B�b�Y�y�i�z�02Sf�Y-!�u�m0�U�͓=,��upH�v,�)�׍��'��r�&�C�S�y� e�pӷΔW��f'��>(�R3:�w897A�f3_�4���]6��r���|�
cD�~�r�s�Ly6syr&��p(������^�����}�T05N���5mp���.��6�y?�W9	(�`���g�U�#e�τ_9a�d�iDR�l	̇jq9�¯�~Vs�}>y����o��N�w�k�o��0ܠ�c�Z�O��&�
o�l\ߋ>��-���q0}�ʽ�u�W��k�)y�*uh^��I�-�V�j/�M�ޑw��7{���pi�^!ڐ]R]&�V�Vӿ��j��V=�$w2��H�o=�E�d��e�����b�'�dW��>���D�今v ��g�}~ѯ������h㩯.@b�tW!t0{�7��ۿ7ZA�)�O}�a)h<B�4F�K:��x�Nt��b���~�;��i���L	�|W-��E&t^�O�G���tR�}n��Jyf�_�I2�̛����9�Ų^~�4�Xk1x�ey|E�8�$9+�j��ct'5������h���g�	��4\�*=��9ճ������K֒�&���۟Qc�=�7/�/�j�kx��{V���?�:4������\�!��gv0�I�%��e.����J��ƃ���04���`�w`��3��Gxq��gp
��ɀU����9�1����BA�	�dZm�Ά��;,z��+��¦���'3��Ҙ���G�T��)/�Վ�&�� Cp�h��Z��A�E�c��k��v���8��6`(Қ=.��CY0��|IS�%�.B�{�G���e*��׮���!��tb
���FG���y�@�:���f.'���Қ�#��KBGLw(���me����I���*�aM��-ϦK��b2̵tIXK�6�E�	�K�qs��1V� �L�(���W�e�/�zE���V�P��^S�g>�}\GI�������
ZR�k��3��ܺuC5��է�:��frC)�F��p):_J���T� ���X���B4`NI���wע����B�;޴J�ډߧlurR��lig�cy\rC�>i6����ּޡ����[�a���]��H��Ő}иw  ����1ovJP�����>��X`��]}��JP��So�7����N����-�v�W�0S@U���?�H_h�	:ˀs�51�-*�p�\e<�X�i0"M���Gbt�g���!�&[�_�p}Y|�zPY�]�6����������D4t�G"����%f6K���H,r
8����hM�Y݇į������u+���8�k�i��k��	�O9���Wr���"轭oǽ�&\R�G]mrcGJc_!��9�G�T��İ��P��^԰��9Y�Қ$��@s��,��zrC�2uȞ�{�k?��J{�A�⨳l��-e܍��Gl���]=j��S+R�wv��LK{x��^�L�-{�23btS�gN+�c��%R�z�ԕ�_B��WX�Xصdf�A6vnQ)�p��H���"7s��y�?^z�"�܁�g�S�ku,�*(��R~�4�%P�!�� ���7Q�c���S�`vz7����9�/V�����5!t�Ai��e�B��z`�0T��o����x���Xo�	ܗfU+,
B.0~���2>[���4c�9�nX%��h�����!f=�$#K-�l&+h7K�Ｙ�F��J�cf�����c��)U��q��ޑc�`�p��~.,���<��"�pn2ʋN>�j�)r�xϙ�DK0����3p��W]��,��1���']�ؑ7Ea���O�k���24�/AlsѴzU�������P� ��V��[._�-PL
ᇵ��Z��P⡐nVB���h6K�W]��,e�g���א�r�G���1���y8/54I�
lG:{���r�(o4�b����'z0t!�S�H����yO��R	������`G49!�w{�A�Ȍ+�$D+��Z#��Xpթ��e)�A�O�q�QQݯC \��A��j��B̀_js���]A�)��Y���>���@,'u8���Je�:�����Ċ����oJ��_�)$��I�a�($��D���Zs�=0��&o�d�uJ��Q�/�|=���� 5��Z�Z� ��5`�\�����%�C�9�M:@��"�%�����
��L �zB���U���=U�j�^]��.�@�0EN8�/����İ�*B���-��kpG�O��>W��1Z=�o)H�Cط&5��ޯ��`�G@��Ap!�{F�ę�]�g���2��J����#eQ�8$��-c�}`BC��~L���H|�T4h��{Ju;��D%�ْN,�h�p� ��ˣ!����1���WѼ=�/J���y��J�ɥ�Nu`���R�zǳ�� 	�e�Z-� �A_��W�p��
+��z �wL��*�ՑZ�ܿ�Ȯ"J*a��&����fyWC]�ڌ5�a|�3(�(QJ�����r��g�#����ܜ�5"����%pĚ]�^=�Mz����g �5Y�^�ac���<��K��ˎ\��*,�ś)��1z"��Q��f������⊥�Yq�v͏kO���4�I~.��{�};�a9���V3V֦�>sYn�LY4�Ԉ?(���Jl�?�5��>vH�����B�'�����"����&��\Z`�Uq��W�8>/T�Y_�)�
:W���'-{��E�ۯ�-b3���TO,�ZNӨgZ�|~n�� ��$�h�2m̺먆��}>�!@�h��aǀ�v!%Zw�園�������a9�J����to������%��ɋ��T8	Sz��u��1��nԭ�W�!����e��8GHی&S�T�':���"+*��}��RN��	�8�b�F|����-��T��Խi�A��5�!ŵ�6q���])�i�ߝb�?�9蕛����0�j�7��8/߶D�kX�����Ł\�lY�Rv9`�>��x�0�L*h��tB'�D�2� R6p�v�/Ꙕ���VeL����n�5��jkz5T֎������M���V�7a[�$��۩#�����ꐍWpԼ����k��]���T�:Å}t��.�b`�wk2���y��������ge`�Q�7ȃ��e#�ae����/�8_�r����Jf��^^sg,PD)����y���;QV����3�=q�ܓ���'�@FM0.���� E.��(��o��
��Hvsx@>d��i"�>������-'J�{�"n鍸_,)�� }���-|�P����~��eչL1�
o0���E��7hS�v M��"M�]͗C#�o؂�p�%��]���E�$)�� �U�L���[;��T��4j@.��C@��G�icI�+�q��࢖��мX�FN�_q��'�D�H���F.�������ufР߉�I������+�x�IN6vq:4�8����	|_�33~�df��ɿ*|k�
��>���X�e���X5�%[���9U���+�ktV��1`w����l�K��7���,���~-��艁7���\k���2f��֊g:��3'�-�'�g7CǴX��x��3u�eG�G�+�~f�j��L��s��cm��Fɣm�ήq����,80)��B|?I�V���?�w"�s�P�D� R��H���_�C��Sc�&�ԭ����[���%��k��囫����3%s1�j;ᇽ�niǹ͇�v e � �|d!����_j&݌��o��,��l0Tn.��U4�;pm,?�!�Pے�p���7ex�\�-�N��D����n)���#/pI�Q����T͢l�oNd���@���V��G.��{9��\�+X�ۏ\p�w!�N�")IYE	��[`C[���9nw��Vխt���f ��TF�j�ISd7�򜿚R�mҖj٩�vR������1q�۹������4.=o�
U�R7���&R(��<��/��B���o�W�H`���V{���2��ܐH0?)���L뮤�"R
�Vh��@�����`4��~�0N�\F�������E��O�cɄ����^�.s�C�&�5Xt۽k >�ݱ��I��?�Q�y>�"=B��0�÷�sA�6�{�� 0��ų6zf���4��A(ʗ�)61��핟4ŗ{��բ
�m��צAvr��A\��m�Y��LJ�Eg;��u��0��Ԡzu}��ċ�-<���r���������"��A*�G�)�����~�a��-�X���V��a��hBg'|��R�Mޥ�5��G:�}���@ӣ��6�c�E���SYE���4*{��/�|������M��?%߈��ɬ~� �"����%=�^�ţ��[��j���Xq��c��J(���u�v�V�q���y%�3Z�gy��}��Hڎ���x�=�l]� ���΄�×��R��`1��;ƀp����s���NA"a"������p�*�2"_E�:�+X����O=�`E����<o�/ 	Z�$=��˕.,�X�򡰸7М7?xCb����~��"?��9�T�[���Y��`��[��g�NH>��6$"ṉ��&L�df�i��J_��Aet���y��|_�iYk�c�z�q���`�و17gp�r9�,z( ږQkv�L1�{-C��(X�Q$���R��"!��(�}rcjs��cj���nw���t)���=�ů�c$�Bv�9�R[���*w,<B�l*_-���\���a����c>�J�Y����o(S���Z�w�<�~y,n�c�*8��V
(��J��}?A�+�+g:4ۤტ��qx5VC>޼�j%K���w~�=9P-�#<����H��o��Mઇ�`���im`��t����菗�{K
�kwq�O9�ݰ�|!G�*�ø0�}��b�˄���>��|��~��N��|������ȵ���y赏fi��|!h��Ȫ�w��^LI��j�$nHv�N�<��� 풣���G肏�A.�x��)6%ځ�<�n�gܸ��G�0l��G�r�B�~GZ���g��rqh�4�+i�s�}�����6�+�Z�J�C^ �	�1&�+fe͞�X�������ǻ#F<�h�	E�8�Υ@�? &�4v{µ㞯9�o"��ƽ9b[�z�l '�;=�uB�g[n��/p�Wf�f�e�DLA��$�����9�$-L�:��#^�[#+Ͻ?1���.�Ӳ�T�M��+0OМJ�Z���ݱ[�䒖\��e����E��P�F���'��(��\�	0��m�:���|+gV�u`π�&%�%�8��U)y�|�˪&�G�k����,�hy�a"x�g���À@����	�QS�FAm'�hS=$hW�C�G���� �&n�<��g��hhT���(��$��`�T�/ڳ��
V�@��qC���-d��'�Ƌ����ޘ�`A�ɮ�����7I�-q���L�9�&*�ũ��������ˀTv��9x$"�pBK|nˢ���C���T��A̱H�(�ZAܮl�3F�ɴZ�@����t�xu�i
V�;9��y�H� k(<l����Z���v˾|`��tOTX�=&}#)[޴-����	�8��L�z/�h�y�4jڣ2��������x��pw��ȐFR3v�zm�c�~v���X��؞v]����d]���֓ަmLj�a?'�T��,� �Ihێ�/.�
A�����O��Ș\g5j6s��l������Z���w�ѭ*�"��a���}_m��<X ��I���mWǗ�c�n��O4 &,������?6fdy����?�O��T݉ #�����\�n$��vP�1<�P�	��L
�~�d��漤�!\ʽ7>Az0�>n�ĀJ�SGv�6Y��Ɵ�Q�/ED������Z�3擥����ݫ�����Bx�Nx�g��*ѯ��h�m��1�ة�� Z�n6|�����=E��G��DUD�
���&�X�ls���r��l��7�3�xt� $��m�C�wY���Ֆ��>�7;w��.���z�$ew�p��!
���A�x�Q]�\qP�:$��s�C����mC,���k@�%��-�3��~4��n�]���闩����I��jq����46���Q���-'���R>��������RĦ�g�Fg��M�,a�Eqv��cۣ��R��B�Ĵ:�j{��Y�k�/����ނ�DwQy��%k���YE5�ӈ^�9ڴ��%i	�q�ϦD��B�@hTN�<��wL����J��8fg�������<��Puq�ͳQ��I�p�mHҬ��*��g��5���_F_8<k'p8u/��Ő��A�~���+���I�g�ZNڷ� ��ċDD�����(�LY<+(�7��Ot�]�FI�Vm���ڳ�M��+��E���:r�cp��	���P�s���ፕp�o4�;�RT��1�F]�H_�;BmҔ�$]���@T��}-�p$�B皂t[��3������U�o7����9\2���ET��u�/|TV��G� /FfEe:�Z�G���^��j�D�1AzC��d�8����h:Oei�⛂��J�8jh�w�Ꮠ�"��ևN��6*:��U�sʧHb���#�hHqu�D:�ץ�*���Ou"`�r����UZ�W����ؚ_�$A�	D��4쉜#����$���~�t��8wt�&���)�f�d6�>��8��B
}Ϣ�R0n� �W4 ҝ��W\�6�Fȹ����]��Jt rju�$�	>R���>Ur�5xd�N.̼�_ڤ
�U"����{��ae���m��� K�(�K�5
n[��խjz5I��\�
��w���X��n���4T����%���s�>ͫه�PB��cQ8�Ge�޳�>7|N�9��j�o�lm��t�b�ԇq�V���"T075J�joĭ"4��D�*��H���Q�ƗRZr��02Bd�Yj�����h����zH���[��eI���bK��Ţ��>�O[q{���|��(oњ�(v�T����՝�ND�j�9&�AD�����BS%�R����%U��T��[#W�6�)t ����검�X��L�]�IQ�Ω�8+����J�p$!�!�8�k6DdϾ;��fΕj���������Egͻ0��+܊!&!�1�Q��ɫ*� ��H+����Vs10 ��oCW/丂���[���{G��]~��B��q�[�*��6Zҍ�Cz��t�!��}��&M ��~����W ��r��Sq��j�w�#�5���nC�&�$W�f���jL�+(�j<J�9=�� |b�NV�IlPkQ�X�>���xП@���<T��6��T)�0B�rq{�����jN�do��-]nN�� ����%'m��~m�1�3b�i=s{��v�#J�VE�1�d{����
��~��)H	��2�B?ϝ��5,1���\�yG���2��ֺ��0�6ۙ���H�䦱�\r
�q�R�W��ѰT	kQ���]ΞӋ���`kn3�w��Nb�q� #�;�LM�LZ� WB�;���q�ËShlp �f�U�����jm��4)�@i�Ð��&Z����K M:?�6@Ë�#ҙ��Q3�Ƀݝ��N �FQ���� hH�=�B�PU�����}�~V�Vg�������|��E�
bKO��� D�Xnn�<F�����|g�3 4��B��4{@�����zxl���!�`��y���Hd@�Bd�¹g\<��Bl͚��⸁�w��~���4�%��0O��%g������ۖ��&���e�#h��f6�8Ո���X�U��2{Kun-���i����%�^��hƜ9�$��{���Qb��f�gow�?L����`��:��1c�NmQ$+X��Kh���r�e@Ӡ�ɯ��G���f�(��Lp�-��5�],k���Z��g�!�r{.L�v��=@�^F�?K���t�\�i5�a�]ṥ����$�O�Ԁ�[� ^6�����W+�4 >�'�T)�5�'Z� f�㣩D>�ڤ@�	���Y�i�Sj�Ꭸ��n�q���'D��|�Z^q�f~?�opha��#���2wp�\��.g>*�����x���#���=�;0�ݡ��p����Y��tN˃+r�K��8�iC��M��&��]t��=�Ӣ�#�\�"۫2kD�+��������l'!�r<�40Y��j�� e�HZ�G6�tă��

���'v��&�=�H;˯"�ν
f	��0q@IJh5�o�����o�~�u��T�!"��J1���hè�eu�`����5�*0�[����~��Up2[ķr�*����QSY˳솦�=��U}���R�ӳ*��oz�4�e�x^9e2&����^1[,���nmyko��{IeE�"�2��~!�
�������ľX��	�
�PY�*9�--.�������-0�)Pl}1	O K��xY�-2��6h�[KU�I��C�@ebDGV{��Nu�L��G�/�>x�bJ�Ēts�șӣ��u~HI{߹ϐR�+M>)ě@�woe!L�G�z0�"��}�t�u���i@k�^����B�ܔ�¼|^�fy��`BE#�-@�ݣv���ݩ0�R|-'���`顨�o$�vRV���8i�*r(�� W3,���9�kߊY>)��Xyv�c���8,7�Q�����a�oւ�	"*����3}�0M 8R2����Öf�q�"�o���O�o�höx�4����t�e����FQ����#4h�\�/�,�GC9�g��c_�v\��X�_�2�n �ǁ��`^���
�4��'�?}#�0Ne��h���2p{w/����k�k�%�_{r��3bd;�:�����-!�H���0����0�q+V&�{�nC+ G&�M��������V�w�'���%:r��F���aK��;�d]B��������6]ڂ=���4�]��	m�_�]^%w��=�ӑ�t�r6䯥�@
��c���Ϧ�x$�b;iP�1���v<�F,u���$��,T���@{G��Q��5����j�����j�H���"�Ӏ����}~ �Ҏ���}	h��`��KI��) \���(u-�ff-HJ0f��������-�P�1I�nn٪��:!V�y�g�G��f7���S�Aޅ�r�~G�̝8�����ݴ#L����L�$u���1���'�ĲR��)�߿�ݷ����>w�����?@�}VJ�4?��^�熪��~k�����X��|2<��F�[�$�ط���}^<
�܅�����`��V��.�ލ��)��?�趒pNW[�f=|0����aLN	5��q��9���j(M3&�c�W_W�E��s�Ѝ��#䬑柃��O��E�����(!�J=pq�1xit��4��������s����$/��D���C��)3 7���F��"�ב�kG}�р���c|�צ��"��5�X�у��aP�9,o���`p ˽`E�lſ�����s�Ǧ%y6:-���`i�����C��re��%��'����:8�Hc�7�|�ڇd/�}��<�[���'����s�ҵ0T���\4�-R9�?��e�
��Xf]���G�2�A�>�����Z_�#��"/�i\�o+�xD�wB�q����Ϲ?15݌=����m��M���c���r�Bt�_x������}�3F�O�M����B xz�,wog�M��#z�g_�,�nEI3���ٯP_Q;�^�%�wZ�Ea�G*o�,V�|�
xnؓ�������#��ƴ+��#�D�C�#���ǔ;N�n������ުXn�mw��[���CIɶ�'޺-G�oB�X�� _i`�"Rka��3ٕ �#�OL�#���+�Q*�dd�3��&4-����]���b�.��zߠ�,����iq�8U�|��j� M����� pR�G�y2N<6���\D����
zn�5#Qx�3=i�j���wp[^Ye�2�Ǌ6XN�>B��Y4!�iI���t��ɭ>X������QkR�]���a
}��c[Q?#���-7E�����t�Y�*.�{s*��]�IVf��Օ�� ���P�M"8Zt�ڲ�J���J��Y�'&���%D���N
]M���g�W53�4C�cQ��E�b<ύ�h¬�&ԟׁ�ŊI�A�H�>+���;%��9��Ռ�H�:����W��z�>�[5)���+��_6l�KI�� ��́�̋�D��I�UJ3�UW]�n��(a�g���a���TȐ�J�đ�#���,��%��|q'i5����Z�"�oO~�4#ŞP:/.�����y�<�n}%���}�MMz�7n�'����$s�lc�T�(H�\z�Rt1��'�P�C�F,yj����vͿ����������r��"v;,�FA���P�ɶ�T�+�d�1bk.�Pw4DO����!��y�����1'��T��A�u�4Ǧ�~^��=azݯ6�g���S�͊��N_�DPH�J
"��ve�æ�f }���혼Xc?��R��`v�aY
�t�J2�ɳ��^�t@t.�}��u��7)�� K�L��ع�1]��(����*�g��|�\��|Z̝��I�`
��"����p07Q����g��x����U�K5ĉ�y�]`���}��O̢e� $*Q���҇��S+ML�� �kn��s�[�{��W�	��ͦ���������b��� yTh���_x�/������1Ç�W&��Qܽ�� ��|��^{����|��y��q� S���DP봃 �i��l�a��J��	Mqk;L�
[��܁`�7�1������?|Rj���S�0o>Ui����q�Eib��� ���ɀR�-j�6�%�1RD�D�%��[Jq�G�uv��M�;�����o]�߿��t8t��F�!�-<�r=8�A��>���1h�i�b�V�5)Kr�Y6�Pf�3{{�B`�1͑��A�}��w\�w�a�a�4��ˈ�C�b��R�aB�ܔ)�4ղ!m����BLDP�����Ýg����5��7�09�Ɨ{��權Q�k}�kg ����r����]��]�'������^�$�;s��(�J"�;���P%�����U<k��6]���[�����LEl �����0-[($������~�^B4z�N0m�t���p��(���1�Sg����fX��T��
�ȈU� (Js�麋RS�ǣN|��|܏~Syp���!XK��K��;r	����G߳ƭ�}C�!&��8��3z��'P�%<�
�,�/�,��,p;��6/yB�n����8>�������(�8n�;�A�v	��j��5�����c�KlZA]{q$�<����g�!*E�:1�4^6ha��Ō@�V���Y�`�O�H\�c���-h��Kq��Jq;��]$xdH�ȁ-9H� L��3SO�z��l>��r�M�͊�p�t��ν�~����S+z3L;9`��q�$^b;��px?͚���08,�g$�T�t�0(RZ�����Վ���v)�W����>؁��P�`;��uΆ-\���EFE�y?���-h��@6R	a���u�c}�����@�XQ��Jfc,�mhAtߍ��9HX�F1L�	�)�c(�6T��J@�\���0�����W���L������L��N� ����	���X�eg���������޽̭�1�O��/�x>'�eE_���d�����5ךJX��d������e������<
�S����>�5�dX��ѨRi߽>�g��55����^�w��9iٖ���8(�|!^8�A���4�į�b[Uq#k:O�� �6��>��7�K*ɇ���s������W��$�Aa<.DQV��<��"W��q��I�G�r�4�%w��>��ܤ������ԫ����@�V~�=
&5�<-��3"36�5@�SY%��ݲ�$��J/m���8"Y8A����A�h��,��㤚�Zd��o�A���p�=��1M�Cd_��L���t?jWY�[6��DH����� K�{!g����w��Jd�w=�ɒmt�$Z�c���R�i��g�<��%�I<��Y��]�4��|��霤�e H�\��*NK>\;��)�GL�*��ߖ�K҈�1���Zmu�RX |&d�C��ڪQ=2���k�hހ2�C�Zv�'�P������y���:L\Q����=��j#ur�Wئ�?�'4T!��F%��<2S=?��i�z�
�E7��4���J8���ȃ���S�<�v�̞c��9&(��	!�V��T0�"���K��1%P6r9�����h��2�H��*2����}����#��k����Q��#����봪���ٌ�����( )�:���~�:��p�{��M�U�-3OD'�1�?��f$�^�3�j~�}W9��-�.]ԉ�N�/jF�͞/@btgH�I ������}����/�u���/"�aT���T�����G��>t�:5���c|K�^�)Ns��cp��5J�X��1A�:fV8g���h�@f��R]7�,���Y���X!��h� ���׮���#�[�q^��N�z%�ڦ�]��bJ�[�7?YӅ��j��F�{>J��&?�;3U:+��ʈ��xȧ��{�N�Ț��碊9G�,�E�Rt�!N� 1Y��)zPŋD��~Q�1�'ܜf��k+�ű�~��jt��ά����7!�B�����.2��:�
�a�i��}����jM���@D���r�l)��l�s��/�d�J;&��D�EYy��Ȕ�*���a��S�h�	����h@n�_>�Pg��m�1�����^����$����s�ܾ� ���>d���d9�,釿���0t��Ue�2Y8��g�pCV�: FYK'�x4s�7*b���|�C�lC�8y�t�y�z�Kv��/2���O��+�_K���,�Z��wFG//�Sb�3�5j	�*n<�L�k�=!�W[ �� Gku4P���Sr�Q���_aC��!��J�s��ڼI0f��F����fP=��E�W�q(�!ٶ�����A� X���q��_]�� By�����|xƲ�T �ޟzH��V��3ȧ���Bز?��k� wN��Ub���U\���Us��n�4a��7ӵn��h! p���S��<҅�$��S�JI1�.4 ֊�& r�B�F`�C�v�0��@-��3���:�Y�o��3��m+J���у�6�S՛�[�X�U9����k���G^�%H0]E���N|���R��a��q� *�aI�������������_�q�܈��?�a�4�P{�~�hT�^<6x�Ni��x�s)�SE� ����zP�c�>	�jA��p;�(��뮫s���m2�A}D4��&�:�S�������J�DJ��P�D'15����#9��-�g\�y<��9�1��{�Nfk̦��˰Voj��~W���}��K����F�@�|<��dI���S��;��P����ah�[��ES�/�S�dǪDL2��w�E:L�\e���&�<&���m&�&��松��b$�=�|Ѷ1l���(���BB^��큕1��%?-��y�W>��d��V��˭?��@�ZR-���a��w��u���D8#����uAԖ+#�lF@�(�&U�~�t�O�֤@�e���=q���e��Sg�0+P���A�m">�����\]cC��t��W�ή�do	}~�O�g�bh[���tz��O�e?Y�6�8�����T�Q�ݻ��)C��`��3��\BC�V�>0R��	꾀$=H�������IҊ7!4����e���2�$�%5C`B��[��}�����3\?��]�*�#���y�����}�G���NGVCq�Z��Z��\]}"�������Z@+S�����7�����­���lz��5J���P3T��p�5��t�0p?���?[٣�y���*��\b�r�:2w���i�UiF����W/���GO�8�#1�7n���@E�@9���t�a`QH�\66��0��"f~�g�K��Z:�E{G'�+ߺ	�����6�PXwQ�=ʾYN��Hn�;������;�&�Q�i�?����5oƇ� b�M'�*���gb�u?�Gj���b��'��/�q�,?�2$1a���$�ֆ��vM���cY�����(C��]��O��(���Q�f�ސ��L�Wؖ+��t��������:�K��·&CH�b��\ScN�3�L�;v�(����}@���ٳ�� �[�m@Z��%�i�@~� �/����/����C�q=�s�@��3qW���W죄𺳂HD"�\Z�Ҳ��0�'���A!.ȣ{�E�$�g�4LɊ��K����GSG�e��3/��eYm:k#�����5�����2�)-�nY�mNRz������)DS�S*������v����FFڎ�fs�?[cڒ���V�a��e�|�;F���p�W }�9;&�&�7��K@Jp0�H�Z�a��Y�m��s_T�l�$P�!�nb(��[4�����C����ip�N��Ug�vz����Q5IPQ�P�S��ƙ�x�Tg(��x���tk΋qȴW��֐MS����S��+��p��p�p�F-�}�c����S*�hH��1�R�&ls�7�u��M�2���F>��G��>���+\D���
x�U�V��{.!.�Đ=�Z�P�������]�=�`i�D��Na���.��g�������Sb3d� �����5׮���
�KR�n\Qz
[4B�S�H�u�_�
�h�M�Fc.�N��$ex��b�*���)����Y�oOL"p��.�
��;L�}�`��ښфE�ݳ��s6�_(�u�Č�����/�@�`�w��$��8ŭ���Y��t������m
�̓��Z#��|s/،�Yjn/�{��" y�xo�)|vh����
�-	C���7��R�[B��[��^d��f�!P<S	���H����XPB��Gjҳ�۹�p���'�WX�v�J��YL�Y�qPS��r�<໱$)2��ώ���!:m��ʮ\HP�ݐ4r����*�k��iw�w����`�z��lz�N���{��q���t����3��i��L.؝��ڙN?�1�L�� ,kΌg���y@���ޑ�� 0,?s!�C�f��ڋ~�{isf�B��L�!�o
o.sD�{Ba���l3�QJ6%ac���o�J	6YX4x>���& �DmGt�&�YW�X�}�rD��q�w��3)0��s�w)����E�GT���	)i���[�o�O�6���/4ws�$������b���1���L\ ����	U<�>� '>;���O��3�_<k��R⻍�c�� &��;	g�	~��7�L:<�ΑRN1Xeh����I�.�;%��F�d�$�`��!Bj��]�3D�p��|�o���79�q��h9K���� B2A������jA��&�mKh���]0�E����rJ8޸1F�py��=Gq&��1���l����(�U���zdb�kā	�)v�!��:���J�>�{�p��63������!��s�y�K4'�u��Ө��S���t���[Ch!�?�W1����jvkK�3�L�L4M2�V���qx�*�
d��/iB>�|��Q&�z#�ƳWڦT?�v�O�d�&���їO5ٟ�uB��� tu�l�OX�����An=|�3���� �/��f�c����O��w�dȳ���ص������M r֦��k"�誃��'+(�k�〯��<!��]�����c;u+�~�����w�"��Q�^*a��v�lc�d�	=���_�V]�fq�C�,$y̨\�V��:�sM�@��w�����,~do"���e��r^���gr�z��hI�eK�Ϻ�Q�hL�s�c�ko�8Ƥ�K�/��'璦q�m��F%��'P��׃3��)�-�'b!��\Ǣc/����A��*�n'��~��u�c�,�ۅ�(���
���%$c9��f
��G}���rX��)�6�	�߬�BD^K���~T>�/�L�D��Zo2��+J��+?��][,�5�Q������WBj=��<l?�V�;[$Bš5���ۃ��j����;NZ��!�[6lS����P�����p�<Һo�%���s`m�F
_�������	1gӈ+�Teyc4a.��j���E�RZ���Z�f�,_Bj3rn+BA��5����G> 6}�!�3~D0h��
K�wP�9��&�!���X��$�;*�e}�KK����)�B3θC+�{���/:�hG,	���V�Js�]67{�(T����U�4���z]������4u�$$c]��� s��M|{��Ó���J+�4a���V0�2H�@1�)��@�3�[ƒb��(�-�g��G�v	��'�hf�I�n%"u9Hdg��ܿV���˺l����F,?Բ<i����P"�) ��@ͼ=8��`�P�?�X<Y�R(gh�[y�F=�2���ݓ���w�rV���F��G�Ѭd䐏x_b���I�z��5�����q8Y��$��%E%���-�4�d"��Y��>s[�S�O��H?�G��ֿ{�C ��ݦ�8�廇�����ě]7�2Թ\~�Q�7.3�K�M�Sm���TB'kd0/�f�6�y�3�J�+�hu���f���+~�7�x�v:�]O�3��cm�3m�l�j���s����=���2:.�È�r�`�;�����h�A}[�!A��-�5�{��_��9}�d=&ơ�ॸ̰��2{���X+[- U\��c}C�x2�G��$�5*RFe- <u��M�r��L���;[�3j��K�t�2��}"�G�K�EBηO-$P�� �ݓ��NH���.��	�6&�bk�A�G�dK�\�U��	@:���d��s+K�}� !!�ǖ�H�5$w^@C��@���b�E�6���/���wC�!h���M�O�������� �MB)`��/���&I��#I�
D���nj��[2��!^l�#h�����k��imtyq�_��f���YҲ䙿	��LX-5�;�z���G��6�Z4�4	��[D��r*s��7lh,�6�;�ˎPr�Y:n�z��0��e	et��ǜ�g�v���U��N������\�%�ރ09_X2S��xc3~��:�.��o��U�i��%M2�ա���טxQ�2������eU����t|T���Fy�ӷ%w/ێWzGq�ZL[��8�m��vm�Mc�4��)Ge�	=rM�U�|�vT��m���Ia.��]�����~���1����t�L�3�zE�F����;�Io�V�|�<E9���'��s�A�e=�s*�Q���CC=w��j��&��@�Zv��-Ǣ�K���0ExJ�G�9W7��%I=�F$���)ؔģ��Ѫ��F(4�?��f
�r��*P�f��|�]�D�9·3Zz�0���Y8�{�R�3�#��JTC���x���Wnʜ��7/p����^;���[-�#Q�\�҃�}S���}�RGf�N�Ai!��p޽E���ɾ���ۂ;b�/�I�{���1�D�c�s�[���*POW��d�h�<b��im���s0}���������Z�PJ�x����XK|�ai3����J��5-�L��W#�N�Ϛ�����["�{�	���Rz�*)�(�����������W�	f[�dy'4��h���(��탇F��&�Йѷ�n�m{�$�:LLJf�� �:��W�;Pn��F�v���4�j���d7����J��*hNk�~Q�k͖o�Ǵa%0؎����巑��/8�	<Au��^�����Fz����׹�du�)���}#����P(���$�
"��<�v9��g�>5��na�g�[�g����id�sum/�(�d��P%�ޒ�p���A�|�� �V�B&,-&Ox�kZ�B8�BK�E�03�1�Eʖ��]�Uǒ09�\L����WF�u�x���[T'������j
�z��J�@�)؞�Y����4���$!5����N[�ٽ�
�w'�I���w��t�ͧѷ�w�w*�����+,��Q�f3�wS޵ҽ�������G����/RK�#V�;
�<f����PyJF�� �׸�]�ߌ�g=u����/D��r_b
��-��h�
 �X���s{U]���^ 
H��
��ܛ-��a8��5-W��'�}�
���ܤRO�a7�e2�R�R�Z�����}��J�ZX��M�!��臽�jD��G~��{D�_y_��_�ؼ���I�@_���Jt\����+W�R\P�� 6�ɥh�1��Cl�N�55V����Qn��Z��PV���\I��=��y�;]��A���97���V9O;�����y��٬�6��4��,궆KIaýzf�/�N��!Ҙ��(�[z%d7@�+M���*�H����\_c+trR1C�кݤ��C��'T��u�oª��n� �"�Ja�6pa���{$q��'����	KȄcLG��Uqz�OK�*��R��ţ���i��w���{����{Τ�|a�����l��)����Ƈ��]�l��?�"N�Om`
sI8ǒ�>�|�r�]I ̘����V:�pҹ��O�>EWa��H,5�M�N�,�3c])(���D!f�&8i��t��L]�~^}[kuY���e�C�qZ��Mvԙ��a��_t�(��|r��w���V�¦d��P������$��^��jZ��Y�{B��v!f4� ��l�yIQ����DwoӉ�YVmt͸Dv��r�0���o�{9�=��w�v���sf�.�mw,a�����o$䞶�����ww���������rc�0��rH���cb��
�^��'����BS�%�Ð8160 �� l�d<��2��34��fe����
X:"j����$t��.�����9���W ������R�ega}$Q��Ti��B��6�ü��@W���кyi����6�U�=���@�8�-Ř+3�A�{���o� Q`_f�w���}!^_`�.��h:G5ל�1*aR��dq1!�i�9$��aߩW2;�4�ɺ2je�f{X��*�c�z��Ϗ_����K:�fyO�&���̃&v��,�C��bD8.v*���v�~���K-�a:�P�$��/-�����u������4<�����<2�Ձ�}�Ɯ�$޴Աˏ�
����j�+)��eג�����?��(i������P[?Y#Ih�v� #?0Б�,�&����xb�=�:[�`^�R]�Ѹ�~�"���Ա�Hz���|8��}@
�\�g��T�}4?���w�7EϦH�
R�M}ĕ]8���}4�-����e��3�!Q�ne�^2��1��Z4s���d|{cd�%��vxS��K�OO�H���
��j}�O��J�1�<S�x&�
�-L�n��w-�@�����kvs]��Jd�a$nu�Y��v(���m��v��e5�f�ܕ�Y��g�H_�i�+G����L�fς�E˭:��S�x��m�I�λ�7v��)ɡD/�6a6+<#,ٚmݮ��&�x����.U��V�D�ܓI�aP���>fF�Y�et�n�S�F���v�T���
��K����u'�X�#����. �q����+,E���fۗr��kS-�=�����s�YԞ9w��KS�|�Z�P� ���S!:�a
��ES��^Q�CC��C}�#:�f�$����2��ԫy��
d�e|(R>��M/�\�.D����ʄQG�Ӏ���D���A��jhxqg�0�S�����t�x\۰�O7�Uc,�/@Y��1}�w�ߦ�u�y�n�����j�-��c��%di��S[E�2E\^z+o��ͼ�N�]hDC�ߢ1�������Z@T�h�%&�y��Z�N����@|I�ʪT杏�����U�1ڻ�/`J�C��J���],���FQ'�Ylz;��H��TU��k`)�ּ�	�[�b9�At��?u4�v���Hb�zT|��G�m֎�=�Y�y$]̟�;jKt|��5/9~?Sp�34�kw�ƻ�@t ����MV[X�1���8B�$�1"�n�b�G���nj҉��V�cRU����;#�&��)d��@����p�m���H*�͑�8Q�X4�B^�U����}���d� ��U7��MȬ����:'Sm!x�G���ѓ�X���[}����%����J�>!�N�
t��X��ϰ���(�B���)���J#�Фs	Wď���쨙�s��<չ*�zd�Bp�q�(�fI{�2��o���|��{mU�=�