��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*������j M����J����Cw&�u����Dg��>_�,��o��3�9=]�sn��5���A<�-��Y�,���AU�G���̻N�	�Ϩ�g�ϵ�w�Ω�k���R�9HO�o�u�(v�W�T�yVL �q^�Q�0/�����)1�cڵ�E
�W�D�t/�Ș���~x��R�X7�]0|��?ͭ�m׭��e��%\rN���H�i��8A(_�P��0];�ű
�0
�@�=�eH��j��闶�|���v��U�7��P�1(��M�[�d�Y)/�ΉQ����{��4kTj:䜶�ކ�+i��ֆ���u��OUgnJ�=��N�v�m�"�M�fe��7.?F��e�4���o�I�By�Db���.۩��-ņ�\7�L|�\��uQ�Jv��(�����yi*��C�:ϥ�u��D��S1�"n�ı��
k��-��i0;XkM.u�!�6��XR��Z+���J�)�lq��c�QS=��*�I�d�V\�b=�[��
. c���Z�%���
�"������P~���V�WAQ�?\d4
\V/E�?B�{��ҏ��J-�S�5�Tr�-<o*X�N��{�\�:	�3��hi�Hu�4q|�|�8��R$�R�� �wayw�Ē�:�p%t�;���Wه�-��8�ո��f%�uޠ2ø�����H�@<+�ҵW���Y��������H`ahN��Y����X��:;�M���Z���d'Ha�^���^y�hnO&�O�&��q
���X���'�R鶰�RQ�J�$W;���p�ps�KE�Ś��(����8��+�m��$�U�Ƈ�A��S��W2$v��Wg��y���2u�@-��]��>�݆q�j'�������LZ2$)Hz�J`k��n�ʡTH��KIe�?�\�+@%�3+L��������G�h������O\��`~���/�v�JD��9���-EFw�z\Oy�~M��.���*��&�|k������~k&�7�咭���<��i)��6{�U��[VuΦ4���d�2�@4�w,�R�����p�'��M��7�Y����A	�I0�1C�mR�19d@1��i��a{6�ݔ7��g!�߇�dao�}+���5n���m��-)��^�}� �B~��/�ɚ��̏&�|V�p�[�k���U-��(��f<D�w[����.�%��}��Z����J�?\Bu<>뮰���摒��%pv�QS�����x$(`�~��{�dc�)�Dv�Qn�=n������$�W6��=F���%�V>�)�F��bI6Q�2Y�Q�fX��T)&���~�ma��D޹�:O���C'�k���¦��1���d����\�l�&�-A1�E��Y��q`2���1wT�9T���G�>/����:2�����>^NG�Q��`�a#�Q0���6c�Zi���Aq�2,k4"���3ZW��x)?,j�[��
'���K�1C��*�`DDk���S��J�F{ΐ����0��h$����[Wu�tT)��s�;g�����N���|h�p�	l����H��#�;��j�[��8��\�J�@E�b����(�"�7UY���3����%���y6IC&�7h��m�A�6�|K���B��ѵ31����.�w��ԑ�`�#�:�kO|�Di�5'@�3��y���m�\f�|����E �ע�c/wƾ�ϑ1&��c >��o���@��gL�{(?���CZ�>�z�PL_K�w��]�u���|s|�Ƃ���M�H"3��X��ꬫ�P��/ ���lk��%�6�Q\6h}�.[s,Q����A�W�#�iэ�m�!�0�WO��,M����+Iz���?;%��_��A��VԘ>�F��}D�uW-f,�d�m��ju�B���p���f�F��5������x:=76Yty��C���-�����T���Zl�a��tbC"�
*A;�z��N@l��S�цg����\w �+��9����d�i��cf?�	�ڂ�S��5���L��4K8����^?�:T7�BK`��a�R����]_
�K,�0�)u� -!��IN>R@+�����*ih�
8��潱�r��ٲ���ؐ�1�g9�Nm���>�E
q�~�J�� !qS������+.>��ǹsY�W��J���AQhDf7�MI�X6�Y��\`h�݊�؋�v�B�#{Wo��R�H��罱�(��7��<��|R4�6P�>��ʏ�]h���[��&����ef��P��K��#��?���Hu�b Z��7Q��pKY�/x���� ���[l�������!=BS�c	���w"06N�G���.��bH���9`*i���}���y��[�q�u���@9:�A�F3iQa�r�V(<��_]���E�Vp�-q�,��}���zP�P�÷����V*�wtN+B�}��4�f؁*��*s�h�?f��f��D����
#N�f!���x���c���؃���ȑ�9���33X��_bgJ�����RW�%�b~�EM�֖�+仾q��v.!s�� @=��+�:z��P�Ǿu(緸�8�F�b0ȹ����@�����'�' 1�m=>��Z u�0SrE�	e	���H��,WpR=h@�?.8
��bJT�yRZ�j	h!�Lf�s5+��A���d(��8����4Ǖ`s�P�E3�-�\�����p�Nc��*�A��GZ��qY����"�k����������kd���L���QF-���\�Q�7����>�s�>B�y���h��'�8R�x��9!8*F���(���cH�C9�@��+ET�D8W�D_�)�͗�c1�Ơy����g��q�`��P�ԊmÐ
	KP�y�.�G�M I\����v�ڄ�����9�L���ᒘ��H����|%��J���w��]��?Z�"���$���2j3r���L����]\�+NM�U�T"�7�2$x5�(*ݥ�7�1]F��m��d���D�z돺����>ljb>x#�[@��\`9y���	���B���E�*����6Y�󏌏u َd|�[�����?RN6<	f�|"��s��x#��)Q��X�#$w�?����H�|#ʩ��WԩƲA: ��Y�{=�����h?��x�@�1�_ ��#����{��A�%|	��f26i��.�>� ��k�>pV��JJ �k�ݚ�������v�&"������55k��t�E@��אҼ�,�&�S�����鲎5Q�]��;t�z���i/��	�aS*�Ss O䯮��Kn(�����r��>ˉ�_X��?�1行~���9���;�x�jX{�=�b-H0����� BwxrT��>��o mػ�*��z��;(�UtZ ���}J{9�~���GпHr���fG�۬j	��V�c�HS �m�7�T�4G�g3���a#	���Z��{�����T� 8oU��I
���l�(�t�ӕ@{��Cu6e����ǵ�����7Yj�����Q��1X��Ov|� U�GS��>�n徵��u7��<�@z�9΂��	���Ǜ��M:Z�^�v!��(Wz�P֡H�&���6�f~ ��^{+xuc#�,~��QZ��m�|)0B�k��	x1���R���h$2���=�>�[A\�k��������*����)��ԡ�M�x�d��/c��Iz4�S�-wN,X���&��ۻ�6vx�q�>�Sj<�|�;���>� ����l�tUT���2���.����s�]�vPvB���{y&UE�I^�kόK��ܪ���{g�(�L�'����Q����*O���3`.u�e{"?�(E�O�7xM��0$�5�w���Q�>�h���A�\�dO�$��Q�ſƞ�5��vU�����7;v|ZQal�N�Y�����83`>�^Br��o/P;�\q%w/��b5�W�gP
�S�Oa-p������R&�gl�  g�G����{�����N�Geu��/�-�]�d����@$G4$�R.��������<�L�Xԯ�w\�<{�VX���K����j��;I�]zS1�zc�P��K��8��#�;�ύ��?q�{�ȫ/��7�۷�W��U�5��G2�F'm��, ���G�D��L��!B�L�25��uҸ63i�'"��������K�%��64s���g���'�
&_�oX�N��j��`�l-8z��k����H~;j7�}�2�� ��v��B��Iv�J��W���Y�a�%�
r$ yo �^��J+f	 J��>rp�]��ҽ���j���j��K��5vTmٽֱ=2�:�5�>C˪��׎��Z+����I��ت>�L"*�_��&o�����)�v"�=����ӏ�"]���������a�\g�Ĳrg�!�w�~��6��U����}��
��?���1���:���Ys�S��*[��fgVH��&�KTG��TF˪�L��|m5�q�"�-B�J��WQ�9���P^�Hb�����ֿ��4\�����O�d�l�#Ύ�ھ���dZ0�)���q�Ć)�D�>8lI�q���J��W2�������pg���0�	�&WVA�*^�BX�!Q��z��-�"C�� �2l��gxCt Oby�a
�u�ƙ0�t�U�C���mqq�
�I�����)<w2-�o���������~��V��v�l˚�/�6�Dq8V}_�w[:��c��O�v�7� _�g�\���XY�`N��m)�x� �a��M����0�Jj�7Q5�!2�H�k�fV�>ҩ`IP��gć��[��P���J�VW{���Xo&�o}rt9K�MM�X�B-n�4az��,�� �0m����[�]ܥ�����s�F��Ʋ�J�h1��1y��sߛ-1�U�*����}�ߖ��s������K:r���V����[������)�8�ēU�(w�IT�"�/������]2�P�q�ԟ�'��f=ݕ/�ʔ�lh��O"��M�d�C���c YI@*L�ތV'ۍ��'������Z[H<D��*��©�6%���Lꖅ�ncO��z�3=��h�)`��Q�F��7�8⾁q�φFKf��(���ꪌ�ف�F� H�����t����V��@߱��\c�m�2g�PI��6xx��q_�@ד����C}Q 	�A"Q7d�PD�u��킫5�����'��)l�.�|���^_����y\�o�lH)0}V8��u�c�)�ܱ���z��a}98��*���I�6��n[��(3oL򞯃\��Vo��M��K_�Ap���~IC˛�Ha]�u�!����q�k7A�y�]���5��[~��Z}
�}�F{�\'r�Ik�y��-�k�C4 ��z4��]�鉝Jz����f���F�nyVK<2�=�~�s9Jy�yػ�o;�^�>AƧ:�g>��JhZ:�i|b�̂�?�ro��4�!���k�(����6�M�T_(9�C��y�x^����8�:B�Fz������ɠ��r�%>�1.h"��hr�L3�_ƶ��L��eǓbc!2��)�T��m<t�Oi U�"��-���%=���Q�Ӫ1^�7g��������?b�]qVK�M�[3�x.I'���j�R��1�Ŵ=q���/��h.`��`b5o�8�~���R6��U��e|d�킴n�������+�.��= �y�`��|��FLDZ�����j�SQE[�g��\�Sl)C�W&�7M�9���^v�"�4��嚼�m�/L$)@d��Q�ʑv�=ﮛ\n�]���������x&6�ı]%A%�?�N ƃ-v��K�$�*8*�6�Սuf������iՀ�]�8*��8Fo����E��fX���߳KJ��X�������J�<p�t�d�IF)Q�
�����~�1ԣ�j��ó(�����(/hu�VPl�a���td��SOb�4����m9i���;|��]����é�K�;Ƶ�JF��aWN<q��q�r ��(�_���>Kf���9B������9������Y�CTɢ$9|���Y46<�f{�"7Z��V]�<FxER�5uc5�(.�Ir�V��=4��� �?���f]n���;Ԧ���q�87j��=�����]k&�ZO�Y�_ҹ�L�K�R�����/�����f1�׾-� �iW�gQ�Nƪ�L�9x�DV����&��HFw�j~��B���$pU��"t��t�<�h������7'v����TjX69�F=��
�*Vel\����m�p� �3�=l^��Ni��w�,��M�O~��Cξ��=�"���Ӈ�lX(�?X՞7��_w�.��o'�4ǧ<���~�ǀ�)�:d�h6g�i٬�^_���A�O@�Kt�㥤3�ss�џ����9�����^!k��m?J9���W��� �j|�O\���
:J�]M$í�*s���V��L�Bۭ6�O�Ր9O�֠�~v*�A�2p`��T�#���:��e�vEJuh�C5s����:����>���YY�\�l"��L�����<��ݗ��I��&NҘg�GU�D ���|��@����=�J�w�R�'�#mv�{o���=av�x��Q�g�64C�e���`���}�\#�RE����R% 	�g�y�M%e���#U�����2Wp����`���� �H	�,e�������b��aB$�^L�̭�L��w����{��A/i.4`�`Ea�")n�VxΚ��#(P�0��|�^�G�/7�1���Rf�;�"'��Fg�hH�DR�@��'�vBJ�c�'7D�7+X%kƄ
 �v��m,h�X�Ǿ��2����uxX:���S��9[�O�<%��2^�F�e㇟c�H��=,�Ku��H+ZL��`�m�'0���O Sx�֐�8ߗ�䔨%1��V�A��*���89��@����~p�;@�U`M
���į1�
���<�� �1u^�r��l+�;�I����!�_Z5�
$��V2�p����8"�)?�H>��o�Z0�s��擏��B迧Ič��u3�@�X�Ņ���ϓ�	��%�����I?d60���:D��|��2��С����Ky���[g��_����&� k�&<c��h#RJ�h\��\di�`M�0�ꙎR�����I�b�Y2�<":��~ԎIPF�p���0��h�͒Ր�v/�S5�`� Յ�*�I�g�N����u��K���$���v�^A��z���AJo�G�Y�7蜤�v9M4���6��I���,~�L�̧8T�q�T�)���T_���T�1���F�����/�\S�G���[���mI��� ���t�#]�Rjv�?PA1L��T��w>�;�����n�Hd֪	s�%�Ћ���o��]k�0�Q2��� 7��/����2*��|(Up�����#���`%QR��O|�Z�]ĳi�h������Xm�����Ua&��E���.�*�_	0!�0��䀴IbԖp�*c<��w��&Z��y^/s����*����:h>R䗒��O���� ��^�B&�e:�g��-0D���5�S5y��K��ozU�]F_�ٿ����B�~�_ZE6��T{�=�Ga�5Ł�Z�N��M�J�dQ���2��vvd��4��C�H�{S*F��h���1���>4�P0��|�N�O9�l�ʯA� �ul�*ސP^ �`�ta����D�{ռn�l������`q�(C:��s;��n	[����~�NK^w^SJ��툡�3�h�B	!n�����K\�ijG#�Ւϓ�&C�E��*Bya���(��;�߸v�Vǣ�o�d6ո��C�ɋ�.��� �i ���>���N�.�>�����ΜS�;�Ħ���M�c�g�Ӗ��Y��s>��W7�z��^���[B�:�!�<�3�h���r�����"