��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�J��"4�=�7(�T�JѺ�ő��,\��s���ӣ�F�؏7ޑ���L�v@`oT�8��y���3��8S"�f�a��Ib�Ñ`�I�� ���a�l���J/��)��H0oz�p�Z �AJ��G7�%~�!e�����Ws�̝�ql�#�C�h�ZAޏj�-Yn%�U@�U8(>��֧��|]����z�g�G0��0�Fw���:���vv���CX<Ė7�={ġv�VX�c��:&Kl���r�e8����� ̀�L\�� 1r`D=���y�/��?)�����x���%ƞ�Y�@FdB������`���O[�~ �aϺw���Q�2c�������ox��'��n�0ngGW����)��1ˠ���˧J��-�{b�H�����
�e��q�H(���^4��IC����� ��ɡ�@�wk
h�ɵ�
	�+<@�;{�i�p�����f��*�z'l�����
�0��"���gߍe����7�U�tF�}����"?e��%ߑ�UH[xr��5K�QZ��
C.a�m��i�b��UyX@��D�����F�K}��!����AQ�y-��6� ��4��V��U��bcc��E��d��V{�?��ܰ᠁�T�8o
1�FI� W�U�x�2��#�7�G����� ���J�݌�f���Zy����,'V��h�]C��F�,Q�P��18s�%�^�2���L�U�}~h��D�G����ct��x:0���n�1�߈ Tj�E���������O@o�>�G����E!!ew��r��{��h���0gڃt^�<P��t6�9�$���s�wOL�������\ ��$�[�����q+���费�p�-(m�'������Й���e/u>`Vltqs��RRg����*��z=�.�z�r�|�en��U^�l�!jۀ���:�U��1�E��&Ǔy�R���f_�c�E0P���蝼�s�ĝ��iZ��s���­���2�U3�e�-�
�,8��&6ڱMym��O�'lh��	������'~�uټ�R#|ɉ����^�L�M�a�WI��[��J�)�V���Х`7�|��(a�h�8��O���ݮ�2R*(�c�0�K���T�@�u���(��bm��o���'�~�grb�m=WB��H[է�2�:؁�����V�Ğs��`�HG�&�ڪ�Lu�&�(����Z�%�"Q���7V�4�7�m.�p6��O/�ܳ��$�5
����F��@@9���
ֹ-Q�dYd�WB��t��<-�<�%]�����P p'�����X!j��6y���';e�bg󃰗�k���fV�5�gD�=�Bf��o��Iu���1�Ń�
o��ɥ+xc u��Ըjf,���� 1,�9���(%GPZ��i�tnB�pFfX��an��s��Ed��_��U�el�������j_�~�ņ�D����x����p2`���w�*hP��c��et ��8r,08��/����ESj�	�B:��m�?��4ٵ�)�7�A�Ya=*֍oՍ$$���A%i���OsH&�fQ��׳�>���y
�R- ��L� ��5`Р�hZU>�Lz!w�b�؀A.�����4�D�M���$e��"��U�/��Fc6�����i|f~�r1�J���Ț�26�r������"�I�Ji�A��A���&lz�e����vy<&���&w�ȭ�&)kLcjs��p�Bw�{L�q��L�4��������lf�7H���2#��"��U�.��S^�3�|L��.��\���n*'�����+Bj�P�g]�wMm�c���O��cm�8lҤf�;���^�GA��Ѥ޻H6B�OKN�O��<�ݍ���Q��}z�*�t0��g]&�?.�౅�d�?�	���|0�{���[!v�;zb�:i��d�.I1K���C�x��4�G=�-����g������]�R7�_��eE�\P��y;�R[9�H�K�q����(_݁DQT�����Ϋ��P�rA��ĳ�OX��'���^-��R��y3���]i>wO;&d|�g�Q�?g�t��b_<Ns|�փ'�j�����j�Ϝ���A��f��sʫ�3��H, ��ܲ]k
4@��s¸���!ӁCP�g��S�M�lJm��!�~�i{{�<C���濇"�i���c��D�8��L��+ݏDC=x��t"��h,���
*��*̩kB���o%d"���s6k,��/@10����E���y��A������K �w�P��(�0x�|ܑl�%�������Fՠ�[Azɭc����,�O��0�v��P��[�ɬe<
 N���%)����$u��{Kޱ�i4S�5����=����c��ԋ$-�Dl-��hvJ��Q�<��n�6����/ѻbm��ٕ5������	2���|��� �A��lf�D���h�	�b��zV �z�!^����v���ۏ����&�To��1M ���Wr4 �7ۛ�X[yc�>g����,�:.��!e>7���u�B����2l a<�2����X��9��s���U�:N �虗���d!����tz���V�Cj��Tn�z��ԎQ	�M�N�(��@�x�ԡ",�$�&l�DSoT^���h���J����Z��٨�>�:v����S�q8'�;�J�����[���^��*V: \�|2��HInԣ_?H� �r/4�QLdQ�1q��ӌ{��P�9����H���u>��.\��b&<�=w7Ԏ ��
��ro�m{^u���|�/�r~�@B�ρ��<���7B9��<�mz�+?w~2
��Y��|;&I�]2bV{L	�1���P���q�SR����Hfbh�	�������������U�>��cXI��y�JV]���lw3q�q���Σ��^�Q������;� �i��xkFynk-��Nr����E��lQe�^s!z�1%.�y�*�8_Oc��J��wa'~�o�"�����v��D�8���Ηb:�G�$���æ���C�r��{�sӒ���?!�M{��(V��(��~SoO�^]�����(������-��f|�����q�=�sh��d�4��� b����v�eִqq$�p�!��>DOS�qz,�U����/��o��L�:N`�)G����ǌIƁ�3���WQ�Ȁ������$S9V��tq��O���qz��ޘ�B�$*�_�d�riǺ�d���hي::#����	&}2���RǕ�d�K]]�����e�F�vq�T���߃�*�X0.ÖA�=�)��[�ԕ�
������(�W�#��)�0�]uB%7?�QsJӧnZ��%�u��0� �u��x���G� �2��?p�|V�m���扵�PC3ƟQ��`n��m6�mD�E�ݻu>ь� 
^d���*H��Bv�K��|���� �:f�<�j�n-�Tt�C� ���?�Jh�X.�[8_I�(�FȤ�Đ��Ƞ�?pD&��33]}H��65�%��<)'ܟAl�]�.}V�2�b��r��� ��舺�ē�����Tԍ���īG��lN{�i;0��A[�_��z�@�u��DI䫤�u̓�&gY�U&Q.���<)� ol������E`N{-�w�)��+�S5')�������:�O���j	���?�;b;�nw�k3��6]]���zE6�
~�V��&����
�����	��ܑ���-)�-���bnS�נ-�n�I߀�S����^�S�щ�1��W���"�ˌ���h�O����~��bfj��&ޘ29֩um�S0��: C/'wEL`����K�S��A��!�b�|L�@�κg�r R�X��EЖefiҬ�խJ��em��*Y�*�à���[��g٫�6���ӎy�� �9?�-G�eC��t�U��sP؝�>|������V-HR����w:�����C�$�o�t�,��m5�~����Շ�L����r�2z�3���|K���{%t�PEκW����d/�w��8v,6ʦX��M�����7����~@��99����֧�P��InNХa��yw~0�L®�d��<B���T�{�rW��9�Xm�7�\��Mtj����KCP��|���=m�r5��Y��K��8�S~������m��Z�F�=�5�!��h���8N����s���IV�Z�I���[z5t��ɪ�j?��
p��k�k^^��-�ZBja��q#����9 �/��)�0�{؈g�5{�+ǝ �������fa�A��`�`�*�wp�����F�q4����۫4BoϞ�{��
�G�F�E��V4�KM;�A:�� |�6�ա�P�6�r��2��L�m��7�m�^B���+�+�)�P_�,��I�=P�Y��)�/��#��+���9־��϶��˩�^�q�k�P��'m��,S7�\��>�ZN�<᱕���F��t�7���-T�2o���C�6��5�C��Ss��2өK樴��Lg�HM����]�)�q��L����>o: /O��O�N?�ˉ�I��+
9��l�K��r���V, �ktɩ-�;-�gz^�V{mT��@E�Щ��^cP}3�=�� �?�؏،!1[G:�qҁE#7� U��Ң�IݸW���R�t(��)�0����lc���� 0�9DMڕ��i��c�n���E)?6x+;p��p��iV�9{�,Q�Z�H�Dt+�	f�[��6P��@�k��#6S��9�Y��!�����=/-l�P' �`ǀ��kR��d�1a&ޑTNQ�.'Y��>�����!�f�Q�=�=�-����#"�`�S8���
��� )��;6�zQ��xk���_̻a v�޲��n�y6�z���R�=A����������Ǘ�w�����9��2��m[0�$!�kw_�qyk�����6�W׎oE.A��� {��b�K�H�EwE�ƹ���T��n�Niˡ�V����0$ص���^{ZzB��ҟ���/W~|,��²�Mc�g�K���ܝp�pS3��SFY[�lo�8y�Y�;l���	�?�cV�ÛR�3CT���N�����
a���"�����
+C{�>��k�
�h�WU�7��r�	P�~��B���'nd�b��*J�u#G��)�(<59U%4��`�W�<ȵ�x�}�4�p�8����T�Ӟejҁ�̘PT�#��i8��Ȑ�T���]M2Xc�3��dEjQW�ãPׂ�����3i�Q�R��p�X*��L:�*��B�,]�/�ڨ_���)({�c@I� ; ��3&�y2[#�����&"*�{Yķ�xa6�XU������b�e��Q�b�&��!�\Q�"������2�W�"����ps`�����F�W�i�Nڼ���r��s�{@glM͘�*]��r5o���	����������$A�V<�\�Y�ɇ����_�E��MF\D�+���p�oxəch��s��I]�C5ԿY]����n��ߞ�
͆^�μ��TČ���#c�qj�eƙ.B��NG���>���so,s�a�6߼�/ɉ$�f3��߁��_h��2 �&퓺a0\'�U�S�Hs���3|���΋_��F�D`#*��l��G�g��>�@0[��}w�OF)�n��=;$('gGC3����=0��>�9�Sk���hp8=5l8a<P\�#m:�Ȅ�n�A�wN0���?�O�L|K�)�\^�>�d}v'_�B��%H�Ǩ	��\�Ec9ʚ���.��KH݅��ɖ�0�o��#�(�hmV��j��(���_4[�
I�iѸ���^�Gd]�vZ����g�����j�f�[e�1�R��n��t{}�?��PJ���lZP�"�ᆢ)畸�<iw��j�u�K>)o�z�5���ҵ
|��x=ľw��Q��.��}�O��Rd�D6��!p�uD
��.���wZ���hd�/�[ߣ/J#��D*���&!�����R���	X�W����H���q��~��;_��ʵ� 2��< .��>��������A��9$���?�8�yP�]��=~#&$������*N�v�~�����Ǹ�8�o�	�{�m�w"���l[�IOˈ*uP�J<Ǯ��煢`n��ؤ���;Q�ʔt�X	bE;],�����:N6js:HƯ�8�/2YFY�z��mrM��x�G)NUR�A���l��N���օ�@�4�!%_�Ɛ�_W,��#���X�g%w��$�Q
���v���՛8�O�������m��S<dv}�9O]#6�8Sk�����b�v�� F��i����U ��ˋM���(K��.�>�'����X�.��v���������W��ؐ9�=��y$���Z��ʃ�ݒx[f�[l��R��_�:��^��fzf�އ���n�ʿ��i�σ"�5d��4���Ѓ�n0�E܃S��N�+ū:�m�C�I�dg�g��I�L_{��\,�޸�5-]��f�X�?f����EO����G��,gpOn�%H򿛌��"4z�W�Yg&5�M���]��k8�)��%'�X�{�1�O��b�P��F7p�u7ԓ0�n�IGO5S*��-*�^���B��5[)��-�@�*J�ye�cSo�e+	kH�{��ٺm��� k7���B�܍�6� =ʗzJ9�'��γ�tY
��SJ��?�����k	�L+������<U*t��R�I�$���>_��Ia���o���Me�5u�YV0}qT
@�'��|1t2�����,h���y{�D�	琎�3`530�'��Z�n��bIF#����"��͙q��58�U�i�7�+N�>\Ϋ8%��V�3jlF��z��y��ф4��؃
��*�Ck�g���&LM(c'�+���`f-C.yDU��)E�
�f/���������dy"(����Zw(.mA�gP�@��z�[���4t�pr[2�����A̙�����~�;#S(�s����Hb��0�@?�3_*ߣ��n����ܪ)���_u�����w��U�j���(+�1�$��'�ђ���CR�xa���^��ڛ����!-&'����PL���΀��b�z->Yv�0�C�X��޼�	��f�[��a<s�UGb�+bJ��3�O,,���2�y#�Z�Oe/��YTo�J JXn��]g�DZ�M�A��2�hZ>�3�.%�j*�Ld� 3��"DG��?3
?2�T 	`԰���+,
�/�
!�D���JW}�N;��ý���u%��<�Y��-6Ntux�ܫ%�dA�ƴ�Ϳ���+��=>(�B��;�LS?H_r �i���Ny��?(h�IeO�=_,<��wa/"�)}���;&�-�%���A��٩҆����D`��ߢ�߲R��k([��O�oL�Y�l��	I��$_K�xl�������p�� 9njúJ��#Dۤ��G�	>'�Xό�,����-��%=Ҿ�0�R�@�z�R+�5���z�AJ
�eT	"��ww���i�̈�R��zi�y��D#�OpsHïu!����<P����Y�ǷF*l��%�si�FG����'��wIC�����T���(����t������.$��}���s�tW4~%�s5�ML��6*�|`�E~����vn+���1dA��
<�ꤍZ����ٰU���V=Ad�X�`��8��'��U��C5������К<�fKm�v�b�s=��]����	}�Y&��w�!|0�ğ;�O����.'���.��f��/���;��b�}���H<ȞJ�h�&Dy�0���|���k���ș}1��IrA��m��n���2��x�}f(^�u�x������R�ʑN���cT�W�=S����c��K,������ӻh�:��-��;�<m�mZ�N'`n��XƁ
,���0r�����"�VJ�ٰ��f�sE�P���p�w���,�n�`���b�2���C�S��KFp���PS^Nm��㄃��͚̂Mə��iw���w��v���']Ay��&��rj����:����άL8�\n��${�R��'��+P��ܟ�������<B)�(��L�!a�o"t)�~���t�ɄOJy�މ#�%��y�꜉��o��}ƙI��#;�
��>h��u�������B���d�RR�A3��& ^*��w�c������m�8���i��b�z�Ҋ!���B����~_[(:\�P�!J�>��+��e�1�t	"��R��J��x�H���+;: S�I�R6����^��z����B�@�D�w��j���~j2C���O�~=*Z/����=���8����Kd�|}f�w�!�Y�04�,�\\�kH�j����6�"����԰��26�t	�y�Q�-�@�����S� �#�G������ ?n�]f��F^�h��B����}=Sれ#3vr?��	��̞�S�ۀ�!񖲢�����8�)�1��Y���1+oo��ެ>��� "[�y�f�׳���F��2B�N> /*�o��4�S&Lvp$���`K��3��[���_V6
�
^�3Db7����HF2��]��Co~ԝ�ej�Ҧ9��r�J+�Uh�Aו5�Y1��w�(��B	�%���ҝʕ�6������c�H�U���(�7�"���Jey��W�,hS�Ih���qz]���e��e��I���'�|*��	��Z:�IH��Jp%u�t�5@5 �^�B���~(��(�s@?������|IL���~���~LL![�J!M�6Y����ֈ��^u�W!bzTp�^7�a�YC�c�4H�T��#�U�V(:I�g���B����ϻ#�5�#.L&}��7�B �a ��V�1N�Q�$��E�\͜B�׫�zM&�^���<1�?*���[��^�HL\��`���)6��*Kж��M`���d�K挒	�]aUzIᔃ�q��k���/��FG��߄8�b�r����i�KmJH�2������~�_8NǷ�G�]v*�:�H7��g\, �ۜ5��?K(�O�͛������������J�-�_����h���ԛ`W�q�O̳g��=ځØY��� ( ��d��ӷ*��h���?�N���m�6m��lT�E�12g�/���t����4��ڳ	ǟ��QK���%EKϝ�е�	�z�Bc�a@F9�%�@��;@�w-�l�0�,b�ߣqt�"��ݚ3�]fN /��ԅt�f��&������nY�|���a�Gi��s�1;L֝<!�t>O��WlT���}[O�b�fhv��k͉��f&�T�����Zs2��O�K��UM�|���ExJ8�mв�K/0�����R�6�e+�-(��_C4��+V�n=\!5S׹�xtr���G��'٥+�k��g �㑔 ��!]�9�1`��T2��]�����?\hKVTF�
��4O���̄Ʊ�8�,��ݳ��=_�l��R����C,�����J5XJ���[*�[�pI��BB+��%����!�C3�G�[Crb�w��a��I�T�Y����2 ����{>�K�}�	9�Ue���Ʒ��d��Qs.���\��[�s��N�������t��.�";7V�e�W����U�[�����R_>rqV�d�J�~��m{i�Ʋ�y���2p�lX�� r{vr�׊��,����R�th��{)���*w�\�����b�Zٞ6�)���#�N��>sr���@ΘCq� �S�EA�4�%�Y���ç?��Wm��/�����9����)�-h�Α�o�q��x��yu>qg� ���	EXX�0R9ܾ슮�9YQ�H�`�u�d�U�Słh��	�H]c�C��\no���tX.�#��p��'�åƖ��MK�=+�(���γ�G�Ϲ�%*���b�kŇ�x�r�wf�.Y�L�lA���H��y���{�K���
ʵ7��\�)Sr�6DI��O��G�x�G�A}2��^����5s��1m���>@��`��4���os��ݏ�w����{H�YE�$Q�ٰ��.�w��g��v/�s�U/���>�Y�GE���:E=Τ؄)Q�8���-�ฤGH|�gW 
+דD�$A8p����,,��s�c��6{�'��������.�U�X� �0�_��!<�z^ ���Q�|�(���۩�嗈&�[�ҳ������y�w�Z��ZI�dQ�
�H�[���G��'>�ʹ5ͮ���V�
�l��z*���䔴�l1��H�N6����9^�zUI%�zn'{��S�t1Ct��1�C?���;�}/4�7SC`�*9�L;���JQ43��&$/��*~)��f�z��kv�چ�y���]�J^��B���R�*9�SHa7c<��(Ͻ5<��I�3~��aA�6�	h�'Z7Q�X0�Q�B}"{G�zL�*���GL��2o��43\ȥ ���W�Õ:*���]��Bv�%Dp
�Tz��%�iQi���`wޭ�j��>G��Emۄ�����]����_I�5�9>J����E���~?=�f�J���Cnh�wϟ�h@�ـ�,�5+\���[��r��3Q�Gָ�33�k��O:�n�v���d�O��;pf���R��3���	tw ��w���]Y\f$���eځ=�o�������U���ĭ��H������HF�=��=�×�x�_Oy�z��F=j�&���{�4tM�^��0W�^�$��¡�_�!��������q��Qu�
�����5��}��l���&�m�r��d�ư�C��`�ڲ����>eze
mڗ��7�m�?g�s��</֠�,��*<�"?"��{�0��Iƹ�$P�8ۅI~�nPuȬ7ϫ�v��h��"����sT�� R��#�o�r���\5g�����n��
��o�'gT�M��KLȭ����P]�zld��Z�~�U��pi����m�fW�3\f-�����-O��k�q�46R�L�T���fV�Dl��
�Iؘ��+Pz�,_����oJ �{�D�1ן��n�lE����6�^��4*ť{�ɾ9�0���Gr���,qf~����5n����F��I'Z؎h���M4JA1�Sgv y@�ƹ��U�g6�RZ^�[����p�1��)*�SxI���*�ݽ��ܖHXu�۞��A�ߚހ���![k!�=�������w�Z��Ⱥ.O�%�.V��%P5z3��Z,?�WoiJ��Ü�,��n^+bUH����|ɠ-�B)�!��h�p�Q�_$��nH毺ч(�YE,��ݸ�:ODe?�����Wv� ��ff��_���G,Z�=�p�l�%n�+�H��:	ф�CU���������Mz;0�V�DcK�[�J�|ڟ�nW˛�G��B���X�ڋ�\.U���1`�8�����V.W�Uͽp��?�`������s���WY���E�_DE�	�#�q!"��T ]H�s��cN�7>��(���7�.%�����]<�L��c�1��J�Rm��,Rnw�п�N�6�4��|XoA�
^�wP��}IF>����G� :�CO&�?> =`���F	�ҹ�S�+B	0�����LZKXǯ�)G�R�d�ܰ�V���d�؋F���S�݊���YAճm��8%{6|�a1����BY���#������ҝ���x���-��&��Wo�$���#�H1Y��& k2�=}5��У��~�(� �I^b�h�A�6��K�эyO���3����_T�H��Z{�H�
u(��I�ŭ��#���c��Me�;���C�6u߼7(N�1���_ДaP����"6M��9v�|F���v��Y�������}�CZU�E�V���Kqډ<Ŗ�G�vfoqC��O^�Í�6OUB�I��KujRutX���.���(Lȡ��0�����
%���ic�=5��� he���l~;[�J�b�z�u_�8+�K��-�b����jT�F�k�uk@d5���#�n�%���e	M�W�;b%�x�Q/H޿`�w��	��kӱ��5Q�?x�"�7kz���k��j�_�^#+�	�&� s�S�|���3K�SsEp� ޲���v�U *�Bs/��R�.��h�@����VE=�9Y�[��5-	� ��:��w�05lP���:�������R&�ׅ��g�#��U��I�Z�� I���Sf=�hoz�[r+�BX�>�����\����vaټHP�����Z�x2LV?g�	����=���Y�\���aA�:}�un,��!AG[C��"�I������L�'����ۨ�|o�9v�h���H�_�C�����cH'$�҄�\
|)���A����c]bH�X����c�F�H�Q���d%�+2�k�+�E�'���@�]�$�ᙒ�F������94�!N{�~&�f�?�z�K��壬����T�LK��2@�%���5���X:m �9�]�P����R���y���Z�U��%����綇� tP�e#��na�N!H��|��1�Giz�7���]�i�{��ۢ�(��a�_�=_l!����'$�*/������v��!��Y�9n�hY�x�I94[4�9Of�t�Ib��������M۲I7l%�<��%��b��Yv����]n�#B��{��A��ߟ�tQ#4p�?vc�� {sِa�v�q �ɤ��8��D�l��"�YE��Q�j�VBLEr:�i%���Y��e�?��,2�W,LJLw��8��q	d�'A��6Y^�DöB���Rb$H��iZu�|�j>�����Ig�v0�3�j>�v�č��i������,:�
�ů>v�7��W�<`�AOo�SYR9��ݓ��|/�\n���P3w
+�s EK`�9d�ߪbW׵9�N�tQ��.��ʡ7���!�Ȝ��C~�.$��wCuV�Q����\;H �X�5��Ƨ�S$[x�Dѹ���eX��Y�z��Q�?�)� J��b�{f0.8�2J|�
	4E�q�t��O�sKIB��A����{���#�,mB{x���*�m��Ul�r�ǅJW������K�;
�����+�I��;{B��oԴ�l��<k�U<�zRk��'�^�����;�,�Dʻ�8�f��!4�n���
��̀�+���-B�~q�� {����a�
D�����}�?ߔfʗ�)�ak,�Q
������&.P�r��5�	�n���#C�Z�Ѩ�7}[�"��y��֟���)00�8�?l����>�u��wS�@�C/��^wY����<��eP�/��԰
���RCQ���2��,Y���Kড͝�f*�幕7'���`R���Z�t�V�2��{�Sx����C��ڵT@�)�6V�,�RH�$�����g���;xJ>�1�����s�c^��ъ}�֐�}�:~���>@3GLn1���N^۱Wh��?μ���{R��"O���]s\!>�O�5f��bq��T�~��l�C�A����S'h\���3��K������kJ��P�?���up9}.����v
�D���d�D��-# !�E�N2{��͏f�����=<?)�^��P}����OO3���i�:T�׈i�tʫ9������IP��9-n�$W��~��E�%��YW�%�Wfx�BU��6/�xͥD6� ��ұ�������e�6@l<�E>��ic�����lP��Ob��x��̦���@J�/�C�Lt�va����#�FU݌�=ZS	�M�&������N������pM,��2��+{�ۄ�b�m��ی�� ^w�I���eR )�]�;�<��&�����rg�w�e�M�2:UI����,ީ�ڎ��}�b �C� �1�)
��H=��������i���d�2�ЁO�&f*�x����A���0w���|�^ҝ��"���y�oL��j�V����rC�"�\����z;��P�\�)����䑶�a/�?���&Γ�5�!��)@$q=�Lh5�kf>�a������Fe��n��£��a)�r7����e�ܗ��y���@�A,���S�����hѢ�����
��JD)�4�%|�HxA��+T�p���i�$ <a�M~��psoS5qw��<��/��ɲ3+��u�v����H��Z��T���b�ݟVKhwTS��}jt�x���fH�u#`��T,c��`7bB��0A�>�P{�O�󻵦2_�[��z�@�w0L8w����i�) ����I�)5L�H��C�8�C�#ԏ����D��3C�������EyN�L'��S��%;4�J7o*ɞڲAl,����2��^,����@4�}̂[�9#�"Q�����Ϥ�aH�<P%��[ר�H+��Z@�)Z@Y�!�iL'�+ K�t��`	��u�����ȦM�rmG��q%��F��n���r^�NX������!����i�ͦ?���A�r=h1��BT��G����b$�sgW(�l��څבO�3ƞ��U���������T־���v2�Ҙ$&�&��1��]xE)�X�_s]���C�N����U�h����eI��!0�*�E�\-9����q�"��)���b�0&�B���#:��'���Su$��;wTo=�.$��@��+�
��Þ������r-��Y	����&p8�0�*ȟ����CR庵�#Ś��G=e�=x���9���� ����ޣhP�ځ��
*�ʟ_���l �[ߛg��	��uJ>*�:n`1�q���a�gvH����Ш�`����s���,�d{���em��c|� Mm	D�?6!^kt��m���7R?J$N�2~\����P��3���r���Z�]+S��ȵ��[h�M���lM��x9�<1�[�������� *oá~`B��|��⮺A��D�\M�?"�<��kmt��N 5vN�/L1�kL{�=FO�r��YE�w�B���+��7�ځKJ��m m�����_�� w�*��3�J�U���݇�f�ܫ�(�X/��*�8xq��C�f�k�Hņiս~C�~M�}V�KW�A��˳���Y�lb�f�a�nL%1ǂj�`:g�W�|V2m�G���}��Ѓu���|���F�ܘ�%_a��K����n��t�d�v����δ)�S{�MJR�>�*$�y��L��"�[#�h��2��^�K/ok.�TݸV��W�<�ï��%�p��J���R���ֶOP��
b�9v4�a�32�pD~�)ա^��¥�Q׿򲒤3T3^~719�E�QJfGV��0��,>��? �%��H14�;<�@Xh΀�C�|�(�9�\���{P����\ӡEǬ������o��6����|[�'��: bl�%!�Nz�0(|���%(���+Y���b�}(��aN�y^+凌��Bɾ�˧S���=h�3�/�adp��{�����L`�oF�&���Q2���>W����P+殣�y���8{	���h�&K�o�F�\�.���X��em��j���/i}��#����B�Oj�o'�{�W�G���K��Zo�tU�;qM:[�Qx��u����?/,�h�(��?�x>���M��7�Մ�p� /\������Uyj��\dp,��Z�� ~�Q�hĸ�j|ܘ~�ʪ�.���Rs�OpE˭S��7�w��b;�>��<�)L%�.�]�}��4 ���ȁ�8f���:f���D������!=a�]D��n2��>A�:g��U��U��: �
�V��a3�V,M9}�c)�}���do$Rոr������I��iH`���ob4�@����$I�~#S�94���ʘ�PB���S�&,=�R��C��җ��/���ь������<Yw�~�~�ِ�{�H����i5W����Z�)�qQ�h���lq������g�)ݰ]S�/����	���U�E�"] ��������|�a-��L6GfOM%TǊ!�h�rRSn�daN��Y�.�6���>�����v��1g�T�O� T?�ߴ�92\��7aB���΄]T�q��>BA�!U^Cֵ�?�jf[���C��w�sH��vo�+��#<��}"7����iFq�=Y�:�b>h���*X�ѩK>��A&'��.ˍXK\�H�f�m��9U(@V?��Õc�(��"ؼ����#{���7�����W��(o���/6*�X.�$��OntZ�D��E�M�ة�S��Ҟ	�����h����Q뚞Ə�˦PAw��	A噹��tc��+�����l>�ݐg�ٯ��bxP[��ੈG����$��B��eѱ�x�C��pz�䍗fqU^��z���z�j�D2�6p�D&[6I�u<
PjZ���	g�2�ka��|����Sp_P�oy�����pňL�������(݀c��=�bȣ��d���?�����"7�R�q����~�Vg��K靑J�-�&Yb��n���u���{�ݣ���z6����塍&TýKh��ƌ�i7�K���%he�;|K���k��?FM�g� Y��lKm�N\A��݋eZj�ȅ������>����_̰z|
8��Z�+c���*�z��2����N��X:2�/�)�/�(�Mv�&��S��4�����D%�}� � ���$q{=G�XV�n˔/�x�kn�>��<Ia9�v�Y��HG�45�]l$I�fά���GIeu.�Y�5�[��e��r#�@R��3.���y�DSΝ�xw}����T�bo@���c*��~�HJ�)�c�WXv����2)z_{<��+n^��0J�*L�Yl�&�;d��\ﭚ) Ē/�B�ju���y����T�'A�mp�%�����@ׅ�� ��d"�,t���(F����o��
����v�h�.3���;�q�Q��-�JvC�r���upؚ1L�H�S��_=�6ܪ�RD�R����Ad�F�.�|�h�eP
�u���-��a"� ���L�����Ŝ~������v�8̱�ȫ��@��[�g<�'#Y���k�y�P]f�vƮ��J���?�5<�p�#�2�CO<b�J6vg���<��Q������_���x�r�&!q�X��2O�T�S�X�,O*0����k(#Rh1��VX*�ա>�������_ǉľ�>�Ɯu�Pa���I�lɗ-{kz�g�K�6��"���[xIM�+ʎ̔�n�϶��U��~��;�ҁE��6��FW�nADk�]}��q4Fh�p����P���D�;q��F����� ��d��5���Z:2��Q=�"f���a��	IbGοp��O!'���1�݀�I���A��D��1j�g2`'�(��tǿ5\�R����k!�*dK�$<b��<���j�(hU�I��KM�T�@�!��T��àg�m�~m������#0_>⯲��Źɘ����W��b��m���E��4���A^�#��|	�C��p�q#p3���3�N-ٳ6$�iS*�T�K7l��*BFHj>�P�MM��^���Vm�'�����mgڋ����]��
(m3P(��G#u�x@�;��Bλ�}h+�Z�f�j�������ə��K� ���m	�|.E�7ݏ��5��8���X�퐩�fIl1�7n׊�-	�!�Tp�T.6&�Mp$=m���B3�վwW�%1��g��D�i�_��#����r���b����G��6Zh3K+X�k�}���P"��ɺ�|X�o�n>�t�pk���ߓ$��&W��n���q�XQi+�۱�P'��-d����z3�H�J�-l���#c�K�ˍ��ib��Ln�u�m�`�8ܲ|�6%�<Hz�{+.Nȸi	��'���pU������hMٕ? ��ʨ��"_����I��	��p� �0p�� m�þ�s�y�>&\��_��"���^sk�~߬-�BC�����4�M�Б�3�I�f��ҁi�K���t�nl��;�.�eDV�I��nC�8<4xmy�k=&��=X�f���1�ˤ�].���+a��c���畯�5Y�-ꜽ��H0�a��dz��#�q�|S_�:q��X�^g�����"#neV0�z�HJjg���L��:;b�����.�Br�a��gF��_�V�X��93x�>���TИ����
ov�q���ȯ�y���O��S�*�"uad�N �� 3활i�!�	1��:"��$\�L{2�5*���Y�݁ �A_��;�R+kt*i���%���X{����?����RfE6�,�(B��*!�b��V�ˌ	�"�4C��6+힅-3t+��(���]��qMa����lh�H�\��%f�fo|��w�e�wf���?v��^W��T��q����,�����9&`<���J�.�Q��18R����NB�T���*�#V
<��c������'cn�1�K���2j���>�H��kvhD�?t�R�{~@�y��Ɠ�Ԅyah��-qM@�tV��;���{@����i�(G깢��O66� (o`s��>��^$������C%��4��m&)�~�4jl���8�0��;k't��
$P�����O�
k��r�/J�e�=�9��C
w�{E�݀���.!�?=wyO�sOz\E�ˊ ?�$D����x���j�žaV�%�LM����^¡é����];]x�q}��8��9�+�TU����b�~���}|@�Ta�zHx�7�:J�Q_�������~Z� g���P�������8����"�:�(�@x$#YҰn�wL�)&$b�K洱�coB��P6`�É�A����$]��2������`�/Db��$��ٻ��>Z&Q�̴�P]��Ǧ�>n��mA��F����ݾ����ɠ�z���ө_g"�$ԡ���l&	��0�Qkh���Vj� Uk���3��H�ۿ���h�>��1�$�J�#�r���8W�Z9�	LB1����8<��9�w72����ŅB�8)x�v�LK0��'v���j]~f�ڒ�!,"���