��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ;l�Fv1�ϯq׆������s@���'����j����դ�P:�Cb�{�'�t�ɟ�>��(Hw-�u�� !i�^lZ��C�{��И���i�-|�|�I�Dd#����i��	�4�@$,d�������v=�3�A�pO�w�tE���M�ȼ{;��?4P:ٮ�7���F�ڦ� w0=L+=~�&P0q[��^�-\ߛw�T��e�z�"�[S��B=q��È��A7�D��]�!Tl�f�+K������<d��\�毙�����gpȷX[���;ފ@n�%%�WNr5��X�hqҶ�=PY�0��WΈ>��uX�+4 ʿ =�������5�i	��,�Hɴ���d��h�(P�pFtk_���'E.ݷ�T�q����l!�&˃S*��, �FȽ�'(�k���=J�?�>:̃�7�\���9����Px%[�C��a�d�%�}�qyh�!�ۍG��x�58��Θ�|l�zFSg�\j=)霃��f��L�U��!�@C(����U>�RRrT� ���X(�A�G���I?�/�I��"�?�Z��E�T�w>�3p�>����G�FJ`Eޑ^��&z9P4��,�N���*�
;�˰d~4�� ��'�L�͛�e��ث
|%��QLZ��s����9[S��ʝ��:W�7��������gG�^:�6���3=x;-��;
�
��_a���-�V�,+Z���N�69"|����a��tZ>�G�.�/�2�7]�Mg�S@~_m����7�ZҫӁ(�,�	2?���G\�^�����c,Sʴ� ���F�g�\OA6��-+���L�����**l�K��:H�\��B��r�A8��ѵ��1M jp��x���?S��p�k��ʷ8ώsr>!w�2�O���q'y,�g{"�b���ipD�L���#2d��!��K��VFha��_�
]{P���(���*8����N}��^�g������ݔ0��]���4��0�F���.tU;,O��w�c�u�>�/��8�cg$ ��Wx�h�G��m�l��S�0���~È�ԑ�,\ߗ��� #�J�!�Ѐ�u�	�h��� ���K�C���Y���BT��KLqÃ�p8��
�[��ь ��cبXK�#N�Jy�B����5ղT�E�N���s�N)�F�b�����V��?2�y���͏���C���COR-�Cd���U��U�~!�o���N��D6Ej>_�R&!�xUjAڕ�ذ�p�H�p�< gh��?%;�t�_���zm�&�.���a�o��n��$AJm��Ԟ>F"���K)m;�gPQZ2�3D���C�d������:S2
в;�P�~5�a��N�jR��Ff)X�^a+�(a*�I(��4: .y{� ���|����|�	?��m�σcgr%���{�L��+.�8z����7��|�)Aj�򄧃�*ٛ[��';������$��g]����6�鵏�hi���)�������;U$�೉�i�t�����!� ��$ ��`�R� �l�M�Uy�՝�U(�F~��:�_��p�Z�!��<�Ǝ0G7>*�tT�\«� U̡�l�8�wQ�S����1���8QOҕ�K]��W/eM{��~d��D�f�U߇V�Ռ?fpj�)ۚ��e�������uQ*�]�?��?~���f\z�-Ɉ�OR|z���>���ْA"����P�x}oz��ۘ+�w?�H �vv7S: ���}�e1\��Ƕ� 򳉱j+x��y<ڈ�u�%^Ϧ_/O+<��9rs��� ���Lk^� ~�����A⸝'e�L���T�M�5|�� X6���By��{�ׯ�:X}0�%J�W�2��� 7�?�gB-�t3p���w�y��.�=w#8�M������=p����ˋ����>�i�mzϓ
m�q�Z�N=X���W���-~�z��}���?�6(x�w�l��t1�����!'�;e����֙,lk@�(O&�C$1�q#�����Q��x�V`����0��jd0���V���"�qt���:!�Go��޴��q�s?͉��@�bjP/�tL���x���~�k��K@|^��x`2�`��'�T$<>^���fJc��å~��b�j�9R�$����w���ۆ�*#�9_p�+S�� 6q<�H�y#9�>��D��T<�
�|o�t�#�8��^)�����Q��]�Nz��.����u	���@��q�.��;�aq ���f@cN9�:v��q�u��$K�R����2'��(��m)�*�2�ǆ����x2�W,%:3-#t#��st�5��k��Nw��I�����<ae��wxk�q����V��]�0(J��ͧ��a�:��2I����	3k(ܯ���3��V`��
�?��cw�7�vꯧn�h�9�y&ߋ�'z��á��e[��E���Yʘ탊���T��U���~-
di���ʭ����V6޺�������W6�?��4*��Y?sj~A��8nm���F���E��nջ�cy���;�s{�O�"�v���43M�Sm�mK��V��������x�ܶb&n�H�	���q�b<Q�'�\t�&�(��v��\g�5�A?�ks�!q��a8�35��oa�ZR�aBM�A�$ꠁWa�����g����|d�Ɉ�6�-�G�,Ew</Jr�6�du�UL\:�M5����dX��]�h[K5^�����j�QU��k�a`���d�g�P���<@eIQgZ�[���	-�pߛ��70ā��j�S-���(Lh����`$��IP����3���h�#DN2R���Nn��8@X~��KlPHE��"�����Z8᜹� �ޛ��z@Ǖ�u�F�;"-X�^�oL��9Yső�(jP�B�TҠX���5�L���G���]��
�ǖV~�Bb8���ht��L�o�9e�ꗻ'�9�Ʌ��v���q�R���>`�4l����^��S��[Z�_�?��d�G��a�К�}��o��6��i�J�Ud��8�N���]~`�����"wTv$U�QKG���Ɩ�ޟ�_$���sKZHߧ/�^�bF�`�[ws�m�4�dA��}���4)�t�Ɵ+�R���x��fGLsXx��b��/���h�וu�}��n)� �X�,�Oо�
{L�#� ~o&`L�@d�p���v�2őM>WNxw[Ɣ�Ŷ�S4���"�Zj��|�� �K��x�� �X�a�6>��O���N���N魂/F4�S�������m�����vhe�apqWPK`�a	D\���+���/����`i����<L~����^�p�Qjyc��0���ud0��g't���p�/��X�ǚ�$\qڎz��=�e�i�)4LsX�y�D��!���?���R!сy��BP7r��Or��b��O��I�_����$c럊��H� ��u6��̍����!�x�=[�� ��`8<��?�:�o�hd
���� .�p��j����ѡ,D�ػ�s.(,�]d��-֔��J�y������8�O'|��E�2����A7//٣��dﮈ�#� 0�����:�i��"���qyC����:�O��0���u��\9���r�`�]Y����a�o�OQWג&�)O`.�]G`;/���v5b\���739���?D��~�qե���\qs_	ŉ��;�Y�V�P��]��I2jCId��2�x�K
�:Vگ�:��EM|�'�������([ �\S���Ԅq[E�<TE1�?Aa;9Ut�����x��93�=��7�0���*��k�5��vZ���-��	1��|6jg���{�B&_z}:�E��b�y�d�c��RQ��wX��7�)�*�A����N��;O�W���r���a�B�d�F4���^���4U�a�f�����C��<Ƥ5����X�D���	X�M�L��ֽ\���0t��8i��<��i�_$T|C	Wi�.U�/9)�Lɐ�٬b�%0忲�tPs����;���gۜ�x]kQ��n�&H�� ���y}<�2��3np��bث�
�TKf�i��;��� ��U\�B�]������F$k��7�5+��l�R��q�.�O	z1�.I<�U����z�Y��r�	���5��/����P`��.8������=Y\��C	��fQ��ZQ^��Y^��Ʊ����p2�>D��@e��׊�CQ�ͯ��P�^8F[
?��)��Z^�<��P:g�:ސ5]m=���ײquN������:�����ku5�bw&����U]�]@u�~�:v��lMJ7e��2��i��w�2 ��u<���v�:5����m�x�I]����=t�N��l��S��	q��^����@f��@�K�w"0��Li�J���d�Щi���,Q_��N�Y:��w�(��Ն�;�]0Cp�i��9�n�9ΘW1���d�s~�����C�sNH}k6��'Z���9+c$�Ӆj�� Ŋ���nb��g�dz��n�Y6������]�^.�S��%$(�?� B�H��G��P�<�*�Y�f�F֪iGNaq������7S��Xe<yI[����n�M��T��0y����SX�'��pb�e�W���GD�a�&]��'��|�H�J A�y`\�M�m��T3�|�xckצ4gY�"A`Z�80)o9M�=�����!�ٳ[Q�J��M�ǒ���U�۵np*a	3jҍs�8�؄kh�F0Z�-�w�A!���j֨$�u��q	
�P~�
<f�"]�[
��zh���}�}������8
��<!����ͷi�m=�]�j��Zׁ��j�R)^	7�r�>Zu��m7��]Clф�`|(`w�;G*v.f��S(�Kq*��$+�8𷫕�,��#y˓�Bh0��Yy�o$��q��0�:0촦a:a�Op씰Q�c�ibu�.'�I�~��t@n�m�W�ܑG�j��V��8����7Nw�j�b�R ��N�@a`F!�Ս���+��qŖA��Z����iL%>���#=��Q��葕U���+0!p�Ғ���|0"�n�@A6���jY*I^�OS�b>c�H��������$o8�ꊘ�pOlI�~�;0A[�}��F���}߶iPF*������`V����	��|�n�-���~>�d=�m0}#D��,y���/ GK�ǟU���B�Q�o!r�f�6/�O�� "�F�$�X=��U�
�q
T\�#j�@�
>���$��K��>��3�*yvFC�s �i����0��WW蹘�yfę��ʊu�A���Mq�V��ɏԛ�w�{;(v˺��.�q��b�Px�0�ԫ$4��]ݜ>k�<�$��a(N�va��lv�F"�$�@�7J=H�I9�+��~ب���u���Z}c��[XB	�y��Ն�xwfk8�J���'Eəe"яY�Q@�K��Am=�yf<���-,�7o��!����74K�<0�f�>*-XV��@�mO�T�U �����i�y�7��!� {U�0BxJ�;�����u'/����+p&2��H/�)�e�Ί�����u������^�&ޟ����iY����O%�Ɲf�9�g��J+����0e��p���wQ��PUM*ή�=?<Z�7�iI`��2|V���^����i�<싆˾�3(��0�O��_"�n1=�S�c�^���{��R�GU�9?`��r���}\f(��^ׯ�2ΎL���h> v;�-р�+~ݤ���a��'��k�`����!�.u�\�?{��+j�y/J2����&��n�S�l
`SM�}��[�6d�<\���@�����.��N� Kυ���Ǝ�MS�*���	���@����I���߽B��P��Z����u�UZ9U����]9)ĎN�M�|b O���8���jFY-�V���w�=������3�Frż�qH�v�{��?��C�m���ű.�7�u��p���h�J�Q�K3���r�6b��q�����\8e��嫊�~Z�H���W䵞���_s�w�_[��b[�.�o�J���RYX(����"UUA���٩��=��;�ޓ'��^��t�є�-7�w�<���u�6r��ח�m�H=��oi���DjP�'/�a߾���>���H��&@,��mjL��#�ˑ��?�i,$�N� Gt��N9�"$��s��̆(��W(��Ĥ��& 0_D�a��{��S,����ok�V!���x��g������hR�;E�[i�V�����LWF�E��3�@]�	KL�g�>ߦ;��~v�aX3��2����#��n�^�<XF�����;Җ}q#T��+X1LO���*~Z�T�t%���5ȯ(��"�G]�w�"\s�8�����_cS(�)���b�HJ��{�Q��Df&�5_���Ï�r[Z2V�H@n+@܀6�޲"��#���r8_�2}ϨZ��M�Tt�5�KI��8BxLׂ�É_gn�&�
 OT�Kn�ýf�_䏵�81,�ڥK��nˁ_'�o4��h˩(P���_��  �~qN%���_8��_7�+B�I-`���;�C
7��O�u8�x8��������򛒭�X(�����8/8� �4A�4'��%x`fݴ|�+���]L �*���_��>eq���<��,_@l�&�5a�iފh��Ri���x����,C.Z"��}�u�eRQ�̅5�`V� <��9Ypycc�n�wٻ��7V��ꏠ`��!QFゔ�ɪ����G��MF�m��������m�.�sAs'b,��e�E=�i|U��z}���<�Pb!��0G�y8�*!��Zەϳ�ۑ�+�=$[�#SO�OXk,!i?�4���}ZF_"&�D{mxَ;P�UǼ��.=��v��۪��7�yW��_� -�IʕyD|7�� $�9���},���		��+��x�#]���t��ke��ij(rk�	���yͣX�krH[���[��7�]�E*�c��f';�Sx�XOH�9�u��Y��ęЕ_���	��}�o�Gt�<T��˓ł�*n��k�z��N;�D��G�[�w��0C�M#2�4�m�ִ�x#uj�O_O����Ge��=�� �~� ̻T�-tf�u>;�c�e1��Uc�|�� ��)����̫�'��Ǩ��z�f�\k��	Y�� S^E�:�Qi�pT�/���|�9���c�V�ʽD������Z��d=c-���z׳��<(����ZG��������i������*��YظI��$Ì�����;JC`���Ǳ�S���td��e��v�:)�jM�R�(��u3{!�ךA�TAQخ��g�;�����$H\�|m����(�XG �b��Y�V�S��<�<<�2jP��N���{ ��"V�|Ӝ&�����ȵ�Qz�yt���6j=�,�vA�)og�;�?0pJ
����6s���m�H&9�Fz���k6�%}��k<m_�6�V�Fg����G}���)�w�ȺW�O�B?��`��' ?�N���s�M���&[�����޸&"��v���$�O�U8v�|*�&�^ot~$��/����K�]�<|j�VS~�V{��iV���h��6��������n�z�}����4�@�;3)/q���k�;����2޾q�%��䵯b��%�`	¤�j��I�۶D;ʓ��6M-�^�ʭMRï�ufԃ}��c��V�^�s���7�|�!�W�Q5R�uU���KO�;���kt�	�n�_��iJ'2��$��[�A�-'�O}������L��3�2�
yb���-���x+�N�B [� Y�+n�ͱ 1�=75���W�Ō��d�p�C>����󔿾��p
D�3���o�A�빚�1�~Vz�B��"���2�����G��#��k1���U�ɶȿ|J�gfx��:V���Jd�Z)�`h�_�9��!	1�d�UuӅw�������,,H�&�O~6�`�;����'�6s����<��%���)(�����>ϯ�j���:f߳�p�)�$Ƒ��=^���t>x�z�F���4Mm���.���Ј�uj�i`��a�tNS���4�<D^!�*����Y�o�}"��ۨ�c�X�^�@�^f!J�V����w��	���?b�!��o�T�z��d
B�����s�_4��G&��	�4��tŁ�,3��[ % �����r#ٓ���X��5lI��R��t�]��`֘3�3�Y���b���0�l���U�V�U�p��桼j`E����jt���k��6�
(��a�J�[L[���i�,
z�+�(�vj�$5	�}Z���2Oʻʪ֧�'ø��w��W=G_���29l�}w\u�9��)�9Oh@�|K际�{���dࢳz�V��bvL1�����j�Q��\��˃
+k�5��K����p
���� ��1�>�I�j�e���,��拡6��B5�>��)���������b����p��҃�z}��F�2��, �������*�/J��F�p������C�X�/@!�S���
�&F�>�޶2Nj��ϖ�3%~���'�a���(�����3�%v|�0bzCE�rO���#�m
�B��>�1̄���r��3Dx��&�Q��9���I�H�C=��J-``4��ɀ;E�;�����~j��C ��~
1d�Sҧ�V�p��j��Օi߄��J���d���R�J�2�w{®�v�ޙ�	���pO�%�� �Ƚ��I ��U�v�<x2N��@1�4�B^G�"`Vv[�K�DEd[���L��Q_w���"��zH��Vb�Π)�=R�O�vB�@�5������iAF^kC���_Z"X%D�c�<0�Y��^����#@�����/�1����}6B�z(�q="E{:�n��K&-��5M���P��xo6��+���|��*}���,�����s% �B;�-���'h���Y��BE��i�ɲ�.�0F���
ȯ}��{&���O ő��0m�pM����"���V���uO�����Š풂3�5,#�6�~��>mߔe��.�^H
�|ߺ� e �<+ݼ�z?����,�suVCN��i���Xb�_�}�e$`�bY8�#5$�w�b��<�~[5�N�ݜ^_�H-�@��0Q�}󁭍��Ewo~X)�V;�Y��l(N�������W��9,�����Z��w	�T���s�-?ޮMR��"/�C40���U�"/��[Vi'�����z�L,Td�v�b�Mә�9$�1���Q�{���3�p����lgG�SR0����_��&�>>*TԐS7O��:�J@�^Ӣթ~�/l�w:b�I���=�e����*O�?�De��&o�\d/G%�g�j:)�EK9 �Cv�G�D��mi)�K�}/�/V�nX��O���N��@�i��o�}jۼ�t��`/�e�tŔk�abR�#��,�[}����9*r^ZeUlRk`��I��f[D��óN�.����Y�6��0��=�s֨�%N���B�{����?�K���y��[C5O5%~"�f\ ��2Ep�|����Ҵ���i��	�*KHO��<��z9sk�jz��Y��le� �<!Z�Z*�Ge���9A�ǿ5#��(Nʧx��> ��-�h��׺{�����_��GP>��ns�R-��5�|��(������H�i2;�w���*v���p�)փt��n��s���~��c�ip�YURNB2a� ¼��j��%�ؤ�%!2�L�!��eK���M ��|��2�~�ѼY�I�I�����g�H��:���q��?�g�6��b�2K�"�h:����HQ�e.K�F=ɘ�dC@x �޹�3>L�ݹ�+/��n�?U����3�Ǘ��F2���y;��݌	��5>�4�E�����.wnYA����Z�B/�#(h��V4�������k\�L/f���\:�&�p���o�-si k������k:��QV������Pu\��_q$F=N>� $E��X���a�WY���5�����󎸵�ɚs����u�q��$Z-�щW�����f�ە�mW�.zz3�au��	S���.-������o�D�y�hXn�_�@����1s�@6�j�������Օ(gݛ����