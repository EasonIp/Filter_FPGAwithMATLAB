��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|����z=+���v������P!��:%G:�FiC�T��zn��K7x��8������pR7�F�'2�L�=����X�m��88��!��DP�X�˴�ELQO��]���״ܶ�d�{�,N8	"����8\Հ��M�42nzm�D��ˌ��2�*I��j��{�̀˼y��q�پ��¤x�oaL�x\(�9�P�o6�׻1I�Dy,Q21����(T2@(Tl���1��;��!�Kf��v$�S�Cn#ͣq�Ü׸�rkp�ᗓ��nN���Z	X�4_V�4pd�xQ�*5$QU�6�-����g��D��-s�{�C�j7���{�R��Xo$B����fŬ�$A�L+���7�H��*l*��'���ͧ?~E�|�.�8x����F��O�=V���ș4�*1�\���&Wc~��͘@O	*gI1��_Ct���.�!��1l��"r���A6t���i�[l�E�т����x��e��d����t3V���].�v ����ӊVs�8�/]oI��i�v������/f;�ԩuc�ҏ��p�����C�ɟ�tU��A��[�$��06u�y���=Pz��:.\�yg3/9����-9E�7�ê��ߺ�b�L������%�&sZ
M�!�,:Ǜj��Ǔ%���~���;�40�������V{�W7VI����[�[�{�U�Ƶ��b�wO�Jಋ���+�膒�r�6�`�D� 6�=6a�Dc��8�L�h5��@b(�o+|��� \�,{��|�^�@�) ����^@���YK�(�+���)�ew�*�4�1F
��꟠դ<a^��C`?�����9��h��ČH�@�1�Ez�5���/���q�l���s�a�CC�w)��ğ/�K{h��8��=��RB)��@9jH���U�PL�Laʻ�e1��nĜst �g���*D^�)|���k���H��ϫ�/\2l^�����ke���>�9Ѫ�_5�}�3X�)F�MF˶����M��?�6�@�4a��QVi)˖M��`sw-��g'QkrY�?
l8m?
��E�d�=�#QEv�j��c��o�����:I[��Չa����,u��PZ�m���ѩGE��Qp9O���?paH�Ŀjd�hE��Y�5�?)���jEQ]�z�6؆D��V�Ԥ�j�(��ᡥ0���W���ܮ�1��x�D���^jj@c�rK�}7
�/�B��}�&x*s�=,.-��t�J�V�Hre�������VӔ;c�f"(T:7{��.20���{d'�����o�Z|>��t'Lp���)�B$�Ѵ�e���:Ʌ��Q���]����ʝ���4��߳��vU���l�y��'�ɯ*z�h���z~���e�Kb�XW����z�t��R��Y��a9�QZ�w(E�|���MH���D�a"�c+�t�í]����2�~Ǚ7�h �n������Q8�w�9�.�9����z�8���ȝV�熣qٕ߾��*�V!�@3ygV�R�l�mھ	�(P~ִ�E0�?�%K��[�c���~㻺SE[9��\��s[U�t��j	��y��`v�w������#[E��cY��N2�|q}�M��X��a�u!U�Z:�.�y,d�ŗ�W�6�Y�*���`��)p��=p��S� J�|A*)aN���3i��9M�@]~����T���TH���P%�L�h�á��D�c�Ɋ��G9�qc���B��\�����Q	�]�Ό8����=V�$��ˑ�`o��4 G�G��ժ���K}��������t��ծ�t�e�	��fq���8^���pq��=
�L���#P�@��`N~[����v1��|��2Z(�XlU�P�D���,���׭�*+k��~�kGѓI*Lmڪ|9!oV�ܵ�ĸ��X�3���n��jpR��3�K��o�B�]���IE�K(S�%� ]@&jN`5�	�1LVEs	zJv`9��0Tu!��Z l �][�ILM���4Us1q/�S$�C>��?�^D��ytc�|L�$�@����5~�r�F��q��,���߫g	���Ѷ��� }��Ǧ��a[,����ll��vw� 
�@� �5�=�����qR��w,.��E��=���U����b��n�,�ZD>gN2�g�A���:���q��b�Q9A��j|w.�B�!!Z}����6v�=
=�VV	�.�e����M�p0�� ��Sp�N	�u!&�I�W��6�X�f�r�Nг��t5��=��F	�8�ӏ;�K8�E�� ��4�t�Z��;��GV�F��*}�
r�Ɂ* �	~���d�A�T�$�%�{Kl�rCy���ɳd�Ѷ��?�_�/�����*O"N`�6��83���(���;"	�u���}���*O��o��V4�� xeM9K"P_�c��L�%q�$�|���X�2��*;�.6�2~�;y�Y�r�����<D�Z��Y���;oH��@X��l�W��!zN;5�߬$dk�p͵�c��Ņ��꧑�$�z��NKȐ[_�)�7/�	R^g[֕�6�H���Z:�*ݥ���]a!gb�3�V_�N�8�}�,5w��o���u��p��1�(���k�n�b0�fn:���8o���U�h@$P[ƹ�9�vt������c�]R&��_�ʩ��L!���TO�,�}o�]1|/�$O�>+:�њ(��`m�$��{	8T�1�!����Cj^�i�,0����`��ߪ�0}IMm>�rX�e��	.׸�<X[��d��L������XU�T�@��:�+�n�z�B�V�[G���ȯ��ȣ�G<�1oJ^��U-Ͽ�K7��;oLF�"�a��
�in��K���v�
}%����ŏ��լx*�~&V�� �o��\�lU!�!�;6�T��YDm��^Q/��Vk5�ƏI�Zj%y6 ��ȻPMd`�J�#��*i	����B��[A_�H�I����8��gJU����	�fǽ�X���M�^����ʍ/-�Y�O��v���C�@�1 �en�����Dk"N��^�KuE.�nvA{*ج����� 0 TsAF��՘��2��h¶U�#�N2�)`^�F�7_h2C�³�@]�\s�h0��6�VE��yE�or-���`kQ�ț��bj2��an&�`9W�����*;N������RTT��[�,�ۢ�P�3�(�H��M�Nz��aJ������<{ݬ죱H ad�v�4�.�1�MRd<�wԵ�$@��#o6̲S��E�A�8��	��o�e�+�D��M�lM����=3�̀`w3�:�y�&���x��~��@��x�l}�����S�-6O�����x�?�[$��b��>�{0KМ�c5�'ԊjC���7a�]�)����%v��ĭ��+ ^��Zɠ\Jy��s�	�{[�0|�T���dFOb?�4q��P��B����y
͞jL-uJ�OhQ������zm�;v*֨+�N�f�eD�����U-��YJy0ȕ�Y��e��"՟����l�v���6�/�7e��m�JݵT��W�Fa�U�(:4�ȌU�'��75��