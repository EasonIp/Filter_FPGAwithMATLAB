��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$���ϵ�׸����^,�7���M���bn�b�o�{�Z���9�C�D과�ZB{���gP?P|��u췒W�m4�n��)�	��msO�@>����}���x1�,*>!�_�����<aG#vUr'��z��X�.�o�Lv�,+[
V�'����Y-'��5��z�5��K_������b�����c�O;��}�����b��Q��+Q��2BI2�Hne�p�Fv	?iVZL@I6�L�2f�^����Zx�\�EW�VN֩Hغk����j��3ב�;�/h����a�Z��Co��Nf�}>��K9���"���T]�,lD��qi8â��(!%go����=��-�F[����1@�%gA���5���4�Ц��/k:J�
MZ��͘��h8Й@���K"7�]@�V����7	�}�����}-��'hBJ;����g�X�;����!y�S���=1�w��Иߕ��;ѿ7��1����,'���0i�6\�`u�}�_z|��5�z����b�Ca���ќKy-�j���ن�3:-�6zxQ��N�+�����O��T��/ ���.Upe,����L쥂 ��b3��l蟙f�҇/��1(Fa�}#�d4h����*��v��ڶ�������̿s��.Gz��v�*���I�9��A�鄮A� ʓ���_Q������l:���?8$9WD4�z��D5�NrZ������ؓ�#-vRڳ&g{ۼTTh�V�� �Q�9X�қ���5�U��,�#h�,F^�i��26�uR�~���}/�ũ(�6t�>��K8Z� ��m��y����ő����n�;�����DncF�LN�,�#�H�[����<��<�v$eލ֌��ݪ�/��'U3j���*^���=d�&G$-��$�O$�# �!���-�fy
J&(5��}A�"��
���}E֡\�z���n*�'cԚD��W��v��E�<��˕����eX#���e���o|a�Ll�ܿ�� ����`�̍�ND[�W�4H Z��M��U�o��U��"Z�Ux�f���/'�@ES��D̆�H�u�o�t�V�->���mgk]Hb�K���eń�8��ˎ�1���ݮ���{����_&~��z)T���0�U�b���*��N��-,x���F�������j�ڠ���ew��3C��+JH��+�<�x>o�������.$?���4����t�f��z��b*p�z�α��c�w��l#�zn:C���h3��L���z��t��1)�ЈV)�Zl���j�Zߥ�#�5y��n�g��P(LҎĕ��� ��B��|���la�)�h/�(_�͋ȏ��?���^�C��Y�I�k%P�Cz�@yL�C;��G��p�}��ݕ+��LQ�o���\��@��w��~������o��L���7M��l2����{�/�cK �R�U_�w� B��70�J�6�#q����鯉��?0v'�%��s�[?�L���X�w=�Ѧ�wI3����fe?u^ro�Lѳ{�">���&�6�������VZ�u���B�	y{�@�[�d�)wl
�I�ґ�w�9�zЩ��1��"���;��K#����c�����L�#���Kjlv��^�af:�N��o��d�G�ݎ�H�v򗌄4Ģf�$��!c}$Ho�����#e�G�#lsR㿧SS�i���h� �䅮_d����3H�F�@���h����R� �W�2 ��N���b�i�����_����0ݿT3k��JV
��7�ngx�QbF�Ϧ�LU8��|�R����g���@�_�L���SF��O�����}!f���9,����G����ϱ��6c��`oX;�C���uf,�B.��w[+W��}������6���u������mBUNd�FZ�l�<��F��G��];Q������#���+Dm�l�q,���)z��o�7|	�cM`c�TD�����,`�/�"��{��W@;bY�{bه�r.E��z�:k+��y�"�Y$(�'���`��U��M�8�T�7��c��J���i=Ы�j23CĔ�.�Zp�*���P��a+�\�u{ ��
u�h�}�c%��2�#��l�X��a	�?�uْ= �T�<�q9#�� ���*j���'�� V��Q�TN�t�"�|������+��JBB{i#]��� ˸���PbM���V�G��ܮ��e�T�~�Ew�C\�
��Z�E�����cI���{�ʛ�����XL>���ӈ��v����M��j����QDg���X{��f!E�d�I~N2��=��x%�b�e�#�#d�� [�_���_�X�2��M�A)��O�&lJ����E>m���D[�Ʃ�<�MQ2�
�"e	���P@'�"�-W@�]��S	�~�͵���.�ȲD,G8�����Ep��[{��J<����v@1�e�rӻh� �W�?O�IH]>-5����?��1.r�;#���#�<�8�+��1z��������L����M��xӥ�t������?p��k С/qO��\���]���a/����>�;`l����8'qRj�f	wG1忸�I�7�~���Yi����T�Y������H����1�b]k�l*<�a�C�[|@�z����SPl| �ɦ�$���T�� �@}���c�p��ڮ�H��/�����P�a�>l'$4�6�`S��)'*�Q櫝Y����[���X�Q+���U���(�6����'��>�/f�1�cW�^US�Z���)bTg&������Ϥ֜�oDZD@�<��s]2�(�n=!0�4����x�ů�Dsݽ]����O�[dp��ba�ȘR��(�ģ�_ pz<C+`3:����X/�%D��OEt
[�v���[�%�X���/ݭv4���*����3r�紉YH��v����rk-(8祕"��¡��n{!C�����B�����҆��6=�g>�ւMT�^�A��ņǤ��&�>�:��\�&yn�;\[�������*>Zz������Y�_	����XWHط����mTн�M�|9����,�Rc��;-�G���1|(���4Ȼ��A4E��=��s�6;}A�I�9�I��,m��zDL��=�?��{�q��E#/��ٛX�`k�K�K����qn���]\���'�m�{ͧJ @�'��ʂi0�j}v�8��b����*�7���M@ԁ('jt�w��\E�NC�D̺|������z�{9�n"��I*uv�/������0��ϟ2��^b{>[W�褜ūd)D~����!�&��{/f�	����o��3[1zlYS��yyQ	������(�&��RfH�Y�;����g|`��v�3K�8�k�=l���d����P���_�l�`�Xɘ�}>*�˲ۍ�s{�T��I�����y���)�'d�1�������](��}�v^�FƉ�N����ؖ��6'�_�s����(ӵ��LZ�J�c��*�G�]E��[���}�/8Dh��p !��k4�©��]qG���z��L���nN��I����5��JC}��^�I�y{F�X[���`��ԝ�-����ߪ�_�΀���#�|�yEf��]:��\ogVCM����ޛ
?��`�lӒ�KϗZa�[�����Ɵ�~��r��rϹ^�F� ���ʆ���W�ǣ�{*�/iW0��fj6�&m�<�k[�]��Ղ��t�u$�׮�w:��Oy��qK�tq��R�:4\Bk!-(�]��ͥ��DS�;�m�P�9����o�P��rAN���)`ٔ�������1����R4]��0���J�k���B�Wq����w\H���ȗ��*�Η��p�K���]����pT��k|I/x]���ԵM��/>W�s"]T�8� uV*E��.=|wW��k��*}��Lڛ�t�&w]��֫�T�<���~�� K�Y��Z"�W��nz׊,����'�sX*�N����������_�ypA�~�,74�5 �M�L3�S-E�,���E�5�8�5���.������
u&	��^����PS�Vj�ݕ�,�
Ք}���?���'��|E��p,�ۆ+*��
\��bF�n�2�E�Ҳ
�*�f2�{A��