��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5��>h?I�D �Xe '�+�*P[�dJ�������ʷ�����*8�����v��	(��������=%T�s֪�������Z��a�� G��3Wn-L��l��f�s�ذf��*g�N��Ђ ���=�G���N�{�$5/������z8Ts�5$\�g���pa����b�1Gf�vj_��4�_�񾀔=�����]�4~0���(�������2���.�I�"��$��c�ӂG�CP`ѡ���n)y_|z�kf�r WI��d�j�b�14�{b@Tq���Y0��[��mK�hQU)`|)%Z�����2��S7�v��s>��L�����!ݪ� f������������NQ��P��ù��S�"&8�UL(N�:i�M���� v�?�_�_�.|���l~p4���{O��+�#��a�x)��I��b���/����E���DJ���q�㘯��%�	����T�x��:�S��I�4פD|��7�6�z��vg���z��p�&�/o���ҿ���'�D^l"�?t��<��)�g��B%9�\��s<��J�{VU����77\��?���O��w���s�z��H�)5aF9�\���#(�|}��!���デ�5
R�]1���а�EH<3��<j�����
X�ߐǥ�E{���7���"���H�DJ4T��Y��C�-�,���"g0Z�IV{�r� �M�r,m����pj�\�KH�wG���ˈq����;p�aͫ}(��@����C������4`�C6�坜Ź�!'S8�!/g�]|R˾�SG�G%��`������؃|Cۗ�<�}�q�x˱`���1)����"�r���ZA��ON��R$\V��Q��M�;jG�Jm�k����i�ڦ̔*��OB9g�:3p>/x�K|śJ��bq�Dt�KO9�S.��!�`h�f�w�\�S�}��~O���I5�*�-w���M#���Ru�|��Y(ޔ7�is��Z�:�X	�W�w-�O�'HRH��P��A������b��^h��-c��=���Y.0����̈́�,Ó���)���sL�j5�gw�0���%�G�K`>��l�����x!k�)�bg]�rS6�����[��a�����:o����2��)g*Z;M@�#h�r3�C|����D�ݗAQ������7ım|l����=��zU��i�Џ�d�6��wFe��F[���ϡ�D������m���P:�Gw�\�^'���	���"D�R%SثWz8y�Z{ ��<�/?�t��S�^����pUr��@�P�c���J����t�q%��|q]���� �}���P�
�	0[&�6�)���>э����GVo����7��H'���0¼��B��u��m��1*`����C`�(����,=�6r�Mb˺��~���ɯ��ݤ<s�I"6��R�_���1MXr�t������C�p��J�8��QCX�߼N���+2'r�㵹��B��$�%z��%:��@1�x�I���v-��������}$�bn���*:��g���'�$Q��Eڱ?^R�c�X�)i���l�����c��s����8���%��O�'5�0(���D���)|1E�|!ť���W�1�l����s����d`��)C�k#�gU�K?f�dެ��t����a��@����(��rԧ>|Q�Tr�9���k"�U�+ޞYU�b�����Uw;�|�P����LYO����txə���' �I����GGNk����S���EP��Q����U�Ox����m{�m!�x !޹;8���K�UhY*�!*���'���s��0\^���o
��K�5�ߤ��	�_�����2HBL
F���P)�c{A��ؕ�J�J#��:ʞ��(����k�E�V;�r�� ���T����2*��u��z7����[g�p��k?q�&�~�nRPоem�Z�"=^3�ia'�jЗ&�uӝ���E�^Sܭ@�Y���E�`�����m��'�=!Mzsv�3j`�`^d�|R�-ϨO�<��u),��G�Ɇj�8hnʨ���LΪ$�b`R�e�T
���ہ���;�T����h�8�{�o�{��'ti'�4�+q���U`N�*{!��0�$����Q��ɋ���ZO�8^��듏'xV�g��$E�n7���j��Y'������1��L�&(||s�O��'���º�l��{��^��eg��*$��g�t��.C�g -��Nߕ���.)�#⾖��l�Db����"�d��T�A�������v=MV��R�ô����Y�P1F�sP�g4�Ԗ �<�B�/��e�ʶO��4��+zk��?q��6��PY�\��uD(ܕ�-��v{j�vH���2esy�	c9E���Q��p�-�fjr�&l����E\�|��F_M�� ������S8j�qb>����r����X��s�&�&��'��s��0�z	Z�����9�I0mCH>�]B Ǆ�A��@;���l���_���1����E'{��q��eiX�w?�O����Ұ�xRSD�U���l ������B���?����z�i!$�.��<M	Y�B͘�z,f� 2J�����yl�zH!6"'�p���=	��:B�X�Ь���E֤-S��<�N8l[���${F� �+0'b�J<�]>EZV��7��ص� �#�t�?am��~��9|i<<�,I�r�D1�껦�&28W���N�P��m`�J���zc�~	� z��-�Pc�RT!̴6(���L|m���u,�
u8Rl}�OvT��O	�:"��Ҁ��絜GB�<�Qu�?��%��-n�0���\\3ʩ�{�s�(��e�<Z��!��Ӡ�a!A��b����"��`lc���&�ŻU���������X�X,*�g�l�������J����x�'�@�eq��E�/�f6"�&)>���J�oڒ��Q�)0!��Ⱥ	Sy�Ǹ�}�\���B�	;Jg>�����̢Ď ���t=��ɻ:e��x$�r���8!N�_вs��(�m 5�%(K⭀��~r!޼'����>-W̹���B*�`��1���#��#�6�b����7���S��.��Dfc�To�U.��?�t��),�!�Ʊ��P�E+ΪO+���o��M���|��c/�������P<ԝ�H�"�i�k(�w�\��π��`n��A���ƞ��b���b\��S��}�/��l~�?T�)弜ڄ�FI��X
TV>R�6�i����{�cJʛ�o��l;�!o�I;+�cl!���%�0� n�7�~?I�!<7S�������7�U%���fb���������O�8�f`���~���EuP��#�-��m��Qk'�_��M��`��+B�����GI-KD�ec���U1�
�##�^v�w�h�n� i kJ��|��{�\C��%�z�G��MG%����u���2�	�_1iV�&��ۘT�f��O�Ѷ<�pRT�i��8�vt-�d��JD�.P��Z&C\	J ���͝�lwJЩ0�4BbA��Rr�V�y�fd��4�ym�Y�4�]�&TEw�s��~,�}���m��y�I���D�����W��"ҥX;�}5����Y�����\���Zu�����)Doo�,�K<1v�����oR^�8��6��>�<ڄ]܋�����z8���#�U�
�g�YT��d�#�:�ǞW���F�-��*�sm:�?DgDa.Rr�p�m-���n[4g]r�F��9ճ#��/	3 GI��U�#�:�v�;�:�Z�(�h��NzfKFbE#�#<; �����oe��� >��S�Z�� ��ѿ�n�������L#x`F7Я׌T�u���7_	[;����~���h[�3�QE���XMt���~�/oy������=I.�V��j�0�-��֋���F�Y~n⊦$����_�sfH�A�з��.�h>xF8�,���O���H���m&�fB�`�$�����Ra�brnR�mo�{�W�?��+�S�Y��٥,I�v�����wϥ�?F��|������ͻO<���f���Va�(IV�@T�7�����������f|��J���~���������9F%f����ѳ7��Ԅ\V=aM�d��l"C(-%)���(��6.W�l[4&En�H�C{_�6��K��z��)�W���P����A��v����%�lu�l�&��~���H�;�� �bM7��P�GC�x�KET ��Gm�DXU��R��ֵ���9��H���]���Ou�E�h�m��_Zb�
[�M��e|k��u�+{�q�Yͮ琌�i%w%� ���O�c0�K�k����驪�[(�
2V"��x�V�u�︰�Vz�"d9�|�r*�HM��a �g����l�E`�����
x�����m���D�R��9�P�B+g= v�y�R�Ο_�v��@I@��
F��m�^��߯O1�h��&ŧZ���[���h�7�!�=�y�H�+Rk��͡|�ܴb� L��̇�*��-��o~�2�v+q�L��:�NrGX�x�e�K�U�Zء��^p4|���ԏH4����XY��I��4�����Ye1��eH�2o��L�#Qn�2��H��F��-+���L�蛕�[Y��~|k�+�uZ�z(�X1N]�V��7���&�"���R�C;\�tݎ�������-U`�� RX��l���uZ�!��BQF�����?�:���o�L�D`:�p��}~�������^n��i4�(���go��&z��\��)A�}#�'��%׬��@��B�M�%	F&A��1b��*���M$�U��$ܚ���b�[|�RӬ-��U��J6��-?`Wx��zT�fÑ���cP0�����z���'v���|Ư]����o�Irn��o����?����9�wz��[���*Er}u������.���0s:�}I+��%�1�zS�ю���Z��X������-%x�i'����8��z�gr����;��!�l@�����>�뻵�ŵ��j�'�����(��\����8"��s��U�!1��c���hZ�����\=�P,�M_ul��Nl�}:#Z��r�����[�/���m�1��z+�V�ZW��+�r%M)�i~%����!*T��F�0jtpm�ɧ�w��v�5=�A�]��w7������׮������=x�HKP[�Z�פRi��0o<H��4X���ԙƾ��\�yb��u�3U9���nǃ���}T.�ܴk�0>�G��a��� ,뮍���Q�>H�W%L�t�m�
,��^]�P��μ�c��1�-SZ(�$1X��>�]��E��z��X�lK��a������'�=F4�<�2���p��3#*"UM�߇�_)�J�M����y�#�ߝ�*T���k�(伉H5����u]���L��C0�G=����W�!wn�4Ӆ8���	;��{����{l����N!����DF[v!��6A�FK)l����<������6�����e��� �4>� C�/���0?U��D����f(J���??cWFEY�?i�� ���j��I�}��%�6��[#4������Ԉ\�H�h$�ћu*�g�|ÏG��躭��.�e�;|�D� =��!mEFXP�v�ǡ�����ރ�T�������սl�SP�X�+�*�=N�@T����H�-#�����7�v�C�r�G*Riz�m���6aU�o�&�?�Ԭb �;�U���^��"��V9X7���K��͞�gDy{e���)�ӣ��)OwN���U�(��{��]CU�,0�Q���0E�ACH�H�H�f�K�'���z���j	���ۄ{FU���$���@���l�8�b��j���-�28P�M������j2}#X�]z/S�,jϫ��ԶkR���q�ԓD[hҡ��V�ylz����X�	�a:22&�8A�q�+���^�m�P��n-h���W������M
��5�ش��hmmx�td ����
`���	Ѐ�~'r����W̒��}�C-��ց��S� 
�'�vd�C�˄�G.�a��C��nU�X3��zf�X⽝�;e�|9F|�_Wn��u�Չy$k�^!��� gᓀչ�V0�Z�?��[��+��+��4��X_�ଽ�
)>� ��¾�{ �ϑ
k*�v�(�m�t�<9Q�}7��m����/�L��[���/��z�;�I��qki��c,�^����e�Y>���E"�!f>|;P=��f��17��e&���#��J��`5��^���HN��ek�)Y�NE{*�$yW\��>���� E��nw�maT'Va�]��A>�^T�)�x=�7��j��̆[���Û����3��"
�x��R�2w]�Ȑ�f�iZC_-N����.��	�wl�1�0No�@����*�v�(���~��1��d���ϼ�ӻ����ܵ�u��I�[g7sxi�y�s�	��x.s^��?"t���4"��c��u���E�2���*��ztS�5E�����Pn �U������\r_B�� @M"�����
wͪm���Y-��cZ!��}Pn�����6F1����z�������:L{�s낽�{�#��6:]W�j��,i�XIt=#�	|*��R�5b�}|+�H��./�ֶ�t��@0���=DR��>�#�0�(@j�N:��Cq�������μh���^t�z+)�8�F�!���l�Q��!*IU���p6ǋ�t��=9�{I��E���@�4�;*�%4NC�'$�G���K�p��̻�J"����D�+.�#�R2�g<��}��)���6㍆B�~(ȥЖrт֠8�|�6xw���Y
�CvTn��$����ג~�-릚�J9��]HC����H7Q�x���*o)���p7g��$�pϬ���?�3� Z��θ��[���E�������LӾ��V�[%D�M�zc[/���r/1���ol�魟&��5�3���&�z�_.VSc'E�u��#���ı�T������@b��2X��ΐ��"g��Y��|��'������t�(��J�P,��O��;�Ԟ� ���2#�^&�mv��
�.�~����N>����J�{h�=��ݧԪF�YAD��]L����p�G���l2Bh�Y��n���;���B�e�!��-4�W�S�u|n�A>��QF�2S�?&��P3��]���x-�޺�$��/kZ�i�@N�=��:�q1�]r��q��2��*�b)t:lD�<	3�[ŧPG�T��z"���f
�_� �_�Ҭ ��o]W1w�K����.X[�w�$����IY�M�,�����{�(��%̍l]h���ɂջ0cgfWi�֔�����_�c3 un@��3%������j�>�1��e_"T�4�����6#e��)3	@禶ͷ5q)ݤ�=vo�e��x�-�G1�foK&���?���^�D�6C	���Y 2OI_<�6�3F���2���]��#���U+�������T�)r��YTX|����`�|ƴ��;~����u4��HG��͹�ڕ��!b�Ɓ�VP��-נFJ.槅�4/{������Ҹ����|�Y��J�x�ZC�6�t�l���-�w� ����b�@�<0��6��U�_$��Nv^�D�/�����!������˄4��,�ݧI �C����?2���t3�P0p�������lݥc�t}3vّ<���&��j��(3K�,O&�8�������{y�Z� ���o�+�*f$���JL�;Κ��	o���82�a�U�x�q8E ��C�=��oq Ս���� �ʣ#�d�6��k��k�v_~:T���T��.���P�8D�¼��&�?�ð�=�δ� ֱnGCNʺ�-'N��\lW� )#�*S�6"{	����,3���po]��?k��ul�@�̚EX�[�f�|�����ź��=h_4��(��nf��ū}�I7���;Zٌ���&�Ŋ�Z&s1�1�3�^V|j|(fF���2r%�ϻ�WT?#��1T���X�5�q�t)����O�rY�����|������e7��ߴ����>O* ��D�FC㦻�ͱC�Žqv�U:�6��ӱ[���W��	��ɿ�ix��, vj�B}�ㆯڣRQa��xT��ἥ��6?������p`W�����T�;�����d��n�<:U�
RV��Q5�R])��~�/5�GIl����&�|��.	:|�i�������RmJ$^�gI�4��U����l�^'��C�~~i>�cژ��Mvݗ��gJ�Q����D�)�w3�w�-Ϸi�j�`~0˞t�oI,�j1;k?�����z�]�\\�����М>�뷰\�v�6__�!�#kb4-}���H;��[y�+� �$ ��n~.�Z$I䢐M�t%SRiF��pEii��FX�����u�V� G�ވ£�@T�=wD�dRPS�� ���Q�M҆{�/G��.��KMyf��ϥ�+ʪl��m1���`.�BǤ^I���"��]��U�le�k'����&<��["�'�j�g����(��m�n��݆��k�K�r+T@-�_jE�߶�Ά�B�}#N�;/�s%6O(�M�<�D[�%����
q��(q�F�*:dH��/O��r<MX����N�03c�7�I��4L/[;Rެ�桪w�r�G�-V��ݵUǌ>P��ɪO���F>�e� .f�6��i.\C������Е���x}*��H��G��nT�ض�-r�DF)�5���hJ	,�`f95h�P^�Io� ��^,x�����ı�,��� 7kD3no�&�� e�������#e���軣ֽ(@��5��R\��)?�C)LJ������Y�jUC��Y��}C
��O��� ?��pj��!}�S$�<k�����!��L�p���w� ����c������T�' �g��2=�Ti���5��^�2S��X�s)�ۀK<J���1�X���G*�>Ɲ52��l~��q�ƛ�r��r�<����q.��
i�έ8烫2@F����<UP�FB� M�,�&�����z��R��b��9����������U Ѻhqm`�����Lu냪A�y.'��`lP���H��[6ݵԢ��uy�z�"�rFJy��A�3�2�!���$���F��?65�֓>,�����r+�v09�?x�2�:j����%O(�g?����S�<^6[�쵣(�����6e�� $�#JS^��n��NKˀ�:�k��6�xż=�8�L��K�Vǫ�A���c?��I*��JF^��9�dȧ�:��3�>!��
��prF��!D]m�{P�nʱ����ҹU%�8�{㯬*�y���drg����\o�(������-�V�3� �S.��cZ�
{"���ӈ5���Ϸ:���~�a�� ��;cԝFE,a��ID_@ۘ�dD�?*>)�m�:i�����#r�KM��_�U��\���w�d�e��J�hs��SaJ;�mCw	��RL��0�K�P�8q�%e��1�`oV񥷡���C���k�W�`MR/,�A�N��.��ٞ��\���
P�,!�����>��+t�lDp$����B@�����^�T)�<%5 ŮC�sll9�}���#���b�yǳ��Xp�	�-%���8m(���>�,N���o5��s<���HK�䌕?+~��ՊEbl6#�=����pH�1o�-��@����,�.V�G�g�@���Q?2��^c#9]c(�
�)��{ˣvt������aK�t$��
�m��0��f�](��~lc�E<
Iu��s^�@��	,�y���1�7���m|��i�&����	nƱ)-�F3��"`	�P����a�准��G�����p��8	^ {ό����e���e&Γ�� ���;Pz�?�G�����F���uoA��eW�>%N�v���A\�~�Y`q����^��-�N�_����j�vI�o͑�|���կWr�X	� \J�$��2����\k�
y���)v������_���b!_����f������;[�ᱰ���IA]�߬�X��Cc_*����I�&�[�?�\Z�_�b��Zt���i,�&�6���C	-�ܠ�t�P+G�|��c	$����QzL�F�����*����l�C���f��M�<��-�\YFn[IB�����`D�8V)�dW���mfr�i_s���v�q}B�>Љ�Yb��i�ڋ.�Y�
B�M�<�0�������M�[)ӛ*M"�nO�Q�S�H�x��BM������#�9���7p�x���ð���]�x#[1m;���BIߏ����6dʡ�^���t*Ίo����{�[J$��ضT�A��p�k�O@XN�]'�)nE|,�\�g��*�>�5=�K��8����|�0"-���-�4l�.�y7ƾ���8p8����H�1�f ����?^d�+Ҵ��K�W�u#����ƃ���z�U��-n�g�y��L`$������Wc�����G���Ā(��/����ָM&���-2��G+-��k%�c�,�5B�D�#+�ڝ�a;�u��eȃ��aq�p�⛵�J6�����]����O�^Ma��P{WZ/�!Rw\�/Q�0g{Y����N���e�)(6߹@ͷl�\Y��4�eV�ǿ����w��?W����4d�Tը҆�{��	}�˧�^(�P���ܛ�r���l���`�@՟HJ(�B�	�4�/T�jM*�0�pv���p'Ie�-W��D�� KR�,hjK���khjd�P������U�Y�C��u�cҠL(��L�/�սlovö��ؾ��qv#[&]M�}O.�`�شM��;�6�1\ �ǟ4�.<�q�;�ԥ~G"���ܴ���	i�3���J����((� ��/��ŇO�-�v-�i}��µ�M3S�ۭ�%�M��ځ���c�S���l�{Qt*��0�9)a�J�J�B�wW ��n���8�:}* �@�,`;���F�?�B�P{�gɠ�H�~v����Q���vh]���v�]������w����g�7��nGQQi�_��>�KWQ�X���$�Z��V�(t�qƁR�4��鉔���֏ Á��ț�N�U�b?^�YA����4�������	G/X���;�MAjI�d�:F��3���y0��I���c�N�p��n�W�{^)c��k�Q�٨�|#f-qz�t63ɠ���i�<\�������6꣎�N�&1�l�Θ� ��xrk!�\{�Ɏ*��D:|�,v:W������$��	#d�}�$x�R�  %��f����I�"�e�b���k݄��_��r��İn���L�3�.�'�7e����Du$���>.5^xO�D�~O�#-�ٿ[s4�=���+
�e��������%m1�|�a!�]">1�}��r��\���,�2	oh�����Q+�B�ݩĈĽ� ��2�r�k�Y;4e�{��69pIY;�wc�]�������&u�y������Wm<�?�����+���xB��XDH2O��X�B��'b=�Znۓ�x�PJ!,pL+���u��q�A��}|v#�.�H�.0��n��.
N���e�$ɹ�]8[צL�D�@�v��v=3�{]�w�]=�5?r���|{��HhZZ�;*�VG���TBy�2��"L�oL�r�&%��q[�n�i��v����߇ĝZG�dٌ��f[�?����a��E�$�n��0v����?WDB���7Ǎ�"��9�I(�oAeg`XJ��Ń"ܹBaHcЍ���h����>�����y�{�i��ޕ
������������M{�qN�/�\Z�M^����^���_���n��N��[�D` uGm�K��%�N|�6+&S]�L��̃Fw�9˄�1��Rҽތ�	�G�W�l�K$�tv�Vx0���g�8������r�� *z�a��86l�4�8���{�2Na�8���$�qY������o��P4��Q��t�����L0�š6	gJ.��uz�����+-�K9},�^��+�C��?��>n�FY���g�}��kMS��s�V����Rʠ��rԶj*/g/�%�sK�X����\���(V��ߦ��&������[V�Rvf�|�t[���̺���õ�a�m�ʫZD=8���Yn�?���}m�ZdW��i���5�^�śB��B��!D}Y��g���Rp��`�O�2K%����;u��L�f��{���*":��$�Ӛ>l3����"�d)��ڿ����w��l���.��<%��g��nX�J��3P\������k�Cbc7$�,T�E|�<FX��4�)pt]$.�@�U'�a��.�v�~K������:��(��庘��(�U���vH�W0��z;
j�J��<שLos�`�3h
ѻ̎�䜫�Y0Q?��{��vJd�6C_Ҫ�0��{�����(�P���I�w,�.~�	gX�l��1����GwkJ���y�X�����_°���zd�	�ҡSd竬^�ݛ�͊�#,�G���7lI*��p� �!�
0��Ѝ���i�M����13�����7r�%�~����jA������?��H����u=n�o�(z1�U��T��N�2���m�L@���{�,�M=iˇ����4�]���4@�v5M�E�
<o�(�(a�m���em���R����ϥ��S����?��wN�p�GX��_�yʇ=��ߩ�,�d:�5f�5+�,x=փ[��d���&yA��Oz�	pa���$-�"N��j����`������LY�0r2�c~�V94����Q%13?X��1Ъ��i�E��,�͑�\�H0������'&���%�KPX�O�}�y�����}'�DRt�/�1�=.,���r��J�恦�|�'T�K��F�W���a��ˀ�*��Q��e*l�83�>@��g�H<������d�ǲڍ��k}�v�
Cw��~V&��]����Tl�BQÂ�F�텾@6�]�V�!�� �K(�/ �����g�V�V�Y)6������&\��BM�E��&,0��I"Fmv���q�֬�^%�H9?�P�)����-�x�8��v�Ȫ^C�_*�R�ba�r5F]��� ��Lk6����'d�s�z�K�3��H.��N%�O@���D��J�L�;�o��+��x�4����U��vl<�m
��g�
�������^�9��	(��� �Yz�g4&s�Vz��v>M�.%5Ҷ<���*����xN&@�r��q���4��`��_.�w`4(�y��եj
ȏ0Z�!	�q��ĸ��۱)��	��\0U���O�x�E,��.��$TѥѰ�'J<rU}�O�(]_�ϣ/��� �BO��۪�*0�#���XM#�m��UA�.�0�:v~b��#�%��Ke���Y[���1�D�%���;9h{~��v�"O�E���N��,���vH�V�#1���}���.Qѷn��-�66�i���ƌ+Y�k~%��m(�B