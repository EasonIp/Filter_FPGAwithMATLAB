��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z��[5�j'1�6$�e���#N?t/y�(*.��#ie�8w�{vK�"��%�F���s��ɰ|b�3�U��@r����@�Z��d<No4��#ѩ"{wY��h�m0��T���K��jش�Y�>г`=,��1��&�=��Y>����S��/֡t��J�R��U��;�i�f���4�J�غ�4t��>�BNbX��;~��]�ޓ-&��7���FN��(w�sj�;��iY{�5�%�ۻE�c�RQ*�����+��zLI��w�	$���V7B6^�tW<q�
�ݐ,��.�LY�f�{W��r�}O���|���;�Kp!��5E{��<]:S Y}�Į��J�_E�k��Q.��̊]�Qh��B�@���@oro�7��ؿ8�׬�%�T�0T���<�>����1fP�s�~�5HՎt��Ef�Z7��į��K�&[��k�^�T���)�8<ԡj&��hK��B.��������H�r�������J��s���}�,���g��!����`i���O Hce��1������T�ɌX�Ӆ���k$ij���*��2){2d	���i`*�򪆈e�OCj��@�N#� �x
���\B�>yq��L?�ro�e���oI���?��j~���5��ia3J��b����.��H
�i�Ƣ�TM���6W�s���!�OgS�= MB��P�N�>�5oI�$�s:#���F�z��1L ���^A'���ڷ���j��i{O���d�'Ji�R�@��E ��Ppf�P��%t�ǖ�~*��B�1��^�c⬨��OV�{�@z�skL�����hl�֭�)�5'�Z�k.�<�KRR4����hrp�r�Q;���"�M��Y�����a�W�دVѓ�)�"*D�P�^��K����:>^����T�k�$p/�ц3{)7~tB��;ޏ����iJ�e9�ڻ��K�UCE�&�f��0�FՇB�%�t�붍Y�����$�0�{��������ݨ�������s���Ӌm���������Q64�8>B��KWx�Q�3}J�#����ri�����K�C�nKTw����=�I��`p�N��g�,��WI�'-�$ٹ ��U��S�b�}�Z���C�Ǧ'�J�˰Çkdw����"����6ok��vR� Dh<5���8\ߛx��FH�>���z�n�|gn�-|E�ms��ѿ�ff��2�i$�ɕ���i�~?�y�Y�[|=��1�W�)��"r<(����<��!�*��㴃2*4�&���� ΅�Q�ʝKJ_#�+����<'��[Y�Bԝ���fߥ�&
��5AB~��;��H�qy����q��q�q\�|�)��(_ t5sr�
a�d���{�[��N����F�o\��i�*"�qA雷���Xnj�G���)ɮG�U8�:2��C"!-5�	��j��L>W���0�6������\��x��9�"���;T�;��.g�nC�o&X��5�<!��m�8xj'àa�ܙ_�Qޝ���U�s�%{���Ep����|��fk�;>��+wg��Ur̕2X��̒4�&�!�8�h�e/�����cǎ��;�YI�K��[l���L��x����0�ݺ0@%���Qni���ܢ�د�V�6roC����qU �X^���K]�[�8a3���HxU`3�AZǣ]�����ΟC�<���eN�������}��)yZ����^[�D����$TR�)��F��M�A5�ނ�p���Q�BlE�q��B9FS�4f��l���B�&�b��Xb����i���*�g-0�뗋��3���Rq�i����� Ǟ�]=4�zpZLs�F!Ƽ
"���y�w$�����*����>C*�����3��$�J&2e2����~_�C8�u�[ ���7uf�57z�+H��\��l=��7Q��78 y`1���u�u��T�ʗs�ꅯ����2�t��;E�P������;���o��%�������Zv$뽏�n���^�����rj��F,Ur�:��bࡄ@�>(UX�����Z�Mz��5� zb�����{@�K��ѵ��(���(�+����p��K{�7�Ƞ����L͑�{�/�g�E�]8��gH%g�9��M��}A�X����0��N��D(!Fh"�X�鎸��f5�Qs� ~�N�1?�#p�[?NL��E<=���'%���O?�ɸ.CBʷ:%��3��j~�h5Ռ�8gK1�=�BV�ܾ����niيM~`_v&g��Y�Tkf�<�ϼ
��_H9ߓ��2�J4�l�ͧ�(�@�W>�9��9�����#���xo�Q�1m���/j-��_56l�	��T~{����t�54d���M�H��wu��������YΡ\��wW�{�\��grw;�� .��k���w�+���$C�_�;�mL*@k�^��j1���) 﫵;p��wD����ժg)&�����$_����Hv��8�2���U*�I�-K\��s,�'�/2�U&� ��F��}�z=�?PG;+����8gr��Ä+,�~�n(�YWG n�� %�0s@��H���@B��?�-���zx	�v�x�9�5������	Ӝ�Pr�E�����F�yiw��V��.J��W+Jk�+�3�;#�&3�R�z�Qg���	��ĉzPs<C L8�o��Y��c�wJ=^��3�L�e A'⓾~}oyOX�����a�6��姲>F�Vi�����4��(7�X�z���F��Y8�R��9ޗ�l��)I�������%�2J���f��3����b�����ؖ���	�7����+���,�k��2~X�ɼ��*�������D����q��U+r�"�{��P�p����.�#�ƺ���C��D�������j�x'��y������\@�99O�R�^��L=#v�����2���p�]	�o��h��o�h9��2I��)T��H��->��V!쏡D�㻌��!Q��M.�*̿
�J�o[tR�)�}��G�A���8ST_^X=��f�T	�����fm봀�T��,F�[��/���QK'
���{�{&վ>�Uȃvݸo��x�yp��#Wr��J��5�svA�|�;��֪��9'���㿎�90�e��T��5���	n��$���I��hW���B|P�DH���{���y�ύ{{���3�a��5Jio~�q�]	�
��>jV�[����X�&��/�Pi�S�4���� ����t�×�b"������p��G�+��|h ;*���sFU(�6�-���f�d*s�d�8�qK\���o:i7Ҥ|Ee���Q�JE��m���o����-�=�lh�F$i�WsѨ��DtyD�Cq�� SG�W�(��CBq[���v|���?����O6����C�z^q�}ۥ�X��i���m=Il���;�����T0����47i�d~re]��M�x?[]=���&�\�l�ν�P'���K)#���������W�g��Ŗ�H��eky�mJ�����m+Y�fu�s����?0�����*�TN��A�ê>!�|72�ۯR[�V���.���_J��w�Rs��+S�̇����V�vj�j���W<{|��������͙xA�0!1��s��y��O����,�~����5��Nܐ�X�������~=����Ӡ��b�j�Zn����g����E|��"��R�|'-*����P��p�Om�e �*oQ��Ӳ�T*
�_z��UR����rF�(xa�m��e�}7��bA���J"����X�G�YjZ�Z`|:�p��LF��F�:P�hP)��_�_��j�tZ��r��^�X��j�����?�=@������l}�H�NmD������pY���E�4����.b��Cߒ�iw}�/�lV�*�[�Zcq(?� W�JE���{SB�ݮ/ ����5�wb}F/��Pd���ύ#d2��I�=7�d��-9E����)�$�l�Wr�l�=���el��ژ�,���"��i$��\�ؤ�����̦~/Q$M�%�I��sݕ	�C��R�N4/B��d1CI.;6ȽsR��W�����9��-��U4T�v�(��&�ؔ��ǘ��ܑ�i������=)��&�MӼx-�j����zu:I_߶.z�F� �e2�Wd��/(����z�%�"��.��.��Pr�w��4)��·?�=M^qy=�LYj2�T�_�U&�ѹ�����/�l\ؙ ��+L�l�az|#u�0����]í�����N��Wl����i ���Ǡ��0`}�
<�7>3�<vu�_�����*'� ]��e	ʂ(�X��7�2��By�E4�S���ã���.�é5駏[��,����d���Bk_X-�RUm�=��$'G����׊�'ء�v�����U,Lv�Ҭ^(8�uL����ۦd5U���+[1��]~abT�3��. �w��zD�O��;��`��/��b	�I�Cj����w��� ������9�u'�7�*��а�bǨ�[�N�y�$�(
x���f��4��U���Z��z��믶8O��y9T���̏�_@��0%�0#�ӕ�:�Q�L��]i�@�ƳW67����;������}����GP�}T��<;v ���@�k��[�=���JqTO��C�;㨽w �z����M�[�?v+�l86����{<�_PB����0�����i`z��M��h���i��o44�O�]d\*��6,�`^@Yց<�1p5K���Z|��+y���yj&,a��#�[�7�G�Ft�ᱣFOk�Apf�JD���5Z���ٓ���� `���i|5@ʈ�j!*�T0���0��;n��M|��6���E��!���Df����q��N&z�a�}����B	j�-����.�Ka��2ӧ���t�9|�b�Q��u��l~_J8�L8�$v0��g2�$�us8��G����Od��K�J����.��� �z��L�EZ�1j$d��.5���|�@�;���c��4w9؎)�/�k��Z�t��<p��M�UN��q��"��e��avjl͝�x�F)���]D��׾x�{Q�$��Pˋ߷�c��U{	�]�Y�f༟�r����4��Wi�_�@T^p���M{$y�eH��a��4� M�W�أ�'��z�����2��sO�v��"\*<�)=S�m-'ː��|�/�WD]M�U�O9���΢�b���
��i#�������4�e-�Xrd���*_x�V�h$��|N<9/�O��@y�q���;H&�h����#}xG��^o�66����O:,����Y?�8����+X����r��+ĆiQ��z��7Q�9�65�ek>�aV��	��(>�֤���&QL����(Z��u5���@/zr���	~ N����=��'�ì�v�T�[^�Ё]f���b&]q	1�8��XtV\pl��A�4k6B��>Km�!�5,(z�a�4Y��\Hc.A"�u����Dj���K_�r�O�AN=�Uy���(�M&��M<P��`����O���Vϗ�Hˈ6Y=�����.Qk���k����t�JR8	HN�Y��}�d�ug	/�=XjR�S�!�4��Cg��f�}- ��ڹah(m�I������n�> eN��ZM�X�k�mS\��nѺ��xՂ��*�,(d�n-�N%�%J�{�4B��Qlq�����+]a��:������I�5��2(�0�j��
2^�����,w/nT��J�V�7��aV���|��A�*-KT�)(�ptH�-V�f�!y��Jh����xr?S<��d� k�J5�Vv0��Ó��ߤ�{a�h��e�V'4Bk|l�+7/����=&�+��b�R�n������u�{�g�{�țr6�S\�q��0�>�2Y[%�X� ��7�k|`	�
�qڡk�B� �{�����9]�q�Q��W�ǻ*X��?����Һ�A�Cu��R�ɷ_�)�?.��G�ͧ_����߾"|�?.�T�}�fy��8�u	iU��Pٸ[~k6��S�@�����t������_=ɾz�7�'Tm98��s���|��h�]侰��ݾ/�.S����)�d ���0����<�荵�v���W��8�S!\<O��i���p���ٱMB)'����%��oYH��ʎ$��M|��2�B��3ӊe�"�1s����kp�DB` ��gN5�ئ��Nߕl��Vy�-��<�v�����	I����7>�g�oJ|u�m⺌���&b�Z[n`�ru㋿͚�[g|D&#�q���.~�=���l��B}S���O�br��hZҔ^�̵&�VX]�e$&E���P �vP%��W��_\U�T���!W:����:����+L���)���=5����7��͗H�ø:�v>}V��x�|�I�A�gF��[�K䳚��Q6I�|� W/AV����I����ȰTȁ�T\��Ȳ��s,T}�2�߅��1�`��z�����`���1O7}j�R-��-&Ew�c/�)��+��M�+�ӑ�4$���R� �IS��}E�>q� �ĵ��j����z��	#��S�k�m�;��3��3D�Jx��Cb�[Y,<��ˑ���[�"ɞ�n�e;%�L�ώ]�ݾ/ً,V"�:ev��"o��pnW�C�Rs;A������`����b��I�C�i��:w掛��t�H�u���
�,�U���ͯ�Ӵ��R���G�.���& ͛ȣd9�Ƥ�B����B�q����6<��%�N�=+)�P�7Ɍ{U���3��1���͟�O2P�&��@�=v�Փ�ޚ����P�ؕcr{�<��F���!;���q1O�f	�b�jB�u"����H~Y[CH��i�1KR�����M��$�A�7�x`6
��� �M@zB���ۺ��^�!³'�[B�#�_՞�}Mb�h�Wl�����x��>�œ�I'�+";LzH>�ՍW|����l��|�I[��Ev�Z)���
�#���;#����gQN���ӯ��E;+�3_�h=�EWB��0s�D塪��L�	)}��*�����'�{���!x��m�g�)3�Ѫm�6��'nܹ;�i�B}gWQ�+�)=�k�sE:�K,G����A�GC �VBs��]�l���`��⩇�Q߯2�ϐ��z|%6����5���l�)n��M�%y�e���b̀T�� S�҂q�^n�bke��DJ�T7X�С:v�H�gA}� X�ш�`���(5V|��	�P�h>���m�[��<r�F��K�,�9Oɝ�Ov\��+-q���!@Q`2&��4cq�{��Yi� �r0��SS(J�mUz�,Qe�6m=Y�!����ܾ!̕��-_����c��H�v5Z�Z��U�[��^'Ǫ#��'���F)���Z�ȣ�/�TЛ����c�X�H�h�/���?yj��5��,d��NߩJ�L:�nnX	��oJj�rÏ��Sz�8(R���0����K2�&�,�ęA��a�|2&F��;������ ɝӨRm�P�S���|*�Oǐ��&��|SC^��wIّ�o&�����g�0͐�(-+\U��ƾ�)�|����2�N:�+w��0�hG:��}��=f�U!������A������o�Ek�od�a�@�7+��M�����~�B|~��g���i�C�;C�J�Ѕ��Ɣ�\����a�n��,����۸�2:B�Ev���#�A��M^�:�,���i��h'�
��j�e��H��YvH��A箉��d|jϐE4��Ֆ��+C��f�+�b����������`�Y����O�����I8�3z�z��#���TT��s ��{Ni<���"'^ڇ��l*I�9=p��敚��tF� (H�8<K�?�C�c��v��:�	`�MH�������r���C��{��_<�:���;릣�P�o,s��Y@F���QO(�c��z{c�_%B�u�"w�!O���2���Q�W_0�tRT��6�zfqiO�dˁ�Ss=n6�zÊD	5�1/�ZŮ��5�֞<�
�#u^b��%O5��z2;h�{��Z:#��"~Ւ"�u�:}?�����g��R�����v�q��JQ��B����Y"}, ��00#NE����@��?r$�EAL$��O�)ƃ08�����2����v���wz��i.�)�M����2�ۤx�
��w\�8�Hk�?!�����GeW5y��U���7�
��|@�޾����]2�֚��c�������E��z�_�H����K�O���ko�MoNY���%��z��.��T��mI��W�a���qnŊ���o��n���^�q�ઑ�5UB��[�����:f�Ae1�
L��G�-�m��亰�QhB��I���l�^��b"�C���� �3����@O�ɔ榞��>G��.qW�`*Z~�y���V��7C�R�����uÆ�96�;�h�$�u1�S���ܢ?��֧�;�_�󨲓�M.�&|K���)�����v�߄�;m��;]���@�G�*	�X�nsۙk#����+�ٵ�J	2�]��"�^�5A�Ά=�bu&Sm2
ք$1ѩ�����Msh��c ���V	 � =,�N������Y����y��C�F�Wܧ�����5w��6m�X'�(kE��WNznۍu4���b��^��T�`�%�ѝ���]�.�&��ޙU+��������O�"k�a����+�޻h�Xe��db���v�ۺ�Y9������Rr@����j>�=���>���,�1�,����l�k����+C�z�`<]��r���R��\e^�v���Љr�GȠ�I5���S	/i�[tE\�6�$"�f��I0�|�%w�w�I�ܥjò�����NkϾW���Ŧ�[WK�z�ؘ!1-���a��"��`�D�� �� V��b1��С�`'U��*=HI�/K�,�����og����	F�ر��z;o�e���$R��1\c'��Pܸc� �H9O'e=o�2�ICG��6:������X�w/@Wj��%W��@�}�O�4�����C6���(~ Z�掳�Z�ۥ�8��g��f?)���`f���	ٛT�M;ȊĽ.�oa߈���3h�<e��l|$;���m?�eFw��D$AeP&�t]=�"�[���P�d�d��/�ۧN�e~9��7��$��eWD�b��4[=���r̆���"vB������]�24�b�c)�߮U~Pֵ%�97���ͷ�{�}����ք
2�XHA$ߠ����b̚8���t��Z9�j�ɛ�C����*�XǱ��ǿ6�5��B&�/ϙM����D�T~�"�w���W`���i����Eh3&i�#��6CP��u.>�&]�"V���F���2�kᅸ& �CA[h�©�-��K܎���mάƌ]�4\�G�yJ1��
��Ͼ�R5�G�L����������>�2�R�8�� 0^�_����:�i�e�p�>	��[ߨ����3�#�����[��`����Xb���1�m�Zd&>�GV�c)��?��L&6'�=�����+?�T�o��l�O�i�iR��\}���i�"�U�.��+3X��Y�@����1�I��V�/�0�@^wa�Jҁ#N ����63���H����Н�;����6�L��%�@]y�]���V�L=_��6�"jQf�����c��d�P΂��<�ȣwƸ.�rə�v�ф��7����}�ix�u?���Yu��u�������d5T$�"b̇��E�;�Qݕ��a�-�r�*�wàx���J�g��%̷'�V�0�R�`�?�`���z���.e��������*��]�
��<�HE1��yx��֌�+�>��j��y�0�[]�w!mٵ̆z7/K8��kNS8�,+�^\�<S�����N���>����Hw��$��$��:&x�ߪ��[��7ܟ�%���N����"sr��D��������3��I�J��i,��U�٨��b�"��e2 �:Z���Y�B�:3�٭�JZ��&��8,��+&��=�-'���ϬA�	x���.O�Ǝ�º�H'��x��[���P�{�ܺ��u��/\��?H"���"f7�T.��!~u���T��A��5M[i)<��g+C�f?�&yƟTg,�w�ڟCiN�8Y��dY�?��N����'�<��:�+��^=�����������1GM�_~��y�g� �����?#����b��� �׶02�� g�K;�3�	n������vsw���pq��4,����-Nè����%�#=����E�����s�E��Y������a5m	�Ҏ�s.�J����Z�����m��7�q	�6�Ϊ�~`u��í���>��ۺ�r�����Gs��(�Yd�)��j6,3�QR+A�D# 0.{ޞ��Y�_�k�m�p-�x5�7hw� ����}��V�8�sa��x0�C�Z_o��ݺ�L�Ld���+5���f0X?'�2k*� �G͙��
�;O��A.M�|��_H���������%vP%��Qʖ��`(\+�Pw�
(!A��s�*�'[㋬�� ������?+e�u�ʘ�}��ɻ4<�:�(�M!�A5/����48q
�^º�̯�}�𬬑1��%�2t���X��W�I��
:��g��zyq�x�b���B���Қb��N�]'=]�N��yr�\�D�9t����wo��lۋZJ��W4@�� bJ7���xqwj�OTK���K�C�q��m��p�=�X�0L(�c�P>9��E�DS��ם���p��H�i��x��)x�%��=k���$P�{'?����Ņ��o3͉H��}AF�)m�%��(��Ql�(��%�_��<�,m��T�Q�?�\Ր�+K��3C��-�y7��f��n]nZ[�	���z��Ů�H�>o��/�±�q\)Ϙ���oyp]a@���&;��`F'��O9d�(X��e�� ,�㦶�Sn'�6�8�bl�?G1���G@'���'�B�B���v��2��P�I���g"p�)Τ���������4�����7$�be@�Јb��^~6V����+  (s����p����\�
:��~�:\��t����%��_,j��H4�Ȭ����vj��n_S�h�u���.rh�������iK��3��&#�w����so���TT-�I�q�e���g�g�;�gEA7������s�rX�������5���kA�e�� ������#���IG����;D\K{ �ܧ�~؁v��簟�V��р뗎xʩo~^��4����U��U��3���ڎ��˕�Gg���d�i�UU��T~I�&Έ$��a � �Y7Q� u��ۭY�r��k�G�GE���FO��u���[�%bX��l0I50������ ���b@ChÐ�3,۶���.{��FC	�͡��7�1l�@f�*1C�|�`�KnxSi������B����ƀ��(Y����bA}t�)	����r�sA�+��ɡ�5��8��`.��ܠp39��D/9�8�-��)S^r+�V5���C޺sO�u����x��֡҃('��"�5�̐�Pn�/��R��_�2Rȭ@<�x�	�����a+�<o&��p��3q}G��t�R��V��-M�����A�x�h%��YPBx.m�W<u��#���ςӺ^��	�\xz7��p�S0Z���� FCV6��)�A4�+vd����,�&�����z����97���D�Ч��n�=��
f����濗�L�pwK�}�[�������L�ozF�.�����e�w���`�ú��D�t�_���}dU��زy�}M�\�+ ����Ƽ��0q�="[@� D;=QyuSw�Rl�\	�}�� �k�����Wmk�����*e�d]����*v;Z�۹	��X���Q�Vav���8O)����T���8�<G,�W1R�#��t)6�bN"v9:Yk��zJ�_5��\Q;�(���#˘徂]�ɴd�!��[�ώ@��v�<4b[OQ��pG�U
ug$R��jDDt�{�����M�EheG�طT�YHZ<1m]ë�
�
��ڊC��,!�r�`鱽����&�7}�ܭ��/���`���e/��GK���?�-�(��)��u�G����#�7ң9��ϫ�,�I	�o��}7~��P���9y"�wݟ���;+>W-���<�ڬ�R3w�|����R����eh%���y�b��l ��̼h��Y#�,��ǿ�ha���駖�L�U�a�"�.�t�?v3�4��Z�"�k��Z��,f���2�����5��z��Tg,81�SSu�(����X;����6��{�,"0�l�_
���36~�,�rj��c(}`E~W��14�s]���"ѳ�����1�&����n\8�n�l6f��ߙ��+y��?��J�Y5���Xn��/�e?����^�9a�U%Pҏ�"R�Y�T���J�뗄�mW����3��A���O9].hD���&������A�svQ5ZM��]ހ~�Ȅ�Ґ�]5�*Z�H�=3d.�_'���:�)���L���e����zf�iQ��t!� �,L��c*���������fpQ�AN�~�ܖ�+����<�@^X�Jy�.J7��L�o�h���>�uA���4)
X����F6P�=��H���ݹ�I�_�S��o��bL|��� ��c�]��`�9���(�so�.Y�3�lE��)�j�͸����)�}e�B�8�H��2^�f5q��S
p���C�6�Z�
x��T]��ڠ�aw3f�aOz�{w���ԡp+Q�Q1R�J�w{�U7z>ϟ�)�b@�#n�w�4�����.;u��$��z?x��Aq)&�{V��D0ɲ� �����d_�I�D�N�hֿ�%!a9�S�|Zv�WǎA`^�i�5P�`/J&��8��x;qL�F�:�3 �I16�3<4F���A��75��v��y�X�5��L�fk�_��bA��~��GU�I$j��L����*t��h-���tN�|�=>8��#���P'lc�Y�>������6}ݣ��u�ꂣW�tap��!g�y��G.O�B�!�����"e=���
�Q}�v�'��%tH.¤�}�~�ς�����]T�*KIS3��׿%�y�0;�b"���=�r=0u�6�.�o��[���֛=�x��"�z�=����R"���#��+~R����c�.�_o�?��r#�dˉ�ش�asI�Xn�HT�!�^�� ��
��[l���ql��Ա)�n*	=`� ��[�O����b�s4������Zn�Y����-�!15x��5�B0�`�{���O�z�#cQ��Y.b��ح.��k���q�fg�Џ���r<�l1�����dF�*�^uC�1��4�$nh&D����\$ae�%�"X��F)h��VuKD�ԿV�
���fa���l����M�|+�8����o�"��|�f�����<�rD�2�Cƞ6�=K�8��Y}Ll���������T�q�w��Ԗ�	p�L)'.ODM��G3t�F��[�9�XǛ�F���L��m��R>Z��j�?���v���r��y$�-ň2��@њ�Tw��hh��Wv�fp�=�̤/�~]������Ue)3�LV���N��~"���j��`�z��y6QĶ��tl5X�t�g�Д"�3��޶wͲ�N?��V4��)R�lj�w�u]T�4�)��xۘU=�v�7����f��٬��Q�3����mٚ��-��v���`8�h��W��oW��9o�7���b�@��cPt����eC�rU�7s�Ӄ�$�Ɩ����M���/+����M.��:��*zY��3��ݲN�θ~�sQCJ8��:�oʍRA,�����:P�Eg*��	�3P������)|�޵?�0z�SC�|2�׷t�qa�* ʾ}ڼ�zM;�����K	rc��L�������׮Z��ede�*t�"#-�\�?ˁ ?�V����.�Ͱ *�ܙ�$�tK*�"	�٣B~A�=��/�D����j�N$���W���������Y�w=w�+n5�Ϡ��q��"��Q��`dEᓊ�M`��opqwoK{�U���`�FeV�QZ�}|g��J-��i5�
��;+6a�C!�������I����?�����ڇ6�L�͎'YÙ/Thg�K��Ç� �w���-���s���Tfg��0U��m�PV��O����|a
�)^(���K�2�،(\>��"�E@���t}ֻoK�K,fT��L�gA�l�.'B��a�b���O�X=G��`I��]�}�c��ͷ3�؄5�aK�0�5̓��F���r:g���5no��\�r��Sຎ�#7��G���מ|ڠ��sO��7�D`@�� B�q|�ZT�������2e}����)�ECE�b��]��x�(�Ry��S�����^�ּe�%�Ke�.�=M`d��{?W��%ь|�@�"u�ܣ��mT��]�n�-4?<dF�\���;��/>eY��{3��g�"��T�n�@��CL��u5���^�뾯�
�w�������#�jD�k}u�v�C����41����t�W=�~�M�ά6��ok�,"�J�?��Y����Gm��Z�>�4y�^X�x��l�����ռ'�@K
Į�&+����N��5����T��T����y�}U��r�Z�ۼ��� (�pk�����
���t���i���.��J�?j��$���c_Y���ALZ][�K������Q��ܠ�%4[��R_Eu_2҃���"V�sH��Z؈0�kr�f��u�2��(4J<ݰ����D�$m��YBNk��J6�Qb���,Þg�'"��ټ�(��-��RƝ:]}dD#Q�)��8Е�q��*!�����l����cSX
����?�:��$?���{����%����	3��N�R��X�i�;�8h�3�H�������{��KyCeEd��%����Wm�b���s�r⬜��HQ��*�2�b��}99�}HT�iU�_7q��-Ɯz ��Ƞ�������NyB ����a\�`>�ٟ��fS���ꃈ���H�{���"�gН��d2�HPH�����qQs�nf:�w/�?f��b�R��b*I]&��vÀG-_�n5X	��E�>���𝑌2��ݓ�s \8�G�ZV�
���>��a+%���n���u�<���()%���\�M�M��ˬ�R�0V�Y�`��^���B[3���%�v)��gc����X��{��4�ٞ�m�S[=lO9g�ͻw?2���L]�@:��W�5q8��ѕ���LK�9��0-��h^5wU�<S�I�U�v9hY����_��#����Z]$�
ݴq*$W��=4���6�U����U�E�q�K���_�����X�Ω���o����!�w��v��O�$�;��"�,Zr2pX��
�K@v�pʧf��g]�لĚ�$�$��-�_ ����j�2�/FC�?)Y�`D�=m���dQ���R��>wA�h���|呴�W�k]��6*3+�ܣ�N�u���c��`oG���(-��ɐ�ap�W8xhؿZ�,Y�p��eQ�<*�~<2������΅Snm^�0�@��*�k���w�0c���)R��,2�D�m�5�Gr�N�1� 7��N�bNy=h;����P:�v�I�az�#`z�b�2���ʽS���`�J2�Ѭ���
�%V��)�1-��3c���$���Z�:��$|��ۉt�c_���Vl�\���5��e�ˈ.}B�r%���;@UW:]��^��9>�BF�P����>�U���.@oW�o��{����ys��c%N������f�hq&Ҙ�{�:!Tc�"�j1r��H�Q������|O �0e�H�ӪM��R��n�\�ڻ����v�ܽn����pC�a�F�DRT/�l����.�ݚ�g�癁�ϗ�m:�>���1����I�/�v�p)�\\�:�>O�������J�2��Qv*]�QA��O�������wFt�a}a��G���������.�é�2��w��߈�k��Vkն\G0�9��oQ�����=���"b�x������YR�܄�F"T?ݵA�C�\r��(�k���NsF[>?9�����������G|7Y�QE��d۸ 1��<���u�R�"���h�Y�Aa���P��~���ښ@V,4D�<�pѩҧgZh%�|�� �Xϕ��SVw�K��Tz���D�VZWy��\��"��?Saʿ��U@�4�-����0ٻ�!��U���x!!^�$P�f���ƍeoC\��.�����H����T!8����?�%'��gq\�`Gu6
���/­2�v5������!g&�DJ@�΢X_��/5����Q�0��6U�J�scf>QR���Ν�r��"T;"���. �|ִ��F��C#�������o�
�p�%�x��d�D5��\�	��Ï4ЪvN�m��ȠX��ei�"$�ЋfY�c��F��ﳿ:���u��\2���]�@�hNh?����j�3��D��m
�☥�;J;��"���u�!엘��SW�K�R�p�W!�|�����51P�_� =Puݵq\}V�>�4�W%���#��:�i������(�p[sK����љ�E�08!d&kG�����D�Q15,e�9u��Y�!�I�����j����O�ΆA�F��-��T�~�J����4���x�4���
�p8����Pv��;V[-ae�4yCs|��T=G~)Zْ=Ų|{�����^b�B�e���;Hۚq�@��<�n�j�g�iծ�$����m �;��fH��/u��~U^K��pLM*@G��m���ύ�rs�,�D+��o�ci^�D1t�L1@�빢�襹i�RJ�g�����ao�h���Y@a"��<�y������������%m
��S*����CJ/�!+�X��g��[%��ӱ��=Y\J���g�z���i�vK~�I�R��SW����6~�9�L$3!ҟ���UO�"��*t�A@�I�y���d��A���=8�nU�n�?�T��32�ZM�'��~�vjiB�P��ON�L���O��������4k�w��6� _�u�!Ͳ�Q�8ͅ�u��O��t�u�_�s�^���]A�Y��O��l	�A;b5PHަj��6�$����ʥ���R.]��=�`[���v����wD�C�#qk��p>1�P`#i]7�O��&�����*�h�״���1��>׼5�G����0z��sB#Z�ˉ����kA������0ٯ�܃��O�P��k��7��M�]�0Q9������4��3BienS���FM}��=a�{��
^�S����d�u�����b{�xtG�5Q��^̓���7�I����Z�g0��mV%s[!����b��C�VP��!���*P�M����UY�s:i�5�T��Q������X�2������a�%��r��-���Ė��6�%��4`��M�=A1���D'���� \w�m�<8XA�L~�N\?']+|�e?���$Cd�!����]9L���e�)�W�|��
�3x_|.�d)�g+�
�ɘ�:!��"둁�t�����bDY��l@3�灗$��c���-*����P���+;������B�x�n�uZ�Y*1J��+���:mV���+_�25v�?x.��ͳ�%!���^�xվs5�-	)��Dg�י�&!b��hj�����L^/��f��#bR���\�E
�!x�r�y{7_G��s��]Xzѝ��T_���g�.�ImI�'��b�ױAl�W��{{�߷�dȕ�k���K�䋶�#Y��8�s�`�,�&�À���N�*�����(6 %%\@k�\�����af�ü�鞠���nx[UMjy�B�4.�ys��&<|�����o�I��B��q1�PT�Q-�^+2�����&r`�>Q�� ��X��G��쳦1a�<;9ܔ�i�$c>!ϊ	�,�p�0gN�����)[���%|P?� ���Fo𞤃~�>޾11r7��`���[�}��+������)6�v�U��z�pfdXP�+ �
���}N�C�^5�:J�b�V�AZ�
x)%p~�Ƹ�l���"�W��n��& >�'4ʽ� �YW�z��˳62�i?'%�^�ƗX�\�tJ��]��Q���m�T �+F��t-Ϯ���8
t��8�:�<ۦ����/�����R ,2F�<C`���芦 V8y'3��;y�M��Iu���^��I�rJ_���rO6i�xI�W˾��<�i�r�G�H淩�k�QNa,sB�)�_���?�4w��"��'����*Ȇ[�Go�!Rh�"Y�Z�j�<r�)��� 6a��(�i��C���pL�=C�l�Bq��"�d��Z�3��к&�A�e�l����q��;<Ո�<nGyl��QZ��jd̫a��l�EO�����|��U���2m^!��R��R�zl�b-��ގ+x��i������9��w�c�_�6B�$���w�8�E<��@���cGv���O4�ͤ�ă��r,X͋),[�*5.I>P0��Km��/p�,���)T#ur-��fQ@v�Tgk�m�����q�ϻ�1�����r���IQ�e�~�rRK~#(wݫxn4�d�m\O���3�<KC0SiK���H {e(©�>f�����o��Y�k/L�ỳU�O�<��b��=R���u�*��B���L�f*�#۟��6e��r�Ic;�Ǥ�m�%��_s�`ɺ�X'<�F�I#��O��$�`m��&n�,��"Ot�iÐmC�	t�}Vf�{4̽0+�b�"Ӹ� ��lV������x��[�-�1�-�TX?����B)rO�Ͷh�ECخ�s�Ӗ>6JyL%���iUR�
��	�����lw����1ZS߮k�����)��֢s�����ŕ&����	����?�,5��YY�׮A(>9���?���M�X`�n���R��TO�u��в����Db�2�pv��F<z�8:��T��$T\=�r�&xO1K������ƑXll��ͳ�6��_?�I�k'��xU�B�b�R��u�M��|����ł�������DѲ��cc���%;�/�2�D@�^�����?�H5�����c�+�K��HM��k������Š��y�v�F�L_h�B�H���H;J{;�+��3����s�k��C~1��X8��Q����Á7�N�'h^��%���O���݊�X�kM��B�cЉ��`v�@��߂hL�P݉g�6�&���2~�Z�$u�]bk��sA4�lv "�b̋�SW$!��ȳC*�j�6�8C%�;�����SRa!��q�j�L�_6�F
�0��~����8X$��Ù&:�"��XT�S�Q��x���K[AƇ�r:%�r.d�)�h� y�����1Ѱ�Nĸd�A�#�ĵ�h��m�s�9�߳�-�O�@���� Z�(>\��x�r�J. *{�9-�x�I���ݽ ��w���Z[��"c3��D]0��L.}�����ߕ���Z&)����I���u}TuZ�kV�tC'���]���t�4 ��1%��e���pG�7��h����rSA�6K
�$�3�%�������4uȚ��n�{�j0�>���*4��a&�j����� �o�/H��i��UA�cS��m�E���ծ�����m4n[{���� `�
rE�f��G�al���tɖ��'��=�����Ta����W:>��7t�!��4�Z>�8�y���sH��0RhN��X,{-�a^�_V�����`K36a�'�����#���o�����`wn�c�IΆ�V����iv��KeZ���뇀5�J�w����k+>�$L�MX祡�48����J�A҄��y��պ"�o�e�w��(j�xw�.�
imJ�����m��ɴ:'�����t���4��Ef�d3ڥ�d	�2t��Q��I����q[c(��P��������u%|���s:�=��PGmci�֔ԇ�A�
y�-�Z�(;���X_G�-
�)�`3��X��z!�-�_@Q
.4�O� �?�Z�Q��X%���0��f�4�n;�@�HVlt;Q�O��'�@mk��҉WjX�
A[b0�ߺ��8V[=A$�z�|�Q�a�=��n/?�9_^�^�W�3���ظpqEz�KD4�L,��{�5��[7�xH)�ca����m�����͸C(2��ⷢ����D�#�oh�E��3[��Rd��~�"�I�D-�}
>��B&���apȵ�Oh�az����n�	{�L]Ӵ�'Ȥ+����C_{���X��<>#Z���i��W~�jM떈�-�H9c���s�&d�3sz8_�*���<���������J"����*�UAܢ��d_���{Ϲs	�K�쫽Z��y�f$�ʙ�`aƉ���[h�C���Y�|*�F0�t�C��������]=��`0�z<0���s�Pg��QO�]�?̉���ɡ���5ρ"�iM�Sc�^�?m���
��]� ��}���H$�VhN"7ύ+W���'s_�A����xwsL�)�f�h��4m�א��4J�����e�� >bG���VM��Ɩ���Qۜ�1p�s�s��X0h�;I|�dZߓ�I���n�:�-�5��j���bYg@bz`�(���a�x�U�I&h�L�W�p8@�@o�(Q3�r�2%r�\�0G�\��]�b*����Y�;,-�Gk�����m�U��'l3�F��]xn3�PUzwrN8ô�K�U^�Ռ�1�Nʐw!�M��s��B�g��i-��i�F��������]M���N���9�='i����VI���/׾�ꝨqI��Z��'���{)
��?������\�w��3k=�Z�y6��	��;-j!��{p��Xd�{�8oI&�J6`�!�6H�S��1�j$�A��d��|K��Kq܉x���(�-N�AG��6[T�$���#��u���e���F��d���fe�l�}���Sg鳣B7F���౶��ˢ!=}�Vpk��n%�S����@�I�w4���WY����9a�x�*�2�b{G9����E���1
�8M�\o�p"� �?3Ē%`M`N�\B�
��RI{tgd�ÍH7l3���k��n�	���a������uZok��FP�k�{�r��4�>m�쬙A:O;h�Hn@k�u:lZ�;l���.p=m��
��O�n�aܗ�Zۤ����@U�:ת�]��k`�|�^���^#Y<������K�z�$���I�G��}9�?`��T�G�Q72F�ޥ�K���@�#�C��G���wS�)�:A�7$��I�������P�6'<����r�$�N����,�%�J��}uǯ9�����& �Hˮ�$���**t'��e��O�����Qw w4 &������]���T��aG'�N�6�c���~�FOi렏�� �41q��&�l5�����[����7��jD�����c;��^a�y��C|�%Z�l��,�a�B䞗	�"��r�5�ѷ#�sx��"߂ߥa�N�.��(4�[g����Y�U'$1*ݣ�Kr���`�|�CΤ?{^��j}z����u��k'ɟ4���A�1�f�z�G�p��pz�\�ԨX��C��]S����	P~%d�W�@��暬=�&��\񂯶��ǝge���7�@��<W�[<�"M]1���1��iFҝ������4���%�k�r�����	5?�l�^+6s�i����D��n�rg���@ct��H��j9�4\�3(�ޓ�2]Q+y�q�}٫�!� b�h���,0lr~���x}Kߙ�3�*���e�{�TÜ���;_�z�5wG�i��
���8���OeZ��7L�Mdc���/6�lh'�r8Jޫ�&)�����;1���8*����R�����BG�̜�h��nX��/^災�s"Q@V��2 �W�Q�~`t�|g79y9�8��yjK�h�
�)�tEA���H����"�Hɩ���%��bSz�Yx�X��&��ҭ�!��=�GG�u�C�x!T"�#������)�nYe=H�Ӂ�??eh��f}���W~��T��ʖ\��^	��k��Έ��Vioa�R�o|A���y���E]��9�&�@�]�03�۸(T����� �&3*�CP�7i��8����ю"����O��-���T���¸���	��K�Ю�I|��fLIbS9�#	I�}����l|�/
\�(���j��w��@o��j�k��Jё��[_��0��B�EWd[>U������5E6hæ���gj0��nH��`@0z�����|6�D8��ծ�W.��i�M���Y�^Kg�G�e�@�|���,��8i�` f����E ���s԰6Z5�LvW�ڒ��;�(yX���D�z�F�����q���5X�BӺ�d�z�ro�d2�
/=�\M\2���1(e������[�@f�Yt�~oz���ک�1�ğ�J@�J��}u=���ڼ5�oK(��I��*�HA������e u�W�q� �{_|ڽ�<�������)7�A����J����[��%�"���E�lp�	!�m��h=�6�0š��{8�ޜ���� ݒ*��^��74������hg"u��Q�G# T��FV�Q-M��qeg��H}����{=�fϨ�!�]6 ƆD�n���S�����~�6��?��  � �t�+��l�p�-z-w4� �9�Id��}J����m.Z�����Q�B�dYl�E��t�Mri`A'�|��y���6��D)M�RQ&t4+���jw�$[Q�w|4~�!�I��<bP���P�Bٱ�tș�W�^�#s�ZL<~�ϋ��.�-5F,LC�y�冝e��g���p�&F�dr���^��j��?�+vśn;r>A�(u|��U�:F���Q鎑X��JȧQ��[����ʢ3�I/ƪNw�����jL�R$˂Q�boy�#���?
/��$m��{�-���5�~-��e�*��;L��b�p�>���AU^�hTH����2�������c3����ÆV��^~D��ᚯ�؅���4��R���\i�nO�d.�K�k��Pa����08���̚�'t�<6"���S.�i�V~�/3�&�F1�f,Ri���Ѵ��.K���R;$��\mj��&�����n�d�������/R9�t�r����֫��c����Ѱ�i��\�D:��W� Am��[�	B��2�]i�������F@ܘ��:�U%T=[���z�LPZAX��f���)Y�r�)`���iit7��W@��2�'�UU1j�B/B/�2�*���ʴ��@���
�Wʦ9�0��2s����z+�<�#ǖ�X��\���ˮ�jO!�m�W���:}�Z�I7-���kdN~�0�U���Y�0h��xC������)P�Y?�d��$ˌ\4��h����v#3m��cq�W^��8\1�?:ی91�n|w���ئϐE�Ч3�f�/�Ǵ3����"Aql�"�ن�Ι�\�L��34����1���ރeRsr�I	�l1N;[_����fy�R w������di���ֆ�Qꜜqx��I���U>�If���N�+�oo.���k]�3�G��}�m�ܹ�sP�m� Ql�-�=�<��S�	x1�ѕ����8��2��oo�=��������O�=���&�G���U��æܚ}V0��C�+��2��a_iٞ���9nt��.�T����zk��|��B���@x_EI���qE�����R;Aa��vE�|p�g�'��h��8q
����Y'��[�S��B��͠�`4{�h,�~�Ӳ(&���&z:*l�|�䴃D���K��1�TH�С�m�'�l�U�4;��+"Z��W.	>��$���(�PY� %e��?n���+�RHB���$ݒ�6��y��$k4�`�T{�=ʍ5Zkk�d̝���4�d�+�M�1޸��!|n=/��k6uSi)�o�њƖNlD-��>�8Lk��L�J���������V16�}
)�z��#�Fy�4`�Ơ�[�)��tk�G��cau'&�Qv�i�00���Ȍ�1�|�
<L�yfT������$�0|<�P�H�8֮~�'��MVS�#�l{xea�5��b�V�oW���q�W����V+L�d��$#,vGDz�ݾPD������x���Ј�-�����|���0�2 ���.��wY��	���ݍ
*^��[}���_A�&O*s�FF������xRO�v���?4�
��
�g�eY�u��JD+*�'-�'OܐܴD�G�����՟o�ȗ��w��K}žL-�,�׿zj<0:���ˋM2�����i�IJ�H��#\�4�'�	Į+}z*������}dH#��ctf��&��,3��9)��w�t0�(p`2B!�R�s3�+^��oג��a_���#a��& �y��J*��feH"1��F�7��5���3�ɝB�
�g3-Q�}R���a2�H�ͱqa���ER��h��B�DAxjŰ���������QV��B���Pe��۽��4>^���(��M!1�h�#��CS���Za ����q� 聼�t�u�+u1��
��{:\���in0=�����sݦ�?�vk��;�8q�;Mb�������s:���h�؋�5���E�,:z�=��i��pM<x'M�b#� yY��;,�$�8�����Gt9l�2w��|���]���+�Q���)�SC�œ��n*v��y�-��o�CV��h�{Q���7)*!����F�0���
��B�\fX�g�R�oQsX�NXx':�ӏ �d�c��� ����5г8�@���e�~x� g��-��~�V���c9��`,�}y=y� ��\��a�M�)�d����b�U��s�Y8n�9z��rD\'#G-�Ԃ+��QKבr���ԟ8��mz(v>r�U	q+��Ai08�|��"��įD�S^,a�rC����jA��|�P�U�b)�w<�?"�Z��3b���+�?_-�P+��ٜG1C���D��58���3=���n�@G�
|��71Z���א؁Ab����y���ס�ڲ�~Q�p�z����Cm��p9��p,OW�9ک��qf������r�6����JZYu悶-$���LH��l�4n����8��V�SA�'۩�k��5�+��T�iX�T�����f&���{3�_�	ta���S�0���:c��|=[����d�m#	�]�)���E�9ÊD�[��f��C:dl�3Gߏ/c�XN��.�9:��	�#J'��tV�dJ�L��h`�[5�~0
��	?j,�i0�'����������� ����-�d��{�k�zw��P��:=W2�?4!��ϭ6���� �gV�L	��h��%����G4W@G2�,�Is�&��@���p�3�� yƫ�pԿ�9����2gZ�E��na8�:�b>�n2�`�$׈��lڳ@Q�y�����mƟIF�vg!C��/��L�G 'f���J3���2N�V�=?��H���LX�� ����R���yM����������������u.#>l�RQD>%���l'޽�hʢ)��w9$�I�|�u����i��/5f�I�t�
r���Aݚ���65n��-�d�\f�躘v�e(��F���� a�U���M��TK��ߖ��T|>U9I�"-_�id$Y�SR`&�����m gg[E�F�^��7&�6���d�<qBauP�i(R�OF�vef����ơ�{�A��`5F�eߖ�[�%�=O��T޹^�F'��/)3��0V_���3o���ƹf�����L6�w�A��[���=nE�$��Ͱ������TʾǺۂ=E:n��)�+���ү�_E�K�4�4�w�]�=�sS�3�S��#F%�%l���tx*��jhKd����Z�k�D	�	WɔY���9��HA�*��iS:�g5������� ��J���7�`ז�'���(^�rwCD�x�bb��.�"����][_�`4\d�Q2|K�`[��Uh����Ҟ�Bך�Xg=���V�����w_�qj��,�RF����X�����⬥>�?4���n�y\�=�^$^��1W�fVO�7�L,#&v?p��O[����\9��(�Bp#�3��i}eZrW�:�:h�!+IO��玃��c�9N�ɺ���M����J���=$F��*D��{�?8����5�B5��2$Đ>�Oy-�9��K���,�4�
���z��u���i�de��陠hqF��G��F�����4LO(��?��z�BKĚ�w��z���F���{	�:��iV�+ �V�$�����Q��
w.����䂴>�$���z�`^f���Y�57J��n 7�u^��y�;�l��?"6��s�#c�)��yڄ���*�o <}PB�H�B 
��"�P�/��(g38���n������RT��7�mͨ�����B�*�k����.�2���Y�x7�{Q�{i�}��=�Kж"-`wˠ����˰`��n�^X�w�㮎�_Z1>q8}80Q!��n?p����B��v2-��E�~K�4�h6�������Hm�o�$�פ�?�����VM;A>��b��eN���x���s�1^�r��)b蟾��j6\�#m9l2ԋ�\j��DL�m�.D��s�lz^�q=��b�7�^RӼ���3*d
���[����8tO�;G@��g�8�P�����H?� z(����q��D<o��I{X��G�`[��uC�S���7���j�W̍C�� �<Z'�Ʋ�<��~�T/ |&�����+��yӖ�;�^K ,������	�~c����=M2�w�����]��_���L�d�a�[���qY����)�w-��� xKJC-l�w:��W[t����y�t��TE��c0��sdH`�� mE�w�&�P=��i��`��UK�� ?<k��߲K]�R�N���Q��w�p.x�J�ϗ�j���T��U!9 �F,B�B��D|��u4U�c <o��E����G��/�~&p����}W��_���S�Qzկ}�����'9���+���lk(��d
�n�=U��W���-���#T��[�լV�-�.��:ICC̓L}EMU6��yآ�."�gjQ�<~�b^MƊ5�������@R7�3j��dDo���+�RA5Z���}I���>��)FPŷ�Ф��18�|���ž����&Y6x~0�#he4e3Ǆ��x%��'��dR=���B��'�]N���aV��򂒗ߚf�ϛ��J�ؐ����0�c��|�8^(�u�B�t�ŵ:���^��=a�'���,2�K�>�`6i@ ��o���*�S".ٺ�).���Fۘ�eڟ�hg��>r<W��*���=j[�q4x=$u��^)�N�7�0GR�V%Ha?�ㄔX�r�O���ʌ��=q�"(sZ�/�q�~*�P�T����F�T���Y K_��i�����JJb�J��O��֪J<�R��U����3�d������|��m�eEA�׎\���������aW�-[�s�?�}޼|V(<9���d�3�g4�a6���\T�j������n��M!��uD���}x�M�x�b�*=Y�tE��g+��RHшΧi7u ���Y���X禌U��P���9��M;�X̛�X���/��붶�X$&#���Ô�?�A@�$��
;� �n�fޞ�I?��$�&Wh�`�/_�Mh
aݩ'�p�a�3���:���a_9\��|�U�En�m�o(X����{�����[���˷-�j�q䄛e�0�n����JG�xO������T���HRJ4.#�"[-�q��c�a잌��$m�ӈc��wZ�i��{����GP��HF����7���:�7�S����%U��	�xě�vS�k������ia:h)$�`�>a����-ͦ���H���(Y$�<�,�?��=��T���̉n�uom$�g��q��O�F���g�K�#cs��}%��W��c^�u��M���J�J=~�b����iGՓ�6�����L��ĆĦ��av����A z1��\�7���PJ0]�E����o0�a��=�9�ă���п~f��-��W����m��/Y��(E 2S��a��-�o�_X¬I
����ݕ���K%���zk���ƁP�{�K�!ft��b̾����m��G�C�Č�V�T��+T�Ÿ��ai�F����H.���H{,��L:�A/����}e����RsR_q6{k.1���i��I44NȦ�2��T��#�כ���P�j��S���R�ϐ|��s���^��xՊ�K!I|w���8W+a���T/��OZ�����$�9�_U0߇�8+�L	�����_�ք��FB>R�����G�la{..��v�G�G*ԿҽI�>� �U]��C����0���ȭ�f/7�~y�q+Ί�@�^��|�h+��]�qto��⺢��U݈,���Nk���>mǙf�C�c H��u����׽Npl�w7�2)U�"ź��f9����y�d��e��F���7��~���"M��۸��9!7�[^|��R~���gv@����"��:��������c���<�]�0��d�1��=����Cm$z7�0����l�z�0$��Ro���fKe�Z:tH�W.��Ր�}�@�s�:�m�ߑ��]����N�r:X)�E�ӈ�	R�I���I��]�a��!�^�U�(�~�.\�[��
"B�?#�)�IF��!+�*���~_ˉ8�"��A�E6�#*��p�3�w)�_���W\W
Rl,N�T�yΧ�9o��n}@i�������3�>"���5����la_�zc/Y�>�o��*��@O�}!�
�Y�hk�ك[�2��j��Q��W�!�͂s�^~y	3��m-0RS^r�s�]hq�^S�?��^A��0-������s A7oD��J5Q���-k]8�h����-����O�w+�w���|@~@l�y�?"�ҳ�1��A'&���Z�3a�a�6 �b^M��t�������M��'��Ɍn�g�v�ٗ0c���hf������Oyrp+�3_<t;�[)E���ӆbGĂ V��8��+-頌��#�QÑ��$��=���&R��2�
v�����P��c��?�x&ҳ�+��0�K	�ZO�)!���cR4>�cC���l����]�`�`7�>ɉAzb(X����u/�(H��f�T<��Q�~��I.;3��"5��6�;%�v�_���^q(y�`Mp�G�w�1Fo�0��������	�J�<_x���Is���tt*�	I��TQKE��"��Tx���Ң���b��$	;<��:#R�9���@5s�*���G��b*���-�F9�t�H�`d�IN5�ɧ<�5
j�.�Q�l�"}� "�c?_�(���h���$��'x���#����+�MT�XF_'�zNl�x�qR�6�V�_�B;@Q�p�r8߾u4	N��[��0ӖB[X'6�.�%�_��IM������7���S#:Z	��ﵻ?k�ӛ6ɫ�͞��1#����FP��۝imK��ND�wL�q0X'�oQ�gLu � �Wmڻ����o�3�J����V>DY�+z0�߂���h�3�U��^��#�����^"G�k
��!^��q���=ݯ���ĵ�q���l[ӧ�Z֝G�9a��|$��/�߯���(S�7����3S\ԅ}Nc���v�}�~�Yqh	���o�nK*#5Ȧ�]6%�^�Tu�K����L4P��W�f�k8��ؽ�ۥqw=�Xć,'��B�}X��F����SCL��u|%k��]���[��8B��yuu�N"Ҟmr5�B�G����=����[���b�;�q ��)g����WI��v\�W|�E�~s$>�;�w���gT$���.�î������ڧx	ɏ˔3�a��m޳�H\��^�ʩ�G4�Z�d�~�F�(ԡ��oJJ�N��f����}��I<��`N+��i;��7Ԥt��S��|��0�z�G����Sk�bB?���W�9�B]���.���(5��q�?�FxV����q�����&��k����.�')���1FY�H���V�9UX�οN�@$B$�a7������ ���sRim&;�2���-�f=�1W^�2z��ܮ��+ڱ�}��6�7�3�w* ���:���9C@o��FC|L8�?r�X�5|���a����(�ߟ�wOG��L��;gL|.mY�es�r.u'��'V�dY�v�դ;�]�wT����DO�nuG�/���X ���1�Ff��氀ɑ�9���\_��?u���������+0�/
��&;A��;��tm�D���1��@2CO[D PƈE˙��X�	M=��%N}P?��<������A��}0T8���oOx �hb�W�6n��X$K܄�I���#�cLG�+>
^���W��Ǜ4]gč��4���9���/bH���1������f/�ĝi���Iń�{Ϫ�8	ȼV(T�*?�|bՁ���]�~��S��(�����EX�݅h����(���[&۵���8��r:b�ٿ��&v��BVJN�%3eӄ#!V's1)ѹ<��_]^ɼf���E�E6��������"�-��^�l�m�y�]q�[��dE������$"�,g���ORWz[����hn+/�qOS��@�{x��#�A�&���B�I�A	�����44l�;�g�+}�Kx��b�{���i��G��e�����RPx��$d��:P�tMk�߆}yI?S<�꼧M/l���͎���_T��|.z�����c�#����Y�n�2��}��� ��aܮ�bf�hq�9�4�jǓ��
zg�@}��0 1����`��>�-������Rgv6r+��	��kH�V��] Z�%�,!bx�~)ˈ1�WAm�VT|�����*�aj��^Z0�>�цŎ~��,)�$�f6��+qɥaT�N^ͷ�es�%���t9����H���a[�r��ۿ�.D�N�xa:pc��jtD^[r0NfٙR�Z��f��E4���������IX�*}N��w5�+�Sgi�>�ӆCe۳MO]�ԊDu�:QLm1�<��9���D`s+/֦�O@�hMsd�`t�lվM��[���L#�)ib6������Q�.�!�as24-¡��pg#n���`��������|�>νN��f�h� !�yQl� Y��n@X1 ��x|���AQ�%#9#5&��P�X�Qf��f�&�&:i��v�{%�X�+���C"���X�ۭ?��Bjg���s	��}:�z4�-���E��#ߔښDZ���:��{0BG�y��{-\�X*KM�oǕ	�SxmG��Ob ˍȲ7���~�`H���<# �7a�O���3:/2{䴍����D��t���l���s��NK��}Q;:v�6(M�B�V�$m�Eצ��w�)���f��Zo���H%SQ�B+��8p3}z�}}>V=C���p�KR�^6o�0ȍj�����P4�]�z�݊��eҝ������"|��p�A>ԧ'B�#?��Ɯ���;#�|�Ҧ�Ae�:�l�\�aJ�ӍMk�A�F'�0Ǳ�� dl�~��P2�U��ض���wJ����Jns��?6mM�=����md�\[�d��;���DMff4EF��N��_-ZvJ%uFk��I��fM��*5�L���!�Y�鬎ւ�%ί�����л	b�ۿ4ӌ9�s����d$º���*8i��I�m�cn�@��oeMLe�S&�?I����&4`sC�[��2O3��اM0�g�8^=�ڼ�:\�z=9�G�g	��E��t)(��j�@t��6��U�oq�_�@S���������l�"�lk{�1���v����)�Ͽ����8�p�܁5h�'){8�v�8C"�+������E.!
���t�=��^،���E�� ��'�s�J�7���ݔ"X�vCjiV\�f�M1e[c�ZQI��y���Q��R62�CJ��-�@uʵ�)��kIt_�y�<M?Ƽ����Ϙhɡ�f�^�����[��{1�U��v��^w�V��#���?�R���dE^���ބ�H�u?�D�W�g�6�M�>�6�rX����԰��忋e��c�k���;�bpET�F���#W�&���^j�"�֋ߌN�_�[4H�'G@�P�/40ӶSK@HqkHz`��?'��!���e������l���/ą�Rs����Q�_�nIO��-������R
�|�V|ҋ�i��[����S6*�{�����k���	D}�Tt'F�B�G[#Ez2�s+8[ ?Vd��H������q i�:="����xj>�]�;�Wl(�$���O�Y�˅2�D���	���D;yb)�{�^9[JфE�,���4@��gn�"��/6����h㢹穳��B�_�J ����1����� ����6?7�v����X��=}��QCwM�"D��'%�ԍ�ʂ��?G��?0�A���
l�����0�ᖅ
Y+�U� Ύ�/۾K$2��h�1}�~�
������L�~��=�Ė~s�gl��V�!����^ǎ�x_�VB�G͹��%rvc%�K�J�Cz�K��|����������B�qX�5%jͅ�^���@���>�z 4�E�_b�S	�T���I}�Pȵ��K���d�GTN�����w��8�~R_9o9���0��6c2�������=`�:,�j�=���ֽ��F���;���9�����&�d�5;����q��(%�mr�Z���Bl@@-D��$����3�}�b�l���5%�r�m#��B�a(�0���5��U!�S��,�����F�	ˇ�,V�i�	}�����k�	��x��r���T��	�Q�Z.7�M���|P�T�Q�m~����+�ҵ�{��&1 ��0�aN���eRn��5�K�I{���d��昋�x�ޛ
���Aׇ�%� �A��Έ����O��_��DT�b��Dwj�tM/��5Y�����l�ϙ����� �N�|n�O����sb���/Z(w�o�{�!]S��J�v��jī7�K�m�$�ƺ�u%�4]a0F'��MR��ʗ��G� �`O��B��KL-.�NS� ��s�]��a��v�}���E_w$��B�uœ����Q�d�?��?���q�����/�	��)>��c]S��~L0>$�#�?9}��*V�
s
V�W��IE�k�{-��������X^�(%� �g�;�n���z�;[g�e�.�u�L�ܛsCN?�O��%W�A�b��i�D*��%�m�đ�z�<�$-6�I"�5���(�C��Ic��zvi@��4��{^n�EJ�u�E�9嬅7)}��c�[y�S�Xc�$^B`E��^���B�u	G���s���'?P����FN$dY=��-¸Er�S�bxh!��w܊�k�mD�is_:�|i.�C��a�ա�M�U~	_~5ҟ�_}�S-X;0�H3�γ13����:�Ϗ$�r�H��Q-�_-F��Ӊ��9������Rr9��y;��PVP~�HdP朝��2IB�<Z	��`��+_��?O�{n[���{�Ծ�A�i��j>�n�q��p��S����J��ঠ�����! �!��≳U�B+ �ɑ/{M�P���i,4nCj-US���z�R��Q��c#VzpޘkŌ�Q�Ƙ?"����x�ھ�8����+_�'j�4��C/\y�y�-�����\g���\��4��%Oѫ8���5�*,/�Z}���P�a�c�����0R}��~���I�av6B�U��m&J����M/2=�b��1�x��jq�2Y���N:�;�YT�C�=1ÿ]�2�w)�9"���QzQ��dȥk~�{�
�8���P�з��SC�x�q,�~���Y�M-}����&^�� 3�!	|�*�>᠅�ۙ[% _�>R�W�}j~y~&�/�2��y���A^����$x�$Nl����fcO̬/��j
�Ǿ���N	���f&Y�'�H"�@$����F��
��+�芴��Ӆ�[�؛G�b'�]��pJ܂���Pu�Be�m%���!��
xܽ@�w��6��12j2�)Å�$/��A�����Dذ��Z�gW��P��,�o,m�9#��eʓJD��d��eR������n�'0�2�F=�+��@G s�!�:�s3HqI��Oh��_i`�e/)����$�î��w?=��|e�KF7�k[�Nf.���;<�d-sN,KɄ�H�s�<�	�G2E��̮����� �Ӷĵ���$��3�q��=�Lק2�|�5U�Q�4��f�J�����P.�V��ѣ^��j
H�6;�,;��^�^���-��ʮ��v�U���~�Կ��-^`@',i�^�4�i�X��'�+���O�!��D���:3Մ�F�L�#|Vw\�n5�HHie.Qo�Cs��?}1���>�(����@�����6=k��\[��G���j�i���3�0���>�"b0���j�xedr��̠~d�K�R�U�v� �����9����E���6]J Y叠���ɟ�5�=�����u���!x�v%��,}X�?F�A��j�)����A��ϰtz�[C����8Q�T_�j��:V�*!��~�qH�Fcu�(�����
�Bkt.H�L2�\�>Y`�`9rᒇ����y���t� ��3M��e�!�G���-�[��H�_�ap�Q�����ؔ�����b���}�����I���"�4W�%��rD,ֶ�O�@gT�oݕ±t�`7��v��We��D����rz�5
]���q�;�޴"	w��Ģ�$���Ӏ�0��K�����@G�q�����lP�CV�k�-3N%G8V�O�����ҳ�*��f�c�x79�*�M����#�M�Xt�Q�����z�p#G��*d�O�������Z�<s���#�Rb�y&��C9C4�����!�m~��m��¥k�����۰��PȄ�nq����=�.P�Dݿe)��b
6n=d�fg$�^�>Km4�5N�ɥ}�T|#p%�̳�B���+;
�X�S�����,�����/(�j����s���1�~�ޱ�C;���g͞�����L*c�	2;2�	�d�@�
-F�#��{֎�F-m*b�U�������S���x�0�"���i�ƯW�d��!hZ�����E�1lW�"\i�|mb�Љ��	[C�6�Y��n8[�NM�U�10�K~�ө�z��6��DUm`w]��~D=!�P���\l�	4��C�bP@	0�+��j,��}��Vf��Z?v�~�T������v+D���棷�}��8���s�c�~$���s�E�&ps4pv�A#ׅ�"��!���E����=j���%����R�J]B�]�_tdh�0`�һ5Z�0���GN�i3��"���a�4�SOmP׌�^����J�c�qm'�B�����b�T�cs<�oe�U*5>�`[�X��u�S�I���Xd>&@���z����G��ф��?��8��q����T	�\�ӄ��>�5¥����/��[d�����O��B�́�����Fl�:��{�i�7R�� `��N �B�x�;����g�R=�@)o���Ͼ����'�� ���pU.2�i�݉����(���j:Q5��%(>�9̮��5q<�Mq�o"Ҟy�UDA?$���S�vc���Q.W�!M�ۓ�ڳ�}|̒a������)Mp����k����e�LՌv���<wh�-Mű�ꪎ܏����[j�@�{Q�{����o
v�lU�:�v^���v���@�8�t�<tF��wL���(���[��ȳ�CZ��'��
�>]n���ñ����4d>�2��}�����`���;�%���5<\���`z������	��n��Zf��l�⅃���� �� R�j�X�O��4�q�Ӣ|>�ꮍ��y�[cVzpb�z��r�%�s{�1�hU��r��(���á�I���J�l`�mV�������2��G�lE��0)	秮���8L�`�~5��fP՚A�tt��xN��,��+������"���&�W��OfBa�aJ�CJ�(L�����/#�B�z�	S�I0E�=�~-�i049?-	��Kp�h.���i�x���uw��M��A�%l �ڐfW����rg�XĂ��	{*f6k�&��	��"����s������:��l͝�iL�Y����P�",3cK�B'���l�['ƈS���d7.Zü�! ��<}�ҫq���NX�A�o�k��CԱ�]�=c�K�[�!�����kj,?O'�K~�F�CӬ��PY�n��	xE�h>�w"������y.���� O�2��`��B9�h|}�r�[�����~���A������C�C�Ǐe=t��u�DC�n�U�6{��΢�������R��/�t��"���6�&ܕ $���v�=n������bfr���m�"$t���=�|����4�{��1��c�<�L���a+j:4��u�`c�(�`�i�h�-� ֣r�04��o�>��x���Uj_�_��)@�*�r�y36F����"��.�}^���\x��7sy����W`�r��ʛk�c�8����z���+��	��%���D! 	���"�[��ݺS�%�q��{5���_KT:@.��K��,C		I�5���	��.�3 qb%)��f�
�����N ���MTA�H|��	�c$���n\nT��4�s0Q�*���>��g�KW�7���\U��
���IgC�zo�A��-���^�@9��)97PU{�(	CQ@]S��8�>r5�%���t��]��`��o��U����e�����^2��6�Cy������,�:}lM��^�)��t9���n���#�����	����0z��N#����>Ǽ��l��g���VD673>kr�r���+�����Z#ͬ��A��VA��G���h�2�p�,5ZB�Ly�2�Ғ�.��M�!	�Z��/\{�x�*K��m��A��Mկ�:B�3"˿�K�݇iR���S��nY׽�fX���m!F�E���lˆP�ЏƃzY[��{L����)�b_D~uzN��W�zD�ﷀT��A�eȇef'���&�KSE��w{ G�'
RR���F9΃����y���N(����xd�88>d�[ ����l_U�������'Ll^��r�H.C���e�\?�^%0��#�4m��lg���p�6�Q��t��x~-u�-+�Č7��PUAm�<�tF*"���m��죰(�`��ܮC�����WjqV 8��؈��	m�w8m9�=�) �3�uX]�2���8,��:�,k!�Ż%��uS���5\ۑ�`Gէ����`3��Bq9k�(��7�7���d�c�J�b�E������S!�j����٦)@�)�����R ZS}��w:�ƣ�>F}�D�O����v���T����la� /�B7�&�|��~~�l����D@~�O���3�q�$n��CU�A�B[YF���Z.�*ŷ$�R$�}�%�ָ��z!���9����>��U����Zݡ'�y��*�$<%O�8�W������d�wiO,:*�Θ�xGh���ɞv4�u�q�d�hJ��C�$�&�N�Q�Ł'���c���D"Ԑr���0`�����{����!�]��,y$�A��2��JC@@�[ee���3��v{���!D� ]E2�V�C��/��w�(���s����7&����27n!�'���'ͫZ�Fb@�u)ׂM�b͏�Vf������#F��T�'F��^��#HY(���@Ƙ5��廻F�J+ڴd�icGh��k��
�U��5���,�O�@�	���c���R��狔s:�
��]��x��m���؍g	�$���)O���	�l�A(����ԯ������%abj�����ղu�*���H��3��R����<�h��1�q��xD�Ê��0.b}t��������D��*c_l�$E
���9�F�N���jJ������Ĩ~��o��̷�8iY�\:���D�E�s�Q}J��PҐ�!�}��n:�B���C��/������9�@sG�����X/yU��
P-�]���;����g0���ZL&�g����y��NDR���^��e�G�%�p���Ud���kE��kn���������辍y���Q������d�I06-�0dk�a�ou��5�)0���Hoa����k�;�d7f���!��d�_�<+���`Ͼ[	�R�"�H��ZW��8N��x��~%J��n�&m�aJ�F͇�=l�u�f$��NEK��e��P�rK��M
�A�/	,DՏ�x���>DUwbdU�#���������n��}o���[R��Qگ)c�/������$<��U a�M�]='���Į��I[�ۯ�3`��o�22�y�˻�`Er��E��k�0_2���/��Kww�/X�vwkǬՈ<wH���i��]�l��%���5��wC}nN%9{N ��Br�k������)��*E��(�
\��/�%&��6�S��ۮw���a�[_(�ly�����������?�O,c�n��cx>b��g�Q0X%���}v~��r�)n��m��DyK08��>�UL����a�e���:�SH9������I�p�Ӗt;ƿJ��k~�NnhD~��ҡk�Mn� ����orٟ5 ���̇���c�1/��jRIjsS�����f��Ý��e�ן_� �4�}⦶�O]��Z�P,=c�\'� ��\�4��o���	��E*��Av�L������E@O�6)�W�jӋ;�I[�`��"�䫗��z�$
C�f!�H�w/���i޳qWp�˪6�8��o]{�K=E�k"��7�\���P���|`����Ɩ�}F-��o��:�������X�| �۷�@ ����4�^�!*E�[q��5u�4�����Aͧ����v�̎X^z7L�u�O��C�-�}S	T�Hg�h�#��Gw������M�W4�nz�'��Gͱ=Day@%���"�?OU��uΆ&���{ w��H����*H����ɟ�!*�.��v9�J�Ţ���;G�}dSiyiԺT�}�7��(�F�sC�[ �利����n7�N$|�T���/3�O{WHz��B}@�5o�r��� (/�`��:�͑:j;lR�z�̾:xKU��������w��[�ʾ}��:���0r���A�		���>h�#Z&iӥ��'uX�4�jLv�!k���8FX'�s�#]���9��]u� 	��"!j���Uj&mq�c��feN�E~-:z��d�A24y	��j��H��c��>	�Ho5�($���F>6���]�)$,6�Q��ĸ��N���ɖ�0�w�=I�$�*�۳��%kU�z��j-����Ms���	��d��VV!0�g��CS�V+�6 ��ز��;F�PbEk���|J.)܁g=rJ������F��k�h��˘r4ħ@G;#Բo���Q),!l5UVk/� =|m�MY���#�QB�Ц^5Ja!�nyP�TBQ�Mu�幽�_=Ƿ5_�>���s �{R�LqHK=�C��eĴ�/�e��.���]0p[���G�V;+��~Q!��/+V8+ٍfV�MGI�$�����ɥ�|)7�\�;����w�Z�*[gi��pnX�"!��,���M;���c~��d��K%��,2y���^��nY�*�e�T"8@��9�5W�"t$���S��1%(�4��N�.�����5d�~���?�Osq\>|/���X��ԭo��\BE?���3>��Ԓ��k�"�NϢu�uB����,>��x�v�0T{V��=]������%i�����k0!gh�� ���Ïk�{t� y��׭j5 7�	����ߙ�m�)�OC	`_#D��:J�2���;K��e�]W3�&���;&�������~_�@����Ci�!�{�,`��s�Q���
�ԗq���"�#B�
a��%S��#�� I��K���jM���!��F�T�[e�$萅L-����\Hq����vv��AX�����]��$���da^ÆF!�+	b)�G�� ���OX[M]9)h�\9�X��DO��
�Zll#����_yg3޹�w���S��g�%����б>���c��z�9xSw��W�� �k��d�3���P��jO�<��W�2������<n���_ɌסAs�'���eQoI�NL��ӕ����#n��{`@ө����)C��m'�ZX';"m"kr�3N�29s��I��.�cL
(����D��\�c�e�o��@�η���`YJ��]9�iyhV)��@8ܯKU�¡O���g�Z���ˏH�ކS*4�b6	{�]�V�Џ�q��-�)�|��$k��'2��l}Ӫ�N�~�<���=oʢ~ݏq��+	����Շ-z|��$X���]��DqG�ݞ�[��E�nφu�}W�}�Nٯ�����$�S�\�R�q��O�ݷ|py�^�����n�,�ft�L�u�	��(P>v̻\����Nt�x"�D�r�ԁ����է �e�]y��_e8�].�f�������5
�����U�cCmV�Hq�mLa�KNƵ�@�K��)�/?e9���&�;���X`��<�����B��ߛ�p��m(��lk��%�k$��p�Ky�	se�2
 �M�$|:S�Hd��qs�[a�2P��� ���C�o�[�cdyAX3��)DD��d��[�;#��7�&w�u�#d:�frzD�n��M�P�[1=�~4��3�!A^����d�f8(\7r��/�����ܲd��+�2��'�n7g���=9ѓ��Ȉ.�"8+�)�("�zU��w�]��X&J(��(��� z]�ь�,HTw�r]g������7�N`Q;w)'�p��K{#��
����,���:�o�5��<*�,�ߨ�����3j;����
+L���֗
���:i���MeB��xD���Eh�L�#��+�|aM�TS�FG�.�*b�p���`�s��/��/�"�c�)��-!c�}�k����}c̞��n}��ڱ�K%3\'	��Y��H�&�>�5��RJ�Q6�z�;ITP\�|�lX�;�*�����0h��L
bt܌%�#){0���D$l�5�"����O�_H<�޵t�W��-T��9N�B�8#�����VX��C�L����Ў~�,�進�6k�)kM��S){�"�y&�8�M� �B��b����'��_��)g���}n�YLƲ�::��O�U���
�):�v�Ә2(�x���ϔ}N52���|L�'��� �]u�N<�i%?#Df����?�ۧ��c�*�܂�ͭ}_�PkN�	T�)���l�UP���❬v��"z�4�r�u�k+N�����G}�K�_�H�7%(K? ������қ�*�6�X�7�0��i�v�<�M�z�"w`�Q�ȍq�a	��RIY͐���︷�+���.Ő;OT��n ���52�i�M����>�����,����9K:kB֘hpl��	�~�~[/�����hŴW1U�&!��>�[����x}�7���@��L��y�mkY��B"_��j:;@kq�+��&�T�w��&Q!WZm
b�A��'Ðf���c`k-ꯅ��+u��7C��:��{KP�QV�#�D�m�������/�-L��A����"�[�#l󡻭��j}*�a�]�*����Էizu��Y�9#�m�	��G8D�N���HZm����]��rU��8,���V�B�C�/���یVC&?tl5"���kUހ`E͓}t&�!�a�~>5@��_l�>���-8��(�" ?A�dU�z��1�B���[���Ӹ_����L�5�`w-�L�=�{�+̤T��{9�d���j�J�[�ɦ@1îNz�K��~� ��C�H�Xc��\Pj�iޟ�sq27\�����䎎4[N�9��z�4'^�C�1@�ݖZLI�z��"���c�I���9ܦQ>����\����@M�8
�rgX^9���϶��������v���-�%�W��~V�Ĝu��	4����l�h�L3�S���TB���1��˒��Cಓ�� 8�\ v���:�w�� 
Bo�q�${HHF�J��Y@�"H�_RL��!�ɸx���T��D�C#��3m�-JLuH�~bΓ�����K5�ڢ5��a:XbԠ��~��G��RQP���Շ\�]��L���Aw˓��W9o���q����pc��Gv/>J}[ث�ZpE�V�c�B�� "
u6ϳ;x�)��4��.��ӝMjx�Ӈsͮ���a��F�S5Qs�������3`4V`���YA޵� h:�>r�3����2��!����"6k��:�%��6�����j�����2�$$�)�H�Y�43DA�8(�D��IV���XC�r�=ڳ�]d��S䑙o�����t�р\���*�������k%��W<v�D��������89���3ޓ4q���rj�I~M�?\7��-A�Ns�����t���O�'�B�Nr�W�ec�?�2K>�|�Erg�Tߤ�,b|x^,����g^)[{�.J:�4cQ�\*�����Ǫ���6�m-m>J��IL�3#�B$�A2���cN0B��>����e��F(|q��"�b��p��`�p�~7~>�f�&d��?#��������8CJ�^�f���2��~�=fܲ���2 ն1ʩmq{

�(�B�w���0Yb0�3�i{Ŕf��,���{h����@G,Ѿ�?<2}봏�E/�93����#��< W0�$���V.�1UjMQ g�y|�S�8�'�[u��.��oO��}��i;���A%ɛn�\�+,gh(�|٭<���*͠ri$��^����ύ��ꤷ�0h9�[�>p pV�+ ���1nSqRH���m�R?Sy]1�ç�.���I7��%͋_��������5Q�AZ.�8�3����@���ڞtE _]���)_D����u��q%x�3F��rD��!�#�|ѻ���C�"�����m�U�\��Y�M���\���|�k��2��*������w�S}�vUYTX?#�0r��K`���_����e� �ZѸ��C�6�RΫٹi'�d\˓E�Rf�6��"��z����Սs�4���+]T+1��k����u��l, �#S���6��Tۧj5U�v�jjZtS�x��	b�<&C6�*"�&c��,|��skQ��!�^�}�~�(�B�)rcW����u�� n>$�{�4�f�Yl4�5�$tvOd�<>ז�����<ӆ�:s��LQ�4lk_b�oo�����^�:N!���z�ܜ�O�"?�T��0���4Q�x ���D�>�}��KYF�q�+K����>X�eh�^@�CI�D�IH�(~�D3	�D�vA@>�;�(C�?�5�c�����=jW�E��]j���ف�q� Hߪt��fL"�M�s[>�j&�ke��R��,\�	zl��'h"�5�ngZ�p`M���r{P����k�r����7���K+-hi>�J~�"X�'�{�%�-O�y$��jv|�l&�	�W���������.���)�)|�:���q-z])+��f���0�lr<,f�Fd��N��~Yr�� 0�纳�R8JJ��m��,Q�H|�0���;�P��X��4w
C��� �<��H����G�B�e5�u�#��K@�#㙑��3��
����H[�{�:T�a7����x�&�ZJ��3J�3.���X�B¸�'/#�F̫���_���5�}���N#��Y�Y��M6�o��m��߲55	�M�|��Z��V���6}�پ�N���l������ǉW��T �6x4�h?��?���נ:�:$	sԸ���d�l��pt�m�cG��,��%�����~f�Q-q���$.�e�W�/od}-.���n�8��o�0�!�V��C:�?��O<I��co��@��*�[u�eG�E5@վԑHsfi ��JI�������S/fR+��x�|ef��\�(y�()�2E�IAڪ�L~��Y)��!�f̕�i����ғ�ּP�{RJ��;�P���	�����Ư��"��iQ	=q�V<��j����*�s"^���)���f5%��~��m%yvw>�}R��s����Q5��\�E�\��S��b�P/y⚛�S/�1�k��!Խv�d]㙫�8��S�s�lAN]S{�n5�>�ˡ�R�Z}X�\ym|���?P���.��Z̥�x��,����c��E���F5�*��Ϙ�>k�E]/��?P�z��s�e�pr���N��� @����%���@����/Q�BcJ�U�X�~�����O�jmx�*�7JZ7)�������`/7(�{���G�W�E�-e摞�a�jv �j�wm�Iӷ6Y���m���U4���L��7GYQ����7y�E����s�GP����aS���E�-MN�Rߊ��bn�_fZ*�U��8���=���h$�xBc׫��[�2H.��~&�l����J�kT� �� ���^������FZ&����ߧ,���j���)i:,Lb�dyp�n�?=~^��'$l#%��Œ��KB#���*6'��O��z����w $��e�须DKw���8Y/ߺ�`ܞ�މ�[��$�8�x���`�����4��1ߋ�lQؒ����I����#{P@~���Wl�Kb"J��ɗ�;�j�2��xI���ʚe�����E�ͪ *@���+�¼�E�RS����ި�O��-���\kM��TX��г�>Sn6�體��-H�KV��0N����@�C4	�;|s
�|���@rw�?���6��2��
�r�o	�~�;��%�t������\� X�s�U��z�5�1.	�e�2�[�[�#�H=�jpܨ�����K�d�+U�<Z�c�E*�	���^��3_^�1]Wp����}�� �	g������ 2�I2Y�^^ۯ!*.t=����M\|5k鳄ҳ,i=Ö�t�Y�sb"�q�wȫ�"Db`�N��h?������Wl}��k�+��ixc����ݵ��k�t�����z(��u1e�̓�������q��~V#
"w����^�(��]�i��sK�;��{V)Qx�_Jcp2ٹ�~�f�h�r�Y����e�Uci�o.�Td������&ͽ��Dk�>��'S[�OW�@����Y��@�e-`q�%�"	+IK��U��U
t���������O��(^�d��������b%�$^�k��6v��9$2b��"-
�T{���1@�~5�lP�X�}��uO��<j�KC�?U�Ci�na�2,;RC)C��YL
c���M��;%{9��;�q�:�>��x��QI��PG.8:䷅�����a��~�UX@�є���G���#��>�=�:G��@ir���>q30x����l�E,}�N�����޸��EW����ݸ�4�E
~�E;&S�y��cS稙�Owk�/�q�\Lkܟْ���D�H�s!�B�3�F�ɗ�c�r�v���K��y�9�!��}YČ���Ã��Hk�ͣ��E�::`��/e����s�\p�.C��pж�k�L���oq?�<��@��³[��AU�]���w;%���L4(�yH���`� d�Y�~j�d�DX�cH�0��<���S�#��[-���F��*��ؔJM?���b�JT��2����e��w.}�l���!���{p�j�	0�L��^J44����mmG�
���D���P�p����$D�c�Tr�*[��{j�-�=���gގ�:����W��u����dn�ɸ) �>�l'��)�mv�֮Q��<<�¥�q�<���
�\v���AI��Q3�=�-�r�&�_�qj�~4�-.`�p[���k��� ?u3eІ�N�JT��9S�1���1���8���TL�<��*z�r���a%��8�N�����!3��/TH�6��iQ)��2<��D��^1�W`|������i&P�^1�o@���v<�Zy���+� ��]� F��/o\�X eV	f]o�n�J�Z1�h�@�@����7GI"b�M���#Y����-w��M=}axWYC8}��lx#������(z�ۄM�O��s��'oC�(dY�A5B��^\��SZ����x*��p���U��;�l��M��M<�q�[d���A��Q<�-�cg���������^b�� �1�P1��I�fܿY�tJ"G��K�B�����}"�?���v۲`�~�YDI	����_YR�����h^�_�F�O�ӹ���jZ�Q��|��2Z/��4�ݘd(q,���h���^�uj�Cme����y˔�O2ig�NR�r!�r�2�1�Ԫ����$����:ȉ>�B�n8�QH����<�E�Y�a��b�4�`��j�a���G���H��{�I悒<�)��N}V2բ���3�/��Y)�-3�Y�4�t�N�ɧM��g#�O�m��W�4[.�NDWh�0��v���]P� ��)���U~�!���*&��+!�4G��$:|}�M���|y]�+G� �3�zɯ�@d�sy�p����:#�{�3��a
83�6l�;w,N<�C������K����Ʀέ%�I�����'����)��f�n7z���Lx��~��͈H�U�_GV6���V%5������!�����v���s�K
:q���N��<��N@�(w�h 槟����/����8�1�{y�+~^e�bFn:�pc��W�J�h�m���0�}�c�H�x��*YQ\�8IޚLJ�xO�DJUF�ǫ۹�"�l�������Ét���3[Ne�����T��姼�ތWԠ��Y��-Z��:mt�h E2�� 7<�r8��~iwc��,�|~�X���`ӳ��ֻ��B튏�����b���>A���\Qm�:n��v#u
r廸��� �o����qg~����~��k8���� ���E���-�c�H�_�o�Ds%�	>��qz%Vvk%w��[$��5��u�g��C���(k�I� �{tv=&_4�H��\g��8Ã}@��h���rF����Ck��1�����_ު $&\lX�X�A�?��)���4��V|����|�W�5�ʒ�_?aY03��Z����â��mWک#ͱ��l^������������4�vo�cwFWn��sM���5��?L?��%��ܜ��pW�5y{�$�"�vW����t�G >��(�ݤ���QU�h.�ݷ��g}��-��dulF������N}ɖ��y�J[���b�o٪l�4�us�A������Z8S[+��������{�w]|ЄDy�K�/�}/ܐ��X*M��i�� ��
��L0ZCb�2e,m�>H�#��Ktf)��Y\�}l�	<�k4�5��j�eن��y0�0^��z���dGv�E�.�����8ߧ_� �բ�d�*+��A1�W> ����+�<3%�O�� 8k�5���f{���r�����U���l姂�BE�*d%s��*��l�H�̲�����=���!��|<y]Մ*?�cR�i V��#�<`Ш��<��_(�L���r�"Q�z�@�a�U֝��7�D�ň���\6>c��y0�7=���R�{��J#K��~ld���bG�Z�!�C
�ȨU�a���P>�[�w�p8i�����h�h�j�1�Ywt�V|���Vs6*�����=`�傶��-'�<���Lk���Z!�J��\�\�����ar?��Ԝ�^�RY���lg=�9����s���X;|�]2�o��_+��o��/�Ho�lU�}]���ܛ�������^e[70R৪ 
 �9��_�����Q� ��"b �3��y���r��<L�
>�/��p�o��LB�V�9�9Q��F���?�~?R�����;$r@��t��N��`��.�;�FL�Ԗ�b�@b��wW" [J/^6���,����R=kU�w/_��~Epc����6�C����,A�m/��	�J�ɻ���#K��"�#50gl 47a�2�^���cjQ�>���1�1�Sm+�8�.p�d���n���#�7���6B��Ѿ��B�h$C�6d�-3r&!����ۃ�J��J��=B$R]{��ta�T��H�
v�r��E�\��
��ӟ>�e�����uD��5�-��#u��)�g�1N���ǖ���e�kR'3	_`�L;@`; 4�2%Q.(��D�ޞ�h�:����洅�SN8HVQ��UH/c�D�VCG��MzRW���)N ��4���3.wg��dŰUʠ���q% ���]�eR%�E��o�&^��(��0�g����{(�A��^�CVL 䁽�f��Er��k��� �	&i#�bh��5��,�1[�\��C��	�@����d�N">�w�@瀨X�H��+���\������{/-��?w}C�a?�|���Mz�:�`������u7�ۅ���4G�ݲ).�i�B��B�T��8��a�JIK�`f"�Г��!��q�+�a�ؼ�	��"��&>��Iӏz+��Z�l���1ߘ��s�˖v�+/�i�D���=�:*paM�OlO5�P`@��|�ٿ��ԎF�]���W$���|���C¯�5�?���?�{ �CV�;w�-����`������WB����x{�QP=v�9��6�~er=Vn}���S%.&U��,�73|c&��L{�#a������L\��-�Z����Kv�Y3�����˴�>��M�Mʔe��E�iu���9-��w�g�v@�#u~����ע�[���m�V��_��0�љ�6����T'�F1�,s�Bx�ߔ�	��Jx�)�UCu�@1�}�.ś�����ӄi�1�IeGs!�i�~e�9�9�@�.��1�MRѺ.ey�C<Cm��}EѮ��~�݊�y e^%&D��%C�A|ͨ�iT��D�2u��e�*Ӕ�gMU�r��mt��΍�r���ʃ?��h,Su�ddMk)�/=��[r4��ב¯�5�S(d(?,� 8���lcEd�qp(pu�lŭ�M�ݦ�ofd�=>��2`.��W)��\bq�Z�3_��3k!D� ������_)�|�?������9���O�[�A{�:쭁	A���R(�TЃ��B�;�"��.Z�F�}'J��a�	W�Q%�� A"�4対�NZ�� �\s4z��W��:nPe~��c.<�Y��0����i�m�Ta�b	W�x��&"�jf>��d�K&>�mG�@��^W�9z�-W��`�<l�4��~�z�^����F*��0m�G�� 7���C��j{E�;��(Po}��D���q�Gi�R�MLX��_��i��9��V5b��Xo��U��L����E��[�$SrҘÿ6u<rj1덾���iЏG4w�vQ���4'�=za��P��\�x.��h�h�Eg���͘�}>^i��ݹ��o X�9T)�]����&2%Zܺ.	���C�	�_U����3$�o/�"���%V��}T_2�C�!��z� #�#�VY	�h�WcNC���F���艗=3 �7�"��?���
�Q:0��3iY2�9�|��쳍��f^����y�y#}�:5���8���j�3r�AB�P�K��O 冽F�6T3>�v2�0����\ƻ~T]�xyY�G��A�qV;"qE����p����y��3�F�Ln����_VW�i��w��XT&6I97��e(�|����k%E��`o.<cH���#H�v�XI��Nhc��}7���M��/A��&>�nc���PF�����B����@}#e�r%qw�q�̆f��eܗ�6�?��Zy�HHXg
�e\�l�.ο>򙩨��#V8EdٺI+g��"OY
��,����_�~�6<j��]��]�^��q�ֆ1n?\~;h�'�,����c�K7$cL����*K��~���c������L�P˙���W˴U=d���q��!�ޟ	v�i�Σ}��W>�nc�Ѻ;��Q%�7c����/�R~Mu�u{�-��]�&���W��2
1�������X��(R�H��"���.^�0�)�A�-2��w��m���5z��Zd�/)c ���b�.o�NW����( 	]��%���f��HQ�����!*�L�P�Qi~P��ώ���+<-Жd�K	��;��(��}L�ҕ8:�f~���֙w�\��Ǝ'���<����7g�!lPb�P��e�����'Ⱦ�#�e�L77?��ކ�\���Bc�`k�!��ڑ�M[�~`��M���K8;أ�ZN�T��\"� �� ��r���>���e���Nq�Ob�
7�3r�-D�S�;\����m�O�(H��PH�D,��� p8����Ս6�-�����Ũ�o�%M$�.��$�&������`��G��N
�;4�K ��O�4�[F�e�(���SZ��69��~Q�\�;�$s���W�У��p��]�(p����	�C��
��v��B<INB�K�K�����ʬ7%w3ϼ�����GA�ג:Z�P	)�D�>���!9(�E���͍M^30A@��i�*r��)�Wq1��x�����k}/��gr�I�b����m�x��Kd�󔒋5m�Ӡ ��q/r��ō�S˰*���{p多�s�n�i�BK*��;c�b-!�C���9���CL]�����ԳSs7j�0����ߌ��\-U+��HQ��#������M;
xrM  L�I�n���
� ^W�����\��]�,+L�GS����z󷠨�yQ$מ�Մ�9���L:T<Ҷ�Z(?c�I[�:��a%��I�6�eC��+c�	�]��Z�o�(��@�˘����]G�e�#.�TmP�܏�<��sE���̩�5&�DQcN����PS/8Ӈc����H�Ք���!��b���a3|��ʲO��~��y&�YZ׿G���R��+.�80#Z�ֵ-�3���p�$��Re��y�(ⴋ�7X JY��KZ���s���k]�(�:�.I� T�muS��/��.���Hq4��b��Nì��yυ���c�x[�4B.���iËW�_a�5�h��K�ą���9��B���:08�
����1��HX���/���Kwų��LQ�O[�c7NZD���v�rm�(xد�ᝇp�s��e��DS1�&�ʽ�pm�&�	(�cI!&7����!S�g��!�ɍVNs� ��YuL��2����@@o�n���)8����yJ-��v"�qL�Y����C40/�}0�����"���Ş2~'���Iz���ǭ�:�����l����|�C����A��{��?����������z;U��D��� �'Y&)75��)Dq�hA�%k�{ƛ��{h�M�@J��x6-�g.����Z\�rj�h��q��W�ح}�G������qO����_T�c>�_v#�M*-��c1�3�4����lb�-dx&��ȋ���@%_n�_�C~T�Vߘkzw��'��_Ld��^�&G4i]{ڤ���G�e�X���So����:���&�Ҫ
�ȴ��p9�)h����p�khPG���^F�
�1����+��լ�$�"�̈́�~�����N�;��Խ�f��5]WR�]ߡ��of���S��l׷f�3C�K���L&�����93jѕ���U��]K�IjO�ܖƆ3� ��3����X�߳�%)��Q��ꀆ���K��܄���{�����#B�9��|L'K���P{��9�7�E�s�\�J��-�Hq�V��~nv-Z��uf�`�9;�&��}�y� )Y�QP��^����n_��-�[B���U��J>dr+���~�\��>�e:�ӧ���2��K_ȳ,�<�
%�@�Y�-&<DQ����7�ⶺ�]�'�'�qF gf����Z� �V$5�}
h�'l�OeE��]����[���t�U�)�����.o/��,GR�ʗn�Uf��&b�(�N��.D���U��i	�;#5b"u`YEN�؝^*�n:���T"�ڄ�9�O��{N������<��.�\y4�;�*G�*	��cz)�*�z5;�XU�*ГٞUǺl�0HDC+[��m��@5$jE|� }�'<�S�b�/��1�ܟl]�V��Q��]����|�[*��*a����u���'G�6۟R�7遻��l`2-��"����n�|T�X����Fo�%���2&Lm�}_P�1%#��Y��Ǵ��W�-{;�)�L@�����pZvl�w�B��/,@�1���vk��D\y�j5��w�Cٹ��CQ�������F#�������}��g�D�'���&�W[���'$�0����q4���l:�������5��TN���"�6�2�C���k�0�W��D���fw�".^���ĉi핝�5��>	����a�@�ka���|sc�4�����Ri����kA�o��n�ǰ	��~3�.�$ ��+'���~;[����� �n�U�Y1�����Y�|�H�>��U~߰]%�I�;#iIy4�j���J~�[崱W���c{�ǍZ��}#��9\Xy\NFF��Q��[;��6���!f��<;"=�?���&$s̗�tGg
q�·�pw�.�&��lqs*`��nlq������֨��4P�(��=���$V$�}&�9;u���1�z1�������9 ��@�4��5�B	"�8�v��&���zw��(rz'������Ai�qo��q�!�_�Mv��b��'�,v�ot�V��ge�H9�{u����mc�%P�>y����Յ2�LS �������xm`��u���~e��UF�.	����$[�uס��J{��(�|>�o����ڂf~��V��,�wgbKT����Guh6+,Z��^礢����؛Z)6H+�A��b.
I{�Jgw;���(q,B�^K�<Z��Y[y~}�~�Z-N�Ӟ���R�uiަF��,��~�M^e��|/��f���q��>�B��MW���&��v#�uzj�S�̖��N�c��%�2 o�)����ޒrZ�L���%�b���S>P�sPu����6�����~�"���sHN4{P�|'\/���J�z��˟�W�`}Źv�/9�;��d��S��u9���2��K��Cp��U)��Y_�y8�r������l��^3>�u	Ԝ
ҩ�b�?�I��J��a�9"#:@\��U�ť��uX]�LЧlyS�������Ņ��v����'ϒ��c�j#I�<ZǕj��h���k�N�K2�k��񯧖��r����dn�J����V����e"N>q"n� �[9q5ԙݓ��c;�P��,h��e3�EF)p�)��&��RG��\��a��'r�F�z�?pY�3z��}��T� �u1��~fĐ`�
�sE8a��R��GVߵ�f6�'�a�)��6g�5���|�NJ�r°�_($�z�~��b��{�j��|�sfp�M�t#���Ԙ�AUY���W�,c�~���sD	�rK����cf(�Œ�l���%�E��ڶYJ����o�!?�n9XYr��s�CⱯUᓑ	�u�C4��ے��9��T��f[)�˿�J�Ƥ���J��nur����I�b#ފ�j��N�8�NgC��%1����2oO��WNfH�|9��ɳ��x�˱Q����s/�`k������Zm�}ЇVsk]t2|*n��w7~FGĔU�q
��s�A�C������w��C�o�����N�r�c0�E]� +�o�s.��
�l/����X�p�(�td���a���� �NK�$/�;\�_rnJ^(:@7fܔ��g�2ۻWF��aR�oȫ}�$�<w��1��3�r�d��e��9��/�R��?��e�����\y�yh�AU�hY3�Ɂ�T��O�^�+��:�6��!f�������b�k��v�����U,�{(l��-���pr@)~�?������OM'��o)ϛ���f���sү[L<_N������xB��$M����fUh����&bl�>�����r6x��R`�8�8�j��@~H��S�{H�cɬ�Q�����D!��.�t����ƭw盠Kߋ��&�yn������£{���+pC$����<k�Av�%s?h�����	�{�*#&YBG�q�W����)^g �Ξ,��~� ��M���$��a+ɷ�����:yp��Ԋ�6>�t����e���7���|*躒|*��'��&�0_8T�{��Q��D�}����| �e�@eƂ��S��]�G���Y��ek<-%�M|$��%�ؐ����_�?����ۋ1�L�
�3�s�;�B*07�e��'�ɾ�	���p�Z�E�3�gκD/��Y���\ə�b$	v�Oa�
��ql��~}{�0�i��!;�!�2j�m~�UX�j6B������[�¨$�Q���|�O|ߏE*�C�Ȳ��	��:$�\�-���4�Fi��iw`�Q1ܶM3��W�]�֮���M�x�ٲ���-"��������ErL<Y�X>��)
��I{1�1��IH~@����x�Uw�\�I��YDr@�ȉ��x�=Xݝ��+Ssse��r�E���G����y�K;PC�,����2�����cvք8��f�5����7ӗ�����,n��mb#~�ˍ�|�b~���[U�����w��@Y�E<�q?�V�8R'�UY"���J��/�3��_���S}�U�V�O��+��B��p&��U���'3 �%�B3�Ľ0%����\ -B���2��P��o�>��-F;�4�y�T3:�Ǫ�s�Po`���y7A8����^�ʜ]	#^&,D(y�F�T�`!�3�]�3����h0�868#��O�$��-���2q�Wo�xz�F����h�T�d��������y�i��%Y;�@�L��T�Z��
�18�K�v*i,�B�n(�/9�<!DV�"�����֦��պ�yx�Y/�0Z)��<��;��Agz������f�����l�D����Wnk� ��t9d��,�t]�KW:m�S(:W=�����:ݓ�'��xY��	ībv�S&��Z��<�Q��i@Kg2���HP�ࢵW��tV��6d�������o�s�ʹ�>*�ԓC�;�A�U�{݃n�'���R��~�/L��Ԩ��W�~`�$�0`���
uD=��M�JЫyXY0Vm ?�vs���J���x=�g��;œ��ć���~N��Ӻ	 ֯��5�Xr����t筗c��Y��IHfxG�!7D��	��&Bc���%�W�� 3i?ڵ�R���V^o�e����A!BA���6C���R��3m�]7P$?����쬼 �i�����x�!�%�H��s���!~�*G�0?gq�x�[��������6�<���њ��Y���{�w�Q���p� P�[�u|.<E�ͷ�����cz��}M��9(Z�OE�%�׬R�pt�ܹ�Z>���T���lv���ʗ���Ӯx �2!��ѽ����e�=M��H,nV��0<"u�<̖'`㈥�U�N�߉����>���8zY�P-���MJ��ݐ�����}��bX�9��"�9w�N�4[�j��_��
z��:p��6X'*P�EA�lៗ}&;!�3q;�?����>Y�S�-��赸���x;q��&�^eZ$רҀy46R,���
L��>Z�QPKG$�y�b�"{ęn�u)�{_!U�T�1��?�R�L�{�$IôH�]�0����u#�CܸMk���GvWZG^��:����T�t�q j�~Gf�s @��uP"��7d��I��߄ /6������	�,jb'��M4}Ű�A��:�1�1=B���(�?�3��4�B�	6���}�`۸'t����ⲝ$�*\��_���x��r�3m�YVcjS\��8�&�y�u��u����͘��V�6)�Ӏ��'wV�͒��Љ������e26x���:�eǸ���y��.p�G}I�NwR�����,D@�0vItf��{:��m�f�4��]�ӳ���{;S�(d�yk���Ǉ7��P��/��
8wS���'� �(d%_��˩U^
���۱4)D�+�ÇUd�YR��ۉ�-S��?�O��IT=��T�f&�a��:�K�Ed����Ma`�|��L5'W�S�D:pHT�A�S��3�.d��'YN�����=O���N���O/L�!�O?�] ��ݙ[�9|�0=.OPy$��uLQ`u����pT}ڳn�����}�o�a��#raB+eB\���G�߀7�{Nu,��z�O�6φ�4'X{��:a]���{������~K8Z�'����o>��X���m�����FG����V3�p3�LpE���a>3�5z:h���Im�T^Z%Mϯ�,��CR|E*� 1�[�ϙ��"�B�LM��vc�W�c�g��c�T��LG� �����+b6�Y$�,�2�(��jV?�	W�+mB! f������'{.QK�t@��ռP
�vkUG<�S�yOg��b���h��m���\�	���y�N��������~�U�g,SIq�m�3��0rH�[����7���\��(�.U���j+T�E�J���ƴ,���]�߄�Կ��:��=O
W�6o.�'2&De���y,���ך������4�E�IR9=V( ����?���e��)��-�`�4�`���w����Kh.3��79�" Q�t`߂�֬Àyd�>/x�l/����>G��`���_X��5�SnX�t���ۺ*�w���3|�����\ӟ0��dR'���d6��:��W�z�;�kMfRh�L��� ��1�G
��w�n�<�;IǵO�K�K����E��l�.wţ$/Q��ՖJ:z�q�]y�,�։Γ~CzDR�>"�|�v��񌢫ܷ�%ŷ�o�ym�t�i���6�%�燸��w0�{�J��Ffi��-�\�@/�䋑��/��=CǶ�.ݭ�h+J�ܰ�65�/�h1!Y���Fa�Kd�Wm-���*e����?��!���;)~�A�m���8�ω���,ݷ��`�s�����3�z������X^����2]"''�3�7cf����]Z�]#�W}fԤ��	�3.����"���Z��'
n����<�L2�t�I�����l�RG��(��#�ה	G�M�Mj+����.nm��A�
J4����+-�-W� "|K+�DL�hXpI1��]r[/�=,C^�/k��`j�E�a�!TJ��ϣ6#Ɯ���CD��:vÍ��54��e~�D!l����T�{J�`6�>y��ly��0.E��a)�Ff�s%�6�^dc�<,8Y:�J�֞:��N�F�Q01 ���g�u1MTm�R�����	"�0s|u#xb�T�Vz����ߍ�1� YBV([�s�s�o�EG��/�R�\��M$�A��&H���GS_�*1"�<|�U:�E0_�<��c��k���IY��/϶'� �V-G�}>����t�E8j��Q~�82d{��5��Eb�.�o��8yb,�q[7lk��72��t\Y2g]-��RwP(���������.�nئ�P%� pM����L�y~q��������h�+�-����C�(��o��[�s������ԩmp̺?T��P�D�c�88g��h{�>l��и�����ݭ�f�'Id�;��Ȳ2��4���.N�)��'�VZɲj���׿�:�U�0X��}2t�H~guπ��@��s����9�"L,�N���!����<�����B�H}�y�5H~�<��@ ��&��fq�M�ַ���(��y�.�J'Y�}���rWx��';	`h�lw@�+6jZ���퍮�Œ�w������f�����J�6��,�0C-��m�g���/�z�Nn���淛m=\"�D��W��M��ng;�+PʿB�	��?e ��l��&:���.�aL�,�5N�Av+P3q�����$e�	�# *��N3��foF�cB���t�%�0�W�+�8;?`��O�_Ղ��r�wZs��2�����b�����wc�������)��I�Q�3y@?pu�]�;�����v��^�_'l�w�;�2=p(�Q����2��Rϴ�z���9���s�V��$(�U��Z���q�(@?q��F&ņ��)��9g�F਽�8��"I�N�(��S,��O�gň쒂C�O'���/���SM�v,p�2��p(Q!���u���W?��~%ʨk�_�Uqn�(K	Z��3�6�@8!�-�fZl�m����d����[~����]�SQS�~{���� M=BM�����
�
�l�
F"��ұ	:�����$v����5��I)�R��
�9%E�s� �Ϸ���(|]����Vr�p�~��V�@�HC|�k>��D*i#ƃO�N{�9�5�<���~CMZ��Ӱ�6�m���hz�/I0��u�Zʡ4����r�m�Н��y�m؁���c�y_���C�ܹ%��@Z��a�Lχ�����y�M�`�%�i��9��.�⻪|K;x5˩Y�g�����w)#?�����(��;`�n#�:��2�>s�gZ�F��rؒlhh�%4g�6��DF˦eL�ːwZ�IwK��³�7^�=
e�\�9[�Φv�yK��4�\�1��C �jm$Z�c����T
�ڜ�p'CJ�&vI�y>b���DړP�W+�j��/G�K����m��vӍ�X��4m�Fxd���������wW������h�*�Ԗ_�d���79L�ٲ��ެÐ�a�=,�c���R*�
S%KP��h#cǴ0�G� ��}��W�fR��=9���1=|wÔ�?�HU���D��.v�9�d'���e�h�`�tyL|p^9��Ɇf��5j�|VU�ژ�N�$�a�q.��q		z���/�'��&���cu��o���:4��ZJ4�H<�R�n�;Cճ+������Q��_f�����J!~��Y%�=0�-S���+������d='Ǻ/G�l^�ٽG"�p���E)Z�%Nut��`�M�]��زJ��!�Se�%w��}�<X�o��}nB8�&������څ�g�x����^�R�o���&�|���?6������(/��I�(�|Hm�����L��3"�#��yA+�OOA����:�q�MO��NqrNb�5q�cY����KZߎ���RY������c4���e�hF�Jb�;?)��j�:g\�R��!$�ldhD�(���7��
��X�SD�.�YIj_8U�0�1#�
k�w&�I*3�>�C�L�m�lW��̮��8΋fò+�P��KQ��Y~����}�D�ؼ���އ���6M����{�I���ɶ[,s� �ɤ3X1�}�ĊX��7�έ������QaWf�gu�~I}�Cق�9���ZLM���@��3��ϕ(f5G�<}F�=N4����/�eJ����,�r��k�:�ewߤ����|���V����ЛKfY�!�W@䝟�s��{gu�6c�*훲�#v�h��4j��i3ӕK��ɱ�%��E�K:� [z���s��å��]ѹS�*�$pW�@IACw�A��;�����T��@��CFm�;�� �w��B�dc����53�I_��*�}<M+'���կʋ�"�V��:]�R�I���t��_gPWT����c+(�4�n�g�~$�#����J�\�ĩ�$���
&I�l��An9)�Ǚ����q���EuZ�h�/���qi��e@����`��:����IX���Ӂ]�Y^)�wh}�4��@�~[!�:$6
)�_�9��RQ�O&���.&����kf�3�R��_�������Q��W�V�Q%l����j<��V3YS�i^��D\h�]%r|���#���-�^٢�
/^�p��E�llU���48�|��n��):)�q7ƨ*]��Uvh�tq?��r�����ұ�p7ɚ��8 �%�2��"M�}��v=�_�Ӄ�Q\����®J�c��z�b�F�^�؍�)f���\u��/w�T�̜$�P;���!A:?7���[�(!c��o�~�CtEʿK�4�v�W�r͑�gȁ4�E=��ۧ��Z���7���Z��͋.(x���W^�e赒�y���XO�0Fh����e�p:ň��C���_ZB�W��	{���c���ϒY���M�Y0:�I}_I���C���EQL��P[ڧA5���ҪS\���B�Kc�"�m�҇\׸���x����q)9��70d��^dmE`�a0.���/�O9���D�b�),YW������?�������izh�~�S>ę����[����ϭ�����A�2o~2f�x ��96v�:����PSPl���s��[4��|����L᪜�� t̄��F��u�ग��.���D���'��υQ=ۿ��(�	7�PQ�w��f��n�*'%ֳO��b<��ҵ�y�pDs?Ht��;0$��ت��+�h�WƷX���Ё)�%*`��ጝ��<E�6�3�� z�����8��)�.���p"�%�A���磛N�|�T ���.��4�T�>j�>$6ڙ݆mv;�}u��f�Wu�����%D�8�l&i[��>!�ݚ.���y���X)�t�
ѩ��[�I�� \ψ,\���$G=�ҵ�����yB�ݜAxv���"�cr�����d�	AÎ��������`Y,��v]CT~۞�by�2�AH�3��<�D��|�&�3 ­M��o��G�0�b"�M���x��4�,	�����T�U�$���m�(E����/�go�|�6ܩ9[Egc$�M�}�`*(#���E^Q����^/�M%��pl8��bR�զ��ց%L���q�Ea*�C�	?p�w�L�u� q{?��o��̏�k.��m�B�BCq-�f�F6?�Ţ���h�;��
��2QMm�cb�2�%S�c	O9��7�5�֛�� ҫ�*Wr<�t]�yH/���m1�Lrte�ŃkG�����Κ-m�s<ZP=��I�(���<�r�̻�È$�g�zo5^0o=!D�r:�����\��%"��ϯw���� ��n�w����˜�I~��Ո�!Am��X���!�n��>�Fmc.��.�S���#SԠP�1�~��������at��M� &t�����e���k��#Fwpka1��!��[�T1�;`zGMaI!P<�h<�)�E|�vx�'e�T��z����� 8㍥d�v��dq8ލ	ڪsGR(U?��ʘ��ek�\��:̣��(I�m�t\*N�w��>>�ղ$��īK8;�gf��q�b���<E�A����㉡�)�:��eV��y  Y�u�y�/]H R@��*���S0��08�� ����tU��8�2gӥ���������Sh�
?�w۳e�{��/�t:.9d�؞^����'���C�����Ȍ�Ӯ�۷v�_�����Ew��S2\��D�\�%��n�����ϟ��T`�H�0��'5D�x"�K�iLR�,�ͩ4��Z�:�=�}�:<���qwܱ,�����Y
TmH8ފO1^��z��UR�Zk���A@
�{����z�t*�a�V��a���5�P ��d��m
D��wp'�K%Q;�M)	Va%�yf"������T���u䅵5{�5�~X D�Ϯ':�����ͽmNּ�r��߁p��:�6�p �o�+ ��oC���ܗ��������D�Wq!�C����)�@����K�y$���D�n�PlȰ��F`�1+���1���J�-&Lֲۓ��ج��D�fRb�	�U,�>�{�ۊ�PL��ů��LH�E��BPQ�5���:�����ݒ�>	&��S�ۖ�g�rw�>E[-��N^���E�v��׼l�6	7���ߡ
�&q ��՘h�l|^Yd�#��������3O̔Lt��y���t��O}2M�����l�h�&ٓ��rl�n����H���i���]�*8Ԗ��[�9�-�μ�D�CDm#�H������7�]�D5�43�bs߹
���5
uhc�%bipy�w��+z�x�\�s8�`(
'�ץd$�s ب�=:���l4��d"]"߂�ns%+��5쩎X�;YUGP�2�Hf�I��ݑ�+�cV�r^�����ֈ��`d���q���U�˒�Y��z�v���IXBy.�40_s<�NQ�S&��?����pH1�˯���Cbh��	X�z��w����˄�Y<����rBT	Z��^!�V^#	�����[̻;��9��l~��-!Uir����ċ����G�}�<�5�8���ΖSo[X#P��Kϓ����(��hE�wZ�3���dM�c�!�N}j}�]�m�
�$�޶�ۃ=�:dH�+5���GQ��T���3DS�΁mIj� M0)H�zF�����a�W`T�tbT/O�J����dHV�-*j�YL|��𔥏s*��W!�b[3kx�-y��r,����P�P;�+�O�tK��j��ZK�������E��{���(��|b�qD�&�R֟�C��GiHT��S�����~4�|P
l�xlďx2Ć�����8\�zЎ�$�-	��52�!-l��2d�qĳl*�iK��+o4ӫ���R$a��J�j���dmG-�1�C'4��\� [���J�<)O��Le.�7�10���PT�\�Z�c���6[FL�hĂIB�����?��l�+��
&=1�9�����r���G�j+K��B�1���ϝY��6���Ϊ$iL���{8����)'vU͂��j��Ҡ�L]_����MI�0�&
OI���
et�( ��4��� t0���ǳ��c�f��=����e�?��{����#�y���ͧ.���b��?)�:��Y;q�]�T�Knu���uO*Z��)b�v����&kbBG��[mo`<6���C�r���^�X:A׾�T���D�!DɆ�L/�/����sbZJ���v���&�\�:8�������^zo
$`���H��y[�}�� gz<Boc:aC�K{�׉����l���3Ƌm=j[�{ې��-��h�YBh5݌�Ǯ{ɽ��4Z��iF�6������wߎO�������Y&�n��I��͡wV���8�i�|n��M6hx���\��E���<0��X�=/>�Nz�//Y+�hsu�L��p}�	����@��؝�sy����6-�� ����[�-i����Oɜ�Oq�P��r���:ٮq�uH��h~ј�?��ٍ��y���"%�5d�2�FN�Ǟ>��� �U��z+�����\�r�)�<�o��^9:��vr�4R�d|��mfF�Ʃt���~���b�6$/����B�K��na�g��6]���27W�mv���}�Hd��w _5�G�0�ۋY�p�� մ���D-7�l�)b?-l���{%H&7�X���@�7R���?��ܽl��X3���첻�Ȗk��v�i���]i��ݿ\OJWQ���k/�GMm��;��E�6FwSx)�L�N�ш�m�V���_�c+�1��lKýq�{g���;I;ƚ�>UJix�WVh�d�m���H
����K���ާ\���ma�N�/��uI�"��;s�0$�0ep(@�I�mKH�+Ǌ�ߜZ���]�\���i�����M�g+~����g�����!trvl�R�3V����>�4�=��wU�g6n1&~���뭔vY���W���� ���23<���?����jMY�#�غG�GEx�����W�I�]O�q�@.�I�}�(�R���ɏ�ZO˿��x�Q���� ��(Y}ّ��V���;�@��V��]��K��$J�Y�X]F8i�L��p�袘d����I,����i#�h��I3�e?�MP�l_Ի/M��(]�݊*7NT<����j��s�M���_�Ԕ7��lqn��蛘���k�������)@�ç�r��l�˼)Iv�=��Τ��Ŕ�n~�x�Z�f����L�ؿ�+�s~��D�_�,ƚ�xXp�w�N���+�	��h0��n�Z�3�Zh݄��ds��{uD��-t�Yӓ6����8�w>���#gz���@��(�S�_�(�2֨�ֳ/��u[:y炵n�� �/r�fd,�,ბ����S2�UhB�k\�H]SDM����=��7j����z2�Rc�B��������β�԰�(���`�zf�F=�c��=��ĬX�䩴V�o���2�~�H��`���l��xa�,�@���8�lV'L5E.L��2@�Q	��lY�0�Â��>�|A��2�̵*$�������b�l�Ua�t%��D=�#�U�}3Lz�@�N{:������o�K9���,oHޔ�O�q	)6���;Cࠁ_���Jݳ����DhC<�+�͖��*E�$�7�0]m�CъU-�J�RlFy�t�qC��3S��vc�{Fw����ܶ�m/�@�fԝ��˂mj����9���5�E�3^2�D�L�u����2��mT\��L��� ���;�%8����g*iZ���Ό�񴰬Q_��T��� 1�{S�r�R@y�Q$�ͯA\\t�{MF�#�0�wq���H����9�On/o����������J���,O���Xx�/��5k3���{�
J�q����"
��t>y�G|)� wJ��N�x���gd��l��2���u���X+
����v�mic�DU�h͐�Ѧ�[z@�F~g�R<P��y0���ő%a�|��M�/�z��W����~\���F��2	�D���p�zd#�T�oQ��%��Y�7X��	�赛@|�D{{�DB��P6�2���k�vx�#�Qb޷9b������ �[�97/\�gS�yd�D�[�Ԁ:SC:���%�2V�ϸ����]6�&�;���lc�L`g -�A��ˁ�o�x��8,�cvJCM`D;�4*Z�_��tHF�u�6�'� R5;������|XQo\F�Z�~q��R٧}G�b����%����q{�U�J0��~-/��8�&0�Z�j��hr����A���h(8k�C����%�\p��F�-���LP�+��5������>g���޲ቺ�5h}ƨ��tZ�^QE(��� �6�S+�D�C&�_���i�#��QGP2
-�U� pp���]��H��Σ~U�["�UNR?������r�fr����6�Th���'4��Ayĳz�	���,h�g5>y�,��~m�����]�5���{�I��#4�c���� �>�
����'Vܸ�-�+67[=Y~^��V�Z^VCL���k�.;bϸD���xx�b�p�hZ�{�ߺH"�sC�	gm_���٪�(^�R~L	��G(�2��4@l]�δ^]H��ܑ;?�Z��IZ� �+�;!�����"��ٞ�Ҡ7m�sj�P���D�8a�~�3������q���&\��,|�ٰ���+p�j���2?j��wz���n,��^��*����?	Mݙ�D܏�,�/{��oA�0ݧ=�$�lC�&-;/�,zQI�ρk�Yă���x+|�e�dJD����*�S/T�Ŵ1��ޖɚ����x�Z��18�Ε`����xT����a�^�Ě^������1鿑�M��rߔ�S���Mdd�\�����Hh5{�j#s�g%��TD't(˩P��9�f��]��9)���EJ�ȍ��+�N%-�xd}��m�?b���2��:_}1p(�M(=��.���M_M$�S���*[�%p�S><�:eHy�����@k�+ٿ�Խv�F�k=�ynu�^�n�a��$͗&���e-h ��gHٔ�F��q=��0Œ�RW�+�_Q���&����WF@mad<�\.P�% ��,�E�Y���?��/m)��3�u��o�jQ��/�-�&��<���,��8�.{�~7�Ҁ����b0[��UX�����9���Ɯ+'ѭ8���h�.�0��'�Hʫ59v�,�h�)�vH�r��#�#8���{��)�rU���O����SZ�������B�	"��^��S&b�9 ,�19O?�b)&4�'b��aϏ2��w�vLo3x�S��g'�)�V�7�E\�OR�� B0J-��������E+*'9wcpY�N����H[�+�6Dё^��ݣ�6��G6�5Y�#�Z�`K|rn��(�5�֗���RԄۧ@�߽.�'�z�p�ͧ|T"K�`�iT��{�Al�O��ڔQ���I�+��
�����E�R^�#Ym�O���@Zj����Mm�����R��%�3���)DEz(��T��"ͩ.T����x�W!Xs�=��b�|5��=v	k6-��m/���|�S�lK��?`���h�|�� M<�%EdH�r��,{<�Mi�9p
�D��:�5�������/�����̭o�D IA5mt�:�G��0ɚ�;�\�jr�v�'^?E� v��E�FW�Q`���,��V��S�( @A��>@F�p���-~��/�Įt�f��M��2ZHب!ن�v;�d�\��M�%�f�@��߿V������h�j~g�1F7*F��!4���&����c)З�(�D��ɇ�O��h�L�u�ߡ=�~�2����G\�2��tlo�T+��KT;��^�Y�����e}}Kx6�6�[� ��=#�t�%�z �wm<u���ރ�FS�%EYw8K��$3l�� �4{r��?VH���A�{�����b�(��{�.\>K�yA�a{6I�p���o[se�VU�T�͔���2	h��x�"�0і��d7�]�4��~D�p�,�:�XD�䴐��˚�rB��2��T�p����,�y�<�́�K#�x�D�a(��u�5'U�=��z��qT�Q�>��_9� �s�2�r��F�Ȑx�@iP�b�������1ħǐ/�Z��_�����M���^����T�B왨8�h3�n�9��O��=,�Z#q���,�O���:?H��vy<9�y��%2ś%�˔=HO{�mؗ�W�3��{~�⏏u�a,YiU",�UMH��p����A���!nO���\N&3�O}�'g�oV1���r�դ֑�E�zm;?K-���kcM&\�N�����j��p�֑��_:���X�p"���?�i������1�9��2`��̱����x@�\��p@�6r��h������^@1�%׭��yQUa� wl�q<PSdO�s��j��W��Lo)��F�3{�U�$����NE8���krT�����<���Xb`8��є�syk�3��rY1c��(;U>V���-�_�?RH��p���!��j'%Ń���ZN �R}�\��4>uE��B��;]����0�R�� ��'��Ll�K����/���p�r�@0��?��Ֆ�3�L��FX����[Td΍��{v11r;3���=�. �}l�k|���l�A��,�^��򲈅���fꂹ)��]CpEU���m��؜p �)��x�1hYB�Q�~�f-������S�g���;�Q���y�>�� !��u���cj8���*at?�Ǥů���/��F[0��	t�Q�u��`L�X>���P"�G��?8-d^-�\���C�>��}��]2�r�01�z�:������s�F���B�}��R?xi�9�ݐ�W�V�܉�k�{��@1�7ʚ�1�����d'ڥ'���Bʹ�JfZfq�
�Q��Ay���*;��9�xzG�8�<��4�I�i�\]�x�q�btZJc��z�^�kc��U!�&�@�a� �{o��18ϼ�^��OJ�4�NQ}����M ��}@�d<��dD��)i���e�ξ<����sk%l�"�!-�h��6:W�U<@���9-�B��+C9߲�*��>�qD�3��D3��8�n�"�]�g@��0�#fM^�*I��!���Zq6oK�(�"�Vl��
�ƎZ?��Yn��~��1�u���\��;J��M�ax�'�
#�")�2�0%��.��=���`յ��|��=a�[]�驴3N�eW�,CzU���fRr��o��-��g�5B�<99������aS�|��?�\�.P��?G,	�p�2�	��ͷ�d'&�;�%��a���`B�<Xċ�c����%G/���N 73�A�g5P�A�TG��K��y�F��/��6/3�#�����p�`������Ip�O
�觱��r��wP\�!�C��+R�Z�j�"6&��6㏐-�������o?r�Lc.6�1��7���٦��`1�U��g(�e��\��?�Թ��rҀ��=��h����E.�����C�&���1>�/�Q>���q�
��ߙ'݃%."m])X��������X2)q��if~jqw�f����SΤT�H�I��f�VW1�9���<��+⅏���\>/�(�~!���Rq,;�ﭹ�1�A��	��V���A.�&Tu�2�y�z�B����<�9D(���ռHc�Eب҅��LO,~j��	�Ý-ns����Z�z�=��.4�-A��6>dF�Y��ᕄ#����B���/����vqOJ^�o��8�����-R]�(Q�Rw�
�_v[
�Kc^T'@B�SG�?��+��'�|��ӿ��UF�l�F��Yf��G�F/�?'U��a"�#�d)��_̕o����
H=��a�PmD�g���*��������]��0�Y��f�yf݃��u6Rr�V���x6��3�'\ID�$���G�w���M���O�]#���&��(7\+�������(���ك�*A�����k�������)���9n�/,�S��N։5�;��U*j�J�u��}=��k��`�9!�Z��y�&��4z2?q{jO������4�"��8n$�{���
E��`t���ϴV+ +��:�xU㏛����!;�g�����N(e��'<o�$NF��*���J� �1�-�J�?�C[cO߽�.�7�~X{��k'�d�M8�ѵ�`\��2-j�ۋ��P�!<�1�T�2!D@����PE#-���r�� b�s��3���6��Q7�e���}��R��.�7�vd�n���t8�ì���_�5�p-���B(�>?)T�1Y���S���_���f�A���m��g�(�*���,7tO_��G���#��i-��_WK�������D~��sa�ճ��Y|���Њ��٠�a�8��ܺ4ס�H�{�D	`��^-���)����B�u��*�1��R��a��5g�X)E�y�j?m�$,p��0!��h��;����2������wV��^[���>�Jq
J}%�ͰɼĻHk�hAx.����%x=���1�	곎e@�s_K�g�Ӫ���"v���j����^�Em6���Javd. ��J�������fKt�~��e�a�az�Z�Űgg<`Vfd%����X3X����z�ʐ�.<��M�k�yp=i�![9.kV�Ǘ�o���ұlK���z����4r!!L{�9C��G.B���;^�=� b�1q/�hq��*�a��t#���w[���,��fʿBW�oó����	ћRa��C��
�7O���e��h�õ���,8h������H{%����:�q ����sM�׮�Z��x�C-;����E)���S���Y'iVk���\&I����u�be�	�{��b!�pt��K�]�>�q�t��}&Z����VDnɰ��{`綐�(�`s�[3��S���巬�2�t�OmkU�Z����M���!Q��Z�Y���|���(�|0�"R�k�Y��rmRk�i�n����������VFU$�+_<�u���F�Ś?���>�4���9_s�H��/��U���ܵ{��6w���u�/Ӓ�� W�Y⛚^��k���g�<�J8�K啲cl\�?e��H;NgOw2yz���ep�����TC>	6gW�4����뤔�,�_y�9��	=`�'/H|��ОJ�~H�P�}Ĉ�ny3����"���9{j3��������U��M�Ԏ;$���;H	�0c�%��+�N���3���/?�r�~���r��s5���%6����l��mc��ߎ`t�/����0@���?����~���o��3bB������73w�]м�g��,z�����ɠ�D�:�w�az��)U�Zn�^0%������+q��Z���.�o�� ��̺�FH���	�:�F��2=7pv��֏P\�$%��H:�ni���A����]��M������HL��<Y����"��-��w�֟>	�(n0�~�R5?$G����p�v �ݠ���_]:�ǂ����-	���*��Y�8�x��q���v��f`�`ma�\�=�N�l���7��j�vθ�s�Պ-ƚ��ә�lO\Jy�[֦|F(�0v$B]q�e�R1E���/�kS�<�RIyo��c/���)���"�-,KB�m��F�*�9��5Ƥ�w�0j雏�9I��줣��F�ҹ�H�xW?�����Z�V62G�V(�� c����榲����6�XnP��)��u7��<��6e�=�K�RbA����[h0��fc��e^�ǲ"��u.��,=�y�{���Fo����Uq�����ю�\�m�ӑ�3��A�m/�Gf��1���̐s4o��u�6�h,斓���)�5�����zڦ�9공0���G��_�����	�E9����aQ^��|��#�ɮ�O���J+ٚ�X�����L�
�N�W .�!M�g�*�S�'��oT�i��;Qz�Q�2�$l)1/U���D*�%` �Ģc�*T�+��ԍp0��j�z�$�]jq�I;��ک@��A	t�^^O�v�6��)�X�������P�f��	n�+Փ�0����{Ҡ��E��B�bKR�ʛF�h=���<Ag��`	|��@�c��NɊ�=��_*�����	� �"�h_����ʌ��+0��\N\.�M�E���&m����E�:��H�r�O�b�T�?�|4���z�[�
��B�_l��g'�.�I������8\���A�SHԺ ld߯_iH��F�\�k ��$�|@����HQͥ�gf�=�x�-q����E�+��Fޗ�Eõ�_��O7^��3t�E� 61Vg̚�w^_��J6����B$��ߙK��`M�(�|%��F̅�S��"�tp���@�n�E�j~V�4T��Ur��r�c>p�gO ;���5���v�����PT�ާ��y"3!:���?h}D��(v�a�N)��g�'�{������Q���j��F�ШgH��ֆ����;�Qs�A �f��ҤHǓ���_���Hv_�����%���Әj��+}���:���I�����7��p��[�Xy'���kػ`иI���_q�d�C�'��\�Q��U��KWk����mL�l8�W�]쀉?�L2%��'�uL�*��fH��*=����[��Ff5zf��.pawTi��W�/E��_=��l����O4�N��V�Րo竤R٠Mh�=	� �ԇ� y��h���Fa$��Rٙ	����Z��X�5N~�S���fN�^�&l�
�)�!���%h!/��Q\ɉ\�U��Ύu[������:А�m��T���y������Ԛcv�q��A2��kQɲ����{X�3ԕJ�z_��`R|(�W�ϊ/�_��4%�-�����D�\����O��Co<�l����ڥ1�e�ە~����<����?�� 2�ͻ�&=S�&-*��\�.����<�H����j9�^g���Ŷ���^K�q�	s�?4N��;��ÈeŠ>��?~���r�͛�8�����zo5)�	,�x���>F�!-�~bi��GNq4Qy<�"p��h�RZ
��Ӳ����S���<�����o�����(��T�,�0�nv�C�pd����ox�^b��U��`���&&�k3RK g��sD�֔�H9Qq��c��2S��H��rʒ�<�X� ���x8.HS8�2���	]����=���ZZX���n�g=��w�9q�Dk�	/ �D9b�I����X��آ�þ^ˮҚ)�J�p;�99JF��~+�z����;B\l�%��Zt�S��(��7>�{c�I�N|�������A�"(p*�s��X�2K�]� �7橹��bՔڭ�d����Ԙ��d��t6�VeZ�U�X��XMt�n�*�Җ;ʢ����q��/ēB���6�%%&{�_s��k@$�2�G��@!��t*��v�)d������ư��=s%�_*d|�@>�x~�ZW�eJs�o ��?���A�_������K�#D�[�棂��8����5���Z��qY9��J�,�	h�ۀC�ר��]���`�� �#���aA�
� �$i�{+>��e&��8�C$�d�2l���v���������F8�^�PS�Z��r��C�%�Q������:��]�G� �i�$�z^ю�^<B�|2����pl���Sf켹 _�yƉ��� ~^��o��u�S{5݀�Oz����J�·�e����7�S���}yv�<���J����"jWԀ�G��u�fL�^j˫0�Vk�aj�kK��`Q�6�W+��"{NЍ���+O�[l�������4CS?m��L)c^�����Ő�?���� |���l���K�-����s#(_y�s�,�H׉k�Oή@�x�&���].W���sĸ�yPS�����Pg� �(b�}q̦�����I$ۮ��<,�o���o7��ˀ�Ꚏ������d0���ʌ�e�x�*E{��8�M$��Z8 �����dG�!Z&k�iG0��܉sgc���DP���δ�s:�����A;�Ȓ&�+;j�B������s*�7�'\�{z�I�|�7�UKju�(��
c�Zʩş���W�:�H�F�d!�nm�L���.����P��:�N3�ء�
��1�v�kO�R�6�(�U.�l�B� �\���俳��s�����D{�,�$�^�������\�V5�)�l��vZe�b��]�S��)�f����)�`p✇��L�,d�~��r��]Ɨ���VD�������vo&��/m�8��]�U'2�����	����$�sRKv��7��qt�i��Y��/��,�B)lV��*t���?�;V4�p�R�@�x��4�Re�ƧQ��6�N͸�*i-����0�7x�q�����1g��-��cֲEf]��9jΈ>�ys⁗����C�N�QA�D���P�[7�9�El\��U��˕����o���o��EF�(��c-�y��
N��l��?>�fӚ�3>�E)a_��q=������[8p}�(u�����itڂ�F�L.]�iB�%�y�T*0aH(�t!�7�|��V�	=}y��A��I�=+g�|�f֧Б�2�&�\���vK�?�ur��e�8ʫ�h`��SF\b=��k?��%\�L��T��W�s�g�?T���7!�0���7M�m�����8���q�3���E�waah2|5(,0��S2���O�m���9D�w�}�83����,�|.��%`�����z V
�e�l��)��);�0Ql������ٜ�5��|s�>3��@���`UF������p�6^�����y���Ҳ�F��7mn�b^/I��G�M� ��6��L��I3V����`���4����7�,Uɠ`}�H����	7�&R��\����J���%��}�[�/�t�Za�(m�	h�sZR���Ƶ���d��r���/��C��[�\�趃@�����?1+�%� ލe�U�Xe�9�?���̅S7�z\�ޘʢ�[6-�_���ʹy#Ԓ0�v�H�V�- ����Y��#���ԍ=���g��=��uߝ��*���+G�8*�t�\[a/�8b�|�N��9s�����"�:��4O�I�'쾯�`��CȇUL@��;��2�͞�;��B�I��������̉,/W���].��d3	��90�)�0>��7:*L��Y�� �2 �V��ₑ!X>,�j2����o����N�ݱ�t��s[�h���Ȫ{M̹e�F�z���+v	�~�bJ��6���{DvGmc2��rc^��#6�x�Gp�V���W���(�:4{G�~����<-���s�-Ck"%Rѭ��@�/2��zX|_}���9��3fV~(��H�Ip�?�a�Js����Pz绯$OX��O6��i��c�-���YA�9k5����˚��� ����+�zj~e'm�@4��_+o���O8��[ﾳ��m��������+�P�j�kd��c�0������z,u�"!���z��
��vl��D#���`D,�:��f��	`H��/�C�����%EZ�N��t�*�^7b�ŧe$��2���������MD!~���_��%��um�K��5�_�u�R7P��ml�[^_uڃ�7��$���̦�j�0�X�M��͖��TB3Ϳp���#L��
�Tg���G՞��k��B^W�D���=������AG�&�{���:J'�So�%k�F�p!:�[��< ��~%��f_A%�AmK��3sQ
�����h[x(�r<on���%����nU���~(�3��"WU��������Ñ��ު�G\K���沈=;l�q�R�#u��HۼLq�s�;i0a.�y���)Il��sl�7]}����͌����k=���-�i��ȍ�7����ܔ�a�0i��wC��������0L|rKs��g*P�����zk'ٹ��-�xeP�nч���Q�z;�e-��=�]�ɀx��310Cu�%�&��׿:q'o�U$��D�T3+P]ưf҄�қ ��yl��;���s2�S}
������mH����Dc4�`M�E��:BK����_Y<��p�?>�F�g8ɼ�э�}J�Q���S��݂f)G�<v,fB݌_d���3�׆�Da��規�%���TW�)\^���~����I�d�|���H��������Jf���lV��Z�'�@^p��?��)�ie��Ԑ����謵�,�9����C�.W�\4�P
:��8
Q?�* �=��[�ĤƊ[�m��ص�a{��y�A��QNǤ�
�/���Kk$���s���Ħ�+E�r������p��.�w�^�5�R�8GA#Im���	kw��U��\���R���/ߕ|b���W��*%�Y��C�U��{�� ����6 ����������K�k�x-��;��h��7�s�.%��?��,�L�6�"�:g)H�[芜>��+TGL�&�m��\1謲�A
J��mf��G�?�qmI���o%NN�sQ{������
ЋM������7���w��6g{�2�V�>�|�|��7g8x�T??�3AP&c�)h�[䚟�4���Y���r�z����z��,,N�>�$)��N��2�/��乏E�rX�,�@F�/\���B>K���b<�+���7����@�aRCt�tq�'Q9AE����)\!�麄6SV�͖i���ӳcP�xU���`�<f�-C)L�Zx�Z?\9���m�.w���Y�d�dC�"NPEy�"I�xs�ς�s&ھ��V������`��o̪M2ƈ[r�1y�)�=�% �%Fa0�d2L)i\��B��O��/���.+:������D2L�9�E;g�.�K�Hy��?^F��1!��|D�0<g�'@�f�2��ɥ N������h�[,2��@�Ļ�<;�!λ�i�)�q�e�B���[��4��"K�Y���F��݇����rI��x��G_�҆�̜!��t�f���݀�L��3��Q;�]T԰f��	���1{t�!�g�2�t\�EI��Dm�`"N���D�&h)P��ڽ�PD��޴��b9+�Q*K6��Q�D�N6�-�ت��n�):��uf��y����Y��� qpY�F	X��|�P�&�0�{��U��B@wxp1�l�?�p���>�esSM,q�B+�C�As�ly�F�g`�: �}ዼ��<��M��ھ}}GB��Z�h�;9{� ��
�HY�	��R�Tw��Ĭ�׫�Ѥ���㡡M0v���{�T(��D�=��\��h�$B��ý�\��z�;{���f�	mxn�;�B|	)�ʻ����v#mh���9L�Ή�)!��Wb�V�;�ൺ�g��z`'���l�:�!�<i��Q��g/]o���B�.Q?Sj�G�M�|`����c#D8����o2�F���'_��0�;��1�{�|��q ��	�s���J3P%�-	� &8���#f��Uf�633b��<i���y�Ҕ5ӑ�<5��JЕ|���n1��j�ؑ�'U�
t�
�i9�@��٦�L��>���w�����S޲5=�>���MY7k��Z(?ơ�n��:���Y>!�fȣgN4��^
�"-~5�8�VE{wl��vH,�͞�s��1�	Z�LT�=������.�4�+]���B���<ӈ����-���%!��D'x�	e�g�ǈ�JuC�]����{N9���k�QLOl��V��ZA��t���������N(P��}+T6��/6�q3�!�+oG��mYq��z�_��2t2?[�!t�t�TY4�G�BV/M↮3x�Cq�
�*�8�5��&��xdX��|���"x� h>��e�i>H�9�F����
T3P&�[�Z�^��~����� ���e�N��mRcE^X��"a`U#��2礧G d.�.7��N)=��)&X��Ē=�Go�g�l�S6öm��c�LJ�$!X�\6�͚C�5�>:%���p��y����H��m� �T�S#`k�jv
��D���ßakR�D
v��$ ȸ5�-�d�'����x=~l��F�]!����?��"���HD��-9)9,�F@7#�PgmUV��/�v,���Ա�Ÿb�nߠbUo.��7�2����G�%�}��GZ@�C���r�uz�vE]��\�l�Lv��T-�������@V����.�\A�-��S4�F�}�Е�60d��p�sϓ���0 	%+=zwv��s�g ׏�
Mbޯ:��V��ol�`�i�`���9�x�u-��R��0?�ツ(m�3��p['�	j�c�Yr�mn��&Ơ>��M� AX�&Dq��	�D�\���.���Lh�*\�5��H�ba��=���s���:�.M�-�� �ȩ����͇���{  (c\ƻ1��]v�����g�`�Ժ�@`��\���nubJ�+pC��:'�:�ҡ��7�ƱpHK��k$��M�
������*BC�7K���ldk��*Ѽ�`�tO����V�2����sh4�+���A��~?��<�Y�*�][*���ۣj��GP,$r���Z3A�<y-�!�������	A�U��Ǐ��[����*�Q�� c`���;_���={�2��m,̧��%+�{���⠽����k���R�����s��.�㫜��5j0S/�',a��ϣ�^�4 pHi��֛�W�z���^\�?r�n����lS)Mi_w�.%�عEf���1sT躉E;4nВ"K�u��������׸5�c�F� ��0���ar3�X���0��M���x9-�R� �4op��B
�[����9'e0���>4��=�{�����X��h�K�&i�nS��vP4��ס[N��KiX�Go��C�N�x�28cwY�F��ˆj�߮��n���2-D��+=�4�9��Յ�p��i>�י�Rt�A��4{Ϩ���P*A������7��;r��6��o�	��7����&Z��e�/y���⾖����j�ڀu��$��ڳ����%��a%�L�Hj}�w�b��[ڔ��с���������<Cۍ����gr��YG>ҤP�U�y��F�O�&�ۆ^R����[8Ύ;4����&y�g�²��[A�$6Ge-$D��T�.��{��~a�tZbY�7כ2�y~:��WR�H~����?�Q���ò�`Ը!�����^Y>�����E�9M���v�f]t5u�+D?3{f�,�I��9�tVfs�^[r�m���� M��|��x�\�����	�t:R��boO�)U��ڨ�m�2J�Y?�ܙ�a�����yU:�	��8o0wS��	Z�m�L)+`A��?�(�~=��(�����+�4�$(��"dMh���6�����������	�>�h�j�܍��
P"w ��[�^2	��q@�1el;�`l-�_�
�I�Ӗ�$6���W�����_��囜
=���ru�
w���>�ՂK��#R��[b�-xJ(t��uss�/$�����A{����`����y�\:+�E�9�.��ۉ��,�;׸�'Ȍ�}�Lzj����%bqg}LطT��k�xB�(T������r�����'�k��C�hU��wǥ��?.$�����1<ۑ�u����{r��H1w�3p��q,&�Ȓ��-�[��BB��:6[�)=��zgy���1�o��گ'v��T��ء��1���>iUR?(�����sf��Wj�<o 0�z;�!Y��lG�uе���xQ�/}}b���l�N��Pm�9��:*���*0��E�8�#k�7y'H1'_5�"t�[Ys�Ɏu._�^U���o�Lu�! ��'�A�.�-[�B�{��$�&��"�K�\� ��8��.-k`��k� ln ��=�J�i�QkA�u�:�xWР��}����gP��/��+�m 攵y�Cp����cDJHm��;�2��;��XAQ��^�nHj�d�:�J��I���V��_���鶇�����K1q���%<;��޴]^lda�s�-iS|{Qb���qo��;��w��e�\2�1��V՗T 4|f�/NkC����O	h������-ò���ۜ��U_����+�q�!&�vV�.���.@i Zģ�<�x��Eǋ�7����9(ƌ��p�
�� $��Yǡڑ�nh�&=k�j1�Q\+�������nX�'k8�0b;��L�����Gp	��P��8�d%�Wj���W��۽�gQ�}Nkv�/�-h�v�u��-{mlF���nSCO�8�v�=����E�b��ʞǡ-#��\���	T�j��b���������sc�����K<?<��E����l,iER7�-�W���2�5'�7P+h�5�a�X\�eB ��8�v�y����o���[Ւ��A�X��C�+'�[��B景�w�3A�|e6]v E��U���X�l# '�v����E��p��ib"�g��5��uz�A�+$^��L����hO2*�a�� �Z<��P��E�k��ntI��$}�v̾@R�A�U���������fL:�V�UD���X���=�ݫ��)�DH��2�&�� `s=�O�p`��j�8Y��af̑�Yj�j%.�a8�*`�?D���V�X�I%�N��_�[�5�%,XX�/�6�o�C`F-��u�w.p���=#�3�70= w���˜1�Qđ/d0l3^K����M'_q����/��#�Y�"(?�caη}_G�����יYGN����ܑ��*ٖ�*D䡅�Fk�]��u�u*��J�K�!�:��-�-�-�<�_�	h�'�ḡ�&���俇�v^U:��
�p6�\�A|�f�=�!;3�CE��_������p��&�ޚ�6��pD�8Q��a:ؾ#���R9e8���#�!A�%�[ٺ�"}�EB�Y}F��c�;�6tA]}��Z��ճa�i2mԗI@��x��}�Z��Pj��y�.�N8�QP��e������[I����pӤ&�_���/Y�~I0�S�2��,���8�� �������Z>,y�er�%�6�i�i�o�N�r�U��kuLs���ESJLA��WA�~�xQ�/�	��	G��/�a��O��J ��W]#m�9��̲�Qڂ�Zˉ �M���ZٵH�S���[�j�w�%���P�Q���i:*��f�$��C���I�_NP��D̖<�ІF���5��ր���,�!�VL��9�+�{��$yU����G}��R�T�OS����B��_u�~~d�&˕s0��i<EG��q]�������8�,A���|MϬ�W��7����ۘ�u�a[v�K`e�>���9z}e��+O��7u5a�E�����rF��d�o'�8����D��1��z.�hP��4�x/\�Ӎ��-V�:K�)Yͣ�˃Ra�R@d��d�j���8�ӄ"��|:���ʗjq#,��_/�f^ޱiQne
L8_�	�$ȳ旜T�o�`Z�XϿ��x��X��.�ň�kg��婱afk�54��~V©Mq}�d6�I�ۏS�h!��]Ҏ"�R���aۮ N��ߝ4���|��_9NȨm���h~4㧣O*{j�̢�k��l6�U��� ۀu�y��0�Ͳ5��]� H�4����2df7�\��b�-���ZW���먄��m8��&N�ဆ���^�cD7dT��_y���x"s#e�'������*����>Q`0vۣB^�@�'�l�+ڇ��s���CG?U��ң}/J�M���t�qbј���H��7C{�iB,�Tm��_n�x�α�=�Y��ݘ�)3���4J~�X���ma�e���(�8w�@��$\���z;?��<��5��	�,��q"if¥]�'];�G��e�p��iH1�
е���D�SMi�H��������̇�o�%(oG&v^�8�״ZN�*��uDq���^��.}�3܉a}�P���`8?�)����Q��k�Ѓ� ��z{�]q���Љ�^Y������_�ta�ۦ�Jٓ����Uii�2.3��&^�H=g�um�.�]Х���X�oƧD��0��O�;��t��(����������%��^� l���U8J�E�f��?�E�Ąw��`R�_W\p�����m�hZ���ʆQ�-�z�[�gKx�|�J���㊵~|���mx�xI����.Ez�*)U��>У��Bs;�ge�*�����a&��PZ"�I����nD㎘ �w�L�6���ٔ�g�,����-a�~;g㠜��Tz�V�:���П�*���IacԶ.p�IW�s�˽2ɢCoI�k���q�h��N���Q� �(s>�Kt�j�[ꙛ@v$�2��gI1Ϡ(��� �\�%6�&�}5��y7������nV�Oob7�$�xp6>)�de�|(.m��Y�~�*�'�Z��Z,_8'�{�B�9�AA?$ ْ�u$�i�E_�0K Œ"V5XU�?�:r{�Zf*�� v=�8-������5D܂h��G:��q�@���Nr�c�Jw(B�i�;�v�{�q�]Y
�&T�I��H�Ш�����Ip �L���4%�2(��\���ȀRs�A��q�Q�,��<>48�k %�Z�!�lϋ}���`qZz&%�d���۸��\��!ߑR�"�9bǮ�k�VLq2����׏^��X0����`�ABEC��
������z�E"�lh42G��I丒�Qd;9�"��cɸ%��S7���y�a$[��
-��'��)�7��!�	��D!b��`(�M[.����oXD�o�s=��B��G�b�1u��s��9��@�����apa�*�j�6����8dO���T%��k������Yҍ�v��NS��"�6z���s�h�H�V�4+�-�sm�;�L�˗f��g�!�ʹ��]��cߧ|�\�څְ2��uZ��?�!�Jn�U����9A��F��[S��e�k��,�"F�q��Э��0�F��y͋u�/B�R�w�ޚ�~T�U,��]\��i��5�*�ރ�_�b�O��z'���4l�vO�!�ͧyfs�%omz���[��h^s���F*�%�r���z�<ڼ�}����*��i��y�=����H��lq3�O3d�#�NRO`s��1;k�Iw�1�k�Lcc�K����#�ayS�Ԥ�?|,CJ&W����eu/҇��2!���i`t).����)�����p�g���Y4���W��I����zA����7C�V@X(�\[�$c�p&��#��;^݄��0�KΓբ�DgfX���=
~#Ʋ��e�"���Q��6��a��iɯ�^��s��_H�j6~j�z�_�C(�Ϻ�E��(�
e�j,Wy�O�}ӄ����a����>[vq�
ȭ?�'d�����p3sˊ���Ò�o���V���Aqp��r��j�����������X����O�n����E ���"��@� �f�C�opI*UZk�Ǒ��f����2���s�����}��>s;�����`uy7���u=�h���4�P��m�P�Z�y���pg?m�-��C����z���f�Z8�p����k8�V:��MbL�c�d�x85$��;���W${Uc�ܳh!nVD%p�r�Jd4	K�!@O�����7�r3%��'�m?��Z0b�L�
�0vb.��za3���xX�6M�(�Sm�g\��ha��A�)��E�5��_�1�=HݢRF(_�4�'�/;��C�cE9,lP� ȫMH�ZK��Y�]�to{�����>OI.�S��~@�w|� ޣ�M����@���s�a��T�/A�BBvT�Ià#�$��5�� �"�����BI�r���o��{P���};
�	� �#6{��<5�ְ��{B��O�����<�?}��iʲ&�r�ԁ]���%�Nu�VڍC�
�vbG��M���"u�NGȆ��W^A�ƽ/����J+̳i;v�#��������K������'x�I?��c�T�qc N^�C��[Ŵ�\���.�d�H�k�a,������Ђ�� �^!��#о�����t��~`��r�֜�j��$�$9Xp���Ѽ�j����;jpz��_��,޸�Ar6�e-�s�* 3x���OW�?��ހB�E��&W����'�`K�Ș=N�{�$�O�8�K���?Q��zܿ��^��ЬD�	�V���m
����(��]���?{��m���P�8�f{8J�S�F��P:F��ʌ�42Z�Q�#Q��m>	�ؐ1��A��q��3c�Õv�r�D����)[?W��>�����p갖%�.��6�i�ZD���2{��Bx�%����F��xTݲȔ�F��lf�4?�(*�l�sȾ���XnV�u5�S�6-0�����Q�>�I���͞O?���<zjq��/JV�}a*ȅ��H^X�Z�N�W���`�O�Hm�G3���
���mZF6��n�2��({�2c��Y>��n�L��K`���Y>-��I���������jX�6�� u��!����h
��tB�g�����͟h#7�Π������3QQ%�Ʋ����(���O8 ��	>
�q��Oخ(����������R�?<i�r��^T-��]�����O����=�@�e��a�.��|D�z�HmZ�Sp�^�څi�d?Ir�衣��S�*.�(@�?�-��t�nHKx�q���}�i����c9�6Um[�*�j2�J�v��MT�	�+'$6a�L�2O��)݉��4p���PG���и���dMR��F�6���K��Y|���S��v���܄y�5)Zܭ_��⃥�{������ef�E]�* K�d.*�C[��"��RD� K2y˧��xԞH�u~�
I��������Ɯa�0lUn�ui~AR��&�Eql��k(#a�5�=�'O�=��ʠ/_����S�L�$�S[/!�Q�;�R�l��w�'�	%˓:z��ՅM�P�<�������Ǖ�9e@�d��dZC� �_:�~��S#"�bӝ�3|�@�N��u��:f��Sq>��1��rjDQ�}��
��f{B����&{2�E!h=ú�:��L&����A�YP�{�>1�O_j+]�fa������;��эⅺ�g�4��\��%"P�ZwIXdU�E�( t}�������^�����K
>��#(�)����l��p��r��1�7 N�[�aoFNH+v�c�z| �LG���]��p?���'W�B�}�~g�������{����O�
��I�.U���^'f�=N���x$J��]b� ���J�7�&�
�Z�H��~�=�:d-��t��u`���K�F�Gn��O��S�~ER5��/���Ǖ,@���zΛ���(>��QKS���
I
��mx�5n��e�$�k<+�G��8D��[�I�x���6\]�چ\�u���S�\��/�G�P�H*�u���fh	M��1��?6¥{��n� �"��
�J�#d/�u��&P} Z82�wx���()��!��l\�/N�}�Z��D�'�jo�7���|�j2ӦQ���+F��g���{����uW����	�L݌���j}?�[S��3�ev�g0.��uI� �$�Nrx*��byq�+�'l\�v�T��Z
��@���ˮ�?�u��m5��c��ys��$,
P���_쾼���/E�H�����	�Ԣ��<OՔq�Gb@�Ȩ@v�V��p���̦I���R �/xC�6�o�J*�%���Y��!� ����P��NB?~	\#��U�	ӗ��e:��:8鲏�~Qĕ�K�c<N�8��K?�/D�����U)�ッ�h��A��m����pJK�[u{�kh*������f�����}��fO?�X���@H��n�v�m4�<�΅Ӽ1�!�0�F}��H���S���6�����K�}c���7ٌ�����Rϱ^x͢�*F�Y���<��LEDB����n�>�'} B�^�/|N��o�6͠=`�M��L�������Y�D���j=y���	��Iy�MG�)��Cω�=��5[�J��gqw*�̬�΍7�6q9S>DA��1��8����A^mҶ(��"j�TE��2N�O�y�El���������3��xpް��(�̐�Y��_��[g;	G<��a�tg~�h��D0�>.�����3����؄
%0�c���q'���%���Z��*uL�=ޕ���W-j��h�,� [m^�E��3T�m�C]vFP|������&�d
��	B�o��]�3ٺ୉�^�T��w��$�iA�}�4���hR`�?9��#�w%3 ��<���s@�LA���A�Rzn�ɫ;󦱌�ܚd��m�3��oD)� џ
��;>�/R���w��,�D�Q�*Q�ĉp��ax�I���q�6�Wؐ5%3���͢�2jt��������k�9Ҭ4N^O�=���m�x�p���`!ۅ�~�('d�Ë�KA���^�)4����p���#%3ql$v4	#��z�](���� ���q�|��8���s��v��٥�׾\� S��,e�Q��uq��D��cR-�v���O�A��U��U�*�J���W{kcA�u�W&ZD&G~;����`�u�m����������:�Մ q�jbbz��$����$ʿE)W��D���	�����yMc�����