��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��<��T�@d�Gu�!�h�����j~���C��P�Rc���FfxXs�� PC��԰�O����p32iXA�t�"�Q��&?,P#̓�*eA�9T�x��0�8nVHAG8A��J	��c���G܂y��S7AC����&� �?�,�	�B�Ũ��aU�P�̧Θ꾸^�����\�(+��F�I�j�z	�Ϩ��y�g�8!�2���%Q���_�m�$�x���b3,B�6����9�@fZ{�G?֔H���R ���o�;��Hd�����������O��3�m.��]k<�B��I_"Z�L2��:*p:߶����aȈuJ�L�_&�݋�w�����j3�����:6���Ɋ=�����e������0|)
m�N�|[d�)��H���ڵE��Jq�)Tꗓ&�^`kC��O bC������h�j<��+�E�v�)��G�i�SN�p��x��Ǔ,�z1��@��t�ܕ돹S��Iເ��8�^x�)�=��V�fE�s��a�3c�e �ɢ5xE�'�fr&��W`��r�E�m�_R�W�(�|1��hR�%�O��p�ʼvkn��I���T;6�<���d�Gt����d��qkcR��H�5=�E�zD�YX�k���B��&+8�w�}��3V��Cbk�9G��3�����h���7�#���J���j���d�]�O�x�kk�J�1�A_��,�&�:�C����+S+�p�R�^4fN���U81�{^��_!�R�q�Da\��p��{��Ox�o��,ȕ����
J��wܡ�V �p~�P�l�}8���KP��שX���B֬ȼ���_�R_�?Pٷ�x��4TZU
�4E[vS���J(R�v��3��C
0^��B7��Vc�������Ca�A�΀V�h&���.����ڶ�HD��!u�R��v��=2���r�]F��|�]�d��5�J�mX�5��/�!*�c����'R�h��lyb���ϔO��������*�s��]b	Aq�)�-�v�r�w�N�gU�l�?$&,�����_�>	��BG�X�o��� ֜'8M�f� ktp�D�ޣ�R'�H����,E*GPǓ�I�Q�o8���dk��"��+��i��>�Ƌ9�P9�K"P��l��e�2u���.� {����e+{����uy�낯�[���i`N14�k���`���z� sQ���ʑ�b��cr�p#r���=͝��A���S�OM���`�z�v�����%5��wa��a� dLu�)��&�i��<�+���=HjJ��?i�ׄQ�n��>AE�Y4�}��>F�, �Tk�J)��8�y3�Rso��`�O��э�u�Ț�� O�ϒ��hx	V5w{���mп`�0s���("37�ۚ�a�֫��qΙv3�}����G��~j���Wv��6%pP�����������FN,� ���G���G�[�q\�yY	��O��j5T���MD�9����g�AV� �ȓц��k���������c��b�*�U]_���٥�3�k�7z�m�w9�CAC��nt�p�����$��b�4�V��P��׉��3�OU�A���~�ur�U� 38�Z��}�ÔN�"�Ї�����$�),�,��}\)�"��;��u.���$��FI4��(0w`M����⪞�V>���䶼���צ�tfg#6]6��@��9zyz�4�@�T�x��IZ�����D�W��Y��3��n,)�/�i�R��gd���׀|9�"@�\�h���-��f�h�.<�KU��M�Vx���l�_���ͦ|7�j�ݽ&�:F'�����<�"0����d���^[n�2�s��_Z{	f�j�f-.�bn�"S��eJ(ѧ���sV��wMc
Ӭ$�� ���j3+�Ĝ�A�����^l̃�[�N,wa�	S�Y��N}UfO����	���4egsא=
��Nh�c^�=�5'�X"��r��pux���(��{��C�ĕ�s�{�o�gWi.FyR���Z�8|0��#��s�\�1�I��ȩ�����G�q�'Z�c��|�~F�X�U�Y�B϶2��� ���V)D2�b�B�Y
>�đ40�h��c¡�r�z��{��Nn;�H1�����t�ִ�|�M��!�FT߻6N���#cܪ��H2��
�2g�@�_�e~4�9"N�Z�l��9� ��3��"��~�!kG��MZ̓�L�޳��쎴�||E��C.�nL�$(#LҘs�(�9=�S+\L{�Dt!�}��P�K,Ȏ�1�´}ӯ���k�:��׳�%7-�X��۶�w�^�ȼ�a��V��u񌟭���4�H��8�L�v ~��9:,?��N{�c�H�T7���;2�d{�|�|��s��$y(�Oke��.����aY���s�ɬ칟����^�i��L�l�;��Ej����5pI�q%C�,d���h���(��i0e�:�́��d �C>�&U8�E�c`ޓ/�ԝ�';5�[e;�!1Z8��l���Ch��(��9<��,���[��o(��r�A��Ɖv&�>�~YIK���3>80��R�Qy� d5�7�+��2(*t�ؗ������q�%�e�\E�����}��t|F��Q���VL��T%[b�L�I���d'_�I�kęգj)��Q`��qP����l�VP�}߈GQ�)���q�L��Y$����7����ܾ4�g'�)� pa&f�;�{���4ɖ??D]'�ly4hz�h���,o3;��f8���� )��r-�*���:Y�7�?X�!��p��&��6���<��¦�ꠥ�����D1~r�ݢS�r��Cۄ�FNp��jzC$�԰�[�m�;�J����[��U*�; 1Y�B�h�lX��P)�9�\���:�Rʧ��o�������ڹ4!�s�_mI~��D�ޮa}�	�d�m@aJE+P��f��hBB�y���4�;���ecq=��%X`d�R�gC�D^"����䔲����/�u�{)���	,�}�&�S�@�5	G(�ے~�VF@�����.(��/�ޙj�h��{x�����4�73CuhVV���ѕ�]J�m�qŀE��9N�`��+E���1�p��S�4��!'��s���U�7��
��6#u�盇5�Ȭ4_5����cH\�HP*��R_-��q2��O����@���ā�X��g[���1�ż��:�A��e�EE �����nB�}_�����C}���N��e��X���r��a�x&
�d �����斎����쭎�v�ۼ��Î~�E8�� Э�_Q��(��m��u���/a\�� 5cS�������jZ�1}�R�-n�>���c�_���Mo�������Z	��[��l����]լuIEK�tc[�F��	ݷ��v^�]��W��u	N��`t<\"8�È$A�ZRX= B�;�Gl�$��v�w� <{�{i���R:�3u�﹩�K�)ႛ�.����Y�W�C�����"�/���7_��^��c�� ($r��L,��	�SOH�%� ���E��ݺ������_�_�h�u�8R��5:;t���[s#F$ف�K)0�hdf��%��5�9�lɒ�V`hy_�j�8S&m_��0��O�m�e��@��_J�@��2�DX���J�?O�A� vY[�B$�˓�[u"�.�w>gԿ^,ls���im\7T����L5ض�O t��k�̱�Qg�p��?�wG����u���Z]�E�����z�����\^}@l�2<��1XTz����`D�A/��\P�ABDvzk��rF�<�7�I7��AZ`m2� :ݪ�pD�*�f��w�+�-w����_}���5�1��-h��@�/HV����+
���j-/�qR���F��٧�l�k�
���o��/	Q�ї��dA�U;P=w-�D��#���	�)3��!���X3��h_�D�� �r�(eƒ&A�o�����=�K�	$�~���@x��/��d1y��
����Ft毰S�tӬqs9�3"�ϧn�_hо?(A��Z����W���qt�����'5��A�L���)!v�L/m��:���}+ݍƍի{	C�i�}~��
����k=�[c4��9�͞uk��lF�l��,�6�tI ��|�n�':�V��e�F������1}��������o�� m�I� �q!�Rܭe�m����k�F�@�^RhĶ�|=�CY�94���ډMΰ��~�ۅO��Xt�>=��;���	3F���-OM��Ӧa@���,�rǠ�X�]�[Q��!� `�)��.�|������V���CN=	�t�&��p�Mpg8U��D��3#�1@�ps���#����bG ��X�(����2}����r\��t�b�p�]0��!�:%3�}��+:Xm���Z���c��6�c�@����Ŗ���0
����M{2M��uM?�"�:�"\V��Ru��*�ECO�?�)p���oO�H3����}��\�c������U�'�<�ݿ ����R���qT�-*��]dZ8�8?A���0M@'�~�02����S��6�JZ=5�=�@����Z?�����+.�Ƨ�NW��ݞh�\/3
j*@�/��Ɖ7S��K1(=��[۽���Lz�Ŕ!tn��������ahu����騛f�r�HY'&�A�:��e�8n�e��Z���=A�u��B��x�	썫P�R�}�̅LKՏ�������j���tJ����d� t�.��A����gTT%�>��#z2�/���f�����r	��l�f������0n�u���L"�)	.��x� �(,����:N�X2�3{��H*+Ϸ<����1@+Pet��?�R���,kmJ�e�y�P;�O{�1;{#/����q@3��aD(I`��),�DP�}�<W�h��v��o3A���Ѐ!�0B�IEJY�4&^ׇ����*�ȤYo8#m���J�P��I��"����Hc�{�q��;e��[E��؝ը���7-�s1$��h�<�s�� AOI?E�H��H��)m6F�㨳d,d�%!��C�)�\1<��2���oT�2����Ժ�17��f���&���9�pc��y	���if��C�ѥ߉�>��+*=!��'�UC�è.)`E1/�m�x:�jZ��q���Å��x��S��1a&�fݜZ��N���7�����+��?QS_M��ap]sև!R[����P�j7hej���1&��*��ǘ��.���w��R�`fd
z3^�V��+B�����6��P��M��Z��h�;Grn�C�t�Y[$���mS�q�88����<��/y������o256`]
1���م�c�)�1-uO�q.�pڱs�}c�G��#�xW͡w;Կ�"jG_36QO(-k�u�X!�ǯ��#�ǚk+�\�A�}�%3�אhW���|�/
��^T���}#p�
6��E�%l�R�Pv��H��4"��c��;a��Y����u?��SM���>�a�5��\��1�\g�+'����l[y�Tn~��B�<���� b@�{�c��.��L��F��h�� ��*��ޫ�:�.Yz|�x��2�v�
0�h
BN��^��!��a]��&����ݜ��u  ~����i���7�H9��Ua�|dd���K7���j TP��!�ɚ���ʌ�#,�V����rm,Ε]��K�q<�r��q�����a�$&�AE�/L�8q�Q(x��-��W\*ᬐ�|�Ȟ�Ǭ��}��j�H�W��(Yf��~�M�
{��s OGkKQ#��u����g�[�A۶����Jw�w��4�w=s�q���D��@ӕ�����3�v4-+�XC!�N��e��T��$KX<4�;&�$���d�ǔ7��e�o_��t���P!Be��C��G�>_<T=��%��R8�=z2T�ȁ0�L"� 7��0V|�n�28�'=w�^�K}�4�;c������2YH���<�V#�h��,y�9�d����u�|�J��=���K��1$�;����@B
�6���� ���s>סAкػ3}3�fw���6�$�}u�ۡ2̐�V���Q�� U?瀧U4�[� ?7?���1�ƑP'�w��gw���b�v���0	�~˼3���h���fc̈g���°���#d������ye\jq:CJ�Ǎ}��3Ux�G9w�H5t_�|��|TP�ɍ�y0�1�;�A������� s������W���Zg�g�(��pU�R��s�������KE1։3m+��b�*��&�g�G�a�N�w]�P���|�m˪���[�@�mN���1�����+_�+ƽ$�W �mW�{�&�#� &7V��́zK�����D����s�����bN�U��$(q�Q�1XF����v5����k��	�ʘ�������Z�&��Q\����-��֞e�S���W?/S��ʒM�.V;n��r�N�[ qq%>�+�!�|E����CU˃�W+�1��	2m�M-��t�H��֖���3�-�,�O�l���P�Äy�j��J�ṇС	0�Ü�R��+�$�X��Qɧ�c8�]Ψ5�d���b��4gr��g	^�;�=���5j�%���U\�k�N˖�P��I�H����@�2a��U���:�I]���$�J�wB�P�W���p@����}"l�U7� y~�g�\̤�P���#0ق	<����+3��>4��T	)��5.��L��K�X�,��*�'n
�3������@w'�)�N��U���j]��&�nM#2�F�͢��4t�Im�'�W5=́����9��%�[�����|�E���s�h>�#8�J��f��"1k�yw/'�`V�xyZ�#Z&����#�7����9�Y�`��dy!F˱���c��Ub��^�a��a���֠�s�O�َ;�"��@ $r�;h������/P�S���WYl�O8�y��d��L�x�R�ǊPyH�m-o�r������\2]^���ݳ,.i��V�o;��*N�.���w����Ra1o,���:�5�e�}�1J�?����a��ѵ��G�N��^;sh���AOO �L�;A@G���з'����Yf�L�#���O�[�͔7�VG#���n4����rpib���k��Ӗ_2�樏��WoS�Ĭ6vN~a��<;Z����*�4��L�dӮP(�n�(v-V{|��W��旪/�UdX�Q�5�:\���0�p�k�e����nߧ�kon�,�e�Ǚbl�:��5�FA(RB�����7����2� �ʘ�?$X"E�R+r��e�V� �b�t/����M�|�j-* tF��//�/l,��BA�i�B�_ò����O������@��QS�w���{:��7�NSd�t�@>UJ�}��O]��.���x�cY�|�XO�s�����f<n�P��<_�
p
<��� ������#S?�pf�?�!C�"X��@sT>\���iXD��M*�p!i��V>-����H`{��R>�J���,[=غk�I�3nP'zo-��!�Q�x~��t{� Mo9-��Z>�NHi�8�J� ��a�s,��s�Oȵ_晎�����i��Hm)��,UHs����t��;"�UY�Q�!RPt{�ǝs�h�"�9�h���ܙ��hdC�z�Fv*�
��8ײ���?���zY�;1����v�h�ڕ�𿶔%h�ɘF���J��^�}�?�2��$`�K�
��D�e��xW^�GY�mJ|�S�~����n1i��FBD1겻D���G��r�0}X�#�Wg:t�y%�J/+�����]Y_o7�+_m`oҋ�y�M�L�l�Q���M�DC��yuO�<%ofR�&q�I���� �-y�mC��f�O���F�&����d���p\EX�'lhe�T��#���3�e�4D�k��(GL8�ۨ�2/�3��v�HX�R��|�e�J?�VAK-�~:�c�f��_����̉qe��	���5x�κ/\4���K�SJ>}�����Z�EY��{�7@D��M���/%������T���a'ȡa�f��P'��o.Y��sD
:k+�'$R�!�+;%s6���/頨��e�?��j۽�.��2��+2a�O��3�w):u���rk���:do&�f_��U�ϒ��ଢ[]|_H��Zx֭v�מb'*�p,���K.N`p�=G�VRw��bH�F
�ߪZN+HqBJ�7�H�Jm�7a� FH� lJ>�J��]c�$��*��^���c�q��-�YC���<���Gʜ�����@S@�gۆ�
#];������ڧI@�m����b�$�1�áZ�Q���h~���Ԁ6O�8�h@7X�T�ɭ3l��?	 �
e��(����{Ķ�� �tC*�~����;�,l�J��[Xg����]Gq��Ԧn���DZP$tfzO�-���q������;5k՞�H��n2�	�p�	. ��3(&#v0���΋q��fa�wc[�����3eݝ������:��Fi�^�_z��WyF3���,��ެ.	TO�5��\Ü~s�����=���E:�b�:S
�k��˛��z"烖3�"R���Ch�(KI=S/����"q��Yt�Z���hm��u���o�"�(li�W'7-�Ԓ�htJ��"E�M�4If���`䭡�@�T���Q�N���3��h���0��������"ݻ�����r���#6��L�53v�v�#n 0�����X	����z"^�o���n��}0�W<*#؇[e���>�u���]�MM)�j\�X~�`~�w��g�I���f�p�#�ey��ww_
ɭp�7쵴�Ң� ���q�qW�/H���K����N?�*b� �^dsu���u���NQ�L����q��m��5�A"L��u�A;���� ��dl�@X�L�P��8�8�Z"]6�!.T�I��x32��>Q�q/aĠ�7���V����RذM$^���k(��L�&Q�x�����	��}�fܢ�^^�4[�_
��/@�#��W�$C_��L;�9�� "��k$���2;��~��=#��mOƆ�����w�G����fU:'�YG�"��
"�5"�2���J��\�pA�Z���3�t8�Jm@T��e�E-q����I7Ϥ�L����.���l;��LG9�Μ;U�&��2��s}�gjc��^��}�nן�J�-�5�@E�*���Ui��VRi��R��K��	[���7��}�J(*8KcF�v=�M��\C�0��5	�s���q��?2e�����'���sl'��t�>8����=:Y����92[h{�qVu��
����
&��a�4�UT%��7-�5���*����Ŧ�E���=����_d�O��������<�<�~e(� P��[�7��Ys9�&dct��ߊWqː���_�p��Q��?Z�*r���������;��輠�ܭ�q�lO؞-�	���]<���=ߞ�\�P�VuGWoG����&�N������q�%]���ˌ� R�կ� �W6�rWڮ�B�LNX�Q��h��W�o��!ȧ��G��ZKZ߇`6���񮘠0��%sI��V��kq��{>���Y�qp�%]����L��r�(��3 ��� ,�{��j�٣����{�$Z����� �@-�F(�|s6Wq�X��{n3P�h�{�����}��cѥ ��`���l|�O���[J[<�Nᢶ=������C}mװ2 G������m�ѝ9 I�}`	���3M0��/��zZy�x�zIz}����&���m�t$f�03\�?��q"g���GWo�-���_���|�e�SC1����D)�$�-[K��L�{��*�.XH�W��Q�񳾼U5�Ӿ$�����$e]����1+�.+�%�)�=ن��������أ1�&JD���_>`��s�`��1��F͜�1�t�����f��C���Zr��~[���>Ob^�>���S
��W�i�]���l4��K��m��px��-�E���CX�� r�����Z��]��3'P�pɶ�h���a���N�w��"��9�]�<o������h5���XdZv��Ȃ�0��)���|5�F,u�e�����D�R�c���w�'%»�;�ח����Qtn��]i6䨑����9=��W;V#��"�ܖ�T=�wm�Vѧ�Q�2�5D�����%��^u�\�����B?�(	�eڥ�B�2ؼ���/�Tr^wǴ���C��wip$Ջ|�� �2�^��L��mv���sҖ���+���w:X@�7!�]!��b�e�C�=���@����EL�<$N��;����NX�-��cA��f���J��µq��������]�Q'��A׃��9��2�r�A�'��-�(+l�h���C۩
���d��r�9�^��v����Rfܲ|�������P�~�S\~qhA�u��o8�?%�x.�'�]�M�2��Y >�\ͼ\��Ƹ�� J�8!h�'����lUb���ޖ��US�/q&=��d@K�*lLZECWd8y��$�B����2�����v�\��8�OYŵ�r�d�L�P=޻?��k����)���/%f��\�=��?̝�Q�mP�# f`�dQ�+�N��ă�VNr�����z6X[0)wM������(������b��|a�� �zSmqA��t��w��q�愱g�󎾲wgeYF�U�f�F���Pw�9j�?;��i�~�0R٭�hX5	�Rk���I=�B�}#�U�q�Cg�Q�A ���T����kw��Qv]�b4]AX`W[�����Z�S��dG�-������FvtRu-0�sw�D��H�(\��$
��R�P�y����ND�������q�>�B��H�[��:I�f_M~��e��Qx��q�H{�a˿�$��|��L��3b���],��`O�)�;�<Z��� �NP #1�˶+EW���UYG����h%���W��+K����߯�S�jy�׿�'��^L8	g���*��
�p2  ����,r����~����G�GǮ���T�!�o\s4b�����|�D�*�ā�] ���i�nm`�E����(�3�M-����c,�#R�̳jPR���G��	�ξ;֦���͆oLu<Z�<5x���!fH��" a���R�����V�s4���34�$�gTG�Q�*��f�fr�A�<��H�v_�������w���L*v�-,���
(H���Hj0���fo#Y�`Z*fY��4���6�x��l�z��<c_.�V=v�m�a{+~�d�M�!�8w����I�<y�H�F�(ydV���{�y"1�}��}���t�5�Q��N@�7"BIi�>�!H�11���n�@"����$��m��=�%ٔ�g�C��t 
Y\m�%r�pJ�(;�+'O����MU�i�H���_)	/!��L,�*�	�K�du��Wоv�V��{��-�5�q!NϟW1?(Ńq,����>	���N��9���q��%p���������W��	�U� 3P�yJY��n�#�C�S�Ec����f���{���(m�I�}]�������^7e],�P�q������j�kP�W &Aa;�z�s��Uy�_�g����H赀�%�l)�� >CRr;A(��D��Qf��Z/���}l��ӏ���X����z<k8<��c3I�I)��2�!��9������W����&�;t��+2������x˂�2B��6锼FKF����h�!����R�)�����π���P�@X��'$h��ԢGg8��ּ͆n(_yN�8��4��P���?�C�L��l�z�*�}D�_M��1�\�Ś}�U2b�K�Cx����r�eڮ������Z�h�F�֊oR}�)�9�.�#	(s͠P�M��R>~���yC6�@�?�X��@�$������V�eV쾖�q��^�B=
����*��3�<�6=T�|�g�s��G[>��kl�>rH���a��r���h�r�ܢ'�¼�_I���#�V�8+.���~}ɾ���'z�`�6�a�c� w�pC���^۷���ee#i.���[}#Y�&l�T�k1\φ�Jg�����,�!�U��ht.�[ߕn$9��A��%�V���[z�/[�4��	ǅ3�L���3��xJR�\�u�
�'����},w�WCd>��!��|}���5�J@���B5d
=�́���SV��us��R �$)��4���N����2�v�Ť�,�S���d��z��3���%$�FE�9�]�`��,����˿�Ч!�%��ޜ8v�P�F<�NH��h�[|{���y��QH�IH�i/����.���K�Y�k��%�3��/�����K�f��ǅF�Ql��@셰/1E��@�4�;�H��(x�
��h��x$2�#���(�4$}T+q�х ;Rh6}��˿�l�ث�PP��`�gS��@�:����# ���حV��.������,>i�qq�(|kP^\SF2�nzJ��(�
M���&�2	�(Y���ZwT��J�3�o�`�#5�ǂ�/\V�<T1ΌM �����QX���_���i�~9@��!�ȩ�'6�����M�������"����[��Zֈ=l*������C�aJg�(G��4i���<?�΃t��E/{;e����~VF��[Ç\b���,����3�5�ث���|��9#�W�(���V3�M�����13�&���흻���M�����Mo�E�i���Pe�"'ࠄ"�`h�^�ɂrX[�d8W��dl���D�KD�E��An)\z� G]6�|N�B��il�W�a�@Q'�Te�8�ɪ���K��Z� �	����Y	黊��9-����x�;�Gs�?��eTR��g��}�������F�֎L��-�x]�����r�ZȀ�$K<@�V~�$����m�!"�S���I���)������Ĝ8�#�k���s��iI'��oH�69~]���B��!]D�@�H��Ok��[
zx�Yi�j� ��� �C�����(���-	|`��׵%V�����VJp8��SJ��`@�HݴkL�4Q�e�F/�$E>T��{q�u��xɐ�����î���c+Sw�2���%7]6N"
�I-ɀ��^��,YM�z�1�ΐs^Աu��hڇ�/�I���spY��O���HS2V���$y�?�'���>x�SN&��ցդ�q�l����;k��<e��%����xR�ƃ_�F3�l%�3v���Dn�Ѥޏ�D��A��`q�}#��4�]h�?��P��A�z��0��y���U^.����܀,ЎR� �&�<s���A�!��?�t���a�ݲ N%I���#̾y���l�,�vg��\�]�g��j�A�c(2塞� �ػ�#�F�����
��NZW�i���@��56KY%BNLSA�9�t{��g��w��Y�d��x���H�R�eÝ�������S�:JbQ`�?��W|	[���bd�b!JZ�\ƻH//�u������>4���9u�D�/�U��*���2B_�����\O�XV���;�shP/Հ$*�ɸ�O��i�VR���w�t��!�<2�ՊN���[r�i^I�����-kc�i ���"�u+m��<?!E�x*f2�ee�Z���4 ���SP�'���Dklap�/0�~M9��Y���8_��E�1m���ۏE���\�G�uw]/�&6<�G@��B.t�9�KTsm����y�<F�'1Q������'�:'���+@���IO�a�T��-�;vxt1���.ya��/�� �r�1�4�U�����ٙ&B7�۷J�9�NE�ɂ����5$ь��"z�sD��p��#s����י�OdA�~��G�q��/e(�ǹ�MC3(eₖ�$	h?"�I��7�NP��dC���	I�[�?(�]6�]g���~Z:t��,�ɳ��>�D�W� ՘}�4\�h�9WinQ�&z������E�"r<��K��$[Âv$Mn�x&%843�l�*�� �w�姏Q�׎,P�Ys���f"����?��{C��H���;)i���+P�/����Dk�^Q�L:ީ�⿟b�a���b���xі��'�BU/��L�R�i�;(�R0�Bp�w/�ajO�<���-�_��E�)��!��4da�3X4�q!��i�
�T-�<�|:�j�j�|a�aY�dW�n7��gF.�g��K��05%��AG���X�ܜ�c��o�]�ҦzW��|2_�Na��S��������^K�/����E�3Jn���Ólu�$U�K�����^ҭ7P�ӑV��>�N�V�]����_P����\%�����h�����k���t,��c��e<��%�/E�ﲡdx�Lu� H��B��	����q<iD�l��+�RbB)=�@C$����#�I�V	����x3�G�>�M=��Q�R�?~��m<KM�-���!�	���"{�j�������@��9�Y�U�we��t�Y�muR��e�ܝd���1MW��L!w�>I��'w�6k��p�Xn#��&J�o:��5��K��M��\ʸ�p2�(Q�Z�X�� u$QƈAwi{Q!�H��0�o�E[�x{y,���ɯ7%LV�%��l�FOx�I�wn��F���m<�qB�gQ������� yw�m�0*��G⓫�Ь��M��x�1��)��;�Hm6ǯ�&^�`�!&^��)@A)Fj���>��BV��p膤#k�橡f���B��?5�|�H�
�4A���i�q(��uf�O��1�cC��X� �qe[V	��*�Ύ��:�W�L`/��w"�شo*�A�
`ڒZ���1@�3������ѩ�;�qVG8�Tcދ�B%r�6'4��0�e���� �D�]�T��G��K���4l�+p 5o_�V��sHΑ����ΈE��C�ww!��n�e��cQV���Yn���{
����Eƚ* �1��*9�mj1hJ9�k�}�(�#:@�����>J圼��L=�h���w�51:�]8i©��yg�'R�QZ<9�X0�H�|Q-��7V�1������э�{}�ZPU���~G[4���R�f�E5k7q��؍&�G�k�~����7�.��r����sW�O�3G�r��qGϜ�ኜ�@�'�Vʾu�![�1�L�{���VF��ɲ��8��Z��5-ߣ���=��'Mͦ�Ë��w�Oc^|E�.�ʵ��s>7��#b4c)[ۡcS,#lt�bAr�V�|bR~��f!���U=�t�<J�l���]�y��*$ƴ5)p�k�&+���C�B��_"��6udA&��e���,�ȋ��Uݯ�$�{]��x���fj!�y1g����U��G7��uQR����i�� qR~��ٴ)¬��Sw��["J.wz��暞Sy�i8U�I,b���:�t�}��s�u{�i����
��.J�	�h.8�����������\X
�
 ������m:����o�H8�	A�%��Z	h�^[D�L"��Z	ItN�����%���8�Ai�& Jl��M@E����t�ČȾ4��3Q��	�F�|I��]����}����A����j�����=�������jE:Y;����I�3�x�i=�j�����9hBe���9�����2�L3��\�+�.I�c�&bEt��y��WNf����r�'�Jg�k�����VXpn��g��*����a�4��%����"�<p���x1�+�Z�݄�#?��c%�/���i,54����E�VsiFҭ�@�t�v9&Ş2��,�-?�Gn�e�s�c��U����`k���P��Nq~���6;����BH6P�~�s�(d�<vF��p�H�R�����42�� ��C6&Vh�*;�$ ���M���l)+�1x*Z&і%;�ti��cD��5M�����/�����]DZ���t^)$�h��y}ºw{�i8��d��+��Z��[����AKtD�LK`S6�O�X�`hC���Q0�R���%�PSh������̧'S������.k�MP�ջ�� ��ً7!�G��W}�A��9��N�{(zWc *��� ���0��F�>nD��yfEs���G�4U���g%,��ؕb�S%.��j�_�����_�x3�w�˒LL��O�L��S�y#}AII��{���~��Ͼɕ<�Z����m��B5CY��3��{
��rM�O�֮H���vp[��m���#����dה�vǽ@��a�P��pA	��8�x���7n�v.`�)6�);���z��Lxf����qY0���jS���l;PV�������#0�`�,n9�<������$�]�Э�3�g��9�V��`�$���;4��������ɹ6�R�1��cf�bs�����U���xZ�ɱ˜ p�K����fJ,2q?�*�=`.�K�ww�� ��S��{V��v��>��B�
�B���Uvԋ�Q�l�t��M�n�%�"�^����w�.<3�p���e�!��/} ��K�5P�u�b|Q�g˽����&��h>)�2oc�/$�vr���M#��þ��o�VS���d�x�a��Pi�[2Q�9������L�/����o��n^�(���	��k�V؋6߃KĢ�fJ�oٝbn��d�S��"�S�̨w�	8ݖd�Ki��W��~Lhn��
�
��/��R7���������~��X�a�Ϣ��ƴnhUȻ�|�T��1�{dlU��O��#�"�9f@�À��"6�M�4¶|��Y�2���ъ��Dq@K�9r\�
X�.���;���r�_r3� )^�Q���F��<Z�����R-�ȟn[Q�r�*����*�	E�[oVd,���_�~:�q>i
���N*lN�Z2�l
tv�C_�����'�1Z�KW����7��B���
���{u炀W�@�������a�����_���[�~�q�َ���P����2��ߙ(�_��������',69��Wj z��3��9{�Ϲd�f��=��C_���>t��0�{�4}}+��;�����|$ �L@�{:�A!�
�������>���0x��^����t{�M���k�@�
���g��5�~Q
��)�������;EQ��
���_��H�x�r-CZiWl�[��������K("C��}ՠfC����2�Wc�xi(��,�=���p ݛc^a3�Os�����AxL�	֠Gzs�'�a�)��$����Oc�e?^����`]�*�x�@��S�of� #XYn�+n���z�����]	��T�ŏ6��(%:�̼a���e�<��,��^��)g=0��(��qv�*pX��ZN���I>�F��RJg:l��kY��=�y�|����ԕf��9�!n�[e�'�RQ"~�0���a�
���dH���R��Cqi4ViC )>HfrD���(V��>hX9�N�Er�Kre�r�!"��	WD4��V���]�KR����S�6}*tN��;�%�������'0��O8~4Z�� :?4�~���� 4%�s�K��X�F��ݣA���yZ0���-)f��~UsZ3�ߓk�Gn2k=��ˆI�Έ�=�Z��h�o�S���/��36� [Q
P� .W'l����$�W�q�v���]�e���ܘ�&!��H�-��8Λ=��w���k���UYڲ���N-kMo5h��LjJ�.��Z_��~�ߛ���N@�إ�i�TW��Svb�]I����r|I�ۢ�)�u*���i`������<���B~�Ǿ��kJ&��*���(��*"��� s�HA�2)q����QN!�p��F���P,�xzx�����)�,�O[�	{�l�R�6�흯���4���I���1.w3��2����f$M�B���*ۙJ�ﴋ�q�.C|������#�7gb�B�L��:Hn}�Li��g{����<XH~�[�����E��U��ݮya�+��Fbu �.M�g /Wp�/��79 )�e�RG�>'R�*��}���99\��t!x�F��!�}��������ͪ�n���L�8�
�OO��q�k3�Gh�2[�������˨�D��bWi���hD�T$�OE�!�������G�md�&���>[�����guo⯃@.�>a��Z��b��w�~�C�o���bo�����?T3��q1av��1�X�v|9� ��#Z�����\��KrW�Ճ�6�����ƫ�Z��O�{q.�>��*u��� W�g����Wh�'2E�����f�;9 �#'�{7p{�g�PEt�k���H��9,�PF>��Q��J\!�M�TAD�Λ/+n��y]�^�-���$�IR�`�����!�O|
�E�qc����N!E���>�1 ���J�ܶ�O���ӽ�P�[6㭢�F�� 8��c#k��B̃�R�
���0&���P������n�FvkS>��r�P���n߉�!�A �7��ܫsG��Wn�Җ��*˥�����߱����%��.�->5M����`�Ș�Ls��gU6�C֟��kϓܪhٸ�U�lDʗׄ���_�T���=�jh�_9�hxw�oc&�4���"�_#�&\��E~���W�v#���g�v8
���o-�2az�e�j�˜I���S7Q�4*�-��[W��'+H,� �-i�_U9�����uA�!��E)�;�`.r$�X�=N/�r6�Ry\����g���:���87.��v��,�6&%܉��$�˿�V���.�;ջ�-m�ŗ���v��Z�`ML�c<���?��3���X�bLd"-d���1]M{g/��'�Q�C+��<n�"�@����ܷ���7YϿ�`���Թ{�X֯��ioZ������[q$pÑ
�$ �f���g�3SP��g�Ι �m��wkl^�U�
K%;�D�\�]�-F�n�jf�mz~�-�4����󍝧�ו$"��sn��z��	��a�x�������������oQ���߹��v[����Mk���J�5����������ӻ�(g�&���ĥ��Vn�� �
@@���OO�J�Y��һ`Ú:�<.f$�#U�D��y"٥����,�؅*+�:+CҐ�>�}�/^�S`
����o�S܁2�%3�' �+8�
	$ݟG�-핦i�
�rH���Bo7��r�f�@�L�ݪ�����]r��w�\��B��# ���P)�5���j*Ww K�Z�mi�,f���0N�U^���̓�b���I<a�ˋ�=��f }�⊖�0�}��8��.��{����+���`�"�~���s߾�����s����A_|�r&v�J���m�}�2��!m�D��&����Af���wpNi�(����t�Ϩ���r�bC9ɓ+�D�X~����l��ieX8�Z֣�xs�V�"��G��/�E�c�dR�V
t�����Zk8�S�Y`+@���(�x�ܐb�Lo.�w�E�*�"sv`�;N��d`6��ԃ`�<k��B����Ja:����(�e�K�_IC�e_@��vA��_!����n��d��Mu ��!A8��]�w��I
�Rי]�pi�=q�X=LG�+��VM!#ns������Y-*C(���M'����