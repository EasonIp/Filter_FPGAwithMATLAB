��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ḱ	I*�ox��͝"zܕ�=����T%>�����,<}��r&�:疃�)�1��N��oS�I,�	�P_� ��^����~\��>��[�n,�Uih-5�* P�3����i9t�wK���g0K
��%�ي��n����F<ͿΏhf����B����VO��h�2����Bqe�L����y;g�`�&A��\onǡ��IZ촹�N�����|��������2�����O�O�(�7.X�a�˸So��	���`.��t��(�
x=x�(�r	������0����}�c���g��?�P�&����5<��@���)��c�o�T�J��c��w���MG$�L֯����uS�r3k�Wb��V1T��ڞ�±K�Y�(���'I�3��S�*�E�ص��'tI��L1G��ID����;t��&�[��'�d �e��|/��偪�+7�Ƒ��4K���aO���p�̲�Y��0!��V�!`������dN&�bMV�"�����-��}�ߋ ��ݼZ�w�"���2��8�����![��d�:"�I0��Op��~�� �ή���ě���?X�BF0����:"��af�(�R�0-'��o��	�Q�+����>rC��!�����O��:���K�D�_W�w�$��i�]k�Y(e�G��{��Vk>"�Xc����+�H<SR>ҧ���5�YM�M�	�V{�;OԷI\tנEx"[mkv��p@�!2u�3�i2G;y����q�2Cv3���pWE,Z�;�+���[2)YA�3?����4��d&�؅σ]U���h�s�M��V1*����Q�[���3�ݕ��VS���h�I� ��/-�P���-��<\L�l���T�k�Y���:�T�ϼ�����k�~��L��H9]RTm����Ȏ
����I��Q�uh)�z��Iۭ�x��o��tN�0�����o|R5ؿ��e�#g� �9uh��x��V�QhD'&�0�q��F��V�*�i�uU[��T�<u{OjXZ�S\܄5�)����UT3'����ϼ����%����54V��8������ ħ^[�[[�\M�$T�dӬ�I��QA���pi{ݧ���)�x.���D�:7,� ��?���G�d0�5��%`�j�!��?�犺�R����D5�En��r���ށ����(_�R�~;�#���c��t�)�מ�̝�{�.��D����i�ʋ�z_x�s�H����e�ػS��h@/��ú�����X�(ҏ�ب�׫��^2��2cj�؂n߃&Ly�&ff���=s{��$0����!�n��,���X[�20����<�^���}@����2$l����� s�X���s�;��4�(���̔�H�E}�I瑳�|خs��"��Z�+�C�C��Ρ9~-x�Y���q�JN#�aNe�0�9D�x"6�Ai}�F�S��z��[@J3�j��h��e�t�֐y���z>�����Q�9���8�����j��wh2�Mࡽ����2X@�O�?f^'�=��C���	95��S�x�J[��{P��ۛ��$KHq���L�sS �e��!�k�}�~z&��4\k�
��;�&�������[; X�)��};��\W�a��D�8��B��صN%����_O�n�ڶ�ɯ�:\oFA���	;�{�t5.��!��d���r�qC�x,k3mLi���ƺ���7&��zE����x��f�ww�pY���(��^�B�C%�2r�)Ku?\���=���~��w�l�,r�B�����O��?�'�m���}ɊkC��Ma��f��Ƥ���.�-c\�j<�?��|��t���E}�B7V��Ty0�_h7Uh�T95�˞�3��(w�a`<��y�m�/1�i,?(Z2ֲ�\\�
�h74�)����]�uup0���Mۘ&L�}~]��A��^s7�F�z7��p1V�f#/2̩:ܝ0s����T~�����C�9ρxH�qZ(�)ϐ����`S��N���	v�&zn�}TD8c�����?�����Wܙ�y�\��./���+$�3�s٭1���%�=��J�b6�K���f�RӨ�_�����#�T�d.�B���2��}NsY&��*}�k��T\�.;;�zS�����) ��E�E�h��+�j�3 ����x�D@[���5�'7+(�����~j���X� `Q���4�ԱqG��iE��9�c6
b���<�~����ew6;����x�ȳd�0������BAH�=��a<̓�N}�^W��<�uE]��ϛ�	%�hp���OKy�N��?zϜ�Gƞ��-4t�$��Ud�9!'�h��9(U2�Bڀ�zנ��Z�k�&v��ۇ������t��QE��nC���������7p�ۿ��6��h�h�-�D��G�A� ��#I��i���2a6�{�O�DƂ��y���Y�Y_�삳vm�eyL?%<��?hv�[�|�H$�5��B#���͚�.�a|�g��W�S���7q���޶�w�W���5�;�����]��f�o�b���P�沈e6�Y ���"fD���`��Ӏ��O�"�E.a{��<O�`GBgQJ���਋��Y�Ǹ8��0.Y��զ<�is�5/�(#�W@Eηͯ7�M�̑��Je�0��pk���^��
�Xxi����x��Oo�Q�ٹ/Vg������!��ң�F1��'��I��j�B�<���l|���h�Ѿ�W���Qp+��yeCUW���A\3}����\u��>��;"]��{p����&�2k�}P!9��=dcԕ�y����tض�1���Pa�Xo�I�_�����J�aۅ����9C!���2 Ɛ���iڶ�cs�<���a��վ@Q����c��OS1�r�1�뵓� 㔨6#y����0�͔I���o�FA�*ԻZgZo�k�7�ۼ؟Cy��؄y8s/x�vp&[����gf������dF:�g�	�{��|_x|�-ȃ�Q�΁��t(Tb{�pf�b
���	˳-N6o"��b��
S,�:��_"c;�3�c�3����}��!I3�XQ�X����<���߱8����@�.��~�����o��N��L8���*S�3KV����ˤ��f��-��`m�l6�ݔ;J��O�P(t���b���.o�گ��AWz�w �ࢿ����1�Z�7M������(/�[z_�ߗ�]=�<��^��h����2#R�K�m�0��2��/�YA:%Wc���	i[J5:a^��Ť2�f��-
Q �X>:ԗ��Ĩ���#�سk�k�ѡj��9L(
d��߹F{�`��h@:�I�[���Ex�&-��n���0k4TX�
]������v�`�jPl�Y��,��6�ĥ�b>!�nH&3ch��Y^��Q���+��*�-tI��mGhGYYr�?'�Y!ď�qT���S6��ޫa(�ݝ
�{戇�H���L����@?����Ҝ�E��s��t��wf�5�bq:�5���P��q(�*"G��I�4�KA��%j����hc]�+����!�9U�xS�`K=C��,M|H��@�����SNc�q��O͸�V�(�������pɮ��|�i�#c%�pL�XvL�_�On����~��I�H_~;��x��|��Ŭ����4:�X$5��;���ߜ-I��\��+n2?�?x/� =%�T!V�
Aw�|���Pm2z�r���n�Xgv���nF?�K�q��*�tg��dұ�(��}P�O�Ǚ���q����ָf���s��ӊ���#�-�._~�Wݘ�?՘��w�AZӎ'�ƓvE}��NK�B��$˿�P2����ͳ�|�J����=���0�D�<��y�Ӟ�';*A��3�5́:e9�}N,�8o
��F�6���i��2�������<e�g�G�B�ag��W�mL&�A�(���]B���X����r�wCO'}[q����ݣ?�)ڹ�������yҳ�Z��ϳ(���9!,��7�GY L�#�Y�(�[��,�~�s��-��������q��Uw��qϨ+!oR�"䨀J^aUR�o�ס_��y��i〘S����,�"�	��a��\ 	�} ZN��.f���"�O�9��p�Ηi�l�-}����/X7�y�~h#q���B�bo�(�}�$�V�m]��&�{qC��L�Q7{�����R��Y%�o�Y3c�g��@��_���2�[h��5T��yyjZ��{��tgb|�j�)���Nm���g���aɬ�����T�3�o����z�a��w>����پ8�6-~�Ij=�ɾ�j������ 	��si�����XB���IT���[fz�6�5\���G���u�Zl�9~��^��Q�Φ��Z�5z�a�8I�s���솝|��a�4���Tv�rގ��ȿ���ֳ��y�o�'�P�H�7��~xӽ&=򆄍�d��zV#ۀD���e'm:���3o�i�Y������4I�����kj�g�> �����C���!�����q�Ʈ�9�7gy�� �{'��FT��Ft֚���cyҔ>_�!���+tªRMdb��v���/b4��H/g�AeT�xd�Զ砨�N�"�ݳ��Q��8�������TY|�.�:��F��Ѫ��f~����񈏊���S����t���|\	����lǘG�v'�8��O���w�?�M.�JE+W~?�Q��ɖ��T~T�� [�/"�V�̖�mD�-i��R���dFw���Z�A�</���I��5.%7?�N:�\*�w�+5yxѣB�J��"���	��/��#���w$UY�߹�n
hf��Ve,oy�80��p��w�ˉn�R������>��CF�[A��ǅ��&׈��J�	&�&�55E�w>��p�MQ��������r���!ʶEȬ�Q���,� �brRϦ��|����F��5��՝t7t�ހ���w"3c�����9M�1�q@^HMj6��J�B�\�ĭ瘯��YU�W%�"��NZ�9���q��g��t�m�!m���YK�i?'k�p���E�ZX�݈��.zJ�Tlu��(� ���o���� ]+S�q���o�1�Q��Eu�\QA�'���
D�Z(YI(U�8�w�3!
R��O���}�wk/��	��XX0@�Ѳ�:e�4:�#"���K3��Q�P!q��\x/�Kz�ua@ȥ0O��=;�����1@�I:$F�l����KY����6'0a���t����Bm�y<�Rۧm��et�1��r����q3����p��C`�g[H��n(�.G1�����`� ��⋫�����ix��,�yL�������m��U���ʫ��@o�'��}2ñ���
����Ox�"���#Q&0�@Z�EA�0�gÐH�F�rsAca���ڿ	�]u�U=�Y��c^pr8�H�p5H�J��e7>����rLhiʬ�c��������n=�&�L@͕Ӯc�a��g��\V�����Z�nq�c��`j�0�Cv��S
�s�D�*a^2��y|�;!j &�O���Ħ.�G�YX�,`�p ��ӵK!�M�0����I:v�hO��lՊP�)�W���(V�QQ7<%Ä�dL�����=Jܰ�>Jy��T��Z��M�>�~4Z@��Y����U��^�:NC���p꽉'?��/��2��^쬥sfJ�����j���V� ?F".Ni?7g�E�z�.5hŲ��ֈp}hՆ��-��Q�q��]e(o%�.|d^�sAg��]FXz���CgD�D�B�{����w.]9ܦf3�nk���:��C���m�f���x)��{�;���{�>�g��"�ݡ��+*c5�sU�lve���DK�[ �`���l~%d}ga8�{��լZ
�� �j���OK�d����b�06O�S9:2�D��s�l��$rG�n_���v�[��#tb=A�pI�fl�)�VA������y«H^�a��g���L,��؋���]p�@ߵ2�J�� ,�P9Z3��Wyۉ+��;-� �d=t����5���N���V�t�>�maO��e�[}[Æ�uKH���3����~H�{���\�_�ag�|�m����j/�װ������B��J��a�:{�#v�[��P�+m���@2�tok19�Ⱦ��_���=�-{AK�(8���[��۽|�3�~��s�kߧ�+߾ ��y^���c.�ۚ"`.E! {�$�����+	�ޜX��k)��O�^Q�G0J��y��ԩ-j�-��e*�[�oiL��-�r8z41/��4���-��}�>���C�ƍ(�R���h��m�eT콩$�jqL$T��5����Ԭ����rܠ%o�I sC�E�fr�A�k����|�
�K�!�^���䍻�.u *�p�(����8e�~J��1{��	c+
��܂��ɢ��߉�F���C�H�oʬ����$3���.r�.G��5�1�uj1���Wf�&o��5�~���޼�a]B�n(^'7JXyX`;�e�(�Xo�|&��0���H;����ec�3Оx9�>nYS#L�s1�f5B�N�OS��(� ���
i�������`���׺�1���Y�@��rן*���k��iֵ��@����^��9��R��F|�4��2�**�L�6�}.;ϐ�+frkf�|vX��e2wF��nWr�EO�=Wׁ�:��y�)�`���-�
�N��}������H�b���WWZ$� C����̗��'�2ƅ�4��8S��WW4�	�����n����!�����[�[̱3��lT?`%?�ak�1dm}���R��M;�#���h�^ݩ�d��6�X�H���{5��b�+ wc�br�M���g5���Y�%��q槶`~~)���m*�щ�F8�sK�KI�X��yx�>�e1\�ՆC�7{��9=�e���Q�7ң�Bh���g*z��Cn8)�*��e�\]Z+.�إ�2��otҳ;.w�J�&}#q^:��`J�)_�#˽�o�BW�]^��ˊ#�9ÞM;����o`.���Lws��
�i�u����&Tv�f(A�&Y=I��~���y���`:=;ħk�C��Q�x=au��[�ěmN����pu�`�E��|]^�D��\�Y�MPΖԽ���m�_#��F��v��9f����S̘���i�kX�\�y��c�qG�A�j���B�u�km������H�E��*J�>�ZZJ��J��R��d\2�H'�j��Ǯ:�L	& ���\G��uY�bή�d��B�W5�����X���v��vQ�JSR+</�+�t���l�PY&�(�>b�4�{/�ӣ0 "�����+|� j9�)�����*�*�2���c�%x��Th(D�Mf��#������N�8\'�Q�ȸX�3Z���M��S"�@��>4:V���
��ތ�;8b���Y����0�]f[r}�?UZR}����u�r#8��@�>���_�jR��3�:7�pn�D�p�^!Q[mVr�a�Ց��	��(���Dl���Rae��!/*R))T��>�L������H�R�O|mx�$���ئ{�����~��L�v��B�vh�5�Dgy.���5��u|�FX��Q(�fQ=��͢4iH�Y2�WC`i��|4>����_ğېxwlK���39n����O�BmDF��'|�X߫z� �uI)|w�<&�l���R��+�~�̧���/�:��G�C���D���;��_�B�`b:x�ؽ#�bݜ$���G�I��L
��Raq�r<;�P ��-õ��"V �,ԏt}x`�l�m�OkG�>{��W]� ��v�i\M2[���Qa��������6��ݞ���.�0s�ڇ��{_�l�*���SGP��.���#2���Q� f�5y)�/`�5/QEpg��G�9���c�z=+Wr�q^�79zm�R�Hg���Zpݔ!����K�yӖd&ڈ���cj�+nv�/�����<�-"����HoABD����IG���9�?ɲz���oӛ�{�@��u^�-NH�\�涡�:J�w����
�ɋ�,�s���%�8��c!:s���5�h�/ |�IU��������-���t1:���p�)Eq��	H�&L�-�6�D� �/��͢OU�������/h�#1N��B�Ӊ.��K�vV6�?�J�gy���L~� ��H�-�v���."���A��Ƅ.=C�o�k��%�Q{]�-c�.�f_��X��b,�5���Ka*��$Z>��D�b���R$ %%�X�^ͬ�Rn�-�_�v�8�R>wL��kG.�dq�J!��$��͘��w�� �u0��H��J�k��w��!`Y��x"�ô�{���Ӻ�u�F0��t�#j���S�Zl7<�%Yg���x~�7���b]����#^���4�Ϩ����Oȟ��(�N��)�\� qo�������(3B�����R�٫��E9I5�B_��GhМ�񒳓Wp%�6�8�Hl+����l�-��z^��,��nP]ÿ�o����B���q����jV5��Ͻ�y�@%g_��ח��n�=ZP�g!����������ee�\0��_I���N��R _��t�t`�L�ݎ#yhO��eX��4lhYng��}�>���B��!f��˝I=J<�!��lW f�E'p�'��9ydΪ%�	��fȼk���b��*Ud��)��N�}F���֊���c8CCk�j�Ard#��ܐ��U�2M�|���͉ܲ#0�@�˘ԙ��8ƛ��I�GZ�W��ċ�AZ~�-N��(�ۼ�	f۰�e�4\)�S��Zz��~%y�Ѣ�+�	K���Tlh�=�V�Q����;H*o�D��3���[T y�3\M~W�L
v~Y[=���=pve[���I�Z�̛�����K	�N��f�-AS��,�G !A���%���V�b1h�~�A�1��ÛZ���t���[�(:}lm�����W,0�En4Ŀ�7�=���!�wt�����I�,�|�`5���meU~��yV5��ja�㱴`#����3$<�����_p�K���NS��ZM����B
� ���tL��������V����Q,F���dVE/�5x��	��J�h�/b\{�v$�v����q��R�Dx�kl'
7���\�KLM2b4�?�'k��֯�!����WV��ɁV�*��$�4Y��3x��;;�{
+�`�99���v�Z$���=���	�ߟ��ȣ�4]����v��fZϽR�#d����VWc�s�-�$7��>N���Z�.ߐ�$���ݧ�s3N�����/����cо�6m����P�պz�.!&C��q�G"������(9�k�x�`ߧkJ�+�������E���=�EP{Ǯ�&�ٶ"�:0XB6u����vm�M9Ⱦx����z ��?.2��B��ST\���4[ʳ�͍����~�"��`�e4GҖ��.o"mp+���`q��?��{Z7t�UC�BäZ�o7�Ʈ5�7o�*���d{Z�(�E��}�ފn|~�7�=�hA,��Ю�\�R�4��O��7O�ڍ�Z��:���tH��т˫/�̉-�\�r�._���aV��,�(��(C_h�FM����տ	fn��'h��Z�OG��(	-��I(u.u}O��x���J�������ѺɎ� ��V�	� P�����E�m������w���x�DN�_ٝ���eH�o���W�,�C�a\��g>���>�l8x���hG:�#:�f�e�)�C�}��^���<⭴���ɺ�Q�&����F�2�j�酳�[g&�c~��c}鹵ң")�e}7`���;�&�5k����E]�Ap+r��.��L�Z�1�SV�X!q!�q"�*��,�+�����ˆ�h@��dW�kM�>��J9��M�����iP��;��=�f̕���\���s�nG�0�@f�,`z�.��@��o�����V^%�;w	,EKt� ����둮�Y^M Sݫ@^��~*�t<���#�.���Av��zA�;���G��B�'E���
�ۙ����ȥ�eך���{j�㎉jJIt��M�"/�js^�ݣ��@��y|���[}��.vq�W�6�t'�y��@��S�˙��̧���Ǡ��5����CR�& �!�)��g�d����S�Gmr�n��&	�
��L�e)O �n�ֶ�p�od��u#47xZ��-�|دثQ�g�&6�Vv��C�᧟B|u�j��>���V3�QL��)�"�t��^<���*��K%6G����k�e��W7�0��8���_@�-�G����~�h���z8�9 �����!��w��@f ��ꓡ&�'�i��<��L��F��-}K�������!:��vri��\t�3�#yoɒ#8zɺ�<��'ux23 >"7iw�� ��f����En�-��!PwOI��1t�M��Alt�X��!�iG���z�⣧��$o�R���*�K���D���(-��f����&�ZI����&��vM���dY����>���Q��L�h��`^fK*�ͤ����0e�)��7�-�Z{^���  9[��� ��X�t}�c�v�eI
M�����NL.7� jv돜������:s����WK�6��|;6c	��>�99ʲt�jh<�2�{�~,�Qr>���ᝋo '���F�
��߻���^�$�;޴��R�|bDqx��i���Uh*=�͞��D%���-�؁���c���o��Lf&n�s��Q�����y佂��#03[2�	a����<dZVT�kh�����r�r.���I�#;+��Ş��!��N��}%�܈����Z��3Ø��p��ĲI����m���N�ͽ�ׇ�����=C~����Y�S�RY�5���Q��������`����U�gf����o�γ��O���wU#��q=!���>0�>�W?����3,q)?���b����%%A��0��%�ƺ̖��M��6^�N�V�@��}�^������r&�4�l"����.�n�n	@Y�h��Z?���neeT_����g՝�}?�H18��P�O���{*�4�sG�0j�H)����M���XR{ަhm�36Nn�%���j[ݴ���C��Q�o�e~4_���V)��2;ػ������x9�i�>�ZFf#�_{ݓ��-|֭h�ޔ�]��E�qD��R}��9}?M��ߋ%��r市���Q�����Ԅ%��0Q5�nM��R�ƣX(�x3ׇ�����@��zw��uu0��W�!���?"=9�xK�Y%q�,5M�H���=�S��[`�˘.���~/����Z8���A]g���&�!#7B4}�P�&�܍�?�������7rR�o�6��H�5n!t�X�ցߊ�h�v��`�8`C�An�ϨT��Lg5����`�j� �c��^��.n��������v��Vb��j{J�n��ʱ`_��q����U�&l�_nU
I&��`�,��ۅ�8ɘr}dd8H���]�Q��'߲TȔ�R{�eH5�.a��\����ʽ@��+?����J� ��!���c���e/�6�@%3�w%�)s�T-3Y��E�� �pn\	��pa���B�n6��P�Zԫ����^��Y���}��sh���}�b��
�G]�CNx����3g�T�領MP�]��D�A����$\I"k>�
{<JPD�@�<�����w�_���97hyl�F���D�7T�×�����Gv�1����nM�m�D� ����Yc��SqQ㵩	t/b&�>�H0pJ�]#���x01R��hM��c�	����ɶ�W2p��	�Bl~����~�� ����ͨ����N*���]��L�v�d�I��ٻ���?��\��j]j޷�~����y��V��|�&�AI���~�"Ͻ؏!�l}
XU�Xxw�i?�`�^�v�?�cR}���������-�?�0t1G'f.�S�S����z��oޔ�A����x}s�Wz���iV�"�h).����i���e|U}������W�,Y�x�	-����]%N�Gw�퇁���^>L��[Nh�;8v'�^�b��a��Ϭ.�f	���2Y�2v�Y��P�һ��`~�l��gcN�B��Z��d&S<Oe��F�� �9P6 � ���+�{w@���t�Y�K ��F����D��}+�E�T��5��j>�M�!���l�"�>-�5���l�=H�e�_L���p���Jr�}��̭yq]�.�AG�2V� �b"��I���+��ϙa|V4	sǅC3������#e���e��}�q���Z��{r�4�'k�l��$c>���k}��S����J/����yjT�'�<2��u� <S@�O�	l�V��}hmb�U���+�`RU3g����T��H0���t�]��=}H!��8g���A'� 璽��I�\�)�L�������̌I��$�G0�F�4�$誳J7��(�XJ�q�T��ԃ�s �J0� ��*̮�Wԝ��V��Eh�����ڈ9���հFҒ,��b�������0��Z�;���(|,�v�'�RU/���	iػ
}�X�,���8_�j}�����������10����%z��iPO��j���L*(����B�˺�Ԗs�C�~�2oO�)�?���m~�q[��i����݁������I 0�>�Z�$C����R�7H�|���s�Gw�+�su]�&a���1Dh�=�U�!���C\ڍ���P�z)l�Ͻ8��`!#�=,��3�=Ԝ�;J�%�J�_�:K��_�'�um�������J�F��Y,!�M��m��ڶs>�ԣ�}�4ߔnk�`���U8F0<�Y)X�h��x*�&G��>�����D�_�(��g�}��^Q���M�ȩ"0��1�/y��@<-C�] ���گf�푍y,�o��.�yT��ݐ��JM~���<e*U��_F��M�rz����c��;C��y���@�̞�_�w4��[��r�6A��A����.��~��+S�S�R\�%����_ny�;_h[
 �����ح�ܨdJ��{L@4d��]�%|�J�*ә�Suڪ�N�5��L�h�RU�!7�|�G��`-����Ƒ�_Āi����9m�Ax����R�n��=�N�Nh_NT��pۖ:lr�/�,���н�����%�$Z;<�+.��u�5ku8��r��?^0+v8�,��%K��?���윚����6��37�D����j�x�)[���|_�(�� �1��k���Cnc�p���r�/��z�fCx1fqՆ��}E�z�QE�õ󻕔w�E�ʲ��J�&�Tb'x4Lܼi��A/���Ѡr���́�P[���V�l�-�i���'ͅ�G�b��AU�T���D�D#i{{�hP�����2[_��d��Y�xyI�<GAhG�!w�.�M��{�O�,g.i�v������N��9�м;�]+F����$��wi<}�Yb_�tRcoB��ÏI�I����]v>�in"���$�G,��dhmp�?aY������7�
I��!�z��4�m��F�$�閧�^��kĺh~��{r���K"?r�D��bG��&<p0����\�(�ܚ^r�-0'�]�<���q��ɾ!Z�  �"����z>�?�'gu(Ӻ4ޠ�X���D�FX�޻�������������#9+�,9�*s٫5	 R@����@,M^{_���	2Ț�Y��쬙l!���oӢ�{W�w���h�JI.��4�f�Z�7��h��e7���z�pf$񦥚���������4��e�{A���0��*{�ocGrs�� ��?���w��Oռޑ=�ȩ�F(D
v��jjR݉�4��5�X��,ל(/���]�%�z�#R};�����2p�F��Y������P976L�H<i��$�(�e#���]��A��0�¦���
�'�(89XEc~B!3$q4���\���q��f��2=���@��b����VV���֙�K�� <�-?P,y�f�~��Ve���yD����L���J5���cQ�3G�rv{��B���D�*<��X�]�tuT�?=��l7ITj�i��2"�
(=�9���T����\tZ䴑mb��c%�.�dJẃg5
skD�����Z��q�ő%��̘�?��
�厂PCZJ��O(�A�j�\��4�t
V������>(�: ��w��Q�D�LZ���w�Ko��9
�*"�\U	� 
g(��v'���-1�g���9D/(��G��Gy�F,jJ2<��RFy����ſ�-k+����QvAڣ���	m$S�R��UND��T)G᠅�=35�^I_uC�[����)�j����ʌ°��%)/�X(�t����"&��Q����xI(�u�g�4L�{�5f)Ɠn"�$)����uh��±�g�5/���G�4�+T����9~�dj�hg�JZ��c�Hљ}�l_��D]�%E�j�[G�	a������C2i�=�b��S�Xz��7�\"CK�p�����NЪ��xu�᝖۸��ߊM�<ɓː�q�oMm���=[�	�6����4OC��źUC��&��CbӚ���Y�pi�l=�I�{��� ��������qs�%��9����Y���Kwu�l#[��k�FznfaK\Z:��D�&v����@:�[���X�ԟ ��׀3��>
w�Z�~�L�.<��Uǉ3�.�[.�ګ��c�Vqn�����Ѐ���[�G���u��v�C���"AU��s}�L�}���w�[������'�m�M8n;a!W��j-C���
%�����v���|5��8Kr��t��S��f�Eja��y�!N�v�08�)�]��ro5ե�"J�q���+�
���zn�F8\Z������Ը��brZ	�ִc�m�΋Y�Jazbe�R�[P�eH`�Q�'�_�w��8�3�=��W��H���&�!_����jS�q����d�:X�%U>ͬ߫п�G�{����� ���V�j`��9$�:���ys;kbC߻�"ע�(�u��l"�T�+)�$^i����65g�ٗ!���}l��5�I|�uY��TPD�f��U�Tkk�!Rw����wZ���Mw7�b˭ FSۘ6�Ζ�e��#
�i!��,4Tqu�I7�^��4��'X�32�f�K2��Y�Pj����w���H��Y�iۓ��S�(�㫸�_^�0��Ej@c�^�R T�+��1)A��W�<W�)����Z��Am'�b��|�3��)M�嵛��E[5T�jk�/&!�ʊ�G�a!��aG�,u������di�*���X�Ԫuky/� L�x$ *���0+�2�qg�3�d�0"��}�C�P���:V�0���@���G�%`�H��R%ƑzuZ�"2��V�Y_q��p�u��X{��Ԟ��Һ%�'Cwٚ�(^D�*��ZsU�M����ֻy)�p �&W?cK���l�J8�� K��O̩��s��ȳ�2W�/�2w6�K���IDRH���� _}�["],��$�g]�z�����	YG���B&7�P�U͎1���x�k��\�=q�!.Z 4/��9�@u�a���-5r��4_C�R���o���c��9���;�^m0�{X]c@`����B�/��r�v���M��F.�-8K�x�gM3D5��P�)��&�$`�S=�2�tm}4N胺�MuW$�椋�,�e������Lܬ�&8�<��Ȑ��Z ���]qcڻ"I���o"bai$���a�u��g��y|�ka������������8�)�Aҕ�\��-#���5�;ː#�d��ǫz8�Hf�#�ѫ�#�(��/'"-�p��H��Ȕ]d��
q�a�0��\#�߿K�i���/�m�� ň�*��&�a�Jы���Fr$>�zLW��]Е�6��;����Q,���>���r��lJU��(]�\~$�(}?m�Q�_Є���<��Dɑ��T�h�h)B�Ԓ�UU�8����|�p��s��l�'�U�Z�$M�>���J$@�3W��'��ϕM���[@���X��}��X�bQ�H�d��nONN�X}]��O�`)w3�=t��!�~*�j?tC(+��	��c��&�Xb������N�.Ť�V�{�O�`a��)�Js����[��]k��@����)LHTpq�$���'{��1@��c�&�,����^`=ڜb2Baw��<O���&�V,[�1�� ē�OG`�yN�f��������Q�������#[��}����ew��CȽ��D?݀( *E�Z�|������:������������MM�;�\�غXe#��.I����ND�Xհ�/�(T�$��J�g�,R��bWA!x֨T�U\�z�Z:�ѭm�9�y?%�gEK�e����ULm]�����MpWj���I`"b�%�6���`�:���V��U�/D������������Z��*�g�ՍN#�޿���)pD�'?y�xT��=3����(f�>�3�8$��nۡ�7!�9dt���|$�?"���Y�g��x(W��|n�����DܼI�~��9M�T�~N*c�a�z���c�����C�����L�t�����Z�];G��.��O��=O.>	�{����@?V��'���Rs��"?��=75�*�1u�Ψ�-"S?͓�4�'GcIU�sO�f�0�����yڽ���t^�(]���f����Yv�4��?P0����_���,�瓏��Ȝ1�p����0&�w���z���|�D���K����)��FDK)�M����Y .NBt/�vӔ�+��ۘ�*%8���O���<8�(�EӞ�(� ����.�y�����y�����\Q�D�"����V�
��7�p"���-����!�&1+�N�S�5�+�%������or����))�]�鳞 ��q���'C]�L��b|bEOF�*�q�J���>�q	/��ߣ�V���cPh�I��Hn`���~��<f�굥&��u��t|rέ��K+�5������53O^��p�|���Q�$��p��i
����tp�4�����B����PӤ�ӛ�UDZ�Rw"jb}+��	+�ѱ��]� ��<��3�=��T�#�-�u<�`Z2�!���a"��5��0jC��^�X��V# sYR:��j$w3{v4��#�i5Ux��#����<(�ʣd�R��3�[��\�g���n����힗1yߺqoB�D�����R�d� p���#�t�-%��n�v���b�&� �~a�p��w�
���-c#�aNgd^��U6��*�iR���Y�w�L��+0���k�V+)ү�/T�M!�Ds'�h�9�20ű��y��;����>��"�C)@X��_W����?D���z���~&L�"0��������ä�b傼�2k���(�bBr�7��*��D}���-!���Eki������{�Z�� �I�Wl� ?ON|��\�SjӞ�ڟ�>{rG��7e͜T�9�+��@��T�����w�p+��P�u�eY��pe��S4ч�H�ދ�I)����{��-O�c8�\�?r]թ�P������Aɾ
˴��iO������P�풒~�������/&��O�}��=����2�6g���vؐ~�� ������ά)=L^e����BCk7"�6����������*ː���J���h��Fn�cc?q4T�K�dg�����3}�3d>f�g�cp�F�:���9�������{}��/���e��������P�Q4��	r�d����~�~���^���4=�H��s������SR��o@'ih�eT�a�6�������o釙����7�.��Ud�����.��b��/�y��pL�T@�� cE|�})1�_���{�}�=�N���8�	6�B���7���s��Ljf�a@K�|�;�e;�G<}�?B��^e�%��7#J����h�%=M\�m�A��:.��>��o��,�7?)��~�I�t���ǀ���u#��c�$z��B�r�%]ѭټvp�l�fŵ�"�/ڒ.�"�7��s������30/��<��P6ȴ]�6�˵��(�d�
��9 3!��D�y�Rd��FF�&jJ���"T��\�����zd����/�I ��EGA�:NuP]H��<è5pK��𤋮w�1͛�.��R��U_pFE���@�!c���t�];v�=�d�#� Z��Htu�l�;.w���KO����"j�}C��h�'iYź�M�����d�DgO��L]!��E�^�Js%9����*������˴��F�c��I�J�p��{\O[s?-�ީu�Aa��/�r{�e���\���@v|��b�x�'Y���du�;o�u�'U�}��1j�jt�h��*���ٲ��v�zsrdv�n�s��v��+��4�+EXCA8�N�c��"���W?H��U�l��3��{�]�V���M0A�@���A^""#��U������i����iJ��\;*^Xo��Q.{x���	X��`��x��\K�\�y������@H��X㧔Ԝv��n��cy`R��$Pr(��A��!N�ws.2���PR�sQi�:��f� i�RB`M*���P�_}���H]k�)5_�
�1PȜ�ز>��^�bv ���%��&��|�q9ҵnI��;��V�"�����4
`7ł9�Kl�4rrT��-�#Ϲ�Ҭ�و�d�D�2�c�b"_!��c�0T����M����j�O@�3S�SS���Y)܇;N�NQl&V A>�u&@��
�}s���~�8h>�W��~�J<���
��$�d�e^<�@�FH.�^�,��])�p����.�A�`Еŷs'����P͞��L�ĉ�s����k�&5K�B����ֻj3��j��a�8<�n<�!�m�6���S�c޲YɋV� ��b������i�'M	�E�6�R��D|��m��(����b�i���o��R��ʲ�1#P��2~�6����z�%D�b�Ӂv�!n�fש�6,+R���Y*t��D^�!������#d߷>�-��E����ˡ��U��hG:3����6{Ϟ�Ka�{\l�F���4_���u5Q2��w� ��0'�����4���gP�K��
z�ƘZȐ=��B�=X�]#�lߙ�[+�3l���X�l_͞:[i��f/v�O��3�BZ���1�=�w<r��� M�҂?�T\Zڑ]K����Y�n��֨g.��|4�%e`Ǒc.-)�v���v"�x?���s�����!>�lP����ıf���҆iSHmI����<4D�h�꓃�>*���S�墓6v�6FU�d=Ժ�z���uk@Mt��Oj�����6��TS�E�p����	���a����Y�7Χ��j��~�H*�=���8���=�S��ꔧ�Z�:*T�!��.�ap��	s�_��gM�����|s���N�U�YE��~,G��'��{T�i�h��m�3��w��e2ծ�4�rQu��.��w���G3��Ҵ�&�_"5@�j�d��?��}ˊ��gD2�vܠ�%�°34���9@N�����B�auR�D!;+��Uhba=��F�sAM�џ:��w����PZ��� ��d���@�Xr��h�`��3rĺK8�6�Dp;X��	�q'����5|���-s��`�$���A����'DPK�Y&{��՗�\�[zi��Ɵj�i���F_;�
Z��/��˫���-uX}#��7��!(�?Oq�/模h��Z_�|�2xM1%M�=Z�ٮ��ؑ[L<�:o51����ɂ�푍�^��#��#��4(8���]>~u��֠��L��q(ҲQ�w ��h� >�L��4ǆV�FV({��F���'�p�Rh�����E?v߅1��g�H�ΑwGZ���|��Vj|�_�_
�{���":X�F.�L�����V���J�5�`/l�X��Nf���R��O�_�	(^B������7rk�<[�a�_>.H��Yd��8���%(Yx%*l�7N���,��ǩ%y�-��X<�޺�W��ֽ�Or��Oo��x��rs�g2V�'�F�&��N�m�RLz��<��z��� m�x��5�K���~o�$iC<,9�{ɵ�$�Vӯx�s�8SK�b �@��F������~�$��ŵz4�h;Hx��g�Γ^��7u���}-�ajD�!ټ"���C�.>�L�^��Ӌ�l�B7��#n@�V���5-J"���n�Վx0sb�Z���bv�S�M�{�Yռ4�'"�+l$�O>��cA�bĖc��e�S��M��"��Y�
�lfo�Y��S��O_Iٲ��_��U�wM�Y��.���i����Ǖ�J���[�`u�|p���y)Tq�-�����H����ċ}<s��
�6��̱8Bc:p����Ȣ cV��l�ʍi�@�:��fje'*A�+IQ�[3��{y�Z��'�L��S��]1��`�I��V�#��h�������]�B�י�;,j]!�|(�U�7����+�+������Ƨ¦��z��E�����H��	!����#�e��\��?]����j�"�q:�}���V�TZ�������\�zK�gW9I�	 ߣo�S�>�EH�%�����p�q��U���Xsnº���SN"5TN5�_N�O9ѐ
79�K�b}��1��R�R*E���BTF�Zv��(i�6���rL��9+4Z܇{T����xL���n����Z6!�w���2�� �j^<�VB쮋�k�FQ&-@x>P2�=��K�h���~NѲgV���P?�.M�G�R5���4L��x��t��v���	;�����h���{�6�_�Ҽj=(�X��1���1�f�H�mU����,P���S�{�b�$v�Nx��@��D���iO���V��W��k��oDwN�!������[gV��5�$���Brޡ��K]t�'?��Z̈́�Lh����V���	�c�@F� �e�����c&��jL�w�>|M^q`���W������x嘫>n�@)'���闚_'�56�I��,�>�!� �4��i�IHNIY��=����<�K��3�=�c�x,2��r���χ��U�Z{x�J00� 3bƗ��}>�T{�Z���ș�j@��C8���^�+�N8����'��˱v�&F�P����B<2D�W�CR�!���-)�6��0�d��:���FE����s�;�HkW]I��JƟ����ZNɓ�R3D�v�э
�l�,M���r�1�����?�bqTD���Z^�kr�Eym^v�����q�ͺ����d�LS\X �:a��c@���q%X��-zǓ�A
�� )�j�ޓ�+R����=�Wfy^�=�����ۺ���]�U�3�d��Ĥ�G�<�ժ"B�so�h%�D(H�{b�{��raD0��ZuKw`��~�n�ݖ�r���vg��k(�[$��EUx����\$�M���"���$-�60f�y��tM�{ d�$�'/J�o�)B7��?ϥ"H-K��֩e犢H��:�3�̫�ˊ-f�vM)�N>�-7b��02�>���%��3��E�	���\ɀжKRS6�x!	���wFz�]�����l�RQv��|����2��	tv�/Sc@,��A,C���,�{�~*��S�"�V��6,���o�����\X��������a���Ό*�7h��Cd��%��.)C�����2�m�f�ګ��N�H(Ch�hg/P1��߰�¤�$"}V���v^�6�)�'�+���n��(rA�E�_�0��>�%h7��PS���lz�kvR��"�����:0��Hϳ�AΧQ$1��5�*���m��K�[}z�����t�?�%P�f�w"AX��|���qP��tz��ǌ��z�{E�W��9��X1Fm6��fJξ��S���Te֝�G�͗�i���� ��83�*n�M4ý���ӿ�:ޚi�FG&�L]�I`m#u���#GZ�f�������'sl��YZy�Ӽ�)Vqt��������%3~���AR�b�������9�ݳm�SGY���ϡ�Gf¥R�;�q0Az!3E��g�6����{5����.����[