��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�LB�#q�@�;<t��:�[-���&��5/(���{���i�9�о=�%}�~BW.p~+`�l�`��c�����eB0���iأ��䧽�|��b�r>Ѿ�>���-~�w���o3�[P����S8�%��~<��L͢^h�5�� _[�: �F�K�d]�`�>�P`I��~��S$�����B)˳�\��P��6�����dE�_��[�+rA��Y���6w�����SR�]����.�?qLA����������6�Ò ��\<�5F܃�k����d�k͚o����ZGP:m�Fk,��e��]q�/�~��F�����!��?�� db�T-���Wv�����8��&��BP�8�\�'���"i���1`ݝ��L���ѩg���S("�	�~(��i�;{!�ec�o&a�_P��S�������3`&������g����?����i%��W��*���L��s��2"��,�#���yy�.�ϯc41s�7��O�����q&Ym��Q�E�b�3+�zd��06S!q�!bUDF 4�)F��+u�|QO?�s�|���:�2�[]~NL���3Ў��!�N��Z!#k*r$FA�d^�{�م�Uy�9�S8=&�x9w�4]�}��T�'C+eiE��@�8�;��B�� �˭�}�>�V�
�P��y��#�翢�#�
9���Iw�'cp&)u���D�GI<P�l���6���ִ��R��I��a��j�+%��zb%0Jk�^9e����5�B��-���N���p�x9�ƭo����}��? �i���D�gn�X^K$�������r��)j�o��3���4���q��l�:i���\;�%�����?��.6��_]F�P&����{��;}F2�X.!"���ja5���*@a5lAx_]���G�����L�%�
�>�L[�lg��@�%_�v�kZ_���i��||1{ư�|���j|��Е��;ˣ��ech��@[�����cT���ĭ=��K��Y2��&�e9K����vZ/�E�xR_���0�a��3�8�@Ɖ���eԒ0#R��5�ڐ#��`�T������_Y�V{'�]2����)i�&�ܗ�E# }]��c'zc���@��zr��2�V�|m)�SFYǁLyt��=ȹ#�eX�Vh����� ����t�e��^�Ol�9h���� 
B����J(1�(� �w�����)~$J�hf�g� �7hO*k�����S�#x�/�V0������a�V�=�!Q�6u�r�v��ύs���R9���E�5�
�4�~zj���� 6���4@9�eE�ͼ�5~E�1���c^eW�����6��@O_�@jʇU��P�V��C�D���>�B�_��v�����x��&��x&��!Z"�޵O&���0IFu7�=�[�S��PQ0�����F(/I}�!]}`�4��wZ�~<����3r4��J�*�����Q��rT���h$�p���e�[�͏xTvGH��w)���N7��{�D��͊�|�j͔y��ᱴp	/�d�,Bk��ӸIM���qdӮ��2��[W�6�L���)�;Y��{
a�w\��;��_,/�J���F{���%tI�""n����$~���o�@k�v �ґ���}�B�w@�y�U�w��F*Ǽ�;/W�>%O>	�u{�[%��I�&���/|�H���")���@�`����F��X�W�����/����#�y,��5�Z��¦�M���[^*q�@�4���C�B?�X�������Y�A`��?+�C��
�>q�x#��<R�@�K���7�M�p>�@0���'���f%��m	�(�U�C��S��Ϥ��>[ibj꿢�?�YD���v��j �;O�P���%m�y����Ē'5�O�'T�;�K���4���l��(��T���s߆����w�.V��r:��R���i����`_�Lt��K&y�
�J艪M�����e��Hq!s�HB=O���*w��_�s~.k�D���4<���+_��S�銻�7c�����~���H8"�Ro&ͱ/�D�}:3r��+�M5�%$����HN  ';��n30���I�M�R���|�6��9N�U�(iX�|Z1�R���Y�ґ(�+6�TՁ]�\��L�i@�������x"G�v�e���l�4�#cIʪ����]�}��~����9w�d���#k����)��`��0���Ŧ��UI6�6�;f"\��$N!�5F5q����8��=����JA ����g �g��:���` UEG4r�3�8,�H���*~����o u>d>��e�$pO��Y���V�4�i �M���}rd�K_C�x�x��1���,R�l������Q�3��R�5:���U�0�9Xs+��7�u����l��ʖ0��櫓2���:;TF�ȬY��_�Z��K�xB#TI0�����d�^w������:=L`�����U#�5%Y>e��ϯZs��V���Z��k/������~�~Iy�F޾r:י�$�����d!~$C$bs�Z�ЖG��wt�6�Mt߆��_���j����Uc6Z��ejلtu/ҝ��>+��a0ЋO�� �V�!ip��'kn�fĞ5��� �)�������J��t��yH����~��Њ�r����#�sY�ՐE*�K�=}�jh:��_/�"��^�}�2�]~���9�� M�O�0T'��D��^^�z4�>�#�:C��E�ܮ��
a�'�>aΌ���@�ͩ}[����/B-��m�!�dTܡĻ&z�@������o��>�i @�����)��׵#m�N߀���9��Vam�޸���d�C.��f�ON�r߈�=���ی=Q���.1�۬�;���J^�/���9� ���f�ck�b.h3i�E_y^��L�'8O|�����Ȳ�}�0��,^L���q�ی���	�ϝ���I�?���9�Rs�:Vw�-%��=����B�G�N�������ܠ��١k�Rno䋿t