��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+@e9wR�܄]�-N���w�Tf	��%�9��#�Ac#�3��@���q��#��e3(s4e��|v��A�K���F�!q��À�۱#q�Q��:V���@dn�s�@�֮�}�
8YyS `�s���D%3i�~�#�e�zdq�Y��?8�9�Sa�d�+�F����]���9�Y<����Ċ5%�V��ȣ��K�a,-�q��M����kB7	�����>�ECT��޸xa{����S+.s��pDA�qgY�Vx>%ε)w'=c�g������6
��B:}j��{+/�j��Y��O�K��a[è��W�1,w��p�W{_;�]:��`Z�f|���"��)5dN�(\<�f��\o�}z'�>������5���ٞ+D1~���UY��֒e�]�8������)�X�N���4S��\����,:��{�eu��tҒ��o?g])�-%�6E1��vX�[В64Z��H���[�$eƣ���o+J�v��{�.�N�er���3fL�y������o_|9G���r;��%K2�yy�UM�ʒ,��j)D�X%�)ώ]u�D]�p\>��f���Z�\%Qg4J�u�I���kG���+�I���He�p�7����
(5�zc#m�!�j3!M��8EXBJ�2�ߜ��!Sh��	��H2�P�ز{e�ki���>�2�AO��oap p�͍,���S��)� ���b5Mj�՜*VG�/����k4��I��3���i��K3���,'�&`��$&�E;����8�ۼD��z�#v,^��/i|.ق:��O4+������oF�1L�WErn	J�+3L&�Zco�I1[]Pu{������I���YX������'�"�(*��Ku�$�5B	�G�%����#��H��V��Z$�#���9�NZ�IR��/N}k��ܧ5�0M���SO���X ��u�<Z�Ï�U�~/��u���ytIK%�V���k�K9�@���H��f����v��MEc̈́�țkz��TO��G4v.�u)*�	e��fX&BN����+�Qk^��5��-X	��FP�� �M{-��v��,�g �z�T:�����b�T����u�ڂ�?�S\�Fm�Ϗ�u="=K��t����҉)&�6�ZDb&<��󊰜0��;5N�
�o�y-���禔���+�{2#�3��G�J�MJ�颳]O$�2���Y͐�2�����`��?K�(`���ǚ'a�қ�e/B����?*Ί���d�����'0��M�)yy��3AB���������@�Tm�Ówe�t"Y��_'����z4�)gUŏ@����g6p�O$��s&��}L�i8��߈guM�ޘ�C�Ի�Q��0L����;�b�)Z�#3�-T�3�ǭ�-{6#dP�V��E�_�3
����6�ŤЛ[8&K;*�q�[�Qu����>��1׶���t'X=�{m3/i����9�9!ʜҍ��P5���*�]�ݮB�% �d�e���p������yZa)��M-N�d5�W1`�O�G�����R���,Ƕv���Y뵌�������*���T�v�??*�ʆo�6��8�-��ox��Gh����eբ�<�ʨQ�)�
�G�dm�'�9��SԻJW���5XV�ϲ�̇5��Sx��:A&����\�6��.#/����^$O�M'`�qq�i3�1u�*�({�<��(+�����0V�Y��_]�D���c�*Ϩs~�#ޡf����`��w5+Qb��ܡ.}���sK�	�"�4��q%�ߣʗ�'�E6�ܗ�������6�}�H���4�����cg��Jy�DiGz*mԍ�s�w�P��oܲ@��0�X���=�@��T�\WI6��`��$a���嵫���r�-��>7�md`����
X�!H|����� �ٔ͡��wļ�@�W<_���1әי<���t���|PǤ�t��]�"A4$CFj�<^��VL�	��]�?�l����K�nsV!�HT��ֺ#��o�H)�h�O������s&���7x2�T�����ˑH�Bm�p"� �j�<1/XH�K�0��s�[�3�n���g���!9��o�>�pQt�J!K����4�fe�F����uk}�ӑ	�Q��?�>�!�@aQj��l�ʒ�_v)"�s7�
���x��RJk^�uջ<k�5koebY�Ϋ�ICRn�|1�q!\7���M/l
Y�6�\f��_�k�`�@Ze�67_ӅCG&T�yz�q��)��_��-b�����!�敶`��EٹN��Y����[�(ZY����c����M �|�{(����`�C�(	����a���4���A��C/(��lQ����ow�+pr�
X�Շ����t�B���_ͨ�O1�P���?��)h��)7� K�!+��]&6>r���岠�b��b����+qBt,��>�>�,��h�#
����Q�'ϡ��"�mڳ�N�#j̙zW�Q�� �㯝���a��\��i1�M������́I oPf��V��"/����s~���2	Pi�u2MF8��:�s�5�3�`����=kv��D=�W��kռ=��2�..���TET�G.Vh}��9V��c��1Z�:�z	��<_�ـ<(�+��*��Y�p�2�+��xK ���a=���FV�/���2��xm\G�$�f#3-=6XK�,�qi�h����m)]� �@d�Z��f��D1C�Ʉ<B�3��c^QO}�@�uR�W
ȯ+���d?)A'� )�}�o]�0�&�R:v���)��`���M,l'�'�*Y�]��:G�*���W$9���K�B�c2,�$��Y�Y
�	q��b2�l�x|��R��w���zMD�i�?��B*��O��8y�X�i��u�gG���A�L�q-H��6t���q��Ƨv<��S���*4�'ք��wY'����� ���]��<kp{��\|g�aq���OV]���M���{`��i��8�R�w��K����O(%�M#0-xJc_��m�;�Fq���y�n�<�:�����위I0J��{^��W͛і�{��bl��K: !0�tg�Ω�1p@È���4<�_�����8�*$�U<?�ScfF����H2��G�2�M��]��_�&u�ec7�jL(�"M��'���b��w�=�%r�Q�4�h� � ���D(�~K]^��o�G)f�e�84/�-�}C	qڎ6BG�W�>.e�@������@��0#�>�,2���Dr��5�1����[��̭���
�F��no�������=����r��w�h����v]����0�C�Q�=x����#��;2Qr:A(�(~xM���2�45eP&�ك�Ig ��Q�����]�n�H1�j-�	��by5T��s#�J�uŤ,yKNjL7�ȃ�UîD��\�;KD�K����9��O7��v�d��v4ؤ���r�b�g�p'[��zzgǃ@V��&[��즤xDKX���k]0���E���]���r��يH�+��_��w�$������ h��tu8���8��=]�T��F+݇?�?L���N�ªmU[�������*��4����\X��5 �2T�Z���p��,0]%>jr%j[_s�=_��P�PqF�9j>�-��i��.k
��r�B��!�H�\�1p��Ya<B���;7B����-�m�1�#����tO[�j�[;�^���خLU��� l��/k�Sb�j����ug��M�,��܁pEDIId��f9÷�wS�W�2Q�RA%2~Cxws���!`(���ZE�� WC��aƾ:u�q	ظcU4�����r���r!��A���Z���"=���8�nd�*���)���#~�'�{�P(���`�1�Q��w8�����w�W�WEk߃I��|�vU~�!�R���H@�z5	Q� !=3[�n�J#�����|�����J��HWl_�eM*�*������Yѳ�w	�J�	Z֌NC�����umǙ��f�٣1��CN�ݬ�%)�}�6�Z8�PYXi����I���f��Ҙ��tZk��!�G�	��`n8���ྟ**R~0^���Wf��9!.�U}IXc�*��*�Z"b��y��.Ɛ,o+*���4�^@S�U�_k��&
�mb��j�C�+x����K�qn4?�
�k��X�L���r'[�Vn���i�'�<����wt�qDn*�o���n�]��!��
2O��tj�5��ِg��]���3V[�X(O�p��Cj��G':�_�j��P��3V8�H"D�^l+�
��w=���ky��it}�e�E���� �X��U�R����910D�x(��g��8�n/��Nһ~w�+:�m�T[����D]%Z���H۾qJ[�,��5����Ui�!�	d��%���.�����N�c9`� ��tA3�0~~��<�)}܎s�R�D��B�IM��	��		�eX���]�Ɵy��ӷ��G�_�p�XV �p�ʗ"�68��-|�a��(��y^�Iɬ-�g�(��{�,��2@�r!��X�[�<E�ц���
����q|�_��Cw����ҁ����[���WH�|C����ˎL�ls�z:K]��삘Δ�݄���KX^�B\��͐�bٿt~���,�n�\,U��$�!�5�J�mw�?o�b�����ѥ:�� �"�o2�Nc�UL��D#'L�!��2��e�D���8F���3=�����h��}[y&.R+�F�ޗ�N�,��~��?��c�ҳ����u���2���v�?���_��\�n� ,������x�
���;�u��\0�Db�^��6jq��66�U:RV��,��1jh�'T��liQ7�%����ݳ�m�{�b{oЮۿiQ�xb���k�6v*l-}zZ�� wa�/wl0m:�2�'ҫ�%�}Q���X�$4���7��OL_��m+�Y����;�=�c<��b=i�d�u��k���-ߚ�%�3� ��PM�p,�G�VvuqC��2Բ�WM(���Z8����t����"�[l���f{�Y�}�|>W�3p9]����w�X&doI/}���5z�Hge�.�����q�+�`����b�MEC���s��۸�����	�����
d�.�Uԅv��s�&E��F��4g�e ��Z^�Т�l�t���<��푱K8����Vq`�F�2�JG���SŹ�Z0n�V���HքdeD�M�7ӆc[��l,��b�mБ�0zr�)q�)f�~����!�d~�G�x����U�r_r�n�I�$Gn��V�Y���P��˒���Ve�>6X�
�SS/jQ}�/r�׀ �-�ź)Mد����i[t�l�wv7U�Em�Ptt ,Pu��
՝Δ��$A�	D�����\���P���ha
.�l4~�+�<q��\����I؇�O�_�k,') ����vp�����?9���|6�\7�P^�j��x\�_-�/ �J�?�9����8��N6���7�8 
~@�9g��:��Y���Z/��<�^��gq�8�+zi@_t��ӕ�&��%�S�9����A��??���q��̊�\�6�q�j�;�Z]�]#��m�s��!ۀ57ʚ�Ǎ�-�p&�`�v�r"��Ћ�c���)A��I��G�$u��������	
 ������\W�zf�Ν�E +~� ũX;�8"P�ӣ�iU�Z�WVD�l�a&w�`�z<��m.�<�	r�1��(��x�Wb�s�=ϠD,�8���i��N��!)�j _��Z�T��SL��AƗ�B'�z�*�B��Zα��J����*�~i�]�ʨ�Ȍ�*sYN������<�E�e���):2�E��|q��.#�fF�c�3���M:���a�3�w�.������+�X��u�c�����7�ً�O��LuWU�j:D�m��\	�+��#��N�|[lm*�4����~1�b��h��Ws"�r.0��i���H:@���Ƥݶ&�����c�Ǟ2� ��j�6��u����#�"��\[\3��'�qh�7�^K'3�?ٕ~�>Ns��� �-m��2��܎`nI7�j��7�B��L�{��_���#��wq�q�78ua���Q$�&7�Wj0{,�$�2�}{l�H����1P�i��& n�;�!�P͉����x�\<�1���i��"9ϔO3�$����c[��3�h#�rĩ�"�z�ս�