��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$�ʣi3N�������#UKnT���ҟ� ����Ŋ��H����F(n�j{���W�T���ʠ�� ����*�Roĝ��5V�1೎������Fx��H.Q�v`]���l]�(.��=
M��6GYa��f�6
:i�*�!(s ��j��ߓ�FPz��lg~x?hS�J�@�b��FfABZp_�)�q��L%A��Ps��:��XH�ya��xf��i�Q��c��~�<�
�b��1�Κ�aG�u�@Ge�n!�\@�4�U4������Y� !@m�V��f(�]��<�Vu��}\~~�@��@��rio�[�q���^5Xx��{1I�2�ӎޡR��dV-R_*����9���Y���X�#��f��Ow(�m���=ބ�2ո��5滕ys��ۍ�
�F�����l�K|���j5����E��o�R�ذ[0�fU��f��w��%ښ�����]����RYa���eW]�8u;e��������U�!�j����UrP�
�!�z�@�n���k�bh�����H�g����A�t֢շ�d����`�s��|D܈k���]�:��F��Y��E�-%���{���XN�֖�dt�G�Ύ���х�lG��J�%�u`D��2e
�$�2�T�пc�p��8⹛�|�[fJS��Do\�0�5�2G��xxs�l0�-������e�jW����֐8(��X�G��'������r*�W���Bܳ�l��:ʽr��S��?�`���+ǫS4���z��* (g��a3�`3<mb��p���k�C�`q����r�BP��B*�ݝ�!��� ̈�o�&j��̯&OP��A�F�a���z?��T#VPJ!��\�>Fz"�^��9���L'*�>����Ik�w�����G���EO�38(��Y�;�L���� ?㳵���5�����ب{���ˋ��D�c� ��s?�(�a���{�sOp��o�*G�O�ɓ���>)�3ۯv��*���9xlcT'(���j��Y!+uYg;�W��#:s9�XO���G�S{ZI0D�XZp���ī����*=��7��B���}��^��R 	2-�����|�{#ލ�6�W���ʼ��)��¤�O�8�^2AQU1�?F� ;_�}�P���ϡԟ���4;���ّM�$A�m��-�����n�Ф�F�i���Xr��g��/��	Da;<�}ٸm!�rgN�� �{*���#�+fZ��ߡ t
S���H���Q��⚩��������o���u�K���� ���B��b�pv�ɗ����3K�b�4��\n�Ҿgb~Lc�
�7#��k��� t?��[,���p����a�7���Rr�8�1������I��
 ���'!��8h@4��R;|���M��H�-���d�μ�`��X���Gb!�1���]y�!�xX�{+0�TO��S �)dU���c�4o�Ӡ� �s�֐pD��#Z�z��mS��D4޵@��G=���l9`����Qq�.��՗Q�[þh8�r��X�+���ĆRzi��!"u���� ����n���l&T�F�?�U��9�4fc�1oIp��z5�fR���ϴm����Dz9�! "Y@_C�?MA��/I��gj���͊,]�D����H<ҩ�-���h4�o�r�H�6V*4]X�,�/X��HM]�Rca����+#�Jm��"{A�#O:gS�}��F$�_�\������;M��枳���}��z�1r����G��������힄J���E�D�s�U�M�$0��ky��A�L&jD��\�#��;���Wؐ�x9D�q���Ԡ�����ӈ=���,��P*&è�HnʁY�_��,qñ����W�I�A��x8[��7t:GE�G�#%�<��ok�5Q���<���f�<t٠�Ŷ��^��BF��s���<t�u���",јJ����4�e�����?YB(H0l8y<��e�{�a�S~l��*�i�mK�-"��8�~�m�����r�Qe����kjz!��# �'�&k�������m�32�����q�{'š#`�R��2G3���C�y�p��L����K�Z�'�P�¾KN��[��t!����TI>�;Ò�0ty�����Ca5��j TeA�>+fB�yU̦&�`�c��s�lm܃�X���/ :3j��Η��J.��h
���ܟn�_=������ڛ��'%@���$�e����L�`���i�2%�_u4��Az�O_�C#d0�z-���5��q�ݳ"�!�!���S��u�h8�Ue�&!6��e�o��	h���.��2=6���
��v�m�1ю�������Bv�z�b ��F�<)��wd��j���,h��ln�~�&s`5�����#��2��ne��N4� �0�%6�Ӹ:�s��cD��� م'[���B3�X�\K{uS�Ys��ǝ�7�Rn������P�G�{�8h8G�?��q��#�<�x!���:�|[(_��`*}��Xc�Ҋ�G�k0�˄��fD��a�l��S�r"�d��A��4�'|��秭~�^�4���0�e�lH������d�C�V��#�<�s�4~��k�9�x�"���x���Ҁ�0�2BX��t s��ǂa�#���\\�W����R*ߏ�.Ǵ�!Kv����B[i�<�Vj8����b]3�,r�͔�X�����@��Ӽ��H����uQv��3M��Zu!)j�=��1��Y�tߏK���p�(�UA�(����ԃWіp)���}���e���-�^�/�ا��QY������Ʉ��\UCl��(�pm�3H��?�P�p_9_G�Ͻ;��0"+q�A
"�n�����(G�������M7�A�X����Ѓ�H���*/�8u��
���*�U=���s"_O�eZ-�!98��}��'�=lp'�F���ϫ���B��|vP�1�sE��ˆ�5�H��Yfۛ���4�
����g�ش?�B���
<�r�n�S�r�ס�sT9˙�O*Q��P�9 ���0�cҽ��x7����gp�u�f��;-�j$�*J%5e
l�[zUN�zG7�*��)����->��Y��G��t1v�1��2[��x0,�����!�
9��#
�uYb�i�^��!ن=��j*� �&��.I'eZw����s	�+M�1v �:�7���r$��Y��
�`UR���<�-}�w~l&hyd�"���\���n���$�U>�
O
Y�7XJ�و�Lc�L�7�)�x�A��pJz���/2����O�x��>�bna�;��_���$�%P�$�Ff��x�㷺��	��8������Gp�AL�$��36VuM��h�̿.3Ҭ�m�h�qD�T�2�$l_��i�f��\=��FV��ޣ'�]�6����{���uDe:���.�k���u���NY����j��-�����m2�˫ʺ��7�0Sm.���F����棨�XS	����Qp��	X_v�A�d��e�ʧ�~���������R:}�5vLv `��T
P�?h[G�fi�J�9�i�M����{Ɏ�9N��3�@��YR��K~6���v��I�N�Y���1*��X�5 ܏r��M}�-�9 8o�%	������V$M6p��c��7-�?gd]���ZS����b}'%�������#&�Ԁ;7GE�s��e��z��K�C��vo�,������K�L�Cη�x����MA���C�f�� ���1�نq�??��a�<, ���;�{�?�;��g+zD[���&�`w��(�=V�o$"�Ȗ��W-4�K�ӹ���t8C����'g�=�+Sd��#R*�`��ȚX(��@��5�'D5r��_#`��p��	� ��6���ػ�h����V���琕n��z��*#�=��T��v%���dXM������B^O�T;�ψd�wJ$��|Q	:����77�[�-|�5;߮�V1ଅG�_�)�]C�m�AU:,��(�u��)�)^������(�V����F��N	�������gf��V̄�1"�Vh�����Z��G]�E��Q]E��Rq���Ȼ��<�LwΫn�R�@�ν���|�����$dz�Cd�%:���%@��~A�&A�Iu�[�Ъ.�c_���
����1��X��RZB���˦��z
Jz�7�M}�l��|\v�h��Ro������:���^�r�)}\9@�_�>	��Dv7p�W6=���̺��7��)���یo�1��Ʀ�[ˆ(�}y�cZ�]1��F��ɾƳ�sy0�#|��"�k�Q�Y����Φ��i#�Z��\��N��������̳��B����;q��(�VZ��
��k���4��{�8ƝN��ǔl�������|�����^I(����Щ�@Ҁ��1iT"v�o;a��D[�����|��֧M�Wk��/GP��Œ�H6jbO?�m�������~�q;%����.�7����wc�;�`��t�� �{�x��z?x)�B� ��O<_���N	nL�I�h����;��$�YB��@�o��m��\��є^R��%�<���j��?�oO}$&���Y��?�D����(��Ί�HJ���|~�ss���µdz8<�Qq�l<r5h�#T.�3��(zf:O��bd#1{�
��Z�$��{B�~=l��p+�v��ִ(p�0>?���m��(lN�!}s6�RKG�\V!��в�7 k��?*P������g z�%[��Ac����M�4�vc�
\�˩�]Ւ�A}�r�j�f=��ןX���g���������CJֈ�SX��0L�t� Ϥ)?5���e�B��^���g�!������H<�F��+��w�.G�� ןƮR<���(�+ـ������"�R�0��T�[��VC��^,-u�J��0�[K�+��O)fG�>@��OF���~�����h8ξ3RP�sU&�/jD�C�PhX�o|������j�}�@��r1བ�Sy�6�Ŋ4��Ѫ��HG�������L쥛h��*��#۸�K��y���X�yg�H�
��	�(�ۺ�f���0�t�\U;�S��$�A�L?�j�!�v��4~�ual쒒�Q";�g�̋C������Տ����
9U��6�HD��dF���Q�j̺�nS����Z�?��O�L�C8t��^� �'��-�lW�VE��OR��?B�ϣ�BB牰l�G��0��(8t)����?b�t/m,�L]h	�:��$�~�L�4��ĕ�
4��Y{!�1u%�n�hA�.��ϖ��cu��.����M�O�(}��@������L��o5xƒ����`�q����i�֞uX�.S�S3���q��]���De���:_]�?bH���_�F��R[���<)�����_�*�,���Ο+~u��'�Cz���&� ���;@���Ss�ۓԱyE�����_�P���7Zg1=���lg|͘��xK�:$h��D6R�&7OIB����ܦSM�F�k=5$JѴ����٣kAp�u��Q#�lnG��{̅za<"��L�������j�7 ��1��'8󎹾3CHgm�a%�v��{wY�O�n#���@�Q���x��zr]0�����.��Q�ҁ":�^�/��T~
�K
�k2�����m�y����{���t�I]��L��y.n��K��%�_vE�7��;P�Fa���	����C򶒀Ϟ����|&(���=�qJ�	�S�_��2w��(6���8��`�FW��/~lLx@���0u�դ�?lL�!7�ox���N��I�+��*�m�;t�X)���F�ޮ��A���:��������/(Tm�H�T5'��1w7V4��TxK^�$?&�a��{鮫�es�j:"F������S �$��S��P*�o�� `�<a
lmj��a�Q],4��2��7EE����u����::�vFd�^�d��v-.��:��oUeܕ/�ޏ�P�4����#�X^��~帷N�o��?�ܞ��mQ��`?����i�O3H%R���JQ=����Vu�͌Ś��!7����N���ȩDB`�	˫_�L.d=|7��1��(���6A{Zn!��h�/z�E,y7��l�P�o�����D.�naG�T{�q3�w���EP}�+ɪ=��_�Nma��N�nM��
0EX����H�5J4��!pgH�k����
<��G�U�#A4�0@\Т&�D�h'!݋!�XЍEQ�P�é��
 ���W9�UJ&����f�/��,+m��rOW_�U*��\U|������:QD���k�����&�3I+Ju_s��|OD�WF�I`L[�'�5�Q����6G��B�E�,:pJ[��� �����By�� �.l��a��zm�.�h��Ε�J�"=���f�ː�e���Z���u�'*1�@�ʁ@�2�,� �4�:��R���Ƚ�\&�45{8��#�}?^���?h�>P���\�9����cK��ڒ�����Xuk�i�ަ� �OJQ-k�h��LL����]k����Uj��j�1����E�c���ԌIS`WE d���� 9�LK��~̲S?^�z��/7{I>/6m1�k��i9�1����{!gfAz8��c��3�f�<�R����:��$a�B�Deb���w�)H`��%f��ML���tHq� K�G��Qh��5L���tu������Y���w���Z�iV7��$��[��e-�d�p�fɷ�W�ȋ:�� %E`�ݾ���	<H��蜘�|dA�"��H>�!�Xq�&	�M��7�w�7�o[�B�(���Z>��"(�tb�G�V�/���%6r2��@��w���9r���%	��/^ۮ�)���6��#�&_�)i�Mm*Q���=O�k-d��pw��џ�J���7޼���3�j�r��q.�*��\ͻ��d껒�qvK;��2=i�$a�Xd16 ^M���6��* Q'��Y��R���R'YPn�K���%ANc��w�wM��m曞(+�W�ʨ%X�J�q���B%C��C�޷l����k7�e�!P�R�l�?,�s�� s=��&o8�03�Z�|q�8�*�|�-ǗE^�3��o	���{��}�O���1L�/��joS��|j�:�37	,+i�G(���4\O���=*�Dc���N�OJ�>�r���CW�TC�@����R(E�쟧_ �w�4�/^�L�?�z��#ۛr Û�+��Uk|����2BǕd&�{�[�O^�u�=#YB��O8�Gm�?v#�!x��2K2���_�ލ̭}���)1�ǌ" �ĩ���@���(�QS?��c,����]"A�K�����$0�h�Qt��RB����3$ E�M���kT�kb�q��ǃޡ�_���w��{�u.I	Θuo*�]`X4���>�����������@����JlB�ch����g%1uu����S1��.��ԙ�"l����o]�����E�ׅ�fg�ɡ4��jW���D�Zc�{�~�S[2U����I�KuK�"Cu�Z�e�X.�E\P="SeU����<Qۑ  ��f��'іzÌn�4�z����	�v^��������kx�A���m,I�k�p��5w�ytB�?`}�-�ހVP�W|`B�6��#V�C�R�H�8-I������J����ޚ�z�#v����U���c���&G%�1gl�G؎Ii)�2��;���� >�q��ۓA(nJ�9QB�??6�ڈ�R,y��5�ɘ�����KB	�p�WмG��r���ǌ�o�͕���q�D:Ҹ��@L/���'��Ш۫t�;���4e�Vk�Z�CUĔ�z���9������x���W?��n��(%9�0�rp�{��rɠ;Tp�M����	+�B��=j�q|���X��~f"�A���3�@��xV�h4a�� Gk�Z�����xy��c���������r�3V���R�Kx����|@-��"��;q���<��-\G�䏺�����G�Q(��-V3�긔�?�9�����ޭ7� �! o�!ܩG�Z/e8������w�A�^��y��͝��� �-kL�]��ERX��ʢp*���Y��	�J��A �/HWRZ=�c�֔��sv���n!O�q��SE�H�3���
��mQ���SsL���I�6u��'= ��� �o���p��*2�nE�r���|`{�GE%�0Vp��� �	Ġ��r����kܥ�H�,`Lc@y����TT��O��:2�CFL�� ���yК�EBg;S�t�L�`J������~�YLB�	��Ԯ�~\�hzՁ\#�)�ĳ3�����n;i�g�#��z#��
��5c��5�(���>��]���.0��ɟ+��ҡ�6���VBJ(Ao�D��S@�Ck���VL�~��*]ng��b���P!��-�27� b9-`�y�у����K��AX��_氆*)�*��;$�I-����>>��Ç|�Q��X���>��y��g�[����,�A� �z�\�`�od�i��X��l?���f�����D1����`��f2�da�ћ���Y���:pez3����=�1����C�)y��Ƞ%�peء��*��6ػ��6��m�/F��g 0��n�r�`��%����BU��ެ���l�f��S�,�P�;�}�HI�Ӽ�����=ݘ �U�ﴽ\�yW�