��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��&���i} Ĳ?���3rz��I�{��1MZob��N�X�����0�D�ɣO��ad�U��e9�3�f����Rxe����U��S]#	Rk�ݸOq��CsL<<��?
�[E��G,Q��TN��P;�Xlr�͘դR��[���%�H����RS�u�� iJ�Z�?)B��p�d��@�1�[�R�-;�l?e"�f������ �,��|!�LuB��Sd�i�?B�:�"���kq��V���Hu��j���g���ED���sBV�+�U�1���+Ӎ��(���ޞRD6���4��{vd�Տ�6<dm�x��e��R# !;�3fs�@H�`��@>76�'�H�{��6�$����24I�A�FC�`@ї'�g<;U� �"ǱیE�aR�g�<�;M�l[7��vg��~�Ƙs^&g��x�F�sf�"y�`,�>t�ѷ��L�\�^u3�\��K����D���<yd?/)#?ƨh���Nǡ���ܨ|��V.)Z�T	]'�����3��ZQ�eR�?�_k�/�EdRpJ�ARbp���%�{�hJ`���T��v�*[[�b�cp��<����������C{�2�w`��o��B;�ϔ	�.x����eP䊜tsA���)(��ʥB�VH>#���u�r�>�b�#`?��,d+�T��6%�w׭䛧�4$��6�Ӽx6�ʩ�!Q�uK�`��'ub
J������Rp���x��#�U��f �u�g-�ϋߋ�j��oE�+�:����@\b�Cee��G*�93��ͬF���b�+m&��� �$B���J �M���Ձ�|E�d������خ cڊ}�]tR���x`Z5E��<<B6��l*�<�7T������X��e^�l�m璌c�93��)�у�?{��Ӻ�~� ]p���ÔFyCˠ�P�^&��DR���u'PV;��~���@��	Uo�g�&�΁]�M��_���-_�f�t�������@i��M��n��\���oaZ��HT
$r0�yN��;#̳^ ��4�ހ%)@(�~j&�;�ݳ�����c���Á �a�K����n�b�T8���*��J��D6A�V��-�j}���f�u��ķ��W���~���U�ը�9��� P��A'�o��M��Ϣ�[:W��ܻ���I<#*��L�@7&�Wz۞tv��[d�<���6�����O� �h��?����k�/t\��Z��Z�Xgp�c�'s���|Ό��V}�2�(@]$�簸S�^�W�`��ϕ>���.8�5OA�ۈn�G��Gg؍�|����%��e�����@�.��_;4�zr��Uu�j�-�џ��/�g'����8�]�PU}�|\��o��NT���$W2#6���>(��C�#0����t%��tJ�a�X@ɯ���G� -?2�Ay���l��mL�~//f���s^�w:���F�`㷚�w�������YŰ��\[%�Sچ���1q�����.�tk�;��rW�X�,VTiZ���d1����z(���ũ�2i�_��g�}�}V��b��D·�rc��6+���XyU�47��F9&gg�*��{�&r�2I�/j�r�wUz���d���4�Y��h��M�b]������F=wt��mς�^�u �t3R<j�\�G�|���w��N�c��ȼ�N/�e���U�j%~k�QD��i�G�,I,��
���u��P����|�YEΤ:˾��]�����s�d�	'��H���O�5��fpkE7ǩ�J��۔���Ub�����f�s�U*g�G�#P�6"�$R�qHæ�͢����?�cE��x����tٵ�B6�qh>/F��#I\�o�O�"'\����9{�@��O�������}>�砉�������I�
]��jL钺k<��F@�'d�J8���\S���G��k��ϗI�O��Ǘ5�I��]����!�Υ^1[�y�<���HJ�kk��=[�`_�:O�/���'�N�dà������S���0l-`��T�P�89�{xȝD��9yN���������8&��N(E�!�����ɐy�M1�?L�aIN����[���c?�L�h�ī�Z���h3+J�B�Y����%*^�l�UhHxq��Q�~����	�p/2ۭ��W��k9Z_��<���g"�|��|�����s"�YC�;���W��m��h;�Kg0њ3�0�K��X��S���aF�D2�\Y�<���*�k@]KF��"w���!ָ����t�,�]��l����_�,A��zh�v1@tĝ���C.3ʶ0� gw���z.���7�.��~�()�R�f!��b�oN��Vc"�HWӍ����qD�Z����2\L NX��o=�T�P��F������d�1�I��RV$��U����/ը�R9:�c>o���@��7�G&�us�}3�gi2#��tQܿ��RR�`��z�� �����WÄn�̬�4ē�ڃ�M���=�)W���;��vd�AV:���(XY����H*ٳ�P��_=p5�,#� \M���UCE���i|7>p��c�Q>�U4��&�ϭTZ�2�4�6�	=5,��h(�P�"}慜�慿����{Gҭ�搡���PL������F�b��}q��*�!�������=Y��DS^y�2t4��C��&����L@�#G�7�7�q-E������lx�.Op'b��YDr�����[ U�P��E��O�9l=܎�"����zсH��U	��$YB����v�a���}V��S8N�%l{�'wJ��m3,�y�"�N���3 �O��X,�z�--�<mq�|�&d��q	���A����%iP��h`*�1:P�Z�S��a��3��y~�9��ň"(���a�/nUi����dŧ-7�	���h��� `7_%���'m���p�(����������3�S���CP,�8�z_���v/ht��0#��ņ<��9	�RՀZ&�蓾�T���Q��Sxn��e���7BC� .T�"5ݠ,xm���5�V�xV�&��*��\�J��*����
y�/�.�Pvh�����+I���m��SL$�8��V,����u����=H��ȵ�1ŗ%Z{���J��x(�� ��'A_ƣT�I�3/j��2W��L�%��uۻ�({V�F��'f�����.�v��F���3w�$�C����$dmJG��;�1 ��;7o ����)ޥ�_x-���w1bZ���A�T�����'R��YaL��u%`DrqM��9 j#����K��2�Tߎ��p˜�]��PV��%5�Ӎ��s��	�؍��i=)"�܅��
JQ�u�M�8��;�.��J��g��\���^���a��a��+C�-���r�p6��h��2�����M���0[�	����|7��`���t�����ZݘQ��>�`��ذ�i�s��=�H���cTg��U4�5�]㙦�S��H�� q�Q�rH�v����hкłB��cQ�f�ЖXQ=��9_��������Î����Kl����Y|��k�m��:)N�N �����1o^V�Odf�/��?iպ�е��0x��!�1sy+w�@�K�,��=At�mD{%��֔�+�8�㘨�t2�M�j�bztQ��.�ev��辤M8��rW[�d�[I���!|< U�~�Ϊ���@�u�����<����>ɠ�)V?��߆��p��m"����@�$%�;pi;Ĳ� ��s���v �z��8'�m���	�_�l�\�$�J�U�Ө3[�i�S%L�xny�k9kf�-��d���F� �~h���G?7Մ����)+âJcg���2��dtf:ȟ"�N���JK�LJ�['��sM�̓?�j��W���1�pj7A�]�g������T�a����;���CQU��i��	c�ym`6%U�(fd��������r�k����;ܐ<<x�j$�2	�5��T	7�V@NF��Z��S�60���_~���OX%)��#o�c"Yn@{����G�D����꼜�&N�tx�	X��> k\�p�ȇD( d����ǳ6ǌI�_�NI~����0�m�O�E�J�H�u�Ev���F�Z� ��Go�;��FPKn5Xx\ToaF֊�C�7Z��� ��F$v���|h#@��4������z��{#��2:�"�}7T�2qv�IQy6�肔y7yRf�~���v��;�+z�&+|)��;��Q4�L��`s~v�8����/�,��)�f�;ɰ�fVW���u*�o�HaLN�R%6��o� ύ�+$��Ev�4�G�2�ҏ`�w�����%0�2<\�ջ[w>S���P��?NR�֯���	����9^���]��o�#u�;�����CR�DqΜ�t:t����Zq��I��\��@��;���X2��B^w"[�^�5-��O
J�%gx(%ݭ?9�-�z/_��º��J���@��		��6-�r4p�.ES��n���5S�y'.C�i&z�OL[-�ok
�;�^�I}56k����0|s8���a4�����,�A�K�y��c���|c��( /u�\��\�'�����BG���i�J��&zD��/pT�x�L�r�dcK�
�Nͣ�ά� L%	%�8(��i�F��j	Ǹ�"�fxMo�Uj۳�zIoD���V�ub��py�-��(��i�i������9"jm9h�I��7O�3BN��G���'6��:�j�1-;�t+���Z±�r� ����ߎ�+��$��v���Q���3^q�.��q�fmi�=*��\Ɵ�ʇ&��D�S�-%A�޷m�D��"�/OZ膢>n��t����˗�q�~�(���6��r"�뒅��1�<�C&�����!����W�DX��Q扯�gM���i�!"3��"��;L?
?L���ö�w��cJ.���
����(]�	͆�;zl���r'�卣��P���ydΜ�:*�ȳ���5��S��0�}��B�fP԰�%���MR���U�߳�9%$���.[�3^|t����6ϊ�?���+!���tO��տ���
c�w��	��d��k�S��N�B���8V��LnF��s�hy�᤮4�wt��ͬ�	�$�@z_~ӁX2��%=m�DW���������:��� ��/���X��~!�;F��ג�7���H�T#ҫ��#v	��ɵdʎ#��D;v�mXA1��>_�B�P�̖�z��������8���Tz8�_�)�ߓ-���B�	jR��Q�T�}��J;�Ԅ|4�ⰕH�Q���C��'��0Rj����C�j�HzZC�R-�
�U��_�+�m~N5���0�2�;�Tlx�7��QUtȭ�z��D��C5�i0]��s���s��\�!*M D�U�Ǉ����뫐��^�$ Jh8DT|�
!q<�$ϙ���6+���������A7<͋p�زڇpsٸqj�^��y,#�����h�轛�^��{-��&�2�~���6 �����4�$��R'��\N����k�1?̧��M眰��輿g���p�d.c^8\	D�x����QY�\y�.��x��.}Dk�t��*D�=�����	(66�F��ꎅ~��[�\@t�7IǴ�Z"Fy�m%��񍑃K=����jCW�Ts�4�J%ߪx�Eb��z/���ˎS{6P*�.�1�T80�{	R�w��k��	���$~� f��wEcr�[,er$]�-�i%���ܡ���$"?f́`�V�v��*�E#��ˬ�cGI�9x����K�}Yy�M7���k�}�([mF�\�:�F����=>%r _Ex��>�=�I��ZmW�%�n��Q��\��Aqy���S��W\�D�]��V}+��_V| �Q �iⲽae��3�U��30�}�+||F��
��[�K�;OS�I���e�E�1�!��qa�aF��?�V^`3����Ŝ3g�J'��F.��^�d��9\y	�,1���V_ݗ�J-�K�p���'`�V[�% �.�ޙŊ_��-V�m�vP��T��uA�6�q�M�C�û⟵��z���0��j>��Pa���?~�p-jC����vɦ0P��׼$���T����a�m?NA���ű,_vS/ʡ�p�}
'�U�B�H�2C]d\��46��(n����Fۘe3�bV��*7� d%B�)��Y��{�qY�	!�t��~���~Q�)�gZ~܇�#��uW�]l6Ul�_?
�ͱ�x����e�tՅ���s{c��n�)��+�N���.$��(�;i�����4�f!�@�F���,ԍF�ae|��ڶ{�_�Z�Y@z8t���MR�Hp���hN� !��s�N+���w��e�v74��*����6A֑�Y�Y��i�{�w�Ma"� ѣ	"�x	w����{�
8��0�
]&�  %M�[�e��!��C�'C��`u�y������>2l��8!����n���E� �M��D+�����gA�!Y�e����$����i�̊xy.8 �+b�������c9�;0���hvߩ�i�$8��R�B�����x�,�R�=%m��§E���6�Y$��=��Զ�JﰗJ�a�D���(@C���hL��
��Om����䕷b�6�2�Y���{��\�ʌ��o��¢�o~"���a����UP��tH{�j���X8U�V��`�Si��T�{�;* �J��O���/��=��� �w���o.��eO=!WI����"Jc�p.�P��5������qq�N���\���SV�'ѾU��m��=�+�?CT!�fm��	�!��G/�L,�.��G�zV���8#LW��.[R�DwnF`a�3��l-(X����C0�B��NW���`�5�ɍ\:
��Mb^@G8(�會�w�G�f��z���E��J&�bī����.�W�/p���B4+�����tDA��M�Ci��m.��A0�9��L��Gk #�R��O6�b���M��\�l�Ak���;�k-uEN	h*��S��(<_k,�̘m��$�9f�Ll?�)�~�h��n���颹��O�=W���|�ʎz1�#�Y����g�H;U����h
�O�z��o�טئg���1�?$vj�Ѳ�'T'���@$�Yap��<7�.
����,�z��-"6���/A������������Z�����w����?w��[|�6�;(\+f"9�y.�w�J�3��X�]X������+k���+ ��t&�Ё^s�w'��c�@��g-#���}���"�������W|�?��P��ħ I>zh@ճ���Zq��d#A��Z�܇�-���1�k�*B���c:WG���ҹ�=�����[5k�?!nV��m�8;6���	�wx��K��B)�Wz1����.�-f�������+АC�~�<}Z/�:IB���_�B�P%P�^;e�nЪ놖�jм	���F��Vq���u�Q��P�,@P�i�C
®�D���P�n�LIǌ�h6[���M3��gj�i�Ե�<7��|�z[�@F��[�! ��Ґ1��~a�*���>��Gku���l�<V�[E6��H��AnG���#��^��3g�'��H�C�X���LS�S��D4|�UP�.������
j�kE�1;%9e#We���۸,
�Ҕ���m���fg\�9.D-ܺ��N�ΈID����l(Bёn�|�25��?�P��[��)5��U�U�N�Ȩ�����I2��� �t[��LF��!P��2Ŵ��s�h��5Sښ��J�d��-"�T ɔ	U'��d�I<ʧϬb�Jf�ͻb��H��j�;��L����L�
���*�![����X�RZkf5�5ʗ%ۋ�"%Pbڡ��q�4|���?���T���:�p���W�3q��v�Q�+c	>���(��;��XV�����4h)�Rfe�i\�)�g�K�0�5̜��Wߔ,�+6I��-S��Pӊ{|sb1�ՆgvY�C|q���2��u�*ƹl�s�d�s���0d��<��n�ц	K���B��ޮ�&��
�4'�M'b��̢ܺ��<>"V�YE�y����D~�^�zֳ�w0�\H/U��E�7oS<5��_�t��'��o
W:��x�Ҋ�8���E��<[�������{��+%K<�-��]����v ����ğ����%�V���jI�'�����{�jd_c�1�RB]N�5߰
��V��6�?�n%�w6����.^����y�[�V�h����܆b/ֹ��k3�L����eNk�Fc*Z9/� Qb�YB�#�4�#9
Uͫ(c��=h�[��,\�<�\ׯ��_���}��ݙ�6�ЭQ��F��5e�ԝ2>(��N�%���4�b����I._S	
4�g�dQ��0/C�f֖eP"v�Hxȸ�U��ژL .����(�^�����*��n.AsE�<N����\k����u�:��*qH�������`�қ!�u�[*�� �gM$�1ھf�t�ː�x�s}��6��f�F��U��ߎ=���Pk��I^�^-uyn�J���2�f,1w�^�dȸH�y�;)��b%�bMk1lEm�	���(ҪB��)p��q�����=�n���Ŷꖟm�0�;:?���[^`�`�$��o}8�g��K�[�9	0G�?	>�~�=�+�xK&��3%$���3���i�Jɾ:��쮕��Կ��̷'��(�i�8�LT���������C�KB�(��K̀�e�f\�I%u��+n��hd3b�E転͐���eCh�m->���eỷ�.l����G7n��Y]�#ٍ�3��`�"����}���be%,�(�їr^�毡���Д��Ŏ���%�'Y�D��A�/���_>����OfK��8��0PS�zmN�h)ؓY/�E�����Z�Ω�8��55u̓<�~�YMX�^Ъ�ߍ�p�N�A��ɱ,爽�?�
����P�Z��G䃞�jQ��L�o
L��+�K�@QHJ��b�Û�^�:�hИ`��`�z���#C���=�u�x�a���!�������T���ڌ~8�q"�k��?�?n�I*=3wޗ��06�	
��'�54b�Lr��e1>ϋJB]?��'����4'~��o��:�n��b��Gg	P��[��t(�&�}���v%�
(����-	���@G�=6 }O����(_�#Dt�n�2��(�e������nJ�K �M;N�~�2c�{3�V�\vo{w�ʭ���i�n18���Ρ��t�0��A�����jB���c��a���2{a<ahƨ���	e��D���~ЧJH��������$6�<�����'����GU&@���5����
#ٔA�Las����g��1�tp����R����z����Ն숧��M3�����bA8��1<�9�9<�r\��0Mvܞ��u�p"���@���B�wYxR �b�|i58��.͹�dn�F���ov��%�7�v�1 �krO�3}�"�(��Slxaʬ�'$�w�dx��uO�]cW|܅<����i�-����
�(?�G�odvǇ�����k�Z"ܳ>dq���,��� ��f��4���N��e�/U�f������2��	�܁,L�Q}���e�٢�~c��΁ʀ}�}>�ǧρw�uM�ɐ=��X �6!�Fm�	��dRS�pN��*5�^<����i���d��l�I9�5{v���$(~��'�g�ݼ���妛�	-7�9��n�%B`��6(եc�ڴ
��E�S]�v�3�Oa\�I��݆d�_}�u��i�^�o>����/�ý�d��oUۢ���D���.�����&��� ɑ��x�<$�����)��u�7��e_b�
	�õ^i,\UK�f�r�@��kS'xq���䊃B���������K��iG�%�fф5*}�7���?�f�z$ 6-i����m��[E�/"�NH�~בl���܉��I.L�Q�:�=������C����~nF�ê�ˮ��{M��zuՁ�/�/CEus$wP����X����E1���f��Ea��#Ғ�4kUF�Z 8��l�%O��s\����kJԒ]��@޸��<�{����Oƹ���Q���z�Z+3��~#ӱL]�t�b`+E6����U�R��!��Ц+���㡬��,Ѽ���7=�����GĜ+M��: ��>O	�Uh���3J{��o��#���l߱Ѻ7��(�g�Ҙ�k݀.�*Q*Z�ʓ�*���7���6+
��ո:�)f�p��y��v� �I��|ߢ$�ؼi#N����̆�%4�ȉh2��`;x:0�H�6�L�|>��l�]�� r�'s�s[C�T��*�׈�K!�a������R�n��S�J0T.]�������.x�J�+�B�u��II�(mr���@U�7租ch�^�~�`��6�\e�g�9������{�"�%�u��~��
IN3;�O��tsy@��L50q���j�<0/ʟr�[R/2���GZ-S;!+�Y�̀���!L��{�e�����X]�.Q���[)7D6`܈����������at�?���t�E�58ıp�cs�0�Df�_ꬢ�����:���
v�I�"F}�; �x�s]�=��h$��`p\\Bh��q���#U.�O`rl��U��	(V٦��k��8�Ma�uzc�i�H��o1�?�����iZ��$w���������'�t�4��(�&�j��?g߇r�p�r4W�;��6WzӬa�&Awq�� �>�B��6�����#m�N�jH1S����B%�`��8lk��4�rX5R�#y��T��T����e*�YWWX�Ct�x��J��l����+����w�����^�8{���u�'�D@E(K?�S�����Ƨv�ϻ+���0�De��)�Х5���.�֔�U�Q=R�u���)��L,o�lY>4n�z=����6B�4���x��9�j�,���`XސȚ�F�����ԓ?n���l�@���L���0�.8� B!M�j3h=mP��O�X'��d�S��?dlMk^ck�صz�����BIe�qχ�\�Q�-A��������X$T��S��?��iu@�;�ɜ�G.=�:R��'�?��Z�����3�OK�>y0"��8��8nԣ)N_��Xz�6�@���(D��o����k$�J!"f(/��h�lҋ^nN.#��V|���L���"�2�#/����O:���~�u�dXJ��/K�ꣵ!z?W��
妅��5�a��ć���i��!o��3p%Y�8�����/�g)�q[�F��|�l��ý�D;�6��g2؎�oS���4��Ḿ��J��%>�;�cm�|��	�I}�ԅ��\UXW)bk�]��fჶ]�J/e���@��b3	^��îd����hk����;�b�}�G�o+����C���^��s5"�7*�&Ϟ�C�p���p�i�5���$���A�l��vkw+8�����L7��{��ɣ�6m����h/�<�a���!�������y����k�h(��#�d�/9�F�:�Wny�	�t��	*�1��sn�)aQ��rR��n˕�,���&�N����Rj#�g"�d���j���Pa_C�aT;��0�e�b�Q� ���lW�������jB�2@�H\i�䝒�U�F�J�)�ჴ��ϒ�-�j��\�݃�+1�\�h=��n�Qذ�xK�f�g5mx !铈�Є`Q5@Q&S���!��M��:5���I���8�0�ww�+ro�dEmzW�G#E��Y4��MQ��K����AiQ:8�ƥW�O �m���嵰-��5�79�aY �j�L(n��e6�����T`��a�2k+�J?3�Tj�11l=JZd��▞B\CQ��S���g𢍩e>�r.�"�H.^�v�L&6f� �>�֧D(�i����(/]ˠ-�wx�z���υ�5o#��Q+Y�1�e2R���wU�S�>�����B�1� ��s�(�l�7�IO!A{�@�G���f�3���@���+��̲(łJ_��Q�j�\a�� q���3�6
�C�J4n�4)����=�E�`i����	�lm03�ǖV�˿<�咽�$�:��S�7.>d�E5YǦFB��Mga ܝK
�e6��Tjhe���t�:��8��K~]C���U�(��ٵ���`º�ܫ�и�	X0��A���i����D��R
x��y�QA�Y�N���~�V�����d��/��<�z-|�WtmA�Z�R��
cBɀHy��7�������4��fwj�/Á� �5��ȌJ��
�Kq��"�}�����.�Zb&.C���u��"I�k�9��h��;���σ��T}B�O⶚�%=f+�T��䦳q��n��䷨�ʚ�����aG�D<�̳�an~����m��v5�s��@?R8i?u��M��h�� Y������]ګ��Ls�iͽ�TH��@�!�y�S��&}iz�}i��\�8+&7��|��X?D�*[ֶ��[Ǣ���Z��/?&!��1��n�F�켝�Sz�6:�x�OMr���k�^��}?���?s�ղ:�@�|�s��b�d�h���M$��kq��߁��n'(r�(���wQ�8'f�ȳ0}D�FU��28�4���H<�k�O��6�NHAɭ�,�k�P`����0�;c��/�ݎW���,��(`h Π�S\Խq7~�I�I�����%9~��U($-]�������6��eؙnj�xl��a�w�ι/1�%��d��������$���0|Kہ�#솶�;Om�914we���'�9�~ƾf���?���' �qU~��63z�&LOP1����#A�v��D�?�EkX�b��vf%���u+5o(h�:��IC���Z��DԸ��K��<�����T�pa������,��Gl b��j�����.wI�&%*���\�d 0�W�%��Y�'�D�5íX��a�P��\�Qúʹ�]1e;뾪'��\��3��|��
��ψ�#�'�F������a��6�!D<��2U�R���̃�ͧmE!Xo1�[��t~��w�}7��� ��Ȅϻ�ov��Fw�U8P�����N����3�Hl��/�pe(���Q̣�jX#JJ���t�|[�wLbAD-���sY�̹�PS��wTb��c���4	��1\I⃏����m@�T8�-{�[Q�#��-�y����T��p\�{)�V��g�9
x(3@b���iB�cѡ�DK���k��M�{����֭
�8(u��f�޼?JH|&SF����@��W�� ��,'�<����,ۍ��^c�JG�2��)r@������è�T���]Gd���b��y�m��k�����p�M��VK� �8k�(Q�Z�ލ���am;�qZ���O�ϟ7�$����1_��f �.���?���/��.�TX�4(LV�]��i��<��b�S�Z�x��Km҅N���)����g.,�t+��SV�t.ݯ��;�N%��n��~�����G6���D�������� S(���P�h�1�"]8r"9�ЎO�)�@Co���\���>�}L��Z!�F��������z~WΣԽ�������dZ�t��N�E�3��3�,�o\�{�d�8�x�'i��������.�L0o.@k�ߗeH���(J��\U�3�ag=͟/p��!<�ґ�3K _�c~�x[�k��J�:���P��bPLO:|E ���`އ[M<��J��Bj�����u�4_��3�-+��u�G2���o��X����޽gG֊��J�n��^���/`#-��駗ec���=�����"9�l�q�o�T"h�`��AOs�T���1�bݮ��T/�4�L�����t����W��3C��s�Y��M4SV�DLe�I����P���
��E$}	��@$-���9�?�21[C�Pb �����!ɻ�KW?�9��fٺ�����yC���9�̒||E�xOY8�]���Ѥ��J+�crT�(BIQ�k�����ԋ�M�������1�����M�K�@�����!Yi�4��dJV7d�sQ�4�8����QHB�i�6?oBB.2ѷ,���־G�#�t��`Ã�3�o�u�R-�i��[��drN��ƻ�E,��g��(�nr�:]>'�b��A�>�%\q֣e�e�0_pu��@s@������y�hɚyiƐ�#[�1�?��� �ϙQ�w�( �,���a~$��wgr���,P$�O��|U��9����F�X6�7@7,a�X/�7DuqLx	�n�X��ܺ�� *o!˼~�{o"g���!�O��q>���,�	� R[���>��\��S���R�&~"��]�fk�D��]���Ñ�;���%��7��i�_�@`O����Z�ܐ`3�v�Ye�,���Ԑ �O4�97K`y�G0xP�]�r.�����=��Y��bs�Q���1&DqLKW,hC�&�y��8P�<�v���s<ek��0���z��yo�����2`��Iˤ�j��c�(aҗɹ�
�`�2V�~�M�J�3�c���o��J�����A��V��-��[���a�/D��$��V����`f��R"��Ae�-" T!}�3�&�S�ߺ#n��4X��[�Հ��=q��w2���|Pl7>�c��"�y�S�n]�j�3Jj�y��C��h7^|@_��(ٲ=0,*Uxo��Ԣ��Kh�<�|1H�4�9=B����a��+�D���oѿ�ҡUEA����bY�^� �*R�~�­�CV3�vҿ�aH�Ӎ�wkoH�-Vq����1pA��f��5���������"
u7pl!v+� ����fr!�̓�*yC���u�9;�j���΢`�:��E ;�o��[���`�iנ�q.n
���oe����Կ_��Ѕ�
	�����`�y#r�%����/Q�F��R�>N���R��M:��_���]'5a�
GI�.��
�r�YoB����nz3K ^��������� <�TD&��p��S`mqD\Ș�o|�l.-WoŐ�e��c|Mo1v+���[�Y��ޏ$,�ĩ�X'� �<��'�W��j�T�$�<�qA8s8~{U�:�XrO�mٮ���S���A��=-��\{<���-j'u�g.o��[�dTX��h���nf"���P��\�}�u)ee�J/�qĨ:���+ϱ=r�ɓI�CLy�}���}�#��E� u�N�4DE�[�T�e��Ɋ���x��V�]3�`ZxԀm���Şa�<�o2�kS����*�'��W.x}m+mR����Ԥ�Ud�_?=�P^�-�xo���n��x���]�1��	�6�,`â��+�$��:�������ƌ�&WR�$�]��f���B� �t�����j,�C?��G{��5�¨������e>cb@�4��:��0���=��c�@A[%��B�5�L�9�2���tz����`ҏ�1$�_Yu0<�|Ұv����v,F���;ЇR1��JƣQ����2��W�)�&Η�:`�'������0常������Ē�5'L���)����7�BQ9$@�!O*9!��	W\2�/&���.2�F�B���)�F5��\4�I`/a�u�r��c�YBYw�Yhi&8<�8�w����8����E�*�!7[Wf�Xt�/s�Y-�ޥ\���y:�@���"
�r�/��!��\4�C"J��ٻ�ܙizI���=��?����r0���kN:bv���T�J,��Iq4ҁ�'>���\����r��Дw���堹��$Ӻ1��j��`,�h9]HV����Ӹa7)Ǖ�Xf�0��o>�2r�w����q;|��@iMD��HJ�ٙg����M���%'x�~�C��ˠ���z/կ�(�M~X2�z���4� ��K2�:%O=�<
�x��� ��`��Ph�JO�M#d(>
 ����Kk�u���ֳ~D�����է%�V`�k�C�k�*'Ʒ��R��V�\���_�b�/*��pۇT����m��	��d��қ����1M�29|��[W����W��a+Η[�r��4-5h͢ac��C�}5	̄��u�ؽf��lz�)N-��e��aX�õt���r}�H�˪�9P��$\�J8��q�&d-_veC�ǲmL3}Jۍ���G��u��fg+��G4���TX"M��z4��!�G<ES�`�7Lb��c�l�f�D�~ڍ�{���:����ғ�"?�����݋$&�H<�[�x�K�o�&fV�ܪ=T.���C�
8�;س%��k��
x��R����@��QH�Ǳ����6��|$Ғ� 辇��<φr���%�Y�5���X���qtۉvs}*�~�afB�%B0ږ��8_�̿�R��"�]T�{=����l)I�b:��^�g������N�2���xSG�4�?������K�/���C�@�/ԉ=r�D.&3���_��< ��7�v��BM�#����V!N�����2�*E�y���4�Eٷ��\����a[0��&��S�e��MZO�k ��p�ɴ�%̃���qa@&]���E\�S�pYJ�e����d��m����Az⳵��.F^r��PI�j�+$.�nn�79��6�9��K��<v�t�Xc���{W��S�u�b"�6���g��$��*�	fd�4&�O+�v7d��͔߮�n���0{�1 �{��#�}o<~C@��^���"�1e8�h�w�K]�W��+#lB����7rIL\�ڟ�J�D��5[��F�{��jw��tq_�4��A0X�}{��UH�WF�`VlK��7`�6[��j��5Dn�7n�f��<�����TÿnpP��ބ@�2�YQ�G&+�
*4_�sF�$���<�/B���,
�>}ۏ���<�41!�}"h�2�8�E���Ub�"N�6���A6#κi� ��ꡡp�v���~�Nٴ£@��&'�`k�k�H�R8񿁀��13>F#���N��`r0�u������jx��-�������f�D,h5�6w�QJƛ"�IH���'���4�����ʢ��� }	Q�s�<�E��f�a�M �EִF�	%�z�b[@�Լ$�{����W�&��H�.���{ɯ	~�Kŏ����������eK�ٛ�?]�&m(�"JU���&�`�*9�u�0�n��u�5H��PDA麡�t�F�Λ%�Z�&E�*��N�H�aG�B[>m{o�7q�^�\�|���+i�Q6w���h�7�=�"f�ϙ��,���_�D�C�ʃ�D�7�WAǫ�,�����IH2pۏ�tN�ŷP��Z�~�vr��_�Ro��P��G�L���`�i�X����l�:F��J����D��`"�OX��.���)��s6�-��nZ�ű�D��b�25�T�� M�zR x�H�[}�}eB���o�ܸm����l�rA��4a� �됒Nvl��%��_.�BZ�_�g��[��Y���c��<#'�"q]�*�2#e��/��B	qh�k,E\J��*ri�&r<\|��$��g�E����$�bixsPŖ��h5��]�4h;.�L�(T����:���+0�h�iW�ޒ�U��-��s5��{F�c��:���r`��	�?G�������ד��y��޾�k.L�z�����2�X���䨬��C���5ҾKQ�̯flu�ǂ�%FIo"t�gx��tО�z䢜=�nE�n�]fiEܭ'�:��_cMdH�ɼ���4|��C<	{��#I~��}#_ŖAlm��8�*��HZ�ynq�؍C`g�˾��6��')7�)��H[|a�X��Lzq*��=1`�s!)�M1AE�U �x��b��&�9|jdd�3Jܡ��N�ja�`ƴ���S�ϋ���T$��>�Y�կĊ�`h���.|/�^pp�Z]��o�'�a�-Ǣ��JQ%a��9?����'!�~a�`��h��O֌:U����-S�F�7��bU� hP��Oxg=�޽���2sn�Oծ�]3�ت�LS`Y������㝪�h���<_]�����cͶ3A�?<�G��Z]�/^�Ά���v�����4�C�`�f�7�����>��b�S�\�!�+�%i�m�=Z���,F'�<���.דV��B�<X�/� O���9,�p���>����y��:)��+vX��DH��	k1���}��iRF1�g�ЕW�[�l����L����i3�U����gx���K5ďҵ��Ġ\rq6Vה�Q�[!gfp�IC�U�GȺ��j�s��˨�b�&+K�7Y�K9�(��%��31���E��uZ��<䶍����6{K�-I��e��cL�<bpN5��;�x��
��xX����0B'.�Zӝ�\��D�{{���2��mD]ʌg�� �箃�
��; 2�1���`]����}�aQ`�#[R�5$��綷��b݊�eQ[i� d��d��c4�!A�+������C�ZNm��H;�7�J�m�U1�K�!}�54[xD<���e�S3�:D��cBH��yK%e8�7q���\�v����F�b����S ��OK8�P��F��N�O^���ǳ�eeD�'�d(�D��R�Q���UU���=�����YRN��cN%�{p��~I��T�?��)��I�]�K�#ɦA����i2+���F�`/�W�(���5q�J��Z�;iĶ��k7m�O��-�}��]�$^o�����ܗ+Ѷ�����T�z�,Q_;<��^䧸��p.?�CU���s��|�Ǽ@?P��Ա�(:���?��9�bKk�G�.c� nf��#�Kqo�[�M�I�o�n�'@���Z�ǫ�N4���	:�J�s~�2�=V� t�$��W��w8�+۶��Z��BS�+��M��/n8�AQHG��M=�s";�m@����b��/j翮Lh�[�jf-ť��M+�i;c�WGc}���9����x�k�ܸ�EWSɡ�Ʊn���m�rZ�Yd�;_����bVD��R�J��H@SmQ�Z��%�B2k�����6J�)���K��H$-偘�7y��5�[F���0}6:����߻$a�P�g�2n�u�� ���\����=����K�	[��Qu7��X.[���<��r�f�TH@	M�p#m&r�L��hEd&; lH%�J^��y��b�Z�p�t<�R�S�hȐ�-��F[wQs��x��i���!V9F��[Z|ǒa��x�6�d���)̕��9��ҷ�0by�Nݬe*�tZo�g1=�[�4�g�ܫd��Q����O�m�ez֎�x�O��7��ѫ2��:|��Q�~�qsI�����V��G�'�MK�<�Y�5'�.��=���ve���= Ү���ޘ�ǅES2M����(��:�O�PD��ꡍ��W_R��iU���ېت�q7U*��\�7�3��k��/�����N<��l1f���E�Y#ɋ6bn�!J=/!R[�?*t�_hI������F^.;u�A+c"Ө�fh��H�a����[`��-�{E yi'�?��-\�S�O�+>�S
)cw��o���Ws�[��ڕX/�p�%���{�=/���O�8Z!�-$�Ow�[�=��ͻMo��g'=�p`1�.|����I-�/c�j;�٤}�Lkc6����ޛD��G1r�ATǔpr�i�ت���l���i�W@��/��5�Y��b;����)������K>'���<rI!#�J�şe�:T#{N��Edz��t���(���É��Y�;D��G�m���bƁTw�R�I��8"x���`{�[��`P�5�&�lȼ�; B�;��/�ޅJV�:�ڌ0�w�w<H���s5�z���b�052\����ql-��Z%���A���-�����h�����X�KJ�u��Ά���<��P1_U��$e��JJS�06��NG�����{�Q*���OZ���0d������f�}��N��۔�	�v	f�<�qJ49g<���+���'��Y)�#�
�&��H~��b%i�r;g�i2ã�����V;�r
��9EZ;6��|���H(���x�	`�1����>J��2lst��d�8]2��QЏ�@φ́E���e�!WM(aPv=�DcUbJ�\���B�v@yO\ݫ`]*�n��9%� �_��P��D� ��R���_AM�}�-�&�aKK��o���2L��w�IM�0\G��#�ma��m��R�Zg3����Bx	 ((�x�e�ڰ02�3wt�I#	��Y7�`���ھL8��������lO�%�d��h���
��9���V$ѧŀq�hf:�;!�'�r��SR6h�^�0O����VD.2���|�3+@>����H��|�G�������{����p�F��r�=�b�*p���*�ɘj�Gx�(0�����>��1�&��6�B�]�����?�u��>d�z� \�r�ɼ6�}+�$���ԫ�2K�˦����w�k�m�B�%���T��]{|�~�b	��25w=���K������.�-�wZ-%���z���ma�}yw����2E��\�>8}*-�t�Ё�qu*�d=<fq��?��O��sP���ߖ(Q0�x=x�����K��D�����-9��`�;8��˰=>�R8�{2��_\�<9����N�
&w��=`aa�ꔐ�����hmQtn�8Fm͝ t������֏m�]��e[[e �r��$\Hh�7V,81�uēae�����)9���dM�L��v�E�2eI�E<y��6��Z��� V�C=}7j	����]�b�&ca���`{�'����A�I���(��������c!Y�Ҿ�ڈ{	O]�h>,ptF��y�cAVk��F�+	��<I\���	_�Y�3Zķ3~��z]��'8��Ԭ(���e�h����#�r}�@�k���_��dnL_�8�tQE[X}���zGOn�� x]৷��a��V�;[U�'�^�����ނHA�<R�>�2�~���,������j�r{�E�L��$�,{�V��1��\?�����硗��R��AL'���_N%�W�-�d��V���p.d�ٸ�
wM���}�D|�|��1r�IxTW'�E��&B�8���䱤V�p�}}	f.�J&��n�O�B�3;��;8�&F&'�/\0}֋j\��m�0x�&1�f!2��G���]o6��� �6\B�rr��^/@�es��|	Qo�B[TFTAV������,����!�`���$1pur���΢���*x���U&ʔu�8㯱����!�<��]� �۪C����$�pu�k}�Wc��֝a��Ť1�E�in��u0c Lr��������a�e�p�b��n���0��P[����R�p��
k��0�X�\^��r�ի҈��b*Һ��[�'
U�KYn>��4ͥ�,����]:('5��ct�2� ��h|��7b{&$Mf���'����3�W����W�Qȭc�)���鵁�@�C���$v��$��*�����8on�WP�b��pn&��}.ٷ�; �w����9	�0]����,���̋��p_]�	X`ܴ�Mh�Ԯt����B� �!A�'��y$�|�v�0�cm^d�~��	�;��!N�M�9���S�,�=��%�+ƔZ<)�	��B[�^��V<A�-�`5#�3��s ���Dw�Ӹ�b^�Y>ޡ�J�O�(�
��6��'�3��u�0�
%qQzF̔�q���z=��T}5���u�P������M<�F 	$S�A`��	���p�fq!~���*h�3�$��s4j�v+T���TQ�:@P��~t����c�`�����-�M�K. �:�a�Cp*k�
� H����F�)�W��E���)�7zJ��&���������^���ɜ��@��ʭ��6��9���J�i��.P G_ Y����疋�hH���r"�Ї�씛ʿ6����~�t���Z��H��|��d�z-.XH�-��DƋ�:�{I���xV!�$��o�͋��>0�D]y����&�]��>��ٜi�K���%vL�P��z���?j��,��Sc�w���|3ҷBش0e볞�1���h��9�+?*ξW)�0;Kk {l�x��t���S���ZH�@n����@C����\B���q�=�$߿@�y^Q����^Sx)��ɤO)q�i3O���j�VT_iC7�^	:I��������\J�L�8�ONĎ�Gd�b�5ۼ�q�^w^��&���b�w�ו�M���\�uS`�dA��B��Ě�׽j��y@�n����.=�e��#*�W֦vcF�
�(�<�AM��jk[��Y~X��
L���,���0�&y��
����>��ع��;�}����}W�
��J{� �΅kt�1�/����&`t��:CL�J,��Qn�Qi�H���)$h��{�~Pjq��Ƞ���^�~�cxc�TY���,�R����Ϣd?S�> ����2�9�#@^����k��g��a��J�P��`2Ƅw�}�[��q�
a����Z5͆'l%��"�-i��Y�Av)�OI��3 ��ȹyP#�鮠�����֟��Z"Q&S1�F�RmFT�e%!� Cd�� {~O%�|�e���a���Ѻ:�Z�U:�����9 �^��2�����T�-�����-C���U$�O���\�y�1�~�G�Z�ƥRt̽�L�F��&�P�8�1�[<q��"�hb�7'��Θ�<�#c�a��ޱN����<�-� 2g:M�m#j~�`�(Z�=�I�I^������U�d���^u��}��[&vwG�huƩ���ݳ���?Q�T�tC��̅�z|�kSM��E�u�ȃz'T%я�����ˡ�?�@bs��69�8��2���S&f��r��9L���C�P��,-���*0b��3l_YP��RMʷ
ۃ>�X%j�c�XU@#/~��"�J��� �~�:Y�E�`��/ݕ��o��i�����L��"4�����*6�Hpyy䩴^�`8�<}mN�&�O{�z��{w����
��s*�@�"S=�˖r.�f��@Hcd��(��1��_hg�����H�3|w��¶���ѯT�2()�g�g��,�*&�Vbe���/Lv���M�=-�~�2�=�%�!�N8ov�r|�2���	l�}��Hĝ�HF��6�F�I���yX3Ŝ1���n9`��*��i��E=�0�����"Kɚ"�X�az��O(g���k�A���,2��{�ۋ���P �4������e�����2��C�}��
�>
��B�1e�ʐ�0��qڞ�?e�[��z�tl(�׿�ҽ OpV���SyR�&�R/"ȯA�$&���e�7�0��#�\�}629�}��F�?ť݌�u���Ji
3�_8:���b<IEM�:`�