��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1h,�mwG�� ��q�
dh������n�5ӫ�2
�e?4�K�����ps�/)k޼��������a?SrL-j7%�"�1�z忄Q���͗��2��B; �/^R[����wd��\���
A3W���w2�;�uhs�SE�%�i�6H� �P�6��v挻g��Z2
�*UO?���d0�0B5(5��������\�s8�9���T�����%Ƙw�}щ�$g5<�Ә�V�����6)q�ą�!	�Bگ��`Wń�zo�ǓL���u��%�o<ҝ���;Ss�W5Ro����@�W����S=��6�)�L]iM��)'w���L\�$�1����dvS��p���+}��Dx�A���v)����ⱁ�2խ�1j��A��*<��$8�����p#iw'^bY�z�-�a���&hW��}?�0���A�f�
	�w���Ѧ�2}熷AG��� ��i�(3e����݊�O/������<�V�V�ċ���Wћ%j�`�'Ӎ^u��i�*���� �����Y�2Hqk�0#��L�˞�qj�x��ab\|�q5�������Q}���O��>F�!o�X2Bʼ���W��Ҥ�f��3��r��4���L�i����<��̵B��A�#����c'ش���9LHk�S�3��";���w2�Fb#s���;����|2�%�W��)���i�57|pS���&G"օ��yt�ͭZ�
9�K�����\~PEn���@�%1���jĽծ�6����6�;d?��q] �Ǚ��o�>���������1����4��u‒V`�֫���mrv]�F䵜T�~n�@���ɲ+z�5lg���	WɣkU�DDi9$>�g٪)���0��0,�-;_�m��~�؊o�
8j�?|��@�+K���Q�FC;
8�]ͳooM��J�q�V��h�p��o�7�O��w?�ٽ> k��!�}4�l�������F�)b��Iak��5�+u�.�!�1d`8���y<۽���_�[���D��m� kiV���#¼��_V,	��a$y� \���Y�X2�����n����ϐ��\�*�f����A���4�ӓo���n���N���#��2M�f����� ���v�����إ�p��6��f\&��i��v�,Az-�\PzBq�b�\�"+ȃf����!�ƑY#�2=E��eݤX������]��`���jh{�3�bw��\���U�o�YFW�Ab0����葤.+ӇG	,bbq,Z#��EX�V�'F��;G��HphI�Ĭ����[���H�be��; j�; :�V�'�O]1h}���hh��}�ۃ�m<��J������["E����q���g0Ǥ�BWS��!N�����#K�Ҵ��2%r'�۵{�<���1m	�^
�ߑz�sH�=��O��^D!���}������n��g�Bs�����n��N��Ĺ�݁�i�3�{���U���Խ����3����l\k�a�,>~��g���8�qz�AJw^~\/|�Ϡ��&��ea��h̃-�G��F}�F�0ꣲ��4W2�Ö{\��vX��͇�kԮ?��Y��Z�����(�_	�i4��l��h=Ī06��F=͠/�,CT��[,���3㏪���?��3uh��ͧ�q>x)A�2<�!�o�OU�5�
�Ә`Z�qê��N�^�8�w��K�U�t� �/��z�Դ)E0���-���>L$OJ���	F��NOF��L��u�/�Jр2�k�V���h"���{�^��13i��b<G��^UOլ Nw�#��5��]���N %��h��`x����<�!���1�)|A�Ui~��@r��G*��_�g��Pd�U57P=����Ǯ�甾�p=Z@��%lP�K�ag�~/����՟0
�ܗ�.�6.UK��}�D�I�*�?�t��ddJo�vB��)(��RwyצN�������4U1������'��NŠmu�z(��0���&�1�(��;o-��&�4�����0������ ԓ#�yr�r+z0ߡ�&�E�#1�;��ۢ_cu��Ǥh��Z�W.o�77�]jC�� �X
n ǖ���p򧖒և�^Nw��ov��,q}|=�d�d�<鵓��&�!:�*Oo?IK�:h�ϑ:�.� ��[�5qވ�r������u#zG��G|˖�*�Đ`:t�>B5}�D$X6_sEYU+-xOT�r��S{�<���a߂KӚ!+���*(.��LE򬬧��)�������ei�S[n�,x۲����'����w��\�7�)�/d�ia�ȼ���Z�Y%U���U�Ҁ%���0�����{eq_�o��e;�\���ɦ�KC-��V3pQ�+%Mb"�ݾz�����S�ǉ7�r,����|� b��>X6ꝷ�h�*��#������R��]WHQ�0�ңQT�h�R0�����Z�z�s4)����.�_��E��Baf�W�$<��9��b|\�/�xxo8��:���i|�y{��+�ߑ��t�p��d-�*��c+X�00�Y�����IZ�y�I�6ǌ ��%SץIƤ<)�p`I�ᖆI~(b�`�bE��n�u�9Q�[�[sB��0P��Q�Mz���:�CfY���[D��-��������aU�m���?0���^zL.,����J�"�!�*��k�LdD���+��G�]p�W�$W�A��� ��_}����DY�9���(��?��L�`������ow�#�GӞ.-�y	9P$-V���4*����7��O�B�Y�CZ?����;;��L�����~�ψ��s�5��H���o
��J��o���3���U:h��������VS1:������eX�'���qDp������`ߍ��*��$>��L?���_)c0,(�����6�ө�H�zb���������Z�JgDR�:�(R�u9p�C�>��"ټg�Ę�]�EpvH��Sǹ�t�ײ��s���ư}�ly�	T��F�ύ���S�A'k=�˧1��Pj>q��]�C�T]�o�4����'���=�b��G<�<��|o��L'(
0�r�����(�8���9� ]sr���vso�ys�I	:q�>�:�`�4os��̱>���2��X�+�`\�[jy�1���k��V����GZ�e�í?b�U��E����=�!�H��!�"T�J���қ$!�0�U�E�Üf�ȓ�S��f��kө���6�@v��*���㼧}�)�W�����=ӎn}U-^�}��J7���T�yh{q�v��u=��+'�PA��Sn���tM �N��>�f'K
+.���#�{�C*��I��^Қc�����Δr����By����9�Q�"i�`��r�v�"�O�Cٽn>k&zs"�y�ܥ} �tM�9�!>A��?��ތR
 \�:?f#����x��(ѧ��~
�Td���C-+g�E�7�98����B����d�ub��_��_,�R�\"k+_�g\U�D�\� �6�̩x��U=sN:��_o�"��<�� �c�+l�C�졢,����7:��ug�Nm׈�G�'J��6,��N�(n�z"��Z`�}#��pB%�@�f٘
�\��?��VU�o�W���hY��*�EB�I2Q����h�{�w˾�ލ�ѳ�(�0�E��@,����P!~ VR$x��%�`�ÔՔ�.h=S�`����j �^��F�a�Y|'-7��K��Yէ*���GT�_�!���LSQ̹fy>�gϐ"-��Ş���w�fq�^�
 ���J�����P���Xk���A��啚���<[1��� p��$\k����ƌ��pG~���,��DSu����X�{fT����P{�gm�\�I��=�0'�8�0�bDm�į�abl�t�� �8ys�/�����[��fLv�e=�鑼59T5t5��me	����r���1р��9��}�O,��7��Q:���=ݖ!���j��mLGX/�F�`���-�M�pwү#rNfķ:i�v��\�Xe��	��q;f�/�[�zv�{��=BX���֓�����s��L�)�h;T�dPf�\�9��~!���B�M���U��Ĕ�cB3�E6�΀9mrw��mqӤ)�NJ��tlx��u��|,؞�`��PU���\��H�!�GK��`����mA���nv�ЩK��խ�ǈ.�gD� �T�ȩ?�~L±v�캴%���mO<�?�hY��^�&�L@�����*ٯ!Qb�T�n��)h;𑽛_�z��~�"�\S��º$&�	E
��˱cn��W�L�����0�yx*�E\f�� �F��W���¶�3�=P��a�5���`��0@�A!n/��1�;��0
�(�I��aq�&�O������6Iˢ=fF�}����?�76�68 ��P)�l|�F�ĥ�J��b1�l��l�8c#��U9���+Z�@$l���r�]��.�ګ�y�݀��Q[�^��!- \a�Kϐ�yp�����_��l�c3�~�����ί�jN��J1�����؆@̍V� �f�@j�Ѣn���<�F϶ҳ�Jri^��Y���?P���m�A����)�L���ģ�^W��i����rz��q8p��,uDLy�D�����8~��UE����/d�"2'F��Ս�Ot�3^Bm�Y�N����c���L�(���z>��<d#4�!5 �h,��P@Ȍ��v�U�uN�N�6����`�y�����4�Pv�~ԯ�\BD��D��Q�����*��봝kB���+�`�U��Vi%�����wM귏8e���y���������G�B=���� �����s��
3$G*?����jÊ�l36W�/�īۿ�z��/3��s�=B$��\�D��Z[j������ֈ�1�`�X�ȧn�'CM���(i�%*Yd���g.T�-s6*"�&1�_$��e�`ܰo<_5�!�R�����k~��~��!�cXT�p嬭p�
X7k�.hf.�����Uӻ��Z�mHI%,oO~zf#JC�!�b$	̻�p���|�1fi���ٸ�)]'/�kbea�������Ğ�04;�J�@�=W���V[uyJB;I�6��A�	��=���4色YN=���W���߫v�+.�V��-[	�ZR�<��@B��"s���4���BQ	�z(-�\jYiVX��!��Ӱ���+��>�Wvy(@�Ϳ8������z�t�3���@�^�,�e����RvM��a����a�)�#�߆�l2�VY�1Ͻ��x�����P�A�����eB�q�����f��t�*�Zu��L� �]���:�ms�m��p�"�E�M���g��`���R������D��\�xf��C�6��q�5��v�"W
E+�;kZ�ڟ�;���v�F{�����Ĕ�bQ��<FQ8��)�c\U}�Y
s25�\w�ffBe�1&��H��7��x�z���-%ҧ�ϔ��M=�
����h
�<��Ö��[�z��݊\��(�`nMY�[�IY����o����I4rq�Cg=$5hǇ1�&��M�(�ҝ���L��yq:�t 
�*�k��W'���
�gX��5U$a��������[�T�h���mZ��$�:�Y��.��FF��N��N?��`T���c����e��!�wR& )k��"���"�y�7�^.7	O�Ƈ��f����E��6��@�;�N��|�t�|E�	�+ZH?F%^��/�܏�d�ጠ&Y���C9.�%ZNG��U��R�e��I��me?�x~]�u��7�[���Q������nZ�-_s: E͠%ƿ�c�6�3��ЕPdS������fy?:�����`'��%�'��-~m#�p~�ԉ���cS7��:�T`�(�tZ��H��F���'��� ����qu��z؟�x@�,1Ԁ9�^���7]/���ä���L��a�s��5˰Y���1m��c�f����/�޸����J,���ȓ�T,-8z7��Y�F���{�8��T��t��.9�ke�ꃨ������!h&~�5R���Oա�K ��P�JL���˼/+W]�	��2
C���i,���Gf:�B̾{�?�f�+b �_QIE�R���i����~Ε�Z:	yɮ��-�҃>x�=�}��¢C�ġn�f�ش���'�1O_qU�Ƞ�$�<���=}�2�^JEl��l	��N'ޮ�B��nsu�I��d�U��{I1����9� �z�Vw=J���(߃�m�Y��?qQ�8��	�#zf)}x0s���^��j�`�0`YAxJ��܄9*Π�![L��Rم7W�NP��0�N���0�K�?�4O�Υ�7�qO�����4<�t�Q\_ N�EJ����PND��X^�Rtk�)�ŧ�+6+.;*�k>j�ű��&p�T���3#�o�nk�	�osd7Y�m�i�J�z��!Μ��oD��'M��Ұ;2q'@�6|�N�&{Y�n��ۡ ��玁)��	谑���� �>��?]l���� �R𜟲���M-s�F��,����ӱ��o[�}n�"Sn��β��q�P��}`B��ɣΊ�K9ܠZv��s ���3��(��Lb�]=$�@H�E��%XR�J�������X^qa���<!��KȚ��Ol���Y��Ź�{q�0�cA
�lV>���2�[u}X�θ"���c��`7\��_���=��L#�0��4�T�D��4�&��p��]i���0�r��9`�R�i寛�������s��"��K��I��ኵO�	=��<����3C8�\��q�����ov׌i�� i��-q���V[��R��$
Nj>{�0 ϥ��|�*�1��Pt���ٷ<���>��l{��AD$|�  9*:̆!�iE�7���To~�QGz���%�5�U�*�b�_l�������E�h:�>��=�*gl����z��a�e"�l	�����JlPVG�,bq�ի���Ow�L�OKV��Qt���Ե|�{x��k|f�L�qf�@�v	�������j���:3m�
�o �; ,�-�6W��(���� ������T�E���Bl[��/����m�(%%�dy� �q�6��9��k"�߾Z�Eޝ���C-ؖv}�a���*ų?��s�
��2�=P��n���@�\��EK�U��0�'�舡�us�,�pW
�o�QA0�e(HB龹��?����7����s�c�?s�.VԆ��f�8��eG�U4v����F��&͘_�-Vw.����Uy��}�D����+�~�ێ�.��=,�~�聇���,��l]F����bn�Ɏ`o7��~�%�^�"�vǁ��u@�D �]��MԆ8�WG�n��B�Wr���J�-I ���u���B�(�%�J�7	<�8�ha�:l�������'Idk4�~���8��݌��4Rv���Tɲ��Ώ0~����i��V�$�m7��_���Ed2���a1����"  FKps	2-i��3���Iц�䎐�)G����S���e�[/M�K������n�dӌƎ���ݕ�/��Auc9�DU';ׯj��u�m1&���끃��1s��}�O����;����X!F��˘rX�<ͭ?>��\�<��fT��l��҉J�22��o�ФϺSW�ٰ�l1�W�1�"�Ԥ��������F1v�o���,��o��*���6R�ER�jp�m�������+�R[�e>��'�� ��ؙD��n��I,;j�g���3����U���˦��)c��>��S3��k�*�1x��Je��F�����R��o���i✴�/���6���!��6��������_�Ȣ3z����ˑ^mN}�Ӊa^��ea<�jF�s��#�ʎ�֑L�7ǁ����VF��]m����	j
a?c)��0�ξ^�/7����o�5U,5�V
L,��$	�t�lAB��1�.\��w�N�Gc��$��9����W~