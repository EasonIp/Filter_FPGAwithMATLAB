��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^���^�F�����b�}�<��S�����h\y�ӹ�+Y$�X5�%y�:�8�����;i�%G���oKp��5�3���=�l���ˊ΃�NA�|Gy�W�6;�E���f9<߄i�XTA�3vv�OW�x"��G���r�z�zʔ�t�A7��myOU�<U�2��qζ��'і��[�w�>\�����	�7�c78�o�N�𔃈�߅�P '[z3��j|��c|`���bo��O�%��ѶYɿO^�O�=-5X��4-; ���^ n2c�瞾����B��?|!�&y2�u|]�g,��|���*�)��}N�;+����'�'�p4�G������	����OR��Ɣ��?�^�<Y��~���`@ke	���+S .��a�5D���Pf[}M9"	�0��j��C�I��e�2v^a���s	��7+��w��[:b���٪�mϾ��H���3�{��H_q㝻�����Rݵ �̡*"��{i=�O���sS��U�^����V�)R'�)�v����Q� p��A���ӺQ�t�,��wR��j<Rl~(��.9")���\��Y�\"^̞��ǲa_>Q۔�<�v$ϣ���U�~kP{N�UZ�P��Ǯ�G�$A��_���]5~�*��b:��nNû�ɤ?���:�<ՠ��S!��Ɋ��&��V�!�Z�2AB�'��1=_y�y�M��4̘Wͼ�>V}���VԄ2w��T���r=恪��[��l�+���\�r�(� �`�p��@�)`���ܮ7g�3�5b���3�;��K�2�lPLνbg���Yi	%oSI�$�a�*<�gb�>k���m��_)-���A��r� ��V��W����#H�:'���ߑ8�T^�K%c~~x��g���l�m�a��x"������ץ�2) F�Ϥ܅@`,�����t�͑ö�w��W_<��bMH��J6+Ϥ�F�>�xx�A=��|b���A�O���brF�� ��@�O��!�"��u�|B�3xK���*.t��o!L���I�oV�~M�~����1�圆�8��7�"Y�ҷ���̞ͯ��a@�b�l��Q&����u��E�����7:2��d�օ�)�O+��;�x�:W"΀��y�I���a~�x�Ѓy�3�f�&[^/l��X�N�@�>��V0q�13��]�_���m��U=�)��� ,�ә<���C�4��'�1XĵeiW�d�4���yNP�����u-],�T���3ǭ8�t\N��t�;��c��VKdbL��Q���{����9W���k�׿e9fSM;�G��ھ��_'9����;%�nfgB�o��C��Bt�����(z�*�~oI�ޙ?N������V.��4��@��uq�9��%F����3��Xy
{X�؃)��J�k>�AϏ�9�$�X�7?-�Mb�z�?\���v��FUܖ�)�%��=b���y���,EJO��u WC����*�l,����:�i�p�ރΥ�TbA2B�ߖ��D/�U��sf/2�*������[h�z�n_n�R�ɺ�trT��׋U�fq��?w7w�ȑ����"�_��%I\��*�[B�2�\ؐ�9�����V�Nw2����WG�QJ��T����G�"U��mܻ���A���_��`�yޗ�'_�7H���qՏ�[��[��&��c��)ה�;	T6P.U�.�=�Hv>6{�y���BwD�~����ff�������(�(	l��h҂�Ư*2�A���V�aqa"E4�n׹�)I��_���@�=ϼ��s:>�M	ϿLg XIbfT�8g��HU�YP��M���E����
*��K&y�}�QEv�SA*Z��f��^p����q����p�eԚ^�qNȣ	�%��Ac��T�Bʃ+Iڵ�S ��
��1���:��YW��\�� @���,1����TŘ�]�"��n<�;P����{�+�����x��"I�OƇ��-�{W\��ez��]������@1BV�*ݤg=�`���S:�aƼ�8��ao��������^�q� a�����b,�l�V��k��Ԍ�9n�G2�rB0�G�7���t0�~�5,����T�R2m*L C9�:z����|�A�ǌA��ߢA�LMd����5�K� ����˛CKｻV��a��~�JDƯ���Y ��]�؟/�������YO� m~n��ة���N�~q�s�Y����?�v�>�;���X��oU�A�;a�*<m!�d�������B�&�dc�`.�x8�H��T���;��^􄮑
M�HFf9�Ղ�n�&��)�N}��m���u��ᕀ�m�g�)�[�>,���������׏08$*d�>&��d �NZw��mW�����G��<@1c��=�Vg�0&�묌x�k�O�%6�k��U���#���.\�C]�CQ`\�Qu�P����#���_oE�m����C�(tKƈ-q�֛�D̚�j���y9I�$����j��Y�n���f2�*)+���X��M*wv�[�t<jO�=HN��1��k�R�1�m��7�W�
x&���#ŀ�2� .p.�)�U�����qjR'��7�<�BO��2�ه�\ v�c-�CS��L`�0��,�:�Q�n��9��~�
�f�XxB/v���O�s�������n���x����c��BC��C�C ��hr���IҞ�%�l�BE�]^����65׼��M�"�.��~�.k��W�>�8Me�A<����4|�ΌAշw���1��ߝ���m�:Q�󜔣>*;Sw���!atj�������m��}h��������S1[��{5��9�̃�1p�'��п.��tT¸�n4�	6sy����zu�������[�D�3��c`KL$�Gb,`������I���˻�z����/2��cX��Y�tH�+���lB��-����)�q��%C༲� m��H�� Ht��mA��+�Z[�M)�e7�F��)��,��J$8��\�r:���ޑ�i»!��}�_�L������!�36r�g�e�&���?�(,x@����l�OԊ��gG��S�k���至\D2�&��U:(����Y�{�w���hxl1��v4h�� C��p���ii�.��$a~��U`��	u������53
 ���S�o]���3��޲���+�ix�X�58G��a.|�L ����fΗ+�xn����N�I��*���7��6�x7B;�#䩄�y�~�a��fl%[a��v;�䣵���	�!�,��	~��Z���6�cn�~�M�����9L�:3�-�$6�/�%��G%Hw�,�X'�V/6��%�ku�Q����WBl�V���D�F�f��rτS��X����<UW\�M��|��쁞B���(��[���|�4���.�`箈;���-�-"&Æӵ<-���T�8F{r�w������6D�8ש��U���f��e�2����AÜM�A�w�,��`b��rj;�I,��(/��Ҿ`_}���@�5}^��zS]u�ʻ��6�d��a���k�܉�=�����{�����ZM��qt�����Բ��f�����ikQ�^WZ��t<=G}$�������xH_�n��E+����L��S+ih�[8�T
�C��D�X�5�be{TY�(���-�_~�}@i��i�޺�NX�[���'��ع-�=k��^�~M���
��-�6����w�����*�⠤-1Rt�O�*��e��&RjE���)���h���A��ܠ�O��:�3(m�wV����cY$p1:���� E)}`^XߋqH4rZn}�^_��G�������-��*�L\��8%�}3�r��x�>R9�;��?2���Ε�9�ܿ�f3k5�Eivk���F
o@��Aϗ��m⅂�G�d3���1	���#)���?��@�*u�(?q5��na�_� ?H�Ni��&O�#�U0��1��H�$���1�;����^HYە�`�<)�Ԁ�	$rG��oħp��%��`WD_^泦�/���~�z�nu�"6_���7� W������{.F���e��K���3 u��k�}£W��}�*)]���=]=%�x�#t��z�+p,���2������= �g8�n7�P3Bb��#1sχ<�� o}���U�\�9!y�M�go��~_u���)6������ߟ5~�rS��.6�5o�z�\��k����Z�3h�|k�3c��� �J,�� ����<�|G��!�o�":F�ԯ�C���?�3�qB�K_Lt^ф�;s?�C\ZI�Nnd�q����c��!~O�p�6��#��Y�r:Fup��,�a�����En_�X�nP(q�#7�2�B����W���v
�?k�q����"�^�$��vKJ�R�]b�Ue�_�h�\��J��yY�k�V^�Uz��/h`��
@ǃ��fW�~~�u
��Ha�T$կ辫� ����Րz�NL&����`z�mg�@v�
j���Uօ&jq�fTB�oG�d����7���dÑ��R&����jAX�|�Vһ�s��l)w=4�ER���{,�*�f{= ��9���|P���ˁ�'��E�J �T�?$�"|���j9J�� ��r�� v!��J���%�ra�����1aW)6tsYW���X,q�����9��|���ycJ��	l��y�R/Շt&!%�͛@:A�����W��P�!2��D��s���,�+���Y��Z�4�x�K�P~���f��u�՜Bگ�lI����Y�����.zɑ��1(_��ډ�`���cZfc{*NI�Z����p���`9����yiPe�ǘ-�ip�*�"&�b�}G����������@MuK��� ���+�ך����̎Yɇ�h����Z����!�wj6��˧3=�عVM�
:�s-��\�a���p��]�C$M��2\D�Nҡ�L��x|S>z9�Ŝ��'#fW��W�w��5���Cntq�Q�9G�F��PKqÓ����J�?y�Q��ڻH��ʂ`�ZH~� �)u�9&M���1F�CԺJ.�y$5���Q6%|�a�Ò ��A�H}�˖�+T��q��쾖��(����X��g��.=�{�U���S����EHi�O26��Z��>J�4-��hyrR��2�Pi9v6�.��,^ɵБ�ĕV��[ ���k 3���3@:Ag���@�}�p�~\9#�:?��C#�<��,F�:-kwXGǭx�Je�Jsϰ�ږ�[C�I;�k����=1`�\�r ْ�b[h���~�?�HL��@5\�f(Yj�/ڒ9Q����)��8�L{�:���Z?�/I�hAqw�ws��8���2(|����fG(F��ᘞ�9)b ����m}16pf���.+���,X��C�ۓ#����ll � �O�BrP@g���u�3^����*-N���;x0!g��P7�ݗ\O�b{I���+b���I"���_�%J��O8���H���d��O,96��h��e��ߏ�E�����s)!v��g G��!��5�!c�h�܌Й��A^�-�m9l�7P��Rn�3�|*#e�~޵C���/��-PUv��?)�Q��r�3c57�u�C ���41���N�C�s��i�Ό��E���pKІ�#���@V�*����ņޟ5��<إ`,,e33���Ce5ͬ����������4X����U��)�n	�yQ���^ʼ�t��'�ȍz*�i'5z�EX����lv���+*<�/��f@J��l�����N]j��,�?I������>d�PiQaJmX/7�� ��<�����X,X?أ	^<��]��P���;��)�����4l��t���/��kr��h/fYU/#u m��O�a^ ;.��f�r�Hkх8���l�ݠ[�#o��_e�6Yp���d��X�Of39O��Q����?�U�r��&�fc.�j~0�z������� e�n�*�	���d�W��zԊ:9Ў)�M���l�q/l��ļ�1������P�T����ʘS�U//l6׌T����?H���m9���1�����B_4o��h�Q�xK�f��LT��H)չ�eEru$8mmBZ��b����д:ɬA�?J�
���;Lj���v�V���Mz�8�pu>B��ןY�������p[l��lX�68���'ד ��2��q�83�G��Xp��}ڸ�
�h��M�{��u�ƴ--d3>O����>;;�F�׌����z:��3.���+��݅W!�?�:/�o}U&�	Ab�sߧ�yT��'�%�L�B�nq���
#���ar�g���d�6��6{�(�+Axy�F��� �����U�0ſ��2
���U��9��߱��3��c�;}{'�P}5���=�X�gl-�v��[P0M(�A޳�{��0���E�"�J�b�s��G�Bg��$'�+�U��=�6��ի�����9��rC��~8�=��3�}�t�:<&\� msb^+.g��?����P0�
{��&c�.{̹긧�(���i�*���5]ۀ�Q�AA�H|@"|׀�&LF�5-9m'�ƾ��Py�	X?1�'����+��-�/b9W?�
0V�ܮ�+�����+����&%�|Ǌ�9�Q�;:��b�8��&n��|u�����唯r�8�����=bGO�ܭ+�_�^ϳ�<��4��aOc��o�~/['�Q�˙�2I�0"����gH֞7o9׋�}W�Q����By�p"�P[:&h�D�A:��؄�h7��R-�j�b��������/�����v��Oj*�v�XH��ekb4�~Y(&��^��m�k�ze��{t��1�����8+�"����0B�<��ɿ��@w��i��ڮ?��&/%Z�zw�L$	�*TFVs��aV��Ǐ� c���=ҥ7HJ�(S�n�E-�h8* :����i]��3,K13E?�:AR'�@Ȫ����'���z�%_����~u-�1NLե�����7��b�A2b���q���{JlH���:+��]�j��B��͉f�<
�]��yn��@�$�7ҌаW�9�c��G"�H�7E�1ku��L)o�7ܶE[�mE�E m�@�6l�������A� IQJ�5S=��4�)��t��b+tӃ.��!�W�_��el��TeѹP���)
TN��sĪ"�*̼TYp�R����V�!T�O��3�+m7�tx�E݅�������r��l-�����\��2�iE��@���[�4�@�����Bb#����+�� ճ�utu�ga�sPl�w+�����&9�K��e������øt����A�}D�Q��Z��R�M�~H*�W).��}�\T-�m	:9�N�}n̂MI9���ψ3���������6qN���1!����Rfa��h>&�]3ZT���U�jU�Xf痉�n�B�(�Vy]x��\p�
��W,+�:��7�dC�%��e�{����\KG��f�k��v����������&�/ے�_���_1��+>�Q�$Ҍ���]슗�Ⱥm�r��P�?ⷜ�q��q����Z�_��8�/�D�ZE��5��8!A:�x,*�5@�?E�swY��t~l���ߞ]$� ��5��рT� r[ߘ��bLt
�A֊X���OaLߒ�&�cc���Z�>-6F��]hj�i��x���LJ3�!~;)�S���c��^��������7N�XO|s�8����;�a�F�d߃�OM��kE�k��Qe?��	ҷL/a�pR�l�-%�E538�Ep9����:���#5�4�~���n7P�||��W�P�/RY����]Z+2r*���8�5�n�<!<�Eiԩ:>p�'_*��9:ĥ~Bzj@;��摐GPRa��\�;!h��zj����+�-���T��}P߾����y�cD�v����_mBU� _Pj7� ���&��&�z���G@%��v.�ڢ����b�^o����`�Z�/�[���a�����Mlky�+���	A�3���aHd��v�������v[Ψk�F�jxL�	_T���	�����;�p^0�J�S48��%׃ݫ�h��3c�t{�i�d��?s��FCb>�A�����^O�uyh6
���ڱ,�,������5�m�9[K��{jF�T�	Y������5K�
oz>���Z�z~�;���1�/bFn+��A��`�q���B`����t��ʮy#��)���|����7���o+ݩK)O��#M�_n��^a8[�yCgvu8�V��kk$�T����r�_AL��5)��^Ҍ"�H��_l��iv	ug?�_�C�wA狀F�:�����w	Ӿ�I�=]���'EC��w��X����9�Φp�!x�?�[�,ٲ���<sn@�� �en� i�垗��gW<�+S2��������Ww����Q��N:�i0�ȍ���;�!%qS�\��^ho@�gٱ�f�*�"��ĝÔ���|�aS@I��.��)� �#�m����?F�+i��Q�f)��v�h�蘗va��^"5��/�2��c��*Q9dT�v��Kq�Z=wG�]�~�x�>����&�N�Q���F�H-l�#��5ڽt�&��	��������E9Nf�v�-�yIˆ�do�~52M����k.���ǍqKI-Q���rF*�x���mT�3W9���@���ԕ�l說h]�#�y	�'�qnI������	ً�4W�\�c�?R���M�l��b��bҔ��e:w�㮾'u�w�b��M���/.{��2�!��2vs�	G��3U��䕖�,���?�l�\��no���ޡ׹��*�d���)�N�2��h��)yF^�#`J���
T9�ƩoD����B��[~���8xp�ET��іRxE�*�%L����W�( �`�ƥ��\Q���˶A���ݖZ����
F@th�(~��聙���n�S����TQ�W�^�;�\5���A�n��sf]��]�a�o��kQ�e5ˬ����BN'�$�pو����yAQđ�`P�QX�R�* Х�1����ա��-qP���|���-�x`�}�J�	Ƭ�&ݣ����y������zv8���S�0�?� *�"��p��w�8n��"C�1�*���팸2�P5���x�UB����� $�Ja<6Z�E%s�+�$����94D����޵K�Fc��](���ic>@��2n���v�w�\E�b���n$�yxk�O'$�>��1\xƋ�#^M%�^�%����UN��.����g�e���x��KE+FM�:mȌT0!�\������t˘.��("jwle�?!�Hk:�"z�	IX���C�	[,�T<��ab��X�(�T�AwP�HmҴ��\��E�'�]�y8n\�5Z,���"���uI�ϛ����:A�s)��������K\�)�ا�M����	dB�ܯR�QBP�$Ӊc~�~+�pɐa�C �@�ӛ&��r��"�yR���K�is��Y��pl_@���L��@�J$*iN�m,�q�D� �h��B�Ǒ�-�̔�!�9�O!�YW�f�/X-�'
@�I]Wz����Ԯw�ǴLx~�B�$̦� S�>KY²1�LnN�v��/}l��vV.���{\�v{O��<��T1,�)k'��D:�a�e�n�d�I�Do9�2��~̂�%h|;�:T���}�u7�Z���d� lg�I�L�K�Pܩ޵REh���W�1���؅jv�W	�yĈ�]���L�ō�g�%k��Vk�T��mMo@��	M�mɗ�P�l6k�BTr��lUs)j�Z��c�[e���;��\��^$D�s[�U�2���V�
�����H������,�3��2s��I�'��ǔ+W��  v�UFV�Ky��'�_]Z�K�W����n,ݎ'^{�7��ǘ[t��w�N�xvv����v?�7=^ ������@�Ӯ�f�����8��~Ln>2Q9�x�)���y
K�G��g�(�h
�v���8�z*�
���o��!>�ŏM,��[�\-4y���ɑK���J��}棍5�U�W�nˑ�2�a���Y����W�b-�7����'�������&2����\=��3Ee�Xc�{�����Bs�v�-����z��Q�&��k���������$h4+�r�'���r���J�����)Y"�n!���:#��֍��lN�"�
���n�ޞ�oK�{��q�U�杴�KAç��+�F�ji�
�:y�L�F����"o~[JNT�H�E��Uf�_f�T¥�1gml��'T�t��������d�����N�Ab/�E̅��T3v�5�\�e�R��:C�*F�	g�.� _F�J��.#���5�2���9gJ�P�ӷ�x�=������zS�f~����Y���F�v���k�h�����q���R���x�,�v.%@��O�+���{��	iЋ�hc!r�u���y;���$���_���'�j! U"������YҀ��YI7���S�kQ/e�<��k��-�F�ݝ���1H+=tiىO"�:�r�?#�+Et� ��h�"\(a�ӊxhV�pE���Kfr��q��Z�f_3]IK��h`R�`:�MR̷E���̒`���j���%�����e������!�D�X� ��!�|�	�f�!EkЕF�4��\�맜v�G*ӹ�o������>Z�t�;H�'���]�w���7�T_������BV�J[pĀ�e��$��p?�<�����r�Q��5������we�W0jX�MB�\z(x����(��0�8�V($�j����wc� �m��#�ʦ-�v�>�r���5Ȭ������P�U�~11�9t��Oz�/�Z}Ǳ��8��.��W�5.L	H��q�/LNt�L�X٨�qsH�'9am���Ŧ�]P���=*�	�1	+A�d�mfPş�scy]�����Q��۪��	�� /��h,Yw?׏����g*�^x�(����S�3c�F4�\;9II�X%��9X�I��I>�9C3�TMx��	BmW[�R���%�t���sף��y{�%���j>��0=M�-g���Li	�/ޡ��^�=�i�u�O�f��V�=Q��_�OAbcIczv#��SJ�:gi[�ՈJ��:<p�I�Z�t�9���U�7����B���9Ƙ�O�H�070	�L��<:��!�(,�<���W�/&P�;'=�δ��\Mv7^_T�4�Yq�̣��4���yvc�S|e�j�T�}^ܴ��㟫@�3�����&��j
zʏ�mw��G���pY�` [���i�<�{�A�h�Y�,�d��'�(�T����t�����݅!���MR�`�^	�	��ilK�W��.���!O�g������˖�n׾���'�U�w���]���[��j���zp!�Bn��)����&��;?��e.�����T.�b�|	��;���e{�PV2�ߣ�L��쪸5�%�ee�����n�s��&���/&�ʩ
v"��`5 �B�r1�rR����Ӗ}�QV��IIa��GgR�V�ė��(���L�o�L�k��j�N�\�s"�l�͸�t���,�5nA �u�xgg^ʫ�6s�tg��|t��%O����^n�I���^��(uV��!����u�����y��w��� �{
�5�Yűj��� _�ݢ����R%�L��˴n0��`��t�f_\uf�N��2lk2���w�49�D}-���{j�NM���A1�2g�Q�Ə�j3�$���[��*`#l�o6��x�	*p1l�;��X��;�j��S$з��?m����ɴ��>B��{l��-�ѤfM�T�`C1L<e�4����O�Tٱ�%��kP}<�^c�H�7gIǌWھv�����M�d��=n3ؖgV�ew�
?Ѭl�ѷpv�_),kcj�?��_��>���'�.�K���F�u���K���ժ�����y(����+i��8 ���@� \�G)U~F������:,z���]P�ƌ%_�A�b�����m�!�p��!
����I���Gѐ�%��V?���^Ph�
�4K�y��P�:�hG�`�#އT0uj�}7��צ��R�VbF��ՙ���&I�L����[��]����·���������%�	7y ���L��:��
AQ�jȺ6��T{ˢ�V{lP��L���Pr	 &
N[fm?�~F�$��y�-p���U��ƄE�'�Kzy��i��h����р��/�T������(�(h�Z6n���(�W_�,�\Y2jZc�bX��䞶��W6�������ɱph�sC��I��+���v�%���}�H���I���ɇSע�������U�����&��*D~���<]������֡�Ȯo��bqeq"���>~4�VvJƽ2+ܴŷ�����Z����B��[jH\���t8D�Z��u���T��l50LaxP�)\Ʌ��Ǿ��5�Fֆ��$��J���%P.>:�R�g�p�=����Ռӛ���@�k�i�r9ѻ��S�|�y�c*9͌����m���!.��)	���� ���x��U�*@�KU�[nl�ȿ��9�A[(��̲�50 s4�3N�y:A���Z0�%X|�Tqh��ܒ�[��f���7D��<����;��c2��PDu7s�A��Xa8Ϫ���d��5�"�PE ��@[=�*��$�ՏsG%���q+JZ�&n�;b�ׄ��O~�Kڣ&���cl��|���|�<���<��z�
�-is�4r~`&����G��Z����}}B��5V�*���*ڟ���X��eS�'Ŧ�ɨ`���ݱ���d	���7�����埗_�SKˋ�M{�F�
����0�l��JA�XE����'*�c�o�,!�R�S$T��,�T��^xXw��ev�ux8�|9�zx�x�+�tT$���9��|�����(�QH����6M_W7Z��zr �H$��0G�K1]�du�^�%�Pu�)�����Em
�XR;����:������9n5�54	�6>ը�c�bFS �.S�Ho&��1�0l�c˲2�b-�U�0����Z��*�7����?�@��Z����o�՜7G�D��%��J����{J�6X1�B�x�݂D���9���2�"q�S5�]�n�W�G����������M6��!� ��L7��E�Eɍ^�5e�e�a=�c����0� 6,0y�0�����2��7H����DY=y+�]e�ի��i�|;���rQ�����)	̲R�^�^�/I�(톜�&7(�a8�d��D��9�����6���T���O]�N�4US|Y��yp�v���Oކ�����;eQf�v���G��� T�Are�& �)DU�7@��4��� ��䟤õ��f=�5�3���9Q;�&�Ps�}i[�3Ū�{�@� �_ܨ�<�E�4���gēfrk��Y�$U�|�C��Et򀴶)9�~�m�1��j#����j�$i��y=��qf�7�!�X�Z���q�+��!mFJՄD=5UZZ�({;��-]�@�>k�~I�zu�����}�u�H�^R�j�ˀ��� B ��`����GƬ�?�`����Y�?(Wƫ�6+f�X�c�:A�2_�P�K���;OW5����W��SO�a��������~��<��ԋܿ_0!��i\Z�Tg�i��Y�6�e�a4:�i�F��(�B���P3��(���T��gn��^)���>����tZ1�ѱ� r�}zt�����9=�Q46�ܮ�Ó3�%?{� �әܧ�lo��UZ�o*Sv���~Al;�$N��Oa�"1��(���ڽ�+��r��VT�2�MV@�Ҕ͆��3W��N�{�����G$#G�l�	mq�~{	��t�py�?O:/Hdw�/{N�����t�f��]��lI�R���u�#�ޔ�/��tfU>�z�~�/$��f��:g�yk��u���/�-wuA;�E���G�j�LM�p��Ĵ�Z^;ǦN7:-�hf`�1~�m��[δ�In]��#e��*��g�x���ɖO�\�]�Oӫ0U��m�i����Y����<��˿}aE��OI�ծ�X?[i'X���Y�;+�UT
7�5��rgF�QXl +���]�����o��r4��fDI[��X#��]N�����9 �?�Á/PpǨ��\�*��H� ���{.K��JU68{�g,,����nָ��s�w���O�S�ȀW��r���HbL���Ш)�ĪF��Ģ�@[?щ�q��^�LG5 ��Mk���ְ���g���7�DG�oͿ�}�O�IG�z�_�I�e����6?�I�,1��tܹ�*�Z~�8�q,�ȉM>�>�v�GX��gn�0�����tR�QT�s�D�����b��v��#v�¿Ec��@�J)�I'��?n�Q��ǣ�l3��R>Ű�B<񤴙B��T��Đ�׿�&"v&�ul�D��E)Ea�<�
�� �����2���H���$j`}
 c,���-Y�����ϏLᅵs���*�b�Iƀ�~o�~�P̡��������ӎ�Q��� �#&���M��/s�mP���:� �=Լk;�]Ų(~�CK�DḨ�E�jO��A ݡ�T������y�(<��*�~
kix+Ä��#��o��V��G���
��Z��d��(i�W��W�w��ǹwU�)dl&�Jq~'ɛ��(8�e�����k���=�oS��Y���G�o��&�(�bϥYe׳-5�Y�2�w�etj��	,|c���ڇ��ߤ��.��\T"&�0���pY�ؔ�<�� a�(ڷ�-�,���b��֬yN�R���pDtyPB��gTf�Wc��l����ځ2vUc��sKu�=I�����Z�Qk�J]P��9Y<�ͷ����G���A�=1�,�ФC3C�|㱗����ǣx�J�un<��Sݽ��Y���{�NUҳX=����gQ<�FO��gL_�!n3����S9
�u������������W��}�T6�Z ��D�o�T"�Q��4_��M��#�߁�]�d�@��lQ� ����^�TB�Y�]��7p˒�l�0�����Ӡ5&�L��e~�D��Bu�ʶs_�Y@o�Ä����5���U�<�T�CbڃV{�s'�z� �@�O��:����0��!���+Y~���%�|1n)\�#�o���bE=���j�Ȧ�>vK�jEݥZll�ݏ�3��N�4\1��{@��kj��!Bx�W��o¢��_\[�DPA��t)�E��w�-��y�Љy�(���k%��Ռ2�4�mfh%育�����]�m`���I��Ϩь�֓�m1m�L%�ME ��#�Iq�4�;�����x���H��i���L٢�����AU; J6ڮ��ض��*,ȳ�O�(���2j�CHwq{�ֲ[�.�v�Q����=;@6�A�ň5�t�_»�YN�}�h���Y6sn�(�;Զ�"�|�C"׆�*_$VԂ�ĭ=5��dD� !]�m_qI�5���X<_�����k���A@���E�K��̵���3��iaɇ�6s֤���H	��3=c��ܷ�����aB�'��M�ڳΖ㗝d���tpD;Pu���2ʒGn/��v	��ce�����G+�tZ�\`��Z��Ϭu*�@<��]��Fɽ���/�/�-�Sq;�]�YW6p�k��7!J�$2�}7#�m%Y`������ �g�'��\ʩՎc���sX��*q�`���؉�c�
�[W�Y�?!K��ǎ)�c���ǖ�|�|�J�@�XrK�AFN5 ,%��.J$�bhڃ��G�%cMc!�3����)�G"K�f�s�������xfw������ԣ�(+j�Ox�B��?n����n�������t�h�s��q��>?�*���Ed��s�2��z�.N�@,0�dh�f�J.l��"4�#��"wϻNl�A\���Έ��@���1�y����cXa�v�j�#��r��2������&�G����Y�ױ��a���[�J-�#E{�X��W���U=^��P5�~�%�<�u	TX�χ����DR�k����+dw� ���g�.i	��F�ͤ��8�b0m��ƽ��#_)�s�c��
zH���=u�u���j��U���J�ݗ���]F�\B��H�%���J̷��LǨk_L��i��}�aE�v�0��)T�v"�CS�7��
�X�
K���ϻ� p\Əi �5pfY%l,m�V��^��<�������'����[6�� �PW�wѲ�-(�Q��4�-��-<=��mܺ�9�f+�m �P S�x����H���xH�?X
�jIH�ɭ���rK�Nfښ���K�����p�X�����z�OE[��E	^<T��A/��Y k��:­'�\���x��f��=A�UƬ �X�1�_=Y҂�M�1����k�nZk�~ s�'�ic`)���w���24ĠR�^뾞2�SG���_9@���܉)e�0�Mr�r*�q~7��������el�]vZ���~���\Ѳq������� ��AK4��&B(Ǭ)�VA�B?���4X��:j�w�+���vo�܈u
z[�����9���)�Fų'�cÙRgn�hu҅��L�(��Ѷ����рm�q��v�*��l�g�Q�5�ٍ�=DE��7�_E#��K	��C!���X2�� �%g�L}����H��������^�G��I_A�_N��_�:���,�4�s�dSξK��^ť��z���e�AG��n]M|���`���>1Z����w�H:޻T���:�v�/��?,"���Zm�mcUT�%ka�^�������,�y��A�	ץ�dLOV��^~KFXi�>>}k�w��h���q�Z����1i�d1�U����>���ߨϪ[G|$/�ؑ���!G_��qr�˵��/����q]E����@�%��2a�;�O�X��G�bU�3�]�=�I���S
��h��?�ܒ_�)�9�����F�����Z�LD�QB��U�O&&�L��o�%;u\Ӗ>��%<~�K�ݎ��Е^gNr�S*��ca]t+�G2�,'u�����ֺ�B�_5c�T��W�[6��U`-~+5�JҠZ�0�-��x�i���Q�"�$�')+�a���iD,��*'#	%��Ȋvi�ϰ���P����nص��w�c����y#)�{�_7�^8Z��X�h�������s��LH��]�ɘ���_s9�e�}#Ր�G,�����i����~(z#��5_�*.�*�^"c��6�C�x��ٵ�L�X9b��f��;'��H��|�o�ⳤ����	���g�wÃ~�U�����c,O�
�7+M�NPY=l;�pϣ��cd��U��l����:�vğ��<(t���7�挆W���Zb��)�d8Wv|��W�����K�4-��>k�Ys�~�&�&���!:�<A�:#�D�\\V�'�א��Ȏ�f�r�;���M(~*�G4$�}���Ѷ	���������4�⟣q����S�v�R�!O9��>K�{�����G7��� �6����.b�1�>3��o��{�$g�����
v��q�U�y��iH�,�� j&���g)x��|�l�\�����V���{��k��n�ToS��.���x��#�	�������i&�1X�2���K
&�96`VGj��� ��a*p�;/���S|U�����vH���u����K��>p������q)|J6�iֻ�1"dP}��^�u�O��UE�S�t)�;+�sx��u�{ڎ��ip���FDA�\H��5�ٻag5L������G��TuŪ�()��Z����M�X�18����-%�5̀֢ᩞA�0�N����(�j\)vH���M�q��B�a*dY����u�	�F^-���h���I}X	L��IH�z/ҳ\��R�{N#��W �L��0��<�@���z�~�Y$��-K�T���q/�����찔aQ�(J��W����R�!�/�*\9j6����`Fqz�T�8�v����D�/3K��yJ��)¦C?���GsS��31*�!��St�Vs�8�������.!��H�(�H?k^���v9i�� O�1��#7ۑ(��c1X��B9z0i��&XBh��p��I|�����r�:|���؂��g���td�A#��M ��sϔ��v��VG&��k�bO$���<<}�0��w��G�Ѡ�'8?�*�`�:��؀��e�[@�1n5��w�a��!w$����EH�Z���p1�`��D��1�/yV�R[�c��>�R�d��� ;�W� g�<5�$���
��'��9Е�Ӟ��&O�P0���
>��V�`�Ը	5�@�o]
��U=i���k<1��JF���p�%��\���e1,󠒝�G����P��4��_��Σ��-#X��失* ��~;ˏ�E�c)%2�a�x�����Y��'B���|"�/���h0e�N��B|w7z��y#�4A��	!y���+��#Oc�����+��v�EՏ�G��un%VL�1��	�ݽzk
2�`���������01�Q��&�RL�lku���/�D�z�?�5-�lY����� �}Q��Bx�� �؄|���J���r��uܛ�㪗喻yMꂍt"�*��*�0�.(�S�Q��n�$ ���R�T��Ա=�\���	O\�v���aC.��=[�|�a�%W���Ys���#)Pd\5^&���/��:�Z���z-��)��;���Mt:A�|���Pڡw7�#�N�@�/Ln���/4~��A'�d�-ƒ�y�1'5�?&$@
*�ƇrZs(r����9� �������|�MЯ�g��Cm�%���әjw�f0d�o[% ��� �%�R�8͞��i-��97�~\�0�N��N%T����b/�121�ۄQ`�
&	Z�:�o�?�7<�?E8BkI�RG��;`Wbԋ�{���w��TF���nE��B�$�j�|�öó��$B^i@�/bG�,�PWz�@��0=ݩ�񴯇��]�@�q�U�4�/�i��E�P��&�f
�DT1�=2Xe��(��S�la�J.)�59[V��*g��+@(��w.�R �J�/ﾗJ_$V~�;����m⩁jg[z�b�'>����^��9\|�+���,=��L#M(Rb�O�K�UzI����z?Ȑ�K~KZ��g8n�������eM��C�t�Z�jevڳ[����R�i��X4^5I���k�5u%o�lC鑽_|J�ί�Zu�e��S��┾�9�+x��=Of۶t�R��]l���9�]{� �'����m��:�"��}sC�������<��/3|IJOd�����ٝv޻�ǃ
���Wr�\�B���UG*^����ԣ��Ά�|��г�h�9���B�J~��=��J��%��T��䖮�%�/Be�F`}���8�"TP�)ٔFb%�c�0a�S�����^��[p0�~"�l����-��o�+w[@A��f�U��ůbx�\3��v���d�l;��4Þ�	MIm�; p�v��Yh$��yU}��HJg_��HV#��*��5��uY�6�Ϥ����G������
�6%�̿I������LN��$�3�r}�$/�n �",/��?̫�<:f��@(!*De�gV�MPCj�X��ȡ�����g'YR��%�*�׃�~����i`�LL��]��[J��~�w"��xK�yc�X�L (��;�%	TʑcY�8wme���y[�٣*��HNo�Vgbo|M�Ii�I`o��l�������3�B䃷$ݍ��>����'�-G���ع�D�a40Vn�f$�"��gk���4ċZ���9V�W?#��VdC8���$1���ʰ�z���4`��j�༚����	�K�H%���L�=�@�܂ˀ�ѽ;2�'�N���UGzN��H'$���p�wغ���*G��	[�~�{G��8o�IꏮK��ј�a�S:I��?{N,93;08l��AO�Y��6��U�nM���;�K��D�<iy3K��.T%�G@��Hg3=؋83f1�#j׼1��o�O<����k���V�P"<|S�Y�Jd��a�V3�4rt�q��n Xi���EQi��Ʋ~�=���:�J�wW�,����
��,mG*���C�}����k+�pAG%�="�:������M�����-Ȍ_>���pD1�V�6����4�#���ֳ��0Hu�)/���<��H�y�t�C��us�w�]��a���8��`��z;:����>�^}|眸KǅN�S#]ϚMo{i�)�}KlD:1���Nci�hδ`��%Ata�N��yfe���9"�ʖ�U|,[aLo��Z����ƏH�q�Xl������=���Ƹ5�0J�x싸K�2��)�(k��9 �r7bpG�D'BlhD������!�G:�#9%rգ頢bÖ���s���� e"*��x$��c�֫اEC������bk r�m*������j�b�Kԍ4��W����;���C9�-�hJ���\Y��F�s^`8'�y���f��0"i���Q�:�Dw� wu�j�9�yxU���1��?�ʇ��4��:ve�A?�L"�e?���<7;�s�"���,f�7�铎��X�)S=��
�)ߥA�'
�BG�{��G?.�&��9���c+q��s|�d�q�M.����^To�!�8���HU�/"G�k@�f}>���7e�