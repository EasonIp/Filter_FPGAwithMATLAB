��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>���q�;�;�g�?�_�q�-�m��5ʞ�œT����
��cFZ��R:�'��o�xE[�I�N���B0ˀ�2|:{4�C[�p6~��n�?�Ϳ����^:٘�!,�i�dF��<<���0������� �Z�=+C�r�.3]r�p0��ũ�VcX�xeQ���t�9�l�~B�'I�q	����{w.��\;�nsϣ OZR�~'B�\��uӉ0�qlo��I\s�$01����?A�V	FV;��06���Fx��<9��ݠ�_$�̄X�Cv��k�Gp�i���ͱ�Uo��\�ss7&�'�"�Y�)���?@iN��>/@����C��/\ ht1R��+[�;�p}��9@�y.������GT�B���+̄7P�����6���ܻÈ#O��q����-2#�%\��ޞ/����Xҕ�b0Y� ���18�
-���j�Pg�c8�󘺸y%�F�hۿ��ُ�'!�����ۛ��l�� ��n�a/�P=L�OYs}؃9�9ؤ
�l{l��V�nh���R��aҮUAI��MS�G�C���#�4��l4<I�Blnq��ܻr�k=�}�1|�H=�#+���(t�񁡢��y��n��Saӂ��d����s����X��M�c2��l�b��7'"bs[���8�Zj.���iS�8��x�4X�1Y[�F�U� ��2�L����uX�!.R�+���KP��3�r��0Ta%�
MB�9[,W0G����%5�J����XnbZxvw���<�Z<E���d�!_����.���^�9ܜ OL!kH�.���U�<m�s'���G��ٍ�ֹfoh/H��t�t������QG�B��C��j�Yh�BJ8�y��?SPjgGMKݚ5}�Ӿ�q�Al�����uS{�j�iP#�芃�+�5�t&iQ�r�o ?&,,������'�Z,�p��[`��gE���xY��H�sAܧaR/xar+��oKy����zE�m�Ǻ/��J���ny���!���B�mp����1��\�e;h��Q\'��A�+/����e��q���]\�`n�"/����${qҤ�� 7O������S��y)f9G�d/,!R��͉��e�.����w�b\)��͸�	���ap۴b�T>���p.o���.r0js��YR�*�(i�:�r��ap^%�w�(��W��������T�1.��0e/��F����ŷ�����]�#H�>�y`3�i�=vko]�Lj�!а�&�'�(�_�RS�a���xm��*�Aj8�5�e�����uͳ|�#vK$����џ�Q���֫����HBj[s-�0�o�C�|F�� W�ՄK�a�O2�Ա�N�ӥ�P�~�qj�J�j����y�&�����ާ��}V�Lo�L^(�o����'沎�l�\�U|z�]��ôd�T�-��^��#r��A�� �]�D�����B$�M�7�MWK���(�#5���0��-�Na��R@+���E����L!���u5So@�{AHz)m:�SO�!9M��b�R�X5=t�Of�;U�O����f�I� �a�lU�&���S�pA9�Oo�˪�껭NA�s�b�; �V�
~����bW10�}������I���Kj��?\3��D7fk����G��FӺa����6�̛�E+�D���L,8Tj��Q���#�Z�;G���ii�����=\�h1� w����
�v��žg!P\.Ҧ����@�9 "�)��P^�^?Q����f0�Ʉ&[�R^	Z3!y�0��}7*��m���]��(�&.4�Q���[�tݧ���L%�.{cv7�̻������8�M�au�����?�O��C����X:�����p;t���ϓ���M�����5��������l��9�ƒQ�n��x��a��A&�t��SV�Sw��S#;�}�L����e�'�5�-�"VXA��p�ʿI
P1���J1��W馵q �����?T	/8�)�sFv��X��=�e����~ǣ�W@�����`}Y����O���A��O\0�Ko���T�6W�[n����N-��\�=���Ѣ��=o��Z� �iǰ��f�=�r,��h�8g�:�ı�(~��M��VT]kk`T/�����'~����5��{�=�,��won�� ��:;���0	����17㏐A��$���5?3��#�4I�M����흱��@kK��R}�ǨG�����|��2]�{줐�r�=12?�S��!�7�F�����O{HCT�%b2��0#h�ʏE�&��h#���'��J��m��Y����f�����4�+"��^#���r�t�\��u!�n���K���\?�O���U�G��B�f�D/wh���S������Oy�X��FSL~��]��A�{�_�M�=�g[#U��	�KĬ���I���RHa�C�TK�Њ�e�R(	�j��s�76V%��+Em����kkC%���~�(v���&��/�C��2�j��_��-b\ 2�+T�����l�uq�Yb��������B7#�'�a?�3�Q�=+��\�;��.wwȥ`��{
�ޣ�Z�~���rj�|fh��,�d�tyE>nJ�cv���@AR�iͪ!��R�  �F�GjH��ޣ�?��m�9�HE�s�!�s�#�v��gE��d�%��2!آ�p\D�n�>|%����pExGO@�;���Xt�E��{Ro�I����W�Uan���*	A����jk�=3����(R(!ܲ�s5T��}gn�f��;�'�o�R�+@L�@��R�����,��8�9��e��2������ꗀ��*�K��z5��7>!��+Dm��i9��}��!��-%6��3��/��Ͱ�|���2��&���q�$�@܅��씾Q����s�fN�KN��V�redĒ!
�Ȭ5[���vDƱ2:��yL�H޼�I"��е*�-�0HM>";�˒�=� [A~>LAʁ���nOz�E��	B���0��nPiN�P��AcU�7\<r/Ǜy���� }W�����/Yh�(i�Yh���C���T�Co=%��J끜wy|�h��B���G�}�RH�P��^V�ݤ,�9��B�1������w3c8�����F�}۷�K���4���']�_�8ȥn��SSB�Qo�{W���9q�i��ϑ��+�>������d�kH��{˰8����M���ɬ�^�t�'��E���oN�[]	�o�ɒ���m�:��3�)�ꪉ�[1��2��/�ID���4a�_-������4u#���Ng�t'L�i����L7�g)�wk;���#�s�tz܆.�Gk�'��Q��'<���K�#\?@~�$�[B��'s�Y�"���,yj��G�����ϝ�'P�&r��� L桯�C�<��L��p�����r��Q�
��sބb�kuN������8�(ͥ>��l#�Z(�A����v=?3���z�s��q=�P�=�>�d}ƅ9��e��M�o�Ð`05�{�e���w 
�������a�vl��-!��� m�.ճ1W�.���H�/��.cat�/����M�\��U���G"tN��Ff��ύ60�Z�wM��-3�]�b(C�=CO�e�s�t����?�22���� fGR��=�K!ᙀ�R4U�^N:0Lg��1�M�Y#.�,uW����A�*�㟽@�;ǐ
�f^Q��+׬ �~t`6��lC�(GsP&	���������(S�Fp���!Vt�q��B��?A�8�8�E:?��2$|%�3��e���L�y��_����,��J��Z���Z�N�0�Ο��W\b�b�`4�`�n?��8)�ۓ-�?83qY�?@RU���p��<=�
������E�F��C��ȸUʚ~mNV��h�wh������uՠ�^iR&���z[yp��ٽǮu�#��9]T���ơ޺�"��D$�$�R�Bkg't�|�y�3��`Llɘ��ٲ�q
��[ߐ����If��v	HhvKEo�K�}�4�{��7�"�Ի�Kz
ы>�EL�Ұ^0��u3Ǵ���f��[dKi�).��2-��:BM;�%C���]KF�\�"��ゟS�ߨi,�W̄Bۋ�AFĩ-�X\I�n����<��{��]H�_�S��v�̛�H���J���Wjŵ��Nvr֤|(�r��1wX�2t��v;o�Ò(���ʔ�GN�Ia�T��ד����.9�,�V��*�	:쫙Ͼ�ʝoY�k�,��S��Ύ�j�v�~Kx�:��,-w��83ϐ�'����!p
���5p��&���뫀���M� ��	�4Yp�}�\A�oG���-�f[n�;]~�#S�Ԍ(`[�tO5���Y��T|���&u��E�Cp�~��N��;�y�|j��f���z�}�]�D>�K����e{��ب���1U�Y
���5��:�������Dyr��XR.�Ȩ��I��9��Z�KA�(�	04b�%���*Q�0+k�xJ���W+b�et�w�?�l��o�$�x�K���8b7�:�o��$�'����5����35�#�d�mk�����zuA+���}�S�2S�������+[pJ�v�=^�SP:�H!�e����9y���	u�����i�q\Ѷ[,\%�?r�,���p�[�Ϯ�z��{�%kd'd2���q��[�_�=Yd��a@bK�X�p�����߂m9o�����<�� M�ұ��X/f��b�E�H�)Bm�X�Ņ"�>**0��ŋTn���Y�h��2��`sk.9����l�LR���Ī������1��_�^C���?�Lgo� ���`6��m��equ��'��Yu���UA���ƏQ�IC�m.�)�g���k ���n{n:׈�ϭ6,���8����9#ݭ��T����Gz���_ή�{���T�8�K��PfƸ��&	�Ƣg@cVN�՗��#kG����4� 456nH]6IS�Ě	^o����Y�B�'XK�d�)�f>�����%^?�$j��1��1�o�Qws4Y��^��R:�� ��%6�c֒�$����C��+��=ǀ1Y4�5H	Cȧ�&�����W�HA����,�" J�"D7u��
9W��x�0w�S�C3Y����5Ѩ�ETl/Rrkvu6�¬�)#}�(J�f�6R�m��?�����5�r�u�W�"v�Mۿ����w4B��r�9G0_5�����AN����\����?HX�I��|_~X�]���pD/�נ�0�E�R�nc'�7eB�?��cB�~��
5�㖦:�gWuV�/2�j�/��.��AM�����)s�>��=4	��ah���hq�Y�G��g$�W~��֭���;W�^囉�ϡ�m������{x�/%e��\�(���|�0��tdb�d	u����x���ьM=�?���u�_p=����pf��7cW�pq�-�<���I]y��o�-K'|���)
,	t�1� g�Z�v��v.����~Z�bu	�E*c�����"k���ґ�b�����gr߅|qA�4hp�A�����w�?�S�!EMW5���D	*it�pWA!l���ÕO��Et<}J�)�{�|?U4��ťV��J�Y\r-�Մ�3ޗ�dD+�7�qK}'�Q�N�A!�u[F��a����s�\{?g$7��Le׬�˶�.$Kع�ԯ��	Dt���r���ٷT�A�'[M�Y�����1K�'$p�6�~8��B��8Y����vB�VE��9���ж-Z�K�'�_�:��v��J�Q�;n.�eG���`-��Ʒ�#��dJP4p�OR8|��Fح,��ƈ/d�.���ʴ��ܷ�,�`�H��r9qΕ/3G?AJ-N_{O(	�j����X��݅L��y�|�U��x�(�CK}��0���������2�Td��0�Gw\��E	:�_F<$���2�
�3��e.��s����^�í`͢��T��\��i���������	��'+�r����s#�K��yr�W��:�p���#�\8�
nk̨�i�~��I�ߘT�����15g@7���=5���h�Dh{vG_��[���Ǟ�P ]�zF1b�!��̌������Q2o8,�o��������21O�u!�tl�Ê��DQQ��є��Q?�+|�����6��'������#� "I�cDV�)W�ہ|:do��ԴS$����Y�k��U�xi5%�%
�^b/`�B�v�y�5��T���\�ֻ�PDH㧳L��V���賗��ƺ�����o��$��R���HGQi��5����Բ>]^�o�N�`x'S����3��{lP�^�o'����;M�������o��[�qۼ�=��hu;k\�e��ʟF@����D�b��[Q�X�Ӿxӗ�%��rufb��9\����R4��q�+�n_�������i�ژm��&�iJ����(���3jGc17�PC�i�F�}8H�/1!�;��� ]�����#��L�k��)1�!H[l�����ә���B@�%7GwK&ƈ16Yc�t�|FRN�)�:��կ��ס�SC(�:��qr'�t�CS�C��B�7p�Z�7�x�����:~~����9m�E�ɦ�b���Vh�����w�E�ߤ��J*I�}|^�%�,*=;(���h�PAAf���hp��M�[� [�HD	O�]X�u�<�������$)5�駟Rf���Hê�E/���s9J��ͨ9����Kͅ���N�'BM5��p�A�$�߉�ev{󴾺g�e����e�$����kc]��iz�~�_Qt�P�.NS�}S{7�6nF�|�#��>Qa��W�(3xi�U��#'� kF.���磱�����_M���GS��[q}�� ��aQJ�e_�������&�S��TA��Ez����>�S����.������ʿ��BbZ|h.=��Z���fnNo{j!��������U�O@�W@t�ԟ]ۢ��S�~\K��\)E�[�"�t�"��t`%46��'e45�}w����S����� m�?��G�B�2�#�6� �$�d�����?45a$~�!�N�C����k�:x�������d�Sځ�����b{B�7Og��孊���q�v֋T�l	�%����s������e�r�+Ojiq[UVz�m���!���&��E���_���V�eF���#�]���	�H�˛*�NS�'�m��%R�CbH���3�c v��~�"l��a�W�=ſ2�o8U��r�P���Z kw����I�I/O�8��'d�C��){�K]8ň����V�����D:����.{����Ռ [e�m�y��M���V��r�
�R���QƸ�H�Q+�~�,F��٠!!��� e�� �X<�gc;��/�"P������i�����WW1�K�j
^x&��c1Z�\�d�/�0��C�s��-��d76#n0���s��V���f�;���b��t�=����)�,��Ϭrp_���g�"���U��4䦂��.�鳰����D�d8�0����q.Ph!�'F@�&o�����!R�%�&'0���F��c��*�H�DE,w�@�_����L��B�D�rz����,�A��&�^�"�-��~���ϺFkm�
q�B�ޤ�68���9��_	�^���O�!s�4���u�%Ǎ����P�r�����Vn�!��#��_f(Rd�-�W��o�"anU�)[-1�M��`�'$~Bj?��Ep���Y�(y��t��˥G��7h)��H��e:z��YXIN�X{]<��pP��GGÛD� 7��D~��Zā^t��XӋ�����Sy��HpR���[9�/�~ȳ�&�&����ev���U�ɘ��]7���&}"k����c#�0
v枤���E����L�]��4UӏC���-��k�('�I6R��k򏖈*?��òN��?����>ohS�����k���>o	z�X�Da��(#�V�?̃� �3U��`��;�p
:1� ��D��B�H�?�,m���f��Yӭ_9���!L:a�zƂ�&�v���!�˼�+�A���y �A�:��::�P�>��f��h{_��o�mQ����E�HAQ 5��r�u�
U*��z����"`���#�
�t��^M�ٞ�A]}`*#-�0�x��\JE��5(��b#y�����)cs@��ßz�;�, �ե�h��Ǭ�Z����_�aɭ��8Y��t&�vE�V�� ���[r���cg�u���%�*[�9�?z��S�X��'%>��:4�-1�����#a�~�む��R��;�2E�E���=��q�������Ҩ�o"��WY�T����F����ҽ�x���M�a5�}O�RF���ŉ3��|Nm?	�l���B�i2�z\OL��ƕ�N���%�c�+_x飈�G%��q�Δ�)&29n y���_W,ŋa��&"��FCR�$��L/Q�C�`n_J����j`���w�:��*�(��&�bC�n��E�5s��WH���=����r�0l첑����~�'��&`|�L�Z���kQN�H
�\�Qg��:�ә�q��� �QT�,��_�E*�j+f?���5��>�}u����d,��9��j�^����tp�qe?՝f��F�I���9�����^�������^-���p��Y<��I:���jD&�jM�nJr�`�J@&!u�U/�.�]a'dd�� M@֗�aô�Z�p#�N�k<u�-8T�/4��hN�0�Z|�kf�\Љ�+T�I��<@]��V�E�r�0n��Lw��JR��*B��Eo ���96�tq SC��Ϊ4	�۹��e�9�Q���P�L�֞��q�.��Ɩ���*zd�"�駏hH�l�<ӄ��8��P�6���B��5���n0*�&��[y��^|{��j��M/���@���6�͏�{̺�9��XET?GYy��Td���׋bS�E�Z�K����.��5�n��� �������'%wC��ǋdFX ��%~���[%&������1����ET mġG�G>)��WfM����CG	�QD���d8Q�tgc8��t��u씽X�EÖ��~�G�y�o��[�:���,5�N3Qvt��i���'2�8�J�C��nѕ4ҴI}�ӧ�k!�&���I1R�6J燿2Xٗ[�	O)X(s�;���SK�5���'}�>�n��2ytdn6xN��"��"9���z�鉴�w�U���؉�����Nb��U'���.�I7�BF�n+?��q��S�����p6�v��G��[CC���J�!�S����{��s�X�@Yi�P�Կ\4u��R���_)�uЄ5q$� Vf�p($P�X�/�*ȼQ�ɡ�� Od�w+�'7�m���V�,��6�w���CH�z�����2�;_�~�{>�^�����2��'��G�P�>�����l)�+�^y%��x��}��>-���i�uVqXl�iA݅t�@��岎�K`/¨���ނ\��EX���:�tP,��z���p���^Z�9��g0vY"t���^�L��4`�H�ɗ�!S�s���
���~�c�
��.��_q&0�Q����l��y
 l�W���8�7q�pw�?
¤1��ޛ?�%g�]���M��~@hނ���>�Gmg���;j�����Fx��{���q�PjJ�������SpF����*x~�>T"芜e������t�6�;����Q�����* �u�xMo���\!��m��jMj[F��!x��ߡ3��̔3A{3���#�$UN�$�۸L���j[|��"��B������Ɲ<L����A��W�IO�,\�b%ي�\���B�����Pl����/��+�,�n��wɗ,)W��kbǜ�t]�ު�	͚���lgɸL$|�Ae�'�?�p���_�}\�=�������L�#cGi��s�E9�S����
�h�f�s�:d]=O�Xk�`G՚ؿWz�	��#�g�#qeM�k�����j<�>�y�am�x���1��9���Ϣ��OF�5*2SH_��ju����(�Ѥ��T�\.3e٢�KL����[���y��u����U��tC!>�|Ũ(�j��|!r��'
����9�����	�oy�؃�6�F�����n4��gO�E��31AH�{�į�v��wI�I|�4T4w����J1����S0�}�D�ݧb���*+U��賉�ɶ�ā��I_y�ۮ*6uc��d-#&�!�4�/�}P�p�]����&v�3���C�#k�~|����6��Jo~��
G���*�-�ְ�O��^�WO:>Ϲ�>��]�2f��u�ۣ�^f����̤@��i��+��a�NԌ���`ǜ���LX��b���2��mLl�M�m�
��~aa��M�{�$�3�#��w��#��+ �� Z�I�,g1�zc�d�@Th�p�;�AƠv�(�^?d���ƿOǬk��ږ͉�8\�U#D��V��o�jRo��%���Ff�B�%��`�&	K��������� �1�fo�P����Oh^����2`z��J�Ei|G������h���se={��&��>�I�8��#.�%|���g�v����,���* �F�]����u�sgo����^�luLp\J�a45W�J�3��?�P��%U��+Q�M+�	'���P~d�k�},Śeɔ[���h��MOð�	�$W���
��'ס�uuШM<-CҶ��I�Csͱ���g;=�f����>Hs�,L��-�a3)7�g���i�as]:���˗���Q�;m<s�ϏI�ҕ�����]l͍Y���ϺXVi!uϔ����zF�7>]������C��Kq�@�XJ𴆇^�l�DϮsf�]D��]ZFn�:�Gϡe���$W�k��.� �j�7;������$ɥ�4n�=u�h�t�9	C���C�B������ie���hc'w5X���S	�N���[����G���~���fG*8�>d��{W Z8y���ż\*�N�O�9����`��)]	���>ļxh�n��3Ԑ6 V�1��W�m�ē�����)�Cn��@έ�E��[��������o���Qp��8p��C��kSKu��t����Z�V�h1�}<����3�����'��i.R;��w+d�=�F��DB�Q��jڲ��nY?���2z�6yO���'���FIzR�Y��+��U�5��1��Չ��M�Yd͜�r��4�O�$��>LNv?�r*򿙁���qp��y���i��̼R�x��<��z�9�z��.n����;�Ыz��.�N�6R�_���A�%�*��E�6��gw��b/z	m��[d���i>�##\�nOη�Rw�U0���v��ȡ]�Z\�y���ޱ�,9�EZ�Q2�!����X1�*�+{#.L�2��]�:(���Y�� ���C��\��BDn�_����ꊬ"4�r��t��8��T�K��9p̂�~�3*�?���Wq���J<3���Gv�k�$����C�6Π�;Q[��:��� ?g[l�h@NdG*z���(��J���yH���&6@�T��R�x�3B)�L��������x��!$��qq"����h'��%W���@U�23[�8���@*:�0?��J��Ќ�%���w�o*��?�d"$��f�i��"������)��=��	��S0ܣ�OwrGszWd��r���f ��y���<�M'J��O��4�?�uf�n�+�a4�?�ơ���������~9�� ���
찺}� ��V���Q=m�����K�fEf�UF^>����s����EG/>"��S���Qq4^�͚�y�*��#�e/3k�����&#�l�\B��*���}o*Lt�������mg����Mdy�q���1�s�t��^:F��������r���F)n�(����3K%v��r�8[�c��l����Ɯ�l]��[9���)Q��$cx9��t�@.��}�+�����W�;�М(�`��/0�%��'�d�v���q�����<MDm�P�KV�=�襻�8�2���E�ά��C�[��Z���i�ꀻ��3�#$MI_���o�ҷ���u{�>��Pts{b���3�)���m\Gzt�z\f��c��-��0������r�a�����᷋+�+�$�(3!}��4�?��c�o�u
hi����=Z%H����w��0�E|�G��,"���)��C� ��p�#��bh��J�>Q���nIit����<DCX���/!�ǟZ���L�0���^t���W_�	Ux$��lR�R���<���nմ����������*���$k�e��5;;�������n��<���p�� �H��zϺF@��ڻo` l�\�Ů�B���\O�b�1���CgT�����͹s'V�:l.x)	�k�eL��&��eKZ'��|���A]��o���Z^���u�#6��c�R���&��4��H�U��i����s?����G��&e�j+�� �T.�[���7HPR৉���VP�AzF/|�RBM��!ڋ����d�6�:���5-����"$��g���=�P��$"�<}x��f����y��.�+���iݜ�����E��<
�3��ŀ�gWfq�ve���sp��7������*�:�*��-��K��{���D4��C��3�	����ȱ�