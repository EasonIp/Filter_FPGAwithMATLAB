��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$��c�\x.-�M��BDO���{�kr"6V���������e�R�s(g3[K�hK!R2(��G���g�uк\�ԛү���?��_L�(n�ù�6ª�+r��R}�0!3�C�A���	ҕ�h0�(��H:*�O��4�Ӛ�I�W}�`�)�d�:U�f�܆�	���3�B�m�h���3`�蝰շ��G�uPH7>�
��3���,�d����I�ă�>ɴ�z	8{r�-��̽Q�
/��ˋ��@X��?��J�r��3����)�k����C�*�
� �y�è �U�+�풠�ҫ���trX�0���@F1��Xy���=ڒ��{��"5�8�rh��a���Ŀ�Ʊg�0rM�Uw��`,�\�AO>�b���M9�2�ٕ�
��ǯ��@��P"첵���^�`�<���f���f�;tW���=g��ђ6B�o�sZGA� zU���P��c��{y�D�&49���(ҫ_b���k�;�9��^���)r��R�$���k�P(y�7���`��P����f�&+޿�f6^
u���'<��΍�n���'�_Bc��N�A)��1���l�T=��N����2)�~�����g�0	�8�_9ܦ�rC@.��i�Ұ6�Ӈ�&b��$>&������|�.E��YT�-�x�L�*V�۾�����_>)���g���(�hp���+H��KA�I)�)��������n̞�����b:������D��y7�{�s�H���
�r���];M��g�˛���a�E=�[�VJ��_4Z7� ��<C��a��ჰf�(�L���I<}a�\�Fh��	��s��r��1޷_?^y��MW(:ab�"/���p| ��nx�+ߔj�D�5s4�2+&БX�L���PG��-��!(1گ�����vn��.dSoiJ�<��A��f�&Kh��%,�ߡ>��Bt��{?�")��~��� � �m���q���R�T���3~��09Qeր�1Y�	Y���͛&E
{��z	� �1��]6������2r�['���ID����_��%�nl�w�@`?=#�Kc"��X�9]�x���Ί���=��k���׿|���>�����3�|.T|`#y����u�n��'C8��Z��8J�{�u���g�=jsCC\x��wH��{�����`S��n���&g�Tcf�òD}��^77�صJ�=�*)뼝Եɰ�I���aX��?�{���Ɇ�%�2��\���Ӷ��ׄ]�����3U�#'���|w�x������f;pg�@A6f��y����*]�w��n�C����Ե��J:�a�h}d9z�Τ�3kEXK�Wd/�J����C����/�k��i �`؀�p	-��n"A��J�ӱ���Q!^B��=��)��� o�D�ca2�sn��Y9�����@ó�����{��'����nFz�^��jJCOY�� ��	Iy�Y���۸`���u� >v�yP y�F�=T_���"؎#�+ݮ.�T�l�"�����0�8j��>���<+�u�J���vKF�n�h},:��	�ɳH1�V�I�i�Jp�Ŝ%}|��[��������\X��*�ۓ'RlOX�tIHb-�����o�2�u�$��h��e���Cp�7�oc
�h�L2����fXS�!^�S�F�Y�����r�=���J��G>参u�k9f=�u�i{��=E��џ��Q��Rx�� |�W6��CJ�Q�m�!I�:^��J�<P�J|q��С������}d�d�
��S�Uݎ�{G 20�W�����������2�5o���"����#S&��:����_�*�ь]�۽�2aK/��f%��&�=�b5O�����[j2q@�l)r�N�r`����5��ڋ�#$��������$�/&�0Y�S=&�����)�Q�q_{��§;��@�E8����%�7��:Gx�ot��v����Z���^��W
��a���$=��t�[c�J��4n��n$5��n_��X�j��!6�{+}`�����=t����+����ms��J�g�!3z�%����d�e������Z��Y�cGˎ�"2=|��X�HI��\2d�2I�.],_��]����>8�Ӽ�	�n�ȦI��QW���Y�aaD�9�:�"d=��Rϋ�;���̥�+�A�߇Z���E��;�U�]�"��pP���[ ڷ�1O��oݒ�KV��o��ޙ�C��{�Ӡ0:�B��V�����Kxz���D��0h���o�܄d"w���!)"��A� '�,��4{�TM� ��Ytk6_;%ԃ(���q����ۇI��<��@�[���M]��b�K�v<^5�
�i���D�!�o#�k�\�:B��MJ�d�A���m4[�o���0�/�7��XZ��ڙl?���$��1��;c^U.��f3�*�>�#E����{��#������I�S���r�l*��G?�E�^�~�їa��O����#��/ñ��� 
<=;¨ S�j�3Cx|*�S�_�#��� �u-��wKq���o�}kZ{�L8�EqWS)Ď�Y���}�����5�Y.��uxS�^)�|�rfy�y3V/���,!�Ճ)��k��B��_�h�b"cm�s���3wV�muh���V^��&&�����B�Ę��  ��M�^�俊ל|��DqO��3g��c�$;������J�s�����G�z#hFW���$�&��"  v�;֍$aj��\(�9�)
9�GLv���T�6¡��w��%8R2���+| H?CA��Ls��O��@
w�;�n��B_�H�,�~R�=\�ݥ)k��˲��G��wW@L���z���)e�*R��<^$��������X��l�CVu����nc^&ЧV�>�`A;4r��@0E�d63���G��SQ[�p��&�m�*؉ث��v�O�'�QWts�njn-�r1r���Ȯ����L��=Z�4~4ThΆ�G#=����ʕ�p>�h��G�����`�& ����6���#��P!�,˾��/9�yO�w�[�b@��s��$l��Ql�=ίc��̱�#�����;�S�u+��z���OO�a�k�N�-2$�R!|h͑��������`'4,���=-��oq�'F�g!>��e/����0�����+A^���#�
�E��]ű,�ɯ�f�@��=Tq��H�`��$S���/P�O96)���x���hH5!Ibj��wn]��[��4}�\�A���r�a� �+B�A�WXwN.������X�bt�����#16F�"������iT@�v`;A-}��'��ǀ�9g�B�(��KJ������B9#*��8~-{!Ǝ�����c�K+@����t���H���͞�T�����C�T6n�#`1����F�G�.���[�p��9� l���kԺb���,��^٨�϶�|&�*.��p��xzku>P0�D��R�ƵsP���2>�%�X��w5܄��Q56�S��mv�49S?����O�-0�%_� �_���k�!;rhC���1 VmD>�.�c=�:B�
��DxĐ
6�:����O���<<�:6��	U2���E���ƆL�D�9���/��5ml�a�p7�ߕ"~�̜�ڃ�6�u�����g�r"3�/2�01]���.�H�yOO.�~_�Y��!%fI��;@6&	�ܥr�j��_�2��$�n�e��bg9M<�~�˸p��;9��c(���SH��Ċ��0��sm��<�oN���F�hN��/�v���Y�D�B9�O�Km��96�p��	�3�y�9!tg�muz$�Z= 嚏��0C���r��P���gܘwŒ�*�r����1k��R^�i	Tc_P�X������(/�~X�Bh63s
��[��B��r��]�dW�T2����O����e�����\3��Z^��|M|E�ga�|Y�T�����A'��\2���TQ:)6'Tv��+\��{���=�+,N�*�!t;�3���\!�p�!V����P�p`!|���Q �	 �2��)�W������M��ئ��<ME\�2�G�\�b��q����;0�ǶRf�{p4�7��܀�w��=J a��/7dǠ����7���N%�����4<F�K�ٔ)�O�Z@8kQ��,�Q�J��Idu�$R|�w�b~k���;$@�2�5j�1�[�F-���h[XG����`2(��Бm���m��"���}�]f�{l�Dd�,/m:W����`&ݔ���սA|i�K�����ZM���4�#��ޭ��bQ�gS1�mH\33?�e_{�Wr痉R[��:�k�3>��YGW����B��6��"��*̌iq
U��cD~r{��7�eŸޣ�=�e�?FOWEV�4=(I��/�f�)n������� �C�(I�Î���)q��h:G��I�y:�1����U�]ЊXmI�tR��㶏��&����
bu�#L�܈K:W<i^I�s��0�8��Gf�����=�58%(�R��~��2��o֕O����"�V��/�N���'T`��9�z�@�T7ޚ��"tR>[��?y���= ����3j��I����0ω�iE��y�؄�|�0gU�]ؓ]4�SW�0�$$^���ZNo�B&K��<������U��ڞ�LБ�1�_ca�W~0����Q1)��p]����g&��g���2BSK�k~D��zɸ�g\y�L�Py��GAt@�IBǀ�VPT3�s�A�1���Wi�U-D����m��rZ_i�*���Q+ZG��ֵG�4�b�d��!�H���DbDo��sG�b��2 _j�!�j��sQ>ڸ��s���F��4�kS���y9��ye��0=4����]S4�����m�7!V��O4��e�[g`_L^	��Ԏ{�1 |��M��/��B5�nPR?#*ba��|��VƱ�У<`I�7���ٴ1�ov����Ş}A.A�;\���U,��Þ(�6�"`�Eh�"���x��q�W/�Ot	*�HT�F�^�hlv�ccE��V;��21x��#X����Rlam ���9��̸�vꏉ��iN-��-�I��Y�MpaŤ݊	԰�g�=���͛�1�տ�k�%�G�i�Wv�0'���&�#{�$�dP�)������G�Qy�s|�X�V��^�Kh�M�)�f&�#�F�J��مӬ���i�8��R*i1L��Q�����pk_gR��\���3� ���%�6�9�x�,��β���3�� FÊl	��X,ȑTȚ���}�۫<Zsl�o,�8� �`T�qW�T��u���>��i�x e�<��:7�΀�����2������+W_�!�����{�+�č���ډ���8���Z�	6�M������-��u��c�g#�[P�����?@���<��N��)tb�y���|����_E��J�弇�ߞA|B� �rn�I�B����yo�E0D�[ q�B ��6@N�"��ohih$�M�(v����)(�n��yja	��%��~/oQҶc&��_���� 9p�iL@�k���ҸW ��
v��<84xp5����F�,������,�W[~¿�y�뾓S~~�{���[���L�4c%�W˭AO0�=��׽��1�
H�n$�<���C�璍��ń.�hM��&r��.,�'��o��[�YoZ���v�0���H���������H+#p���.��o�'r����Go4��O����5�@���&͏u���`��K
��kՄAz��m�!�!9r6 z��[�t?o�|;�.�ÁP��\
�e>����q%=F���<L[�O�jv�>Q���m��BF�%�P��_4@�ٕ�Sc	G҉��L���2�Es�ýy��U���W��/�'�<�;Y�c%f��7X1����i��	v3M*���L	�*�c�gt;��q}��KC����6:�T:'~�-�ƻ��̃@�妷g5!d?,T	;1�n�N��u�H����!�n��5W<d�����M������1��?ÿMTo|�M��[��~��K��0s���C�'�pD��'
��:z�>�r"��D:O�e�>0��c�xQ�6��Q�I�
�md�g���Oƺ@H��4ogi�~[�����?	�_X#�u/��r���d��������>��Û�ᘚr���t|f:�Orf�'���=V����j*k��E�#;Y
�"���s�%�p���f�2gڝ^�7^bD�W���X�|���� RLO 9�ނ�('���B�[QO�A�>�����) "��$��}}����Y��ح��v�I~�^��>�C'��4�5v��*0~휌�}�K�8�OO��Z���h��m��s�<�a�,������bj�
c��j�Z�KG�����e����m_��P��)�I2h�� >e)u��`$�9�6��+�%����!ɺ�-.�®۞�	��;�hbؙ����y�4�Xd�h6�۝]���,]����P�o������Y��!���w���?P~b_%��M��C4ڸ@���t��9*_M
b5���%�k��������X���5���K)n{J�n@�6pi!Æ���������Uڟ7s?�K��0-��H �����=�U�8m������ً��p�@ ����o}VA��x��5�i�!�E�V�KP���wx"���ء�u���Lwc��q���n�>�OZlm��Z '�h���J�,n�!��k�Уv���
˴�7#�m� ��UT�s�r<D�U�nbGA�`��d_�j�����P�(�{u�y�6�����he��������1.Q�Rdkup�:���{M3�}QJ'I�Ǿ<�&�U�Rh(gq�}�kYɴ7|(����ק���q��D����$׀�y�y�U��������}7#>�H���@��U��b��Ϟ�Ԫ�S�Ur5�h,�F!�t��q�w������S��Uh4�Γ�L*)�2b�θ��;/KҼ�+�ߵ����)Y��g)�E�n������ff����񦙞�x�Wf�Ҁ8gQ���4V���t�?H��y羞7���i�#��f�y�x����,��
�q��|��ly��ˁa�mNKa��?T��]^�Q��E`R&�rt���f��~˴m�6S�w��ْ��%bzv�{�P�UV�S��Н�n�li긅~�8��?3���^/�<�����|�X�T�o�j��@2GH�ᄎ ��k֭�~������\�VT�����UKF�9����Al+&e����'%<>�!Q:�Y��C>�8ԅ�/F�a۷	k�s!��֚�wx�5V�zvo��������$hS��w�V��-Q����=����N���@���21�?�4L����;�b^���+o*Kf3'.ֲΒ�#�a6"\nl>�!��R��-�*��M�CC�L)���m�<�y���B3U���ADS�}mM�c5)w�}Z�����N.�'Ҙ��_bN,S�DW�s�V.Gn��޽!u7�GC�v��~�
�#e	�8��oՃ�͙����I�N��ԕ*�a�U��Ի�_K�}p���*�(��ט��d�-�zH����)lz���������~៑�C�(q���n�4�>di�c[X榃d�*1���\�j���)2T��S��9۩�ME��p�����Aq: 9���d�|M�X@h�խi���,s.L�(B�c���<HB�XS{� a(���a�ϛ2�~��>�n����2�A[	5����t�v�t�w���6��>p=(�6���R�|�JT������"c���h��VJ�7��嬡PJ��];��O�����c�l?$�^T�5�q�>!�p�Z���v��t�cU$�H/����T���I��N�&[���\���bY��_���$��
����5V_n)A� �r�5�nPۓ?Yx�����:7`��[m�d�/�<�R�:~�w��ψn�9ρ���.)9_�i�tG������`�I�u6�G�j۾!Š�Ъګ���#6�,q�ö��I�����	l�/Mt˝�f�!3�ɘ�Ql������l"�%�'�
��Zt&����t}�XIYSc�ӕ�ʽ0V����a�U�+F�1