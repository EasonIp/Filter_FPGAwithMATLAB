��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_ �c��2)����$�a<��d�6�q��tӏ�ˡ\s�$�L���Ÿ|^*��g�@U�*2�X���2��^�:9��D<��;�h��É}����a$;��몬g��>��W��iv���o�ăN�G\\�[�4�������W4xl��0�;O���V^��@��l5f+��\�&�7F�CqϮ�Y"�� C�T���/��Ƹg"���l ����~G�_y�kIe�+E�9�>Ǹ=�oWS�|���WV��P����������L��΋I2�G�r	y�i&�l��vЦ5�o�#����T�WrkV#��+�ڛ����C��ɀeG31>�����k�\�%�̶�@J�%A-�@�'2�}�0�΋ha���RN;zy�Q}N��5Z��}L���Z��¼�1<}M�����g�) $�8��Ρ�g���}E����G�@).�b���L��<�1�~:�~"�S��Y�p*-��^(Yj�����k��=98VK�ϲ�=�Zhy��� �#��_���c���~���YƯXrh"� Sao�%��Ƭ�;���cE��:�<:���6��E����Mr`2C���L�g.�T�"/)(dAX �B\\�xG�� ����	��r=�ى��x�⿐�z{�&��!�$�ȠC���}���?pEp�����p���р�e��Tu�M�@(���v6�ɥ.D�{(��Ķ)B0�h.ˢ�ا--��I�OtQ��I�ǧ�b:�ot����'�� �AvY��ɲ��c�Q��h�v�z�Fo�6$�ǧA��h�;�X��?F�4�E���j���X�Qd�i�� �C���¤T&=Ò�z#������z?��:�]q����k��V���=cT 1���A�Ƌ敬��%���f�@_��Gj������?�B�*n�Z�g�:�j�[`�aG&�L�q�O-�0�\���в� 9�n��_�y�ǷE;R�),���>���ɣ�v���H#���>Z�1�)ݝ���9�`q1�y��Ȭ��|� -
��E�k���Z�<��p�|��LD,bۯ��"��dd�t�����r.�]�S�~�ښ��Cx�\��Ե�N�?��Ώ��W���p�>!_Q���A%��x��E���hl�Tfap��W���o���z�1=L��V> �m��ZM�����L��"�K�+�� �~�qWƒHP�fT��	n7��3~��3G� }�7���˪E[�u��
lti���s�?�2���{�C�J�&�l�G��U�n�F�@�A�>
n_����3�	䯅��g�l��VB���2�7o�}3�=!bC�(z����F�F^,1�6ݒ���vU�OU��k��F���Rl,��S�&����Z�{�8m;�D��J�{���Q0�9��E>���_�"s_!Q�|�n¯�j��ރ�x�;N��^�.���q�S��l���/�l҉���3��0�T�!#f�py=)�&9�ez���-4M��|�<�;�2R\���BL�5 }F8e�<c7hy'��9b!\s�9Ƕ�M1�Kc8��/��EH�ε��a�swSª]���7]��T�0��R����e�Xt�:`���,4�J�X�B'���m/*RA��\c9 "lW��m�/�:�1��� v�F��$����@تN���aE�?��%Ό�s��%���t���W�8jR�0��|�Y!?*O�~�rA�PH&z�z���,L�vrӳ�q�z\�����+���"��>��Ѻ��`�r���z�w"t\��ֿ�&����N)���U�^jh�X(��W#�_�.�E�R�i42�o1v��*&B��pspH�\W,[)@�E�Jl&�1`߹����c,呎��5�+��P>�.:�@�Wz�ߐ_EB@�^��#����:]��y_�&W;�a�N�	'F��;ڼYL�nP_3+���'�c����������='�yrNQ��x2P�|b�~�l��%A�K��F�K�%��VmzK��I9%ȭ���J]V/>�j�1��5�h�**�8?���GF\�JG�Oe_ w��C^��쯭�U10M|�t�|��������h�<˿�y�!�ӿ(|oJzH�8�������M3�m��$a����g��t�������O+"dՁ�QP;t��}����m����d���q��hu�e����o�'7 ��a)f�����/M���j\m#'�( ��)��N�y�ݢi}sR��m�Iht���%�P�|[�<z�n�1Ђ�*&��G�3UM4d��[񳇧����ջk
].J-��W����A��	�m�Er�:�'U ���Co��>B���J'2�!gM�q��`�8�kz�\������]��b�Oٝ5��kr�_u$ �t�Z�v�<�΄�J��W��:]P9Z���kR�C�x�_dPtg}r���b��!=��+�J0ِXJ9�ެ������k62-1�8���X�1AX�@���-	U&>D?m6\�c��ԫ[��j	9q��Ӑ�y�2�pS\0�_(1ZS����c������7E�d��0cec�,�������
׌{���@(=��OP�M��T��D�&��j������K��4_�X�=�j����<���ݢ�BJT��}�?�SW����ߕP��R�,i҈0�7�U���b��_l���M�oĉ��:�h���B9��}��A�TQ���v�K���&��9Ez_��͌�]z�ɯ����d�y�M�8u��N�0_�3	��j<��X2�x�K���̶ �1~�em���*:���|	����+����K}ʡ�`����/'��v�52�V�8�'>N�9���-S@���������U��� �J�����?٧��T0@���~�~BUɛ,%��r��1V�ذ"�%[��#��Aldx��r�Q>j޻5nG��꿊7|gPs*a���_GZ��Nr��cĞ�'vz] ��b*��y�5�o�Iϲ�����X���%M4�$6X�	LY��6��)�����m�a���=�� �/�݆I�'��S'K�O�N�j;ŭ�/.�9Wc:��I�r7j�l1�qm�:j�k7��b��S���,�C��P8[�����?���v�"�!��Ļ�<6QQ�d�K�VO�ƀ�����|�k����h��|���{Jт�xtaP5�R �MJ�Tc��Ŵ�[��B?�@.��U�{uL��d�����MR>Ԅ��~�J�zO%�UW�w�A���$$�PCl<"�C��Y�yG�]�CS�S1��0��hT�=%�������)]r	�:b6�i��'����a�=�!��N�/ޞ	��uJ��1�qm��RO�ӆ��L�3Y��Qn�O�	��nh̿+/�z������\<����s�h}P��p�L@����ˡb�c���h��Ie�	��$����#>������8}���8[!-_�"` �L���w@b��"���c�f���� �?+N��>�B�k��B�_������Ê#}��@Yyz�f���8F�`�$v�6�[f�T���ȅ�H�,�Hv
��y��|	���R��6>�A'���C0Nn�|�O�75ICrB3R(�tGGNQ���s2�}V9Q��\����!�D�In�9�\�\�k߀�攖M�E� O�S���_p�˖�(�~Q��L�K�5n���}d�#���tŃ�����$6��܃Ԫ��2g�ﾻD��?���I�!	��a'�*��In&y=�A��K1X�J�g�e����8a�I���r?��V9a��@)ZuM,\Q�Y��i���Zr������-������x��hS)����J?�C,2���y�PQy�Pv�u�*�u��.g��IٓV]w5��(�������l��
�o�N3���2KU�͝�0��z��M�g������V�6�R]^��9�t���?ظ0��f�A�kH���рآ���D�&Z�u�u�Ob\K�I3k�'�����ˁ�)���^��y6'����'�^�lr!��Y.�!:�=�%��c(�4��,��(>ՠ��8�������r�z�Ʊ�'��'45�;������XFEIr�!Jୱ� pI����"���*��\���d�=��]���t%��缧 �����"x�E>�ko���"�J�`�d0|yS)�v��r4;:uc"�BS`������%,����[u�_l�z����
�S�����%u�9hT�ɖɴ9�F࿺)�:��(��m�w���*Y��@��T��H:��SPв':Iv7�L��W���/dS@��R�}f�����u/�tȔ\�FF��X-Z����������I&vM`��<r: �����FA����t��)R��L�T�K�����Ђ��"���M��!l���8���m������`yr�jq��?�7'����S!�sX �U=:g?wr;�r��=`XN�'4F��c�ɫ�C}P���o� ��#��}����`˥�[��taӞA������ƪт�Y!c�r�K������ҟ�`u�'k*���7�q!~�v���]�Ǫ"�?�����	�5����2A^�sTA�?��F�#�W���E�8i���x�NDr"���J��ݭNXy��d>@�+ǋ��/�:�.�.�mD�����8�"0JB �~=?9^�����B5��b�X;�Z�'<�N|m]m{Ь!m�����H�MĻ3��~4��9�Ջ\Q@��������R.$d��t_���>X����U@B�wNq��$����(���-��H'��KW�c*EZ��e�Jf�+1�.uݫ$�l��P;��[SD�~�[��� ���_�**��։��O؟��e(��p�[
"L�) ���J�襪����}������$O�{���	�l���J^F�"(Yy!/T�vy��s~�âC���}������B�Չ�3���F7�{�)z%9r��5$��;F!��b��1�:��0~��ߋb;q�*Vo>�@�HJdw�po�ȓ*�v�N^���:�����iMō�J�H@��M�$Ra��9l���oM�|ye~�~�,��s��k�	kFҷ�t>�NW�t=���f�2\w'�`ƏRfϑ��<N�BqZF�Y�k��Z�v<e��
����\_�B�����?��f����-��2+^Fֳ�[]�V|+�T��.�+���'����
~x���Ps���u����e|�CM��G ��*o�N�~��l��&�S��]�!���~��#�&�	�;'�lڧ��9�&���S,�bFY��;hbU*�`>t{5�;U�h�(-��$���=���l�C��V�@.����\	1���5'au���m���v�M"���D[�u����?7��P�ҩFx	��&Y�.x����'mCx���<��cO�#i�/ɇ��y_���j�����!�JI��w�RJ"���������T��,�=�����u���#԰݈�fjDt&G*М�p��%�*-d�����%TL�XjY���a�?
�
��f���3<S�EM�E�m�_��a~�"�f�V;D
=��Ճ!�H�I�����_{0ІX� M�:����8+<�y��$ۛp�%�G�n��f��yz�8c}��.��&Ɛ�q��n�A�ǰ�T"O��m�{��C�O5�]d��<