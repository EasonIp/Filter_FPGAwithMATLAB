��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$���v�4y�ߐ�΃����0����n:�4Kf|̔�\.��K�#&�7�W�z϶i��wD��0���f�6�Qv䉅��XL����+�OZwv#؆�.U���)`����n���Q'�
�Y8��-,�(:���.E�Q��bN�^O�
�g|�W Q>E�r���]bg���9�ዊ�����u�2y3�n��Z]r��K�&FU��ϝ"Ї �P�X�����?Oj���`F#5��8��h�+�W�gh�"IJl��Dz&�J�FX��ZI1��>�--注��V� ^���Q5�Pqm7i;��ޱ�t�u����]x�t�J�[}���kt������_�0b���'�R�rΓ��}� �!�VP�?��t^Y�f\I��'I�1&��I�\��m�S�_�h�t��M�� e�p0"���A�0���>CJ*�G��P	C�m�T��"��X䢎��w{%���~}�,Z'�E����{������v��;v�E?}����>�bR�h�D�Ro[���7h�b�t��8Wz�~�|\��Gה��G�;����
|G�����lz��7��L�sY�R�&q��u��|��ȺM<b����7f�Y�A���ve
��&�J�'��I���6ēb<�bɆ)ɐ��j&o�����Q���M'��/���&������e�b����a��º�SQwH����>l[.M����?��
ʼ�π���c�ND�ծ",<-`�=��8œ7fj�){��mS��QI������HPQ���D�4����v��$�P�ӓ� ��EVL`����)����i��l?��zU�|/�_Ճ�4��W�7������%"�Vm�'mV��.}g��8��J�-5z���a�=!_(u7岻�n���U�=�3��7�M������l���~���%~��Yw��w>�>�+���ϵ	u������Z�J����𦛆�=��x�Ϫ�������]ም�5h�8�����A�S�K��G�)<���;�� �[{�~�].0���!i���I:!K�NW8A�B���T��)pu�^�1l�����(����~Y�����A��-�U���.$z~���d$�9tRփ&�"B�$H�� i���-l�h�I�}
h�EχlM;��|���HzJ�K֓5P����3����Z,�����&�Eɭ��>`Xa#K[a�ֳ��)��^)3d90Tn�~v�p��S54������H''�����:3�?���خ�J�{��|������VBUo1Aga�oBZU�; =��4�ŕ�O?�Бj15�Ƣ�z����D!�=6��Eǟߦ��{~��ȩk�x�x,}͡�AY�S���e���[�����ˌ�t(�/��-h�יH��H�c��b����8�'/&#����LG��hxxG����qK-�{
�ޔH�Fd�$C�ux��	g��|g{����N#�-��xmكfm�V@�<���{��N���6���B} �(��ʅ��=I_�(_v-0AR1S~N��P�;^�2x~�|o^��*ߵ"�����R�Xb������/t)C���&Ɔ҅��a��y֨i�c�r�K"��s!��3�U�����������i�>k��ubkS��A�����,Y�u`;B�9�v�hN�}����������6�Հިz��vd��m��'���(G��5�w�̯Ʉ�b�p�V� ��8&$�����a_fg�")0r7�����~p ;g!���5��� ��B(⅄��������7vs�*GfS�+ب��+4���H�$��O��/*�������=�f��;�l���F���T�gh�����⠺"�h�8��j���*��LX<��pO*�i��L��C~�ח�|BGP��(4
���\�P����Y��P?�Y���e.��c;�3����̏���о�*!���7��9��1`�JI��0��.3
�&���`��-�m�4��Nט��\�m�慢��c����W�-%�_�u�*e�W��XI�����L�BB��*���x���:xŤ;F+D�p��N�ZB��g++[R2����B�h���=����0��~b���	��Z�0��^@=-�!��8���M`��Ȝeb����l�_�yFיE�^�jP1�vDkp?D�Dr���Xgp�Tr-���:J5~kď|Q�j���%X[�c郾�O����l�o�1����d�G��v�E(j�ت�~d!����z��T�6˙�Ι �ڜ?�l��ɍ��R��s��=���F�6���gq/�Y�0����Aڠ�������V�A_(G8Si����;o@y2S����CH�Ћ�*�a��}�zY���ZM��8L�R���N�5,�'�'������r&���d�>q��I!y-j��-L7ܷ-�1�5�-w!��
WΗD�4n�`^B#�X�x@˞]S��q�V�폩n�H6�Avx���~e���A�qp�u�۬7�2o�h�ʍ��}��M�1�o�� ��x��l���k5wE�ؒ�*L��9k �����[���H�Xf�D���J���ڃ�\꛼��@��7]$�����fۡ��E�Z����#�Ko���6E��i�I/`3�X�~XD�����ul��?z�?Z��
�h�f��{�]�v��P3���_�zȊJ� u���
.P�J#zYXV��б۾�$F�b�f��k�gjL�ƺ��ǚj���8�2C�&!����a��b��گ��?س�?����p$��KW�`�����O9�zj{@�7�@��݇i��ŐLn� �,���䂩�
�=,1����4����ſ�11���������;��b�� ]��0{*N��%3���؊!���f݇V���^����v~�|��83�����]2$�S�f�+���&����\o =�CG�*}W��)�<l5��� �H�I���9��օN9˧Hइw-�ҽ�Eȱ6�-���������t!���l�_�� ٥
��Y�tb�C���<~��z�&�E8L �d	�����[\�����6G���V͘�LH�`��+8Sl�z���,f.��7����	l�Ne~���j:jj���
���P%�;g��$��G��� *J1���Rk�mD@���ܳ��ǩ"�&�!��`�a��M�>����	7��SC9�d
&�6�gT�I2>Ʌl�>��l������1�~�(a%��!�Ibeb#��RQ�[�>u\���y�Tܚ�
`����y�m)�a�Q󝓷o����J��j*.`ynTPC��пHfC���3,ǻ���&��?ʔ����r�j�6g+hl��[���ͮJ
t�v�8�[xW��2,�7	��IA�n���ej��B�� ��D난��S� �@��Y�F���F�����'c᰾����:��ͨ������ &*���1x�6B�φr��IN Kd�2ӭ,"s�����z�P0�#	8�a�d}�,D��o�.3�������۽��|��R�ƪ�[F)Hg��7/�6́�L;�{�j �F./���h<�Uw;x>�w���C����.�W����J��cP�t1�:��VUtGз�P�~Bd�>j$��
~�',Y2%�6*H���ևc�ڋ�|uWe2hV��m�DTV�rYxr�-�l><��k����4]*�5Y�A��O��|㮳QL�֟��rY��S)��[�Z�E��Lc�g����h��7��p�������˅�E	�J?��-��C~_�ꭅŰypS�(���~�
� ���"q��FIj-bӣ��WeHt��'��}����:边 �M�*�֢4ybj�%pw�Zf��Y�˲�����ߘ��h�8o0v"%"���!��եu�'������p��I�_�g��mĉU�%�s�B���[qD��K�5!��W"�����2�8��&�yBo��`�'���gg"I^�R���gr=ؕ*R�2��@%X�؃�M8��C��Jb"H�ӧؖ�t�1�Շ!�7�C��?������<�74����Mn�I�
���8���z���[f΄�eu�(<���U�iP�c���1ʩ��KqD&���e��w���n� ���9�����B�p:ʋb?�Cz��������-�����{ud�^��.��_���M�pl�AJ7{��
��������"ǳ�=m	W���2n/�唙�x{Ol���z�:�_�Mr�t/��O�б9B� �m�2��si�:��E�Pzf���	�Bwd��t�̚bݽBB�ԡi�.���؋��<�ɺV�	_T�D1JlU�1�(H��T�=Q�1�!����x������1�J��2SB�u���ʿ!h� �_Lt��J��Ŭ��tV�����1��-3-��h).�C-C��o�M]��o���!PC��GR]JS�?���,���K�Tqm�E{�%|�%���! ��?�ݩ��J�$�2������t�}Wm�4� a�	o6��UX�j��z�ooʻhRą��w���0}3� 2R�ԅ"��"⥑C��%��ͧe�r�:B���g|��\���U�	�p���i�K�՛�KM��>����tN�%�t�`���;GJ��s,b�4Nٿ����t%���RZ�f���Qd뮘_�w�ۿyL����hF�;3r�k㞞/�`�%�=CW
�o<}b���I�Ƣ{ܨ���Wk��0�'O��]�x��#}���<�)bR��p�ے�����:#��l�12k5*ۧ���Ȝ:KWP�.K(�-�I��i�f��
����y:VEq�~=�i�K��7��)�U$��5�]�y��2 ���e�I�������M.��+���n�_Oj) PB�����=̠��`	!�;Jj@[o*�|�LJb����^:Ӆ0IpంOn�C? ���U_��7���u׿���8u�9,�a��̄��f���.�T+7�~<���0x��U���ug��n��#��;���ҿ8��P�+0�ґ#�D��l����Ww/��i�?tW���T��9�}d��H�AH�m ZB�UGIJZ�'ֺ�����`��+o��S�h�=���k\� ���'�;RR�B��&ԟ����Eʝ� ��Me,�M���nn�B"��|����45��0�I�����  ��F&�/%�`��%�+��J]t�卷�v�x���sE��1܀ ��fp2_��LQ�1��]��D��>H�H�wKJ=��=���p�˟�$ԃB8A䈙�5�E���ksk9'au�N~��g��� x�jh�Z�?a-����-#]���1Э�Ţ�ߴQ�i{"�-]�>Ϲ��ٶ8��^|�3~��
Y��! ��m�>�pL4��HF�\]���*9i�b�n�B`pGk�K�Yڙ���)��/fW��sF�v���3�?	6����V��J�V�+�F��}`f;��M�Jkaw��%�>��Q3=��vj,��M���5^k�O2�gMl�Ҡ��Mͮ���73zlt�E�w�*ז
|v�qH5�U��䨛��J�	�����w��I�pə�tR�	�`\�����c�b��=΋c����QV29�>�~Нҕ-���.E�<21��!�y� 崬����.p��ۖ�|DZ����Hy��Y�"2��b^���
C�+�����sm5�àx�VP���5���d*�9�-���MN�n� �U!�z+�/��%�,�D�r3�n��',6;ˠ���$�K�t��ۇ�^��@3@���l�34��n+�e�8P���Ņ��E�R7���yD�ݮ�e>�h[%_�丵��y:���K�Е�-��<ON�N���4	����\į�۲�e��ɕ /¯_LŴ� JG�y�bLW�ܽ�����Ĺ[���g@^(�)a�a<�[��KP��5�fcy���'	��=*tM���Boic��4��΅v��_n���C'>Kf������r�0�1�d7 l3E{\��4 �
��06�
���&���c1�Dq�)Rj�"aI�?
2I�~z'��d�j����K���;��q��t�R񱽙U�"�x[R`�!�.�Wm����Q�~�$�xT^wa�,��mU0pg \�/�=B�R�� ��e�'^x�+Ij�m�F��}��4��a�NOg�q1�![�֩ew�Y���»�U,1����MK���r1���3�ϟ:qWA��9e_[�lW��EͶ��2�`1g�G���Y�t�;0�s�>�v5��|�"yג�.�d���"�+�l#B4[M&;�ܾw�Un�������n�RCy�4��[��Nv�A����C��D5�Ò�mO� #I`L�*-YGz�E6�qe�X�X8!���hg��У�)�&8��{��e���:���]�0��=�}E��?u�F@c��U������_ƃ�8�`����#GŐ�B�vV��#f�Ȃ���>�u�_�n�}�+e�F�
�i�c��ǊჟC�����⠛��UtO��ʛ���D��Ƚ�e��<���/�y���MP
��,��|5KW��[!���O�R�pYBH_Ӆ�a`�V�«{���ū�%Q�����ƈZ[���������)W�V&�9�ס
Fb�9�(�9��HqF�ܨf�������t�{U���k����h�7���m@
FGc�r0B�#�~J ���le�#S�h������Sl�%О�S�����C�~��kK��c� �<����`1�`�D݇.�L��=q�la!�f�r�ǒ�g�k�/BN���کs~��_z�%����"ȳ4�ү�0�k{�*��&��B�a�zW�`��2R�y�[#`w<ٰ�f#�Bm6Qg>X��7����+��Rs_�
"OXT.��D
�D5j��<��P��$��4�^��g@�o0��t��B��'�p�@)�U�&�"+\�3|��V^Exl�N`�2���0(�R�O��/=�opv�yN	We���-�-�1�X�	t��A��lsq|W�R���SL
�!N��������s�؉�掫�#6|��:K�H�)a��o���A��a*23��$���f��Oj�f�ѿ?�,Qt=W�L��
$?JR����WP!��'�B���ch�t��������3o��G�=�������"chˡ=������E�����m�a%�h��hl�*����-�W�D�gp��kwPp#�o=�U�I$����͇�wqp~9wJ �~�<�k�p{P����y��E���#�8����5[���&�2��%a�釆MStE�[�m��l��鱓�0�Xvܼ��4T�p�>Bl���G���T>[��-���gJ��q��Tf¶�w ��D@��پ��Sc�Y&t�I<�Ƚ�;M�_.�.�~�;��+Ҭ�������|�F$ȥ�.������u�%Ow=�'�
;$YXvXMK6ʖ��%<�X�<��md�W
x�����\!��-w~��m��0���YN6��04	���S��p��y'��%c,�S�:[�\�({��2�y������H��^��u�� 9�"�����)8�6�rzԻH�i���ƽY:�[_�� �{�;0���#uL��x�ԵD�A�S�Od#���P��8�W�g!�N�I�"�a�l� ��c��詹ApM��)�ɒ��z���r9�����s �A�-�b d���2H^T��$�ݥ`�]��OJ|�6��!'Ȣ�����u<��`��:�~����f���B��,!�0��mgAXm�\��vpO�=$���p��+����n���d�o��}_:���\������j���8���XC����19�:��#A%J{�Ez�<IҰ/~(yպ庥��խ�q%և��6��?Q'���{����'�3��08�z��Ƙ����d������@HK����<q�Q�ĚA������qv�*r���n�a���|�|ݬwl�߳2��ގ�[�Ô
�7�y�deN!�*G���OR����/pӸ��e�"m�I
�q���4����y߁L-R���ñmb�Z��������u�|��"�Vnӹ��A�Za��NB�%������t"BO9o����G�3Q�q�Sݮ��^�D~�1��'� 	�S��w`�maYG�o����	L]���"��*�n�߃��xG�XU"����4����:��t���W�4��E�-����꺭i�`�-�����o�*�a�9�� =�?����D�p����5�QF"ӧH]�X�#�����p/57G2�1�#9o��S���vL�٭)�ۻ����TO�$4��_ܿg�俊���n���%璉*8]��ۛT��uN+H;�J�Ԉ�A�]���Y�U�%C��99����?���M�Q��C$F�<�vnd�2�k:����~n;����f���]�( �V/GC���Y��h������	�	]�a���!�A��F�[E�L��=E�][��F����iϰ�v^���Mk�qsc�y/���֞�qTS����MPhz����Dn94�t�b����
����-S�6���%�
�X9���J��:Ue�s8�؉��8;P��Ä�A=w=���13�_�V(x7*��kX�W�43[;����ڳ��8��'vJ�+�|��k<!��z�	�K!_Ժ(ěw|ِ���F��_��q�J�h���5����!��Q��@��%'��4�9�98���fy��O<n�� ���g�kc���㔶���+�叚?a�1�߷~�|%�ُ�J�
��q�	�}Ų^X�@���H����f_�w��{L�s�{���?Չ�� 3�.�a
�HB�Rt��Z�6�
I;q3���i�x�6�Cْo����H$�����o?^��4l?���� ��<f�z�>�L��������X�f;u S�>���������r����d�q�q�� ���#w�Fp�Gx�.�O�6jt�x?r৊.Xʙ֋���5��c=Ա�hKi+��1�B��\PϽ:k#xތ�[��Pk�Q�Yީ���2��%,�-J�~�[}�q%�l���dQ�ۜ��7I�\U�4������'P�܌@0�n�B�7�wI>ZؐZO3"�v=�	��l��{�6L�f<r�DSGwWŜ���G��B�L����4~8]"(Òc��|��^k�5l���C��՘�慨R�J����N��]=���8�qg'O�!�����#�����O����)����Z/�n�vB|cU�a���rsI��f�{d�G�|ma�xƭXp��B_�a��_�}MFp��O�\1wO�ٖ�H
��Z#'�3����qB��8A�`�✻<O)�n�������)��e�����s��(�9� z{������x��i�]����X3r��Ӂ�G-��/>Q�i��&���a�H�6z�wi��Yv���M�u� RJ��T��T�X����T�r���N���.u?�M��V8wǤ���I|Y�=��>Z�C:��}?!�s�֝�Ϣ�����y�ΰ�>&ջ�8������.�O��Q����~ �����V�k���Ԧ��>��U�5G��\(Q���$o͕���5��@ z c\q���ݤ���|�&;UU���CK�"I�@��x`��0���u��-�� �]��>_3��l
���Q��/9�&�Y�����v��s�}�>ǣ���vU��'��o�>h��<[���I��&Dv��a�r�b��Tr�_Nc�K��j�"�^A�s��jO�,�X0��Z��L��Ĕ�z�PөN�S|,�p`ڛY��{aN�����m�pJ�ctM����X��M�fȶ�TLdK3�~$1H}���z;�\���wk?h��iI	m���`%�G�5��{�+X6�1i�4����q@�j@nH��{d\EAOs�b�z��� Kk��A�\��o���N�J�]|��<�Uף�g�ѹI��^־؆��H�+Y�2��Q5P�H'#|�V!I�_��Wu �����hX�Ց��1N������Ę#��r�:����MNl�Af��"�`�E}У+�v��0�X��&�m�$��8;RE7o�+��S�~cICf�Wt-]�[���uj%�n�
N?U�85� ��Q$~i�iN��Mn������zU. � �t�m��2Q	&�\�W�b�ۡx+���̦OǼzLK'!��"��u�1zľ@�Gy�hej~�\�y��'�u��[D�*-1��f�k�*�N��5eځq5��
�#]�[�R=�D_�B��ꈲ��̳���eDm��z�����@y�<�;3��39�h(�~��?E>�<E]Ԛ��Lӵ���ьm��L�������r�(����]�O�P��E&fAW������T�*�i2#���`�^�ʡj��Tn^�d���R0SЦae����i�È����F�S����Q�Hȓ�C�j�&]4�,Q	��N.���������0��\⤌.\a9yH��r<Oס_J<K�ܔ!���y�:T�CXq�4d�C��2i���p1;��7׆�ZH�fL��Y��*� &@���&���	!�R���zWD����#osyI��U����/ ā�b8_o�}� >TҿP�MH�*�����5��i��G��!Z��\Z �K��8ݦ���I7���l���ɅC#{��F�@�R����V}��u�Vo�t���[��TZ�4�#��L�� �?2��2��[�
���+�F?b��݆�`�g����V��p��L��#ش�t��J1f�cG8$��ѣ(5����"�O>�#6.B��i�?�C4�����P��$y��X��XjeÉ�<���B���=��1!)Kz�F4g�S�;Gx�|�hDո��C0��mۦ��������jrr5HzZnn?��4��j�؄�O�Ԯ�UR͆���^��v��������t�7�Z���#���U@��Z�ڇ��I�#e~�����MO�g����N�v�$M��)z]��EsOquY��H����X��!�.�J0���`d<�����k��Ď&U��v����Q��������I��o��~��eW��xxM�^�&�9���^<��`=���~G���@����D	�O�q����.s\ɫL�����@э��W)��'�R�"|��K��o;�oH�(�[M�)@���EVݺ�L2�����'A�Z��M|�ˆs�]�k�q���e	�X	���!��������v���p���c�u�$����Dv��J��[1*U&��>���@KU�s1E3�q ?�>��pP�/k\
���; )k�Qt;9�-��חч��R�ۥ�������u�L@�hX]�x)�k� �QYj]���>�v �2��ģ�)D�G^$F���g����!��)���BLqxDU�m{����%�b���,M�~��YMF�_�tlM���0x�Jp[A_�S|s$���ʭ�F*����h{{��?���d�kIt=��sD�J%}�xGt*}�� ����HM�;k�O	)Qz�0��>n���ŕ���C:���U���+2 ��U?�ue��A9d�rUZ��`�b�የN��d������𨨬nsß��/�I�4�j��/���w7�B���uZ����c��u�b�d�a�o��G��w2q�y�c�w't�bT5����ZBG�PT"���<��VmQz!B	1�k�{�2�gE4��H��0B_�1������<B/j���p�wKֻ�`�n����#!�����^H�/�&Y{��ZE��h��W�ױS.
��+a���)C�a�ǐzR�����o1X�Y�M���W�z�d�4}.�6�P���Y/"����2�,�`c],*� �BJP��?(��N�2��=g�mj��V��[�k5O]&�{�'���J�_LZI�����	��P�*utr��C!�
X�2�.��]��%����2Fu�A�ZG�)��������̲���P��k�$�493��Yk�9ףT�Q]J�@0j���ߍt���`ꡢw�I^���s�o�4���6D���HE]
��A;�Bř�tv{�m࿰�ūI+{N��g(yB�w{G��O]��*���}9u�����Xv����x���?$��lx2��ߜ0�sԮ��*|����������s5X��zI.���֔P6����U��.�c�o�RA�Kxm�L�f�x>��9�=��>f�sW̨W����a��V�\��2R@�(�d��8."|;�5
[zٳ��� �E���D��"xj*�/�a����m��͕u2-|Xc���zg���a-�Q�G��S���'��q�6��)�8A��`�]�|3L#����Wt�ao�Y׹�g�qN��G�>{���4�9h��%�?A�Τ�0��0��艺�ȏ�O�����v�����Hf�O���m��S������Uࡪ紒�6��dۙ���F�K�ui���Xv1���9��N���y��=��_��+ �V��a���-T�z��qm�j���k��i��Ֆj���.��)���_��]���T%	��G�����R$�7���4}כ{�ڜ�t�T�*N13�.�l�N�.�����r�t/�Su��#R��Ī`�X+���<�I8��&����8�v�l���ʗ[bZq�� �64x�K�������&�o)M���Iǥ%0?����%KtN�[<,Ö���=!BOy{uuҪh�eN�ha:z����M�˘B԰�ޢ�քz�d�H�<��ٚ��mo���Bj>xo�Y��_S�2�������Y�['���#��a9�Ct�#w`̤�
��|���P��0Ir��j���5d�L�`�Pj� ��~�4�ַ����z��j;�@5Z�H�2`���Vܫ	n<e���s~�o�_g�b9.�O�Cы5�滪>=}��P噬ꛂ�I}�!��Åi4���%c��f.�ޝytx�rR�+eɡ�ɱ�w¢>�wu5�(d۽W��N�E�"ȁTk!H
�>H�J1�q�Y?%sOQ�)U^�tAs��T�q$׈��x����SV�0W���h�W�����7K�%�����0���~5A�����â�C�eP��!�F�%bW���&�I�)��Dt�&��'�~�ǻn���Z ƏW�+f�Nllv�_e	�T/Q�9�N���n�&�*�N 
Uæ[��'�ש��^c�j�%�j�ھ_Yv��qL`��MHP��>=�:�K!-�_�nh�H2���a�̬(J.�ʬ�W�i!Q�V{��rp�(t��s ,���;�<�2��؂��{pr�\zW��VG���	���;���no"f��p�g�
�6��M?9D���t��eH��?�f��]��:'��P�Lb��8�g�-���6[<z:�?t��#�~-ڮӆ�>�N��޽{���'𢹓)�(iӻ**�e+ܽ Ptw�n�	y���,�F&�eJ��%��π�������C�7x�0�.'V#k���|������,2g��T��h�ږA�ΓhRG��q�G����Z0o�2��U�+\��q�����Mh�7X�D^�H��Ȏ��23���A�Q�<��ʿ�4�������CV&�����Cՠ������W뢡�<��-EW��R�}�`����v��B���%1��BS@��j�d�
����y��������56s��5*9��?? a{+��b37�e�9�G��EK-�L!6�K��׵S�}����@��.ɸ�LWop�-S�7#w���Ry	,���L�q�&f��e{�� �\����U�a��k{��ea�إ�������=$�@������_Qn�Z�Ky�a��>[�8�b���5�Oq#ۉ�R%�.�_��[�|1������Ť�X�*K���of�3j?7J-�#�h)�ȃY~����5���Z�e�&W� [흌ks�s��$�f��"�r�cj_	��i-r����V��s���$�.�{Z�?_��E-����|ʵ��P�6����8�h��dh��H��ZF�2�M�����>���A�^~�U6��L�ek���9T~���F���$��w��]
�e;�lz��Q2��<�h��^���Y3!�ͥ�Z����pɺ�-��"��'QC:�����U��tS���{�f��M{<NӎDL5*� m��?3�#{�)z�m���\�߈\�Rw���"��������*{G��_^�K��W�CRXG�����>g	�4w~)YX��a��&& Dd�[�U�+���Fr���j|oA@�Q���L�z��ϢfV�.-M�%�^��n���A�p����R6���r
Z�'E<��K�i�>�sKf[J/�j��$�$<L8.����gg~E �
Z�J
�X�_IH���6�u�l���OA֯�ȶ���cs�*� {���\F?��O��V��1�0�4@��#𐩥�{-���I�%�W *r�<+�.q������M;�|���:��w��w�+9C����f����@؅Z�[��Ty�}�
3��Oe~��z�é�Y�T��?O��}��ulu�m`dOçu�3����`_<܆�2�C�Q���d��^��E2ƪ��`���B�pWW���֞�)K��d�Ծ#�X<,��ι�+:�ǜ�1�������T_2ʐ�L��"��!������O@|���8S0y&��ţ�x ��b^�}Wf�ABe~�޲c��]S�����k̛�Yl|��^<�����+t�֪��T�a�����E��2�7�?"n��I���U*�n�v���~g�.K6ߥ	��&E�J����e]9�Y��60�ҩ�F�r�y�Ǹ��ؓ.<G�ә)�84K��`��t�^6Ǉh��b.B��-��g ��ڔ�ʑɸ(.��| �6j�r$�z�ɌM�N��5?�؃�s�3z��eo�tb�A1�������`��n��牳����:�+���F�b7
��n	~j�1�߾Z�V2�T?��$0J��^O�����r�F�,�nq4�:tk�^Z�6 7�KXC z�SU��F`@�'x��؁�\��MḴ3�F�I�4���*�H����RL>���Q���u�mB��8���:wdou�r����g+��� �}���d����"RRY=�<$t��	�6R~��r�ƛ@��:����E7�l�	�[�T��7�pğ��M�y&�����@�j��8�?QP$�z��+q|�c�dH�[�w��F`n�gn�7n���ʒ��k�'�G��C��a(�AY�a1�v:�y:�F��V�s�.�{�?V�op��D:]'�<aX�*��#ԗ,Tp�NEQ�T�(]�_Ա0r���53���X �!�Z_��	�5�=cy���l���q��iv��3�c��T�|f	��̞�ʞf�A�tQ��:�-����zw�v�z�kև�������P��B�2��dH��V�w����pB;�*�
��Tq�)�Vo�t"X��\���@q���N�]��}f�1s�j-hQ��
��7���/�̙��+�~N����n�,& `�/�՟��z��ħ�:�31��<�A�Mx6�G+���"�(V
�~�e�%*;q��0M���N�Pğ��`5J�Y�MI����c��^��2����&���jae�ȕ��&��z��)�&��s3���5h!N�xh�I�6{�D���X����;���C8`
[�'���62V�|���4���L�K�>!����d�D���X뒒?��M��L3}~V�ӻ���+�t,
1��z������d{���I�.�p�19 �]W=������K���.eU���pggw�p��ٙA\�_����^2WX�7�(Ms�6��V�'HMOP՜���-���HI���n��M�^�qF��G���2��v������3z��@�LL'�rj�L�ך�|O������7��-;�!vD�# ��H���t������~�૩e��9_�V�@�W�d��7;��,��"���B�k��ѕ�T� �H�*���~6c�_���,k	��' $���{�K��_��|F� 3�f��[���������+�a$>Fa��,?��J������Ҧ�V��M>+���j�5n �u�h��9�N2����t���)�� ��h����MH�j�'q�7�j��c%�o�dp�<�� 2�ϝ��6�;�0��ĺ��� ��8��|�Z�Tr �xF@�B��ќ���n�a�fS��*4^iPOS�����*���k���%"�.���+��h	�=��bl9Q����V��B|e�܄�9R�`k��z2�Y]���� �\�Nr˺������5��GϹ@���s'�)��Bp���A.�g�>�奣Y���n����~m�CS9���m0I�� ��!��rd{�-�K\�?#u9dV���R�����JgD)}��&��
@��x��m��w B��29�"&�,M�1���s���S�,�M&y�W��G�`����YM��3�6@c�pD��W���a8̀_7g���^��.ot�|y�E�'�Ł���?��Buy�\��7SAЏV�aqA��*���C\��Dqm��[��Qm��o�_2����/��hӤ���%�scn����97�=+���t��.���g�Ip ;��k�JC�AW���������88�V��=��r]�����n
g��� 󶸤�ELm���z�by���1�ߤak�`%�n�m�ჸ���E*�n��Sdԥ�[H\&s�ȣ�����w�����(K}{��w����%��v^s���uR�����������(�?�f�yy����Jq\?x6�1p�g�suLXR����)� �=Ք���:�% �A8��Xȕ� =�~�Lz��gl�1CR��My�-8�1N�|#躲0���/��6%��k���I7ſX�@U�;�/csf��=��!	�K�����&_�()ވ��_�ݍ����(���y�a�ݨ3�\n�;�(�U*���r�+�]E
'�/�@�"S�K��O�[�i�3�͞[Y�T�\H�L�ױ��-�l_�x5H[%���'0���f�Y�_ol�¹3�A�I%D�x�Hyr/��ߤ��~��v�}3�u~�v0O� �}�DJ�syC��u�D�*�0ps�R����H�!*��xG��5� �@�ۛ��BN��:𽣖�ٚ����NsY̿���4$�L�����pY< �Wg�˰���Fk� ��Ig�%����
�|՝�?���1��d�u�6&�(����v܋m���B��-i���-yH��<�,',5��<����fC��ѵ8��p���!�iN���-�j�6יS"�C��T��i�އ�����o��J��BY�U��M�}��Y[���CT�����k�Yܯ�/0PΖ�+���J�j�C4:,B�;���x�XŠ*������в�*ծ�We-*m�\��u#�9 �X�c�o�w��[Ωs��fH�,$E�;�)�p����\}+�������"��^��t5��z�~���))!��x���b+O��͗D��AX��t�5:��/��3;���L�2;�d��Ɓv���W�d��У������3��|%�Y��(R1QX	�w)¿���)`�|��]�t��H	��"~t)ab���SP���@)Ly��ڮ}f���Q��9�>i.p`F�E#x�Y`��$bd,A�{�j�JjŹ�������A��n�o�DF8�[���1#��$�h��/�'��q���-��ZU�K.�%��,�a˒NKOª<��0ٞL��Lh���SR��r7hri&��<���~m/y.o	�^M����t拆�����䬀����j���g �pP"���x!U;�[B�6��'H
�l�F�8A$�9���x��zQ��s|��U�"�,�5����\���42�̙�����r4�"<����N�ӝژ/�*~T1X�Y���<T`������2��M����b+)�V9낛��J�TҵSS���i�
��W�
�� Y�g���xt�h���BQ��75y+\nn/)�?R��Q�I�7
�`,dH��V��ue5�όO��Pau��2��%�F���75�m.D���W5&�┭�Q���/<IN�ӥ���&�Ylz>��,u�ڟ/�����7]Aarqye��ʶ7w��F>�Vw��)<�����y
nw5M�jضϱ"|��ZP��g�_yr{������T����Xݷ��bxl�҈�d�ĳ�Rّ5�=QoZ3�mn����R��ִ��-`_�C1{�9�������f`@ ��冂�)�i����~O�tn��ҥ=]ܔ��PYd��0T�$p�Rp�=���{&b��Yݰ D`�0��C/���]
�8ݽj;�nI��:7�����^��T?D���z�&��z.��!~4\�2v��IEZhUHm�1��m�B�:�eU�cВKu%�'e�S�df"EJ���,�1*
�Wpz����"T�u��,\;��aT)�sJ�t �-���͖:M�Z9J���Q��L��N��MI�S���O1Z��󡘟���gWE��~'ю�B�S��U>���"�)a_��m1?2ٖo7=��S����^�m�up�zRaA�g����Xǭ\�*;�8+�.�-2�]���� }�
Sx�VTt���\!kZ��Lt7�j"n��bݸ_�������#p����2��ɘ	�j捚����[�������B��.�'�muf�z X���$��a˿����a�/��<T�r��&�Un�X�g��G��G��A�6�������ܤ�6(dz��ٔ�ч3'WԠ����`���u�tj�������;�(�M8�KX�V�ѹi�V�|��fe�T�^�U��w�jZG��ojv����$i��\{���I���hٶ����wIf���F�De Q��Y�+���k�.dN�W0y)�vgsB�;�|�`�X
�DD�Q�Wz�l\W������{��k>�ul�A���_�ۥ��a���.01z�\)}�n{��˞������/�s2i�JP��s�e [ؐ0hm��,�e�m���X�dq�W@��n�rŀќ�7(�!oYp��^�U.�yT��jjJރ�y�s.B�R��zԇ�\�m�5&��� �[<��53�B��r�3�-!�;l���ݍ��*�,�7S�;Y=�8=��1���t�I�x�W8�e��۷n�-T�>񔟽�>\%��./�gH�� j���]\�$�F��I�p2��N�]:�5Z|�Y�Cd-MՍ %�/��Y�='J��(�Q��Ám��߱�ef��֦7��7��������'��L��8��r��w�ՙ��G��$�o�Kh��qIo�Oj��80�d5VY��?c�I���}Y�T+|(��FR��J_����!��Ai���'}�91�(ٲ�~:�pqa�9F�� ����;����Q&�)Nnƃ��u��t�ZZ�sSna���# dL���)��~[�c�~�E�������[ߓ��j�Z�r�%D)�����wyA[�C�4Z��i׮1?��#�-�2ƆC��sX��h�c��OB�|�)�a �;h�2�]Vo.����� `�q��O	��G�0J+�<��¼M���ƆRn�,�ə+��)A}@t�Q�ֿ�$`�<f�S�7���ϛY�0J����nc۵���S�ا ���;1�!ᢛ!���j������,$Z�[%Y"Mo���w�x;�Mn�oI �Eф{�iR��k�cZ�׈���6*=�_�,01��Z�+S���[�q����2�(�+Ȧ�kP���b�پE�$ W��g9&��J���%Rx��.�05���)�!'���SV卟6��`C��M��}��/�10��ݮĒz^~roD�E� ��Ti6_�v��>�/Sx�R��(��$}�#�z��$���װˤ���0+��� U�	B�2%M�*��8�����a�����Od�z��{T�lO����Q�s������K�?��9b��@:>�{�V(%^πZٮ�
��=�c��%P~f�J:Y�?�c�xi���V�I)��4�'�&�4GN|�uQ��fqO�����S���FxDD���z/��e�3�Ta{ʺ=��+�Ug�Y��� L3s��g��:���I���@�N���jf�;/D�yL�_d@Ei�|40�:�C����'v��	�E5_;۲H�.�z:�' v!���B%{��(QKI�,,4�)L�rq3������y&�dJ{Uۮ�UÌG1Ϙ�����V��h�OdW�s��bTe�|!U�� d��H���o�b:Jh�y���!�T��%�~i���ɼy���h����0������8e��>��[<�v
��,�F�Sc����M_���IM���"��~|��L��M~���ʫ��LK��`%�5?H�ӆ��w�MS��e��l�#�D�(.��d@��X7�	���~�{�L]t��x<�;-:=�M�P~��������Ng|������ŢI$�!}�����ƚ��?��u<�QL��ÎK|�&��3�Fo�0ec�m�JDY�wu�څm,�d$O�w�a�N��\��^W��Ig</�LB4�t�,Ш��`���y�a�a�X�2��Q�$}Vm�Gm�Ky�ϗjsM�q��p7��a9xɜe)�+П�mvu���F�)�:�֪�怇L4�Q���2Ae3P��g�$	�i�U��Q�J`ۈ^Q�c>�D8@��/�R'lYf�ĩ��4�w
�4�ۂ�E����Бߚ���e%yJ��ޚ(�S�+�	��WV�Х�g:`O��5$]������p�ZCe��|��ۼ�vPs���Ʉ|b�/�L�&����ϼzo'$��������׈�����WT�� m/��h��ܬ䝳l
.�:�GS�z*eR��$��=vmcȎ˨�?���ߊ��M�:�<���#����Ӝho:����2���Kr���#�����Q�m��!��4�mT�V7��=_�턯�0�i������W���UՈ�]lA�Z�����o����;M�|��[H�!�3�ycg5ۢ'��J�uj�NŘ��#}7!�D����h�R��M��T�_���e_��������vT��`�J���C�UJ1}S���X�[ɷ�m!�#���X��N�f�J ����DŚ�!�D�H�薑]�Ro]�|~��C�u�:Ƚ����AZ�}TWR����φr��m�w$��Z����:�c�YJ	8d #����̉�q���g4��r��E��ӈ��mk�^�qH���)�ul���|m�����b���,4���q�-i�} ;=�P��=�{i.�;A�U� (����\������q�AB��?uL��¾W���@��Q�+���1����mj{V�Tkg���DA�o�LkT��4n�-9�}�k�y��e/���ǧO�~�N�f�<+���]x���RR}5�%�����[w^PB�����+�U*����_^E>�%���Q��?X�K�A�@�bM'�����Btx�6�,<M�P|)"���/C������A�(�Ч���9^θ]�Ql9��\T���xIB[�>�-����]vgyz�#t�i)�wдyg����G�e��$B�LKI��̡�wK$B�]0�ւ����HJ/U��d�(�:��<�xM3"���H��С$�!��Pju�18&�.�A�U�\�W��ܥ����wW�I�|����P�p�Pi�2��'#�`��������g�������1����8�n7��;*�D~�E�.giM�j���,��5��}���Z;5�'��L�!��k�8R�Fש��X��0׼Ċ��1)?z*��Ջ6'L�ކL�F�����6}����q����fit��r��v�,	#\2Dw\�:lV	��C~�698#�j����߼���2e|hu��j�y]�to!�
m�Gr����)�r��IKП,��!J����y��1Bn��u1l������M� j	pa�<>�N��S��(���͗��b���}d�1wLAlH��b�;U�!��n+"u��;�`��_��)��	s���@��XPP&�e��&�����_���xkGS��J�{(�!�NK�yV�w��@?R��z���N���CLO��ѣ�	W۔��D��x���]7����3yU�k1]�e�=����;�k+�����	Aʒ�RMF�4Ԯ��}�z:�A��D�+i����wn�~2ΆύuI9?R'�b�X*��a*e��#O�&LN�z癍!��Rl]A���|n�![��}�3>L��QzoX�~�W�='�/��4��_�Cę�}u�̱H
��"Y".+2���_u�/�Ԟ'������q<�)ajx�>�2W_�aP�b�* �x��ז���4-W1�]m��|�]���R�nK�ǎ/�A�m�ѵ+�R���?s��6�A5g��C_�c�[��W���Z~��,��t�YL�B7�! ���[�[�����!��o���i1ȴR�W�m�햱Z8L2�3w&W��&�9d���[BJ��9�5m��	~h��s���2u���lI9�*�� J~�����>��c���ɚ��Ul*�fٯ�<-^Ƌ&z����75&Ws9����k�E��Q�Y!.�io��e&՛���#_�9W�X�0:��!���"�q��0	�Q��/b��;�΄P�k�C�)��Ҕ\���|��z��+����Ӗ�:+���u%��-nL_�?V\�w"��d��P�����Aζ{H)��M/Қ�q��>�і�[���У�o���-�-OE����,Ⱥ)�/��V�\���*��UZH崈�!�����s_�3�`yD�͔�j)�T���>'�RҒR-vg���
u��X�J&B1K��Swū�>�pIp���`îs�H�X�.�s�j���k����[.��o��~;�D��"7*�XÍ	���AnLJ������EcR�w����^�p�y#���i��{Yx��O�W>��=�m2��H�E�KT)��9ú��Z�Α�4�YP��{Sd�⺾���ƞxM�1�8
�z���e����)�b�9�U�ј���Y�`���'5-�A�F�Iv�����+G���K�߸�a��̰�J�绳<��^��DO�ry8�<N̍��E��	�(���aL�#�:��J�����8 F2��ʬW�g旃A&�� ��ƽ^�x����&̀�R2.�Aj�������.	����co33�sk�k�A�������?}����"�M�%1�Z̐[AJ-�(�˶��=�'�c�AC0���Ƨ�R[f+9٤����Ѝ��������ȏX`��8
��6����D�i%q�њ���-*�U\0Xq�?
��Z++��c�FYS�eR��(8��T)+	w\�T7(U��@��4����t=t�8�8h��n�G�*`Y��IzG���!p��$��9��7!�n*RJ����m��y5��$p1_�U�V�%� I99�L��[�/1�
��v��X�`�����3�`��rt�ĂQ���0ٺ3��c=�V�>p�j]{;՘GI�i+ԏ����B��>��Y0����K��e6;�՛:l%{���8_�xD�c_=�8fz7�Vt�3&�D���*�w��6~����a��}��pL@-)[���(�9����-�������ʬ����
$ fR."�;*�v�ب��5x����b�E;��0�>��gR�N�W�,���A��ZҌ�3նL �Bq�y�S�C1y�k�%N��`؝sGt-��nAb(��i_��Vt�Vӹ����M�Y�,�nǊ8?�S�sB�C�%QNS������b��g�Q�4����&�_��aI��H�'�FH��޾$?�C'0wh>�ǒ�$*� )B9���Y}o!n��-�"��������J��' t�㕸��EI��S��8$�Q�dC��Ψ�֭n�FZ����%�����Ҿj���P�����7�Od�E�:��q9(/g;@͏ٜ�A��Ž�!S*�6�ÃO���a-C&QG��U�Nc��}�~�"iU��� 
��a>*+~i7�Q%�e9�(��W���*]�:sB�ݖ�5�e\��)�q��mHa��c-۹3l=���l�F	�!��L3:�#�Ŏ�JU��w[q�Y�������R��XM�?�p9�]x�Y�e[�{>�!��-rfu�L̢���������٘_��d��Y?���e�JG��%
B&$p��<��\A
���C#�ʝ_�E�n���|]�z����(HÓǈ����I���B���s:�|��Q�Pc'����c����L�1��t2wC���.�x/���������^�饒��_�)�y@Bv��Kސc�ċ��RyEVl��g2��sv85�6Aa�czRs̼�F�o�{����`.Ց'P�롟k������=}R�%H���l��fl ��� ���Q��q�
�SQ}1�v{��eԔ�f���uˆ�?,�������NU�P��h_�iL���a��H.�(�>%2J��9F���*G�Z�g�����:J�Z�)d�"����o��ppW�ț��s�+��}�bN��Mp/!,��UTl����o�9"NY�AF����6o��ߺ�b,E$�r��1?��j�9�K'�6�2�P P��:4sP�+�W�]PQ�p+��H�~�v��0�Y5��x����}ت�R�ԟ��ri2�BT���	�[6���j�U��������#�Q_�.�_^D�g=���U[9�f_����'�ĂF��Ng����W�h���D��H�����a
�1�*;�3R)A)�����9>���T��FO5ѝ��>;J�@�O�(Bʣ���:��<!r��sTi�L$��T�J`6R��Bêh�9E�4��.-	Oy�c)�`߅pN���걃�}��8b�r�_��cƴ�hzAR�@'�g,k�J�t_�(��m�I��Ҥ���p��X��G��oF13�V1��M���e'K3�{v��
o��%3��m��r�`�g6�4G���"%���U��"+T�f����C(�
ןR���8{m�su�!5O����tb��b��%�	��C���Xq�Lh�)��� %�:e�h���6��]�>9ɪ��wC����P��Exo3W�X����,�ʉE��՜�z[�Nm7��e,�׳B� ���͡xi%�K��2W ���/�i�W���c�[�4��z�	�]G�rU#˻���L����Y7c��(���tzV����t�{���Fj�]$F4��e�e���,��X'��H�Y�����?t���޾=޹�,]����҇H��+��.Z� ��<1l0g���k��9��aPgFj�dˉ~�8�|y��g�Rc��Ia��4�tiq����w�@��yP#50VQ��U��N|�)�T�ҀwD���6�yA�+[�V���\����οR�b�C!�Up�^68�]rb�Rۏ3�%�;�����q��Qw�ad��t �����G,7	�8��Rqȶnl��7߄
K!u�1K��d|��K�����N��9�Ǝ��8���J}V(���:t"Iq�~��$�[R����f�jSN����駮t�F��$�\�p�ڵ���ik�fmf�aՓR^���f<�[���;8��Z�zf��G������C���J�_I?Qc�Ґꛐ�C�P���]|��O������s|�ڦ�r���$��V������7)��uC�f��ÍW:>�/��L'>R�Y2h�_��䲜�anl�\��j��/q5&���&��O�<���Q�ʺ>_f�ǎ�a��ge-pH:�Nz�"ץS�����wWt$��=J��@�4!�����I�s¾��2*G����/ ���OS��7Fd�J�OY��$1��`�I;�����`��I�H��S8t�rOl�Iη���M����Գ��o��=���0��#-�^g�g&I�42���jh�����!B��[?�ud��:��佺<��A�{�*\+���aĎ���:�����@��(�Y��eV�6��`Z,ק74R�lJ�Ξϋ��U�'�������1���A�p���(���}��[4��H�ߥdߛ2v�P[44�<�J�A�P��c9��-g��@������"��g��?a�)LÖ���\������O��&g-Y�2�"\�ퟌ���,�x��	�ko��m�c� �{���$�awR�/�Ϸt�G���#����N�7��ͨ��U���w���M���kA�b홌}֍�<�[�.�f��.8�-����#k�C���ZDP�
�
�Ns��%��!�p���pX�L�^XR��&EϤ#�w����u�/1�Gʸﷆ&넪]	_��"��W8:��>Kj�Z��j���b��;��
}MB��1o�}�fQ�e��$����c7���������]6Y�=��ӳl'ηw����I��r���7weG.--��;�t/�E����顗������D�^��#�SK���<��nMa��>�����&ӣ�z:H>�7�� "C��Ǥn�Q�a�B\0��
����[�����Yf�Qs�jtϥ���"����@����x��7�]�*������?�j���'Pd^i
��v���}7z���p��c;��^)�jR �)���u!C�tX ��.�������%� ]�OmY��H�ni��a
����+���ڂ���Ot�$�2N�J�Z�?�D��-�WF��[�-~o��Ӿ���q��>A�frj\�SzL<�Ŗf�s�ۈǹә����C]<w�J��X�o�9A����X|��F����R��&�`���M��qE4����^5����M�(�$%4�&�2�Of�����7S�6f%����]}HA�f��G�1�%�_D��\��t,�M�S���T��s�l���JB
X�����'cƐCax0�R���y���^�1�ڨZ{%��m�T!����b?G&��Ewج�\�l1O!%�x{��S��i�-�4�,@��:іo�fg�u�N����S�'Ws1�'NAP.X&�gb�:]Ɛ�����K�8�3�u�$�8�/R$Yo���6�!^�;U0f�Z���!ۅ�A��xƨH�����w����ƻ� ��:�@w�-*.|��b_ex����eeE��7K�����GK}������3���LE�O�S�J��װJl�Y���3����=�u����<����̓F�d,��[�B=J�R�}�ɶ��� ������
9.�8�o�D��5�~<F|B׻P6��h�S���w����h�c0)q�[��X��P���L��i�������Ml��І�*@��g�����s��GC�^2v��;4����A��ܝ�p��~'�H35 AV;}��(��^y�r=���9�O�_df1�*�9�����sT���e����Ib�\����m�^8�e�ʲ(��� ��謪���)���LS��W�u$D�F�
��/�~R �Mt�ؠoʠ����u	��ĕLR����{F�̹�>~;v��K���Kw$j��Z�"��M��Hi�5�E�׉��ޜ/yv"k�M{�̏�`�eM� 4UXB*��;��W����
��T���r%X������z���E��*��>$�Z!�c +��y�J�Y��Q&|