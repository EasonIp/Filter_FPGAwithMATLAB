��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
N�m�H2
��j�Y�?	l�Aō4�8�����>|�f[؁���
Ζ{�����0>��������'l�d�b�%#T���QOo�Rh��&42`�-�R3Ml]�Gq�]O��ל��J���('���Q�5�.����p��� 6�	J�/FM��8���b�)f�ĐI];�^�EL���j�����D�1�5�1�K%M6P�]���*"&	а��u��~ٷn$5h����k��O��L���׎D�y6"�  UD㍺���"O��ܣ2^ �4"�.��d_y&����V���k���ƭo����`���%ȯ��e��εA;�3Yй3V��l%U}��N��������aUiJ��������X(7:�_0�Ah9�[��=�2�5�����,�_���i+���C�m���K-?�qi�b<�-�a�!?@�3��w"�[^�J�������+��A��W�P���
�sYy�ŏ7j�S�����h����nK�L����E��#��-�\�9Ú��U���-|{s֒Ѩ�y0z�]�C �_@Jn b�K� ��A��a/�F�B�!�Ma��Y'�����G������]�LQ���|��gE���,\6���Պ�E?��d��򄻙���R88���Z�c��5���G��{,]n�M��������ܵ�l�{h�W�2;��+p�εn���>"q��N�G�T�����o�-�m�%�xG
�o�]n���	l��'��a��qB�d\|���Yc�Z�t�x�塳Lr��X��/'>]��59֥�'�w�ƣ����2I~ٺ}���Mw�q�ckg�<�B��<�� �b��ű�G̹�[�(�R����Dz��#hu ;��9�`6.z\��".����X*Q�dP�So�4�K��z�~�n�^�a��W��3	# ����k%��t��S0��9����N� �o�����.�Nj�z쵱�G8b�1?�v~�W��e�POOs!iъPU1��� ݀���e7��o��^�]F=c�59�s�+7�ҫv�J7=���z
��_�σ��y�\���h�_��s|��Z.����*ô�XE�@�L��:���e�P��E�U��2���Ἒj��iu�*�9*���^�y�Y��ja�3����qL%Q~����P�l8���Y����3p�V_�X��U��2�p�R�
J��p�ӥ�-�؞7�;���
����ԃC�B`)��Ђ��#�L.��FbOx�4��w�6�c��Y���ia�W�le�\�L����
NBR��@9��+����dϜBF�5��q�>��&�.{a��n��k��/|�i?ڜ��J���|�pP36���ҕޥ+�ϻC=�;7_!�g}u_�]�(��1Y׵��B��r����Z���aqB�������_��2����<�g�$��mִ�Ga��)�f�"��{(�3w>�R�5��D���t��8���A�����VkQl�"3����}�� ������z�����T�Q��@f,�V	�
�ib3-m�''�)5�4D���{�c�+&'��'�}9�5P�g8�����-;iaJl�$��W� Cǳo��zH��%N=����Iq�>n�0��| �H0�,�X�RhKM�Xۇ��tQl����Ge��j*��x�G��K.�"�b��.�o�\�����Kg+T�Z�����m�Ĺɤ�
��ó��&��)5�&�+�m,5TPY�Vw�~%8A|��=�H`(���JآD�ދ�(�K{B��ҝC:�%X�?� #�4K�������lTH�C˴�t�ԕ�(�<tۋ�$�� �?�R�o������|����O܏0qt������4����/a�+&[.b&����	�Vo�-�0�,�ɽU��-A&4�#[��u�d������y�e*��]�E�����1rGz�D�b���������?��C`�� �̲�	�Į�j�>|e@�T9�K�q-�C���7���C�kcn��DqZ����!d��su&���������}�1i�������������>a�\�۲$���UO@���χn�%�G��Ϥ�@��`��pE���C��4V'����I
�)��_Q�I���NA���,�~�JX!~�.���0�YwfX�20g����T��J�#�ݱ+�����o�'�a։[���������� \aB��7j�v�� �� �>�F��3�(-��=�Kz@������m�S��赶��G`Jv�b�BT��re�=Fx�W���6��Oc����s)fA������9���t�Y��A�b9c_[+��|�ы8ő�q�d{y�:|���25���������a��t��Z��\(� ��N�r�oÅ�
���7�==�	����t>�w@�RV�S��,f�=�utf�*_�ꢕ�®d�?䌺�@����q��i���W�����jD����\�#����%c�D��ܪqV��0�ܖ���5{	�\�*�hɀ૓�£\�p�N���S�)<�H�O*9�i��	�1��ZF�����G�s*p�������H��$�ʬB���o_.۔�D���J��jc(��'kV'�
������Ƚ��܃)�A��nUhp�@Lb0�-�Μ��Q�Ϲf��[8�$��I��/e�T���6V`�/�46}|_��q�ϙ�5�(���o��ٲ<N�SB�R�&��w�L2�aP[������tzz�5}JSj����3�h�|��H�G,�`-|���J��LV����{vo����O�R���R,x�b����g����!�]���Z"e-�C��k7:ZBl��E`��:��������˼V����6M�J�[;=�vQ؈�U�{�c��T�#��$p�����X�Î�A�Λ��_&�÷��r����z����ˤ�lg��Q�HX�C�i�%�4{}o�B�,Rph�P��r�����|�2���|�[����?�y�,l�}�T2#{ ���l���8��c�_O~H/{�u�-N&/%��a���p�.�2�HKmM�A�Ћ�9�ai�^��O\%&�6P��{?+K�l��U���_����Zj!X����ف���up]l3�Sꏲ�CP>&da$�1��	��m3�@�����t�]r�V��ӥ���\-w�mY��;I�U���us���N�������P>UY4ިI����c����EM��/�G<�6o5u�ˊ0GCZE��r1�����'������Wj����ߋ;Y/K���؋$�8���a�������Iӂl���:Mnd�d�0����f>.	�5ZHE�����q(�s�̯�v�I� �sK<YK&����wᇬE!�|��C6��p�E�?��%��`j�N��l/��������ލ 	Z��%1.#�%��EmP�X΃x�7��8['|��@l����lo/��2�Ku!�m$��Ro���3��B澼q⽱�o�TqƖ���"��>V����ck��Y���L󧅡~W�##4ݝ~�^�^��� ��u}k�Q�ݗˀ~���+�Q�H�tߐ���s���Ry��,��^���5���|	T1��+�H=m�^djx��xl���Vm �L�gmt��S`�����~�Y�A�Πiք^R�� �*Z��g��c/����]���L|g���������[iE�<�DB��p��� 36�*R�X�㚒[��߻iX��UW?/��ʙ�]5!:�S^֞�Q3���wZ\_7 �%]�"Y3:,PA��O$�i���Ԋ������)\�5 W5��/�ے��V��%�	Fd:E�e���f�z����C��/eܮ&�g��s1�b�9�y���s�@=N؂Jf;�E�T��W�U�y�`�XmԤU��}�;��Gs���-����8� 0�!���$ƕ���DTm��)q��"��͖d���ڸ���J+���Cn	������R&M��� ��%�M]�pD��)� ʤeem����WM��~fY;z�+�s��7��bSd����Z�z���Z�=��7O �,^ᥜ�U��H��.v]��'��㜯n����d�\���7�؃6f�ٺQ �2��X�E�L�#T/��9�8)ͩ���}�.�i��O֡���-]�P�ԥ����Ņ��;�/(�8z�e�i�ã<r�ډ���[Ö������6�P��ˊ���D7"-}���F,�G�O�?�P����_Ъf1C�{[����s.��5f
捼M_�7-�f���Ϩ� ��6����Hr�(y6���z�%������2�o�9�BmL�QIU����>�oXf����� ��y�GU�
������F]�u�?��J�M<��ا����>,�]��l\ Qw���}��\G��ݹ�X��F���1j�����Ӏ�Y�B\1;+dݠ����:
�z��Q�!!��Y�A�+I�*#X�.@kdl��jŎ{�D�֞��)[�2o/��$��o��I�,��'����W7�*��bI��(ly���*1�	Q�ŦoS{�[�����~Q�	�j��#_z�.o��H���&���$婙Lz��R`�J��*D�(p-�[B2
*��¯���X��b]ߛ�@�n/�h�*i�[n�%}�辡2?}]Z����F|�v��d�F��w+0xϛ�@��=w�r����К}}���}��ax(�8{���^��:8sAred�0����R����-h����%:ܔ���\�f���:��|�E�t�	X�Յ���Ȉ�13(��I���筣��:S��h���7�E�1.����%��6g����+d~[�t�%҈����������+��6<q	D7�Rh&= ����Ћ��y{��p�\��3���-N!��NX1υ�S�B] ƴ${!�L2���tN�K=2����An52�ު*I�����RC:�	mHaK�/Ղ���Oy���y�KH2D��+�>�,��r>4����c�� ܣs2��7��(��>�QQe��Y��	|���?(�		���	�pŘ�-����E�(�Y����&\rmg�������w��ǳ��Id���^�S��oB���7Yj�U�Zgl���nFL�<�e�x�Ǭ���&I��3�|N{Kp�O�;����E��Uc�6Ķ�!>����۠ߥ�-���X�j��gx �����O�U-�\s��鏀���X���g�l��{�%�����s���W�H��P�L��XC��#�Ѭ�}��C�s�N]w�����!�Y9���H�4�%/�qǐ�^Zw�̘��R��7ձ��R36&.��W�Y�>5%���%���t��r�<W��S�Q"(K��ذ#\�(�,Y�8͜�y	��I��p���˲5��Ǽ�9+�R2����T2���pue�=a����������le���/��i���Q��w頎2����J��ݘjw����ë��I��~^I���F��$P�ǥ&�"<� f�{��8
�f�P��>T����g��N"�10�r��]qЭ}�S%�^��T �*���]���Pe��·�r�u{�E��Me~�O�W�cP1�xy~W\���+���7YK밸��1�6q_�_,�/w�R� ��Ս���R�?V�A� ;��(Ѡ�;e7{�U&ج͏R@'�SoHmGa�HtW`X��)ZO+D8CW�G=��� b�N)6��f�fɝ6��Z=j���
J���de�O�b1���b�N�D������+N-L݃S�Q�k���Ͳ[�����<jKS�yB���ft��7b0���|4 ���X?|^�=��:V���<��b��B�e�E�G{(o��8�1�>��;3�W0U������!��)�a�o��ႆK��6�i��צ۶���n;b�����_9auwf\���x! �g�v���Q�A~�R�r@�T���r��-�T&տ�����*�Sa�@���s��{�V#�8�ZqٚYk��Šlw���
id`-ˇ���s��C��P�h�R�џ�c��*d�H%�~�?�.�����/�L��x�k���=�t�V/�JA�}s͌1��k�k����^��������x��\Sq�6Z�A�C&���|��b�'SNZ6��Rq�^�Y�U/�KnЊ��n	|�V�];C:���`3:�<2/�t��D[���I,D�j����̇�qs֠P`I��w�5�+Y��-�U�(۫\�����?A�X�"cX��{Կ����u}�}<��?_EUxYN�x��X�<=K�Q�'4��\9��~p� �m�V.����~���®?:�%�G@�&z��gخ����?��΋�$$�	��C��M��v��G����W���W`���7�9K�"�����\�p�m�Dך!�a�6�B�}B �sˮ�ʎZG�v����1q@�U�0��"+�;����#�hC���6�b'/x֘%���(]
t1a"���m�����������Y�N)ڙv��C�J+$��L��Ҙ����[�z�H_C�|�7{�y�kK�t[yoC�S���O!w[ät��ֽ�H�3�3ּ��HSh�7��ߍ���c>����	D��ف�>d���ܤo�è�L��)Ƿ�5�@���Pe�hv3h{˴�� ���oo�[ЁR3Z@�I��Q�=�2�����DĨǜE��t��><@;�?(Ö��� d�����5��&�Tշ��`������3yXU�N�p�d{���y���V� ���a����IZ�<�
�!띷�O�`�B,�\�S��t���MS�$r�7�3�����*���A�!?#f�=]�=�w胙�q�`3 �;�� a�Sf���_v}T��1���dF��\��� �c�@/��i��훞�x/�C���bFI�=��@�ɬ(>�Vu����܆��(p_j�8]��/���\�d"HbS/�nJ�h$DuB�*]�KB���h���-�4f��U}��b}�6k�p��Q&*���y\��j�D�$�|.l�Т�!�_ �i��7���M��44 ����Kk��w r�<!�*<���(	�M:Ӄ8VP��ێ:Tt+P�=q�I���L�J�!�u⳰`�ڙ)A�Z>|��b�3ӭ<jQ6h&���Ɍ�ߧ�Y`��+īcى�Qv�l�@kP�����	4�ikC9�Go%�%nƋ������sx�f�g3>�������9D9{�\�_��{}'Dt�'���9eFUd��g�t;� 1`�y���rMJ�I�yIE	���JS%ƥO�*k N���%����& jX��#[&� ��\Yo����AFwX�6ߜ����{�)�c5�e�����Y[
�y�$*U���:�O���L�0e������8�Q���5�_�J�K/E��^!^{�Bl�Qh����nˠ0�%�ir�7���|���AOY�l���گ��&8��7����,Rߏ�q+��?$�;��g�x�f2�dD��Ǝ�)ը6A2��$�yy��b�Dnш�b��w%��X1��Q�QL&)��+�d�EimODK�W)p��1
Ja���F�pI�����(�oWw�� 
��M���/ɬ0b��B���?����v��u8�B�S�s!�.j��*��y��,�稃�6��n�/+��
M3mj�{�t3�V�נ|�p����R���ءh��~�GԲTA��Q;\�	�r�8ږ]c�T#��IF{nh��M��*D&�̳��u�V\Ń�))LՎ����$�.@X�(y�����Ul� �u���쭯'S�F�.����j4Y�a�vHiXx�-��7��U���*ll�,,��Pʓ��t�J�}�`�48����[�Z9}&aJTyl2����Z~�-9_O-W4F���(3�2u]9F��ky�%�'}9�6�%F�@E�9��;�&��D�DZoR�����9����"��GVY��p���ɾ�A�?V�:0�@ H��*n�A<1k���&� ��tZ���]w&���&ݕZ�<���b��,��O�~�G�}��Ñ5�����o��Vj�l�<&�?�,BKW�RVK�Qɕ�#<���xs���C&�	��X�v�m��ۊrAD���� �͆8��	�6kי���;ZT��#_�Y̂)�P߷��vP�5��,���YgĹ,Ofk�жh��!j�	n�;$"�R�6�YlpM�w ��z������`�b<a�Φ�L w�(����/��f�3Vl�A�K+'�����H��0 /#%�h��ʉ�T��H25m5��檲�9;	�$��Jg��M]�������q���Hg�qפ�/N��+k<%�9�~�b=�6����+��F�.%B���,�/M�>C�ϛ\E�� y ��שR[C[z҇E�F6�/>�<A��jD�~E�z��LpjǢ+vޔ�F��[�`]�X+y)n`}���D�����͞��N�YBI�%�ǊVȺ+h�R�?��W���̱OT�o����Y�&6�n�������Z##��[m2��>p�
��M� �<���u�� p�o>�K�K1G���Rb(�S�z�B����`�����'��庉�!H��x<<
(;���-ٴ~������\�_��E����������z�̩��d���}�?P�UѦiH�}.���$�@�p�t�(�8Yo֬�bP9�3Qr� ���w��B�f͔c��m퍩�Z���~��gG�p�!:.\I̓(��ƕ/̍}q�c��yP�{�`���p{  �S͸II^��y$���@�0�B+b���B����q*���L���>�~)���T �8as	��/I���&�Au��y�q�}�	���GF��w�̵5��BG�h[l]žu��j��YՑP)t�j�F��A�d�=�K��>Rs'���͹�|~���+M[-p�G�X�"��/]�]���dX��׮����y��ZB�Ӡ�R]�G����ɮں$�2SeB����~���D6P��(�T9��D���y�D��sC�_H�a��e��w�t�P|�$ Q�$���+@8�V�D	;:�+�m�Ұ�M��]�%��O�h����0�|���&��Jz�ټ���܈�4~��VkFz��0C�xk���K��ѫ<��R�4ًY��S��zO�����t�t�s�6�#9:��/��þ&�~(?s��d�LQJ�$��=4����Po5 �%�b獵����a{#�~�� ��;�
�d=��wW����Z֯5������γ���,Rح}kl�#�z�|�L�m��>�s��Śfz��˯ci�E4�)z7\bU�̌|��h"(�9F'��_�6�!���V�/�!����X�)IŶ��t��Л�S1L�1��Z�����0:����o�QY�a�����Q�p�Lmo�'r<���T��l�0����>T�zr>-������X� �+%��c=��~mf�l)��m��p�Z*�|k<Lmrf'X}�k[#�Ȃ�	�m�Wq����7P`o;q4o�H�E��6�0�	����c��-����z������q,@r��˞;3|Sd�ǘ`8:�$���-��ā��·_ߏG�\�(U$A3��̱ 1�~��D^Vp.B�:�[<X�C�a�5wd�zb�n�L�ON��p�>6����{��/뒙�V,�'G�(~G����qG�m��d��pc�f����!R�F���E�,�7�~A�F�p�-�V[f�;3t9Hg���s�pݔt@yُ�堼"�^e��=���<�����,�?BAS�c3��?�LC�� �
>��ԃmO���l�n��}��W��Vh�����O�ˇ�!�t(����i(Z������v�J��z�ϰ�߭�Ǘ{��pCI�`U�ٕZ�)�$��rz#Fs�7�^i8�q^J��n<�}�3����t0�Lɷ�9c-�8�i��b��4QN{��U5<<�!a��-�bU��5�qRC�=���ف��d�@7���m�Ff�Vm�63�u;L*�=���|�R�N�ʾܾf�s6J`Y��ua��S�׆�M��/�7�o���4{��S��b7��
�����o�-J�uH� 콤�k0�g�Ըu��o.�M�$�K�K��PS�=�l6@~W!�r�#�`�}-%�ѯ٤$Z*k���`l;���Qk�}Վ��\I�/�����\��X�X �<�A�j��Qx1�a}��g�o��������'��ҁ�K;S�O��?{�}ػtt"^�e�EqJA����R?X�y����j�1�"l{��y-�����[����lE�=��@��&�^n�+���]�e��6߷����z׵C�i�׷H>JP���;���F�=n���blu�#62�<x������~�Ȓ�@�$�6��4����1 !+�r���}]��c������Q��	G�g���,=�$uF���c͡á�wA1$��m���h�Ծ���){-?�C�N��������D	�h�Gj�^k{����s��$�̨9�C�3�l!M��0��z�6}[9�1�Aw
����ǉ��x��B���A�G.����x��ݔ����Oz��%eXY�7�Wr�ê�~Ds�-�Z��Ivp�+���g�%��7��Kd��1�n��ε<;*���u�)y}�����.�>#�Z��]/޴�W�&L��y��]��:�p/���(d�3����vH��
���:I�t�O�@�5���R�����U�m��Q�i��>�¡Wwa�"���H��,��f�ڑ�?w��t�fR� ��o��9E�0Y�<��`Ԃ���0Q���6w����h���R��)�ǹ��dg,���\U� |AtH��	���E��0;��:ls1��*:�y�����R>���.Ü���ra<��ݎj�e�1A�x��z�� �JL�����.A���鵠_��Q���s1�o���;���Y��8{���F��b�΂b� <��>M�,E4�c�:��(��$q�S�E�N4<�s��8�)h�#?`���K^4�amh�Ϩ���bJXt�fU<0	 a|d�iM���"߹V�0�TԈ��d���-�#��ð%�\���!� ��lcS��G5������c��8>��Mv$�n�\��������X��Eث�;v���~��1@��s��nu��M��/��X��X�5*(杢r�g��a6�����x t.g� �g��!�
w��]1B����a
�Lڃ�G7 �!	k����!�����姱���X������R[����4���^�NL�l�E	�� �R˘WG��/��&��h�燀�@����9!��s��>�Z�m��^���Kԫ>�˩����S�)q�R�x�ٞ��o�9�|�m�ȱ�p&�h�T=�>���!cM�TY��}y$8�x�k��F��9����_&(���^�����T&�^�R����P=ʰiRrrTV0�CnT�i��H�ǒ4��/06�����/����\��c7���~k�-��M� �i�����8u���9U��
����U�PD� AVQ���@�]�-&x�3�����B���W~��?	#��x/D�f�����R���3m(�a��Ѹ2�o���"�w!��5B'���$��j�|E4y�l�sl��CiP��͇v��x���4N����)Л(��� r^�MrȔ\HJmw������� �����o %�q��,ܱ�ب���{ nYF�bc�@c�K@���T�s2� ����Q9Y)|z�`���j�����D��ƒ��ln�#p�2%د� Y-o�?���8}f���50��giQ]u}�%����� m/#d0�˞�=ݜE����X=����	:�x�����Ƥ���{/�M��?�Q;r��i���`�mp�U=Jz�,�F�������N�B+2n>�k'�C�	����I��ݤ�[�{��$�B�f��PsL ����~y�#V�Vob��%�4ѫ������0�_}zS����5B�p~6A�]�kJ8OΡQSlm��'W���+6�8�cVi��r���t�mtݒ���=%��Â�X[�u	[�$�5����q	7
����}�z����oUU��
����8��p+k�QM�D�A���$8�nI�-���/�����?0�z�@e�zN�ǜ�p�c�l�/�ZU�d�Ě��uFz�$��P�/�PA�Rf�E/`���KJ�-q�6�M�J0�LK�������Q� s, ��2)QdVF�>�P�.��Y���χ��1�G:�T8cd���]�$��v�>ia���m'fG
<�{���MS%�AK�|�i��rŢ�jG��V�~pE��v�t9,����ACgN�ç��ͧ����
�~X����9b�#���S��u(��< WE��|��� M��Y�2��-���R�2���	UG}�e�BR
1��p�h���� Vt��p�� ���W���=�9SPV|S��,�K���6Ѣ��v���H��h�`n�e4��[x�U�e^���tۍ�V��F�X��Q�w���[��(�3�J��К�N�Ӥ9����k0q�Y�V]ou�ۜ�@О}\֙5���^��z�7\��Z�u���	(��{Zn���҈�.�h���\�R�xs�@��0jF8��7������t��B��LB�j`��M暹�^�&�v�_L�I�#���b
�"�N���4
�+����5dK���y�x�랂��m#q-�M�ݺ7,C� ���@�U�2`����ߋ�,)���G��+��r[ev4��)���w�mJ�������%�*��P�g�� �?���-r�A�v,�,�Tv�a�~��,�d�Ӭ&��Jc,��~ e�<I�-]���XZ��0��c��� �� 
~��.� ��)XӐE�
QO[����W�j����T:5�=;|U"�m�� ��וb���o�!?�����^���\��;��bn,g�t��x�e��hF�D�pnFX=rb;R��(�)i�ܴ��w�Kh�ʮ-R4Gx�|�MM��S��ϳTz�`B��L� ��)��ի�B��e�߇t� ��YFo������~w�|��ȗ��Qa-h9��r+pj����ܓ%*�
mM�~?�
Y"+jj��{؜�%7�=�E����(��^LN	�,q�i�;\��G5����u:u����:�:�o�rAL��k,1��H"U�^7���D���
�L�u�
�[K�0Ů$^��b~�RI}f�\G��'ʋHU�q�W�&(=�>���UGշ�Z��5J����
MȨ�~�~��w��B��k�;R�'T����Q�NpDXn:�g�E�Y��w�r���!�����e�� �%'���u�/>Y3���)�y����Y�_K��TT=.\��Us�o�G'�A�� �1]!�9f����Ǭ��
9�#���������V9���{�RH���0Ghh�2��#���4�^�V�H�wBJ0�E_�j��,@1�d�O{uxd}�~��J�@�30�1�����^�W�n6Tr����[	t�G�K�ß�r$�5�b� �Z��=��4�p�K7x,��^� ���IaedeƲny�p�;�E���+��_yg5c��["Oxݦ�4��a�� MHB�M�"n$ :�?	-�r��vEf!����?�DL�8��/gc ��hI�b��DۇO��x��;*C�j5��й�°�-���D&�[2^MiT��=�l��J�mËE�P��$�T %s�|��t��s��ݯS��O� Gy���Ѓ��ó<��``D� ��υ�) �˝A�s�֦�'.�����䏱R��P�!��:��#Q����Oԯ"1A��wQ8�;��T�Ne<�])��=]�?0�&GGу���5�kDI`m�Sb{g�55o��t�J���4Z/15�Y���O1*�C� �u-#P�Rݸ�����5�J� �7��a\�jh�ᗫ�&��/��w��>�,%�k�ɴ'��ʴ��f*��r�!ϴJ�%d'�r� �*Rg���2t�S��,-�=���7A�Nz�|HN�]�bw)s`�&�uJ}s�KWT�A�a	� R(0�z4¦C%��9����N�nG�5`\mg��6�*Sg�i@�K(�#� �P�%aVķW��_8$u����+y/l�G2 A$@����X�>�4�����6HU��Y�9�|X,c.w��cX�y-C����WY�#��|[��,���y�Q�|��cPUQa�WM������V���6����x��R7`��Ѯb��0�BkE7���tT�,��Bj#[Y��k k1������+�^�C'"��P��M��9&��~�$�,���Wx��j�ipK'`r��0�V>׶�� �V	$���l���f�`�{Lk1�5sOH��O�|ʠ�q�K�Г���u�aJ8�̇��Z�ا�ˁ���䌠�,�W�o��	�h��v։Q�.�߀������g��B�uݏ��� �P����A�)�ެɻi�i���0DÁ�R�TrM�������jH��/���T5����a{ɘXS߁�3��G���E�9Sl� �F�OJ�j-��}!j��^��&B�������Э65����aף�	"��!��="f�=b:�t�V6�i<�2u�"�E<i\=·��� v��)%�.�����~۶�'l��'0�ׅ�qD/�����Jށty6uO�D���!U��M{�����!��Mtt,X��h�.��J�=t�om@N&r�+31�N>J^
CQɧ�3y�j�X����ٍ莑��hARLx<��ܥ��$&L�*���s�;J�7:������}]A��4��/�ũ�[��v����ؗ_(�L$Boa�q���_&ty�������*������@s�/��%�c�����[)c�(Ր��GE�����L��������t	.?����\ ���nO"���S����]{���7$�;+�� ۈ���ꙇ���Zy^U�U��YayV�Bl�;�rx\yz)��# ������m����k�ž�Q�P*���\FC:
�~�#1]��#;�0�Ia��XG �ߖ�(�w�Q��^�m����h�$Uw�.������;~����L�n�	?�,KwQ��\��2N�P��s�%�W�W񉙯�������;���\��@�
w{�)Ѐ�q�����W�1��<��姬s�!.�~6[˧4l.3w�6����y-i�)`I�;�'nCX��+��J%��ⱁ��ӫ�o�AE
��_\���S>L	��P�dt��P�ED�\��U�?���v��!�qT�8����]?�6I�^��|�Cq2�3�cI PjT�>ɗ����l;����*��Q���P%`���"��@����-(�H��%@�B\ �܇Rw����G�$6~.W+��C��d���9W����к��ڞ �%x��z�Rb�WQ�}~������V���m����rMJ�W �וse��Cq��KE��=~NXf�x�By��s�z����c�"��fB茰�LEO$�N���&77����ꌤ�5��;����G莒�HR΅�gi6�_�d�g�l���T�q��b
0�Ǎ<R�ڭ�Xe�d��*NJ%.B�KrZ��m�Y������k�98���*:����~��an�}��޳�G�6�),^���z�{��״64��Ջ��d�C�[�M>��u,�r[�����@jޮ� t:q��/e�c$�o3�G�|��r��a�g��<GG��Q�^z���[g��T���_uX�G��/W��b�Bn����)�
��i%r �?�$?m6����\5��j��A�:�l��K����f��O�7Q59���9��w���u��me}�d�����\���V�1vS�xR?�4�L}ɰm
O�
�Q�~���i�b�#�l�f�j�/�\1�91�(�W'�~��[���RJ�Y�R�W;O׬�1s*��&m���6G��yC�H�.$+hF�0����13����k8�~�ٓ�mj����K���[��r!��<J|��^��M�'T%ՠi���Ic������~�CZ9�&ZCnjh�-�'V��I�����j���t.�q��{�
�k�4��x=�jDn��6UIPqеȿ�m]����`D��u/V/:�5>F�8��[ݮv!b!�s1P�`Vh��"�|��"Te�����͕�`����4��Q6��;���<�4�N�}e$�� �hu_Ay�k6P�ݹN���og���/А���TD��#�#a>��ڶ��A�벲6h�E,<�ߦ��ج���5��L(cx��5_�)~�iP/i�'�94"n/3�t��_p�+.�JJ%��b��2�o0TcCT�i�!؏�?���%��1�@p`4o��.��,�k���T���>�� �� q��	�x@����	��|�M	�b�%�1|�S��,��3��n2Yd�T�]_�!j#?�Tv�WB��48��0�N��C�C(��bD��VZ/��)�f4&���j��L����@��/L=������@lZ���Oh9p��z1#�`���3�����D�r#�&Q>-,���ٷ*�U���rڍ�Ȍ��n0κ�uo�v�i��'*!�e�+ ��7�W���n��~sR6N�U�!��(�b*g8FC��8�)iN�	��b�$Q��0�O��[����W�������A-� 2DU�Z�\�H���8��(wفخ��-�p �/��Z��ﭦQ������d&�X=#���OT�����H_Ր(�(�ih����4�@(��I��O�NClӘ��>i�U)�:,$.�h�*A��|����K��'.͍�9�rʶ���
�Ͽ/�i��H�_�6�6�;43�����kn���D(	KN-Ȇ��&�$�S�n��׫cr����̻)�O�a������
yva"�4����끿�S��^ݲh�^�25��#`�����0�󟱀�n�Z1����L��a�cC�z�}���\tZO)��ot�N٬�27�,�74�+� ��F��!��~OBlK8Ǧ��Ȫ�L`ߗ9�#3���O�^�צ��U��_����8v��,��g4.��^G�:�?Z��rbU#��X_���y�����g-��������/T*�6K���A{�2SxM.��E�����;� a�vx�W��Hp6��[H3�i�F�����hc�89���]�U��L�e1 �{��&��@�Z�����rF��kT&$���^�P������ҁ{�>�NɈ��\�/Bw<xx${4Zj��5h	��h����2�Q ����q��o����,����� һC{W;�9���T�f��اˏ���q"�2�_{U	���_xb[��`v8u�e^�Y�7��z9Ej�0�j���lu���%Y�^�@���Ȁ(��S�A2r���NC�>gzQx�W�l�.݃�R�E�U�>����$��{��E5�ڻ��I�Z}a�M�)K�����_JI��Y��t�J|�X�H��N�r(ێ/8D8����M�D5�%���� ���Q�"�j?\���\�����z~"[�/�O�`q�Ρ,����[g���Aa�%ǛQQ#���	��1�Dƒ�&k�)R���2�0fD�\�MS�J�5?���G��ɝ��3�h����mM��M��I� f{-�2�7]�$2O�PY����J��YM�+����;;؛�m�A���n��G+���򮩦�CAs�Y���i�)��:Ƥ&q+�c�T�(W�/��~ke�QL��14%��L����z4]4�jy�]�G�^�y�uC6d�F����5G�����."n���4����,�F���$��׼����(~����5�̉�G��9�l�^��wwޣ�AA�d��~_N=���Y������=��^A���{�n�˹���cX���I^����A��mSv�y�"*�8��42���3kY͠����壇K�ϒ(Tl���"-gR�SqU��~D}��O�j�Cy[
�Q�s��rB@��!8&+Jy�۽QD�1�v����<}1 s��"S`���v�Ǖx�$�3�M�f!7/T8:~ �����������C�Vj����dA[��V�C����sD�np�2��&#4 T��?,^@t�L����<�Z�w��H��/+���'��?y����0q�-�	8/$�n�~�z�����v��Kn:��ȶ��'���8k�,8ܣ�:
\��P7�<�it�����,��`��\�	�V�s��b���L�U|P���]h�%S�����O�榎(��2a<%{�����1~��q'�+�M��-O�eР�:OAbH��	��by�7i>h�;�*�Q�����h�mdڔ]tW]�]��4v�ӏK>�5���>Sr�Y�`��{�!�校� Gf5��^܄���P���֋uʍ���+!8*Oj�6rh�{B����}-��6��o�4�:X���JU�
���$?��"�t���O�{pr$�.�M:���P����*�/��"љ�����Yd��S.Ra��du�b�rs�*a�W��B�q��sB]TD%F��4+��&�����:zU�q�JL*���Xb$R�����d����U�L����G_U���=�a�^��lЪB�2�>>�jkU�-����d���m�<�Tĺ}jI�$^�̺_�M��>�# ����6��mI���2& ��b�*V�n̊*e�}#b��b��Y���{!�!"�j��sD��Iل���+E��7ZaZ��@�͢a|p�>Kt���"W��o������;��ntv�@�9&ך�胝g�@N��Z�,xv(D ��8��jh$�ù����z۲��kk����}�|o�{�b�8Lv"��N8)����l���]��ezǕR���
�>$P����<������~L��S���'���m@
��'qL�n�6^�aˬ]&	tVj	>�-/�9�RE1-ꮴ
�[
7(���4�0k2?V�S~�Y�iS�7~����Uk-�<,�԰7*(�:�����]����R������.jH��G�З����Bz�q��ǹ�_yN��1/��o��S�	 �������\��u�Թ����L_���:�☫���0���$��������܄%\��%�L�z�?W_;D��CGlmJ?"X�hnfLI�	�+I���\#r@N�]�h��~��z}�3��v�4GϮ�v�����UK�c�=)�k�$�� �����'��;O�ۮ	Ճ��`u�mtP�·\�s^�;��W�N]���Ok�y��u�t�xh���~X��"*�	@6�c[*
Ϛj!0U˻�5V�v�v�8�g�b���4��y����f����~��F��M��ɠx3�/j��| 0����j١%e�wk2VF���<���D~�$�7D�^v΋ ��>�}�	�{�h6����$a�pW�	�(�O�2����n�=�|7���$L���Ry�Ͼ)����) �Qg���.�m&������s��-��d�@����ר�Q�V"f
D�+���,hK-� �]�i�Q���:O<�R@�}�V� N`�.x�~k5I`v��ر/����-!�ڮ�h���� r������N�E��:i2j^�84��B���K����)��f)�4ʗ�ӧ7"�V�h�]�״'c�GU��^����ZxC9�^�n��H2N��0�Q����!/ʓ��kQֲ��ٌ4Ծ>�>����a���x�^�
���?]o`/��Ef���-*�'��FT�.*�Y���G7#�6�œ��4X��<{�9$z�X@���I�bc@�!w#���n�WkT�0�isJ�T�� ���+F��M�2ËK9�Ah8�I�g"�z?�
�Ժ]|F�~`n�����&�e\ŉF��%�	""V\���,��5K!��}6���τhVH늭�ii���,p�8IՈ�|���7�1wg��O�LSQ�`�U{[Y��0�~l :><!�5�Y�[�tޣŕ�j�?Rv�O�*��.��e�����<��q�%�����&E,�N����궤&&,����/KN�|غ��v�1v{��^&Vk�T��ӊ
��T�X�o��ȷ�#S�k{�o΂���(xae;5�\��"��0�~)�N�묇��嘌G��HG� ����V�q�s�7^�(�k)r�}#�������h��e�Y���S�ʻ�i��IV�V����#D]�w}�{�.s�yվ�R�{m�����9��W�29�o:�-���z#�G�E�g�����x�3[��u������+���LƂ�Z��˿�D���3�L�!.�Fdm@\��0���8��b�k�N-�}��u]"l]+2�X�8}]�-������]����Y3�}a��k54lzCC�����q�bPZmʹ�َ �L��yn�w����K+J� �SNC�0��a?�ΞG�٘��3?�2܋���|��_������?�MWw�Jɷ�����&�p��� ��i)o��*���R�0���3;��y�G�T��c^w܍(���U�ᗎ�y�S����0�w����U�x��W�KL��ρDF�Dy��( �i��P)-�J�s/���؊h�G�	w&ߏc�=4�E���H����P9�?o	C��lɏ����"t�qZO�7ۯ�X2��I��J:����k��s+� )��y��Uk��,h��b��-����:i���8�@7�
�$"���4?��N*j�$�1�e��b2�.lY�``�j�ٝRR��"�M�黇K�A)�Ra �b+�_�1�d"�����=�'��}Q~��3�F���8�fKq�LC�`�e�>iqԔ�t#�>�^�9��҉}�KKk&%� ���_��>`_CV����0 f�x^�W��ͯ�2�8?���Ew���H�nW����$���y�M{��2(�+3�J:f+����0XI4���^Κ�!���ԟ�݉{�����$݄��������8�B�K�ptֿ��r�(�fAҹ�XWR8����x�AI�$֧(-\� վ�����@ɪ���"ty���9`�G��N��x�ܿ�8h�mx�	o)͡��Zu�sWڊ0:�b��m"�L9�fL��Vt2�k�)}��v��x��v�c�+�"~<P�H}z�)H~KL��|>6`��8j2�K���
�L���IH�<΃� 3_,�����Cpɒq��ofg�,�%]q��V۪s����d��O_yE���(9:"E��R�<o�p�Ş,�ǾK��1�ة��Fc!���� �J���H���}�g�v�oɡ:��%{���vȏ���ϣ]"#J'f�-��9Gq�4_��y���u��i�LY>֨�)v�R�A�
<�˴��l�0�f�.���I�FFT�����wD.Ssj,�BJ;¸䲘�5O��K��5�>�v��������!b�D���PY�v˲W �wq��0��VJ�}CIax�0rn�,��aF�{��}z����LF�m��;�Z�v��i�R��Y�r��e+��jq�@ ��%��/�y&�������M蓑>5��ɾq{���{�� a�m�ҫ8^D��A�Ը&���;KӞ��AA�����j���vŶ��>�.�ଗ��Զ40l�1� ����G)=j@�DD�,<ٌ����\we ,d.4$	��cu$��̣'���OJ��O�⭛KCp {J`�w�`�Q?f�[Uy(��R�ƪ��%�v��i,j�X2�(1�+�>E8�����jN�t�l���8K;4�S�:o��:׫�m���@S� /�1�>��f��#�r�7农��0�W�ت��
>�^���\<O�D������N��7Ց�`�s��KE�,"vA�v��>f�n�٪���B�����/���;W���~)>�_/C�nW�f��Xd�R�`O�M޲���x�}PK�����?��%|uC��j�Lh4��L��z�0jn��L��?.Vb2���(�4FXO��?}�'V�v_���ʙ���g�
"��r�Ώ
+�Z]X}��Wۙ��3@ZIj��c�t����:dfX'vCFk�?��P�����e$E%�-](��QSOf��'�V�r�Gm�
�<20h���iػ�YؘH{*�[��k 2��!
��#��l�иU���<�����oxnyG'ۙ�5	�f�eP� ��Y�iB��,�KS��c�M���^���`�wJl�\A��)�A���&4oW�ļD1��_C_��i2 ��E�?#w�wo%s	��䶘��`�����W&v�%�;d��F,�;3���Q!�;�m��k�2��^\˲�wQ�h�\;U���l>6G�&���Mr��"~|�T��]gǾ!'�h�@?�E�W:�X;L#<�:�ٛ���	��{D d-�:��9����u���-���?S�՜�@�ݗ�n|5t�W�>4��ЮW����n�3J���.!���w�į�2j����E �8���6�w����1�ޤ�_��c����%�nr�g�/��A:L�A��~^�e7����R:�c�