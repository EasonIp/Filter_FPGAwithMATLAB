��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc��3@���;��̵*T���që �|c\
��`P��o]L̛�鿕Z[<eLl˭�W?�;���Xo����^����Z�<�F�g\CT���/4�Ǎ�@�����(�Lx)�EF}��N�QÑ�*�����Zf�ϏJV�E������V�M>؆1"��0}��{�ƽ�`G�%[�,s���>�ӹ*����ںA��j�'j��''$���F�Sy�,�v��i^ٜ��/f���.�n���WG_�kQ
-,�.UI��ۉ;��Y��ULCͷ�,lY{
��B���<�����N�CĖ�Y���3r�����M�Y����>c�7)����H+ѭ���h��%nIV���+���tF�)@I=.!�vl�h�06]�ca�+sE��=����`��e���\�i���R� �#-r��Y�Zի�[u}�^i��.�� ck�(����^�]��P�#"LE6�g-��b���j�Z�[f�+!K.�nQF�0ߑ�K?���%7�@��!v7�,�N����y�ߑH&�R���k]��Y�:U%�3�W�a}�P{'O�Cg^��u_KNr�ԼS�q�M�d|>�F�?��ōQ�o&�D�U����'��V���V��c���1�~KF	jN��{�>��Bi'�l��4P��Nl���q*6��Op�4��EN��&��r��5lM6��r�I�Z�1��Җ�R�w�P��U$i���rG_ p�����:�!wuQP��)ӑ.u��Q �v�������-Ra��UI�"%Q�!��°ߌ�ՙBEf��{wٖ�D��~L�p_��+� Z�oZC�9:���g�B�E�E�\u��!��^ȯ�.Nl�}�q��i^"y�jD��1<|�77j�4*�Ygը]��������MH
m|��j�}��G�I�؜�}��*�I$��y�"R�L� �^�{n5�	�/�P���x��ުy,<���0y�\Ѧa��\2 &s4�zi��J�����'��L(ܔ�y�[��P��[�*ûD��3�A�� {��pblq��ܴ��ٓ�R��(X�`��r���>�ZY�ySQ&�<DLTfM�P�����d<+62A�J�p��D���ϭ���UT�(m[�&'i�ٛ�܀�;%����d��Mc7�ŉM�k��R?��a��&p*oޅ~6Wtk��xe�n�W�Ԫ��Z����%T�^��$���b�/II�W�/�����k�$Ry����іeZ���"n�5�5���vG��Ҍ����]�]�Nt���lAc�E�!��|��;
S�Tni�h�**ҁd�="Ҩ��)��۴��dݗ:��V���/J(d����b�ԛƪa�Ai��)@�#�@�#�(��-�|����P1�����(]����
ƌO)@���y�)u�_��{[(�q��m
1����t��@�������͟﹗ �Dz���c�JX�.?��O��'k�ԉ���#2��l��������=9�M�Z��&] �>(�����j�rC��.���_[���������"��|�����\If%y��_�/6��!z���A��0	���ykn〳O�62�f�m�+���d]f�r�+�$�T� 2��0t�F���n%h�C�k�n#=��L��V��L�����_��w��w���$:��	��F�C@1B��R���`���n��ZB<�xq�jX��#՘]&"Ӯ��l2N�g��/���O�(� �h�RYS������3��0�&`�9_*��9����l��79�zaIF�U�b�,�Ą:u�����ۦ3����dUN<���~���f�&��8�P�Z2mm�T��"p��D����:uh�Vd~��Z�Tl��IcW�zlG�>ZK�I�B�Z�yW�z��Y�)���JJj�8�ħ8����dH����h/'dVx?���u���>:R�Q�P�Nδ�EY���<1P���r:��x�x���, c�M�@��]Ȇ�^��z��x
�vh��g�&\���YWrYNPCE��*)�H��ҦNVM&q6FY#%�wlY)��� ���ި���]二�r�2VP�_|;.c�܍ޕh�>tS��A�L!h~�9Yۿ�M
e��IL���z�,�`��!�'�Q�� p4^1yu j��]�=�p���%�d]̡���s�+����%ӻ<���nm�f�xh�	U�c���.����[V�c6�q��W�.�x�r��K?E���܇��Dp>�ׅ�H�]��5N'� �� ��2���haBb� ��JX�P��SA2��~��_g�O��"��g�͝�Y�7#U��g$v�8��:����ʌ�rt�b�8�f�����w�@2D����Ҷ*Щ{jl����4�źԌ���h���ys��1�@�yf��n�}���Jķ$5ot,�{�=3�?���m#���V�b_ ��&�B�z��JRC1$��#�̢���aY���F�*�K\o\��b��F���%�*���G+H�Sv���;d��i' �7̈�}�@y�完��w-[���2�@V�Q%���e"�����r�:)�x����V����*j�Z)VC�GAH�3��H��VO%6��X
w	5z�Z\�<���f<q@yw�8�%U�;�{�O^�^�.��jzO���q���t�c�<Ty������"�ZKKȬy�N�S>ޭ[�Wq�ү}�s��W�2z�ô �X��{^X�j�,ddF��K-R����VU�$ZJH�^Z�嬞�/vW�c����t`�$��tn�����ۧ��B�ݎ�]V1ї�6�=pk6|_�{� �eJG�ȮتW��q<�)�X'�e,F.���}���s��3����.DVg���暌�^�`�z�Ƨ�c�@v5�1jAD"0��E��6�D�R���E���{�yJ�n������RL����9p?hb�9��;m�}���z�c� ��DI�蕀��:��(m�Bȥs���d1#J