��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$��	�LJ	l����D�����*�+^�ؕ�M���[��[��r�;R�e�.3�R!3aw�I1eRjsm�Sǅ�),`� ��+���ߛ�N��!�8?��<­m4��#�?�Ȧ�)=U]������jS�������`�������a��1��;��m��J��'���w�nK��;a�u���hT�?�n������bFA�ӁU�F�ٕ��y��
���yP������C[���T���Wc��5S- ���e��n�4m��r�pH�V#6e��& �hD)����Ds�p:���L�&�z� ���j7�� J�ګ��d/o�JF�2<��4"T�0&L���楬��,]W�G�� �~��0=��v8P	v�o�wg[����A�t�hł��%T�����;�g(M��F��8B_R��bJ؈�����x�G�$��DMy�u)~�����R�}�Φ�~ZL�q��Q��F���QB�������Z�$X�/�T�eb���n�m�{�O�۲�71��ɵ�?{n�O�T��z��ڏ��)����c�:�|���ɕl�鬎���*��G_�o#y%|��ra�5��e��Ϻ�S�Q��6�!�c�>v[�ouy *��q�LMJ ĉo���>�����W
��a�mG�5%�L��6[?`���-X]���.��1�}���o�oE�&�[I�K�O����[+�C��Ӳ�046>����:	��@�;�w�?.�[�)3�hF"�Υ�OKύ�Ad!�PT�O����0�� ��+?]T��5�w��Z��u��+�E���:̙̤MuR���q/�`����7�X{��s�������J��^|5�d�# �������p�V}_PW���O�͏�<�`Y�\�z���i
�@��E)�G>���F!��p��P"�n����z��0r�淁bU�k���Y��Y[��U-��vv��3!<Ĭ��x��%��V�^m���� ������';D��ƿy�������Ѽ��<G4����-�Fd�퇚��'��e�����&=N�q'F	�&)_��^=;n�|�Ȁ�v`���n�7�B�mhA���(=���,�~�"��-).4t"¼�ӫ�ʮ$�5�qf�֞�=y���c�9J\�&��w`�%�i��'��|J?�_��%�Qc��q���>zF����;5y�B���)�_@[�bj��^̈���i�/ªݥ~	Z�6��_�<l����'�aT��ݦj��+��k{��@��jW���gL�bOz�8_;&�P(����M�����U�PTo�_��(6�y$��b��R�|4�����)|s)[����M��<���5�K=O�Ѵ<S�AP,�����
���ίޥ����
\&Ć��]�T���3�gC�M���u�i��?<�"��7�=oP~wx ��7��ت��N~gg��6�½�^�p'W�"LG`���gܻ�5��p��kl�:�y�,��-'AX�����CDC^*ȡ�-�jDٹ�=3y�"�Z�G5�HSi��;��:R�C�V��C�2���I��+(�2��y��	d�M��U��w�8�N�?�S|kEg�uIb�U�NQ{�%N;?z:@́��a��J��ϧC0?��;�L�[_nĭ��>BvO����I� C��mް�/�$��Ke� Eѣ�b�4[��p�Tc���QL$�V-��y��󨋱
ER�nW����;�ۨ�׆�&P&��F�$�$���ͷC����ޙ������Em���H���٬���F�j�i�O�>�v�6���_Gc�H�C�	J·��>�d�����R[&�j��������.�J���^���C����f�%�w�&vs�[
��-u8�CAf88�f���O}�}�?Snq
���hB�(��[XQ=5�v���ָR���
��#"c׎59�q�d����F���)A74���ͺ����{�NY��\�p�
Nݐ�xAyuv��t���[]2F��0! �jl^ �X��up����/�0��ӌ�]E+,.MH����\@����e8�4C��5S����;B�w �V��-z�H<䧲;5^j}uP�<+��+6F�M���*ݩ%#����4 �"�3��A�o���T�g��>���`hY�� z����}����� �눿��u��Ww��4����4��@��/+�=XU_]9��8tiɉړ[D0����?dMؼ����*w5
>#Ueo���x��H�M���ha��I=�j�x�i�MJ(�\Ũ)�"Oz��Vv�O��i��(G�X�b��m�"�������K�N���!�k[8����������tMl����r�D��'�g��L�YV�Ř�7��?����>8��Ev��f!�ߊ"��l#�#��Uf^�վSD�<���n��Ϙ1GPy�x����+u����O�Z!>ǁd.p'���� �Z^��?Lp���\˧3�ߐ��$�zS�rF\L�)$)��zv�e��0-]����ILeҞ�*��#C�_�����W�}D.W�\��V1�S��7[`X���m��1�l�E{�V]��bP�8�������%�y�xje&a��%V,\k��: �ǀ�$/֠���*����鰐a�����N�$�jMx�Z�_� S@�@Jr+�"J�C��!���1X�/�e��Q����.�/�v���D�hs"�P��_���o��;0��;VE0��G��ܧ
�uɝC�����{��נ1�	(��|2E����|�C>؍y����FN�E�P$8R�_������5oqS+l�D;�@N!j�K�OT�T�a�Hټ�� dG�i�`��j6H��4�q6�7�(C�iu�+L��.����"�g�di|�ێS�>�jb��,�V`�^��QB���������A�ӚNY��v�uF8���n%l��1dx_�.bv����=���u�J�uk�����7`�eȧ����q�]���͚�C(q��`*��5�)�s
g���g_|��@R,��q�w�'�W�Cإs�4�W�6v� Ͼ�Y�:�{[0^C�*�flw��=�ff�n!o	q����t�d�,Ұ�Y`f��{{� ~��1��گ��d	���FXj"L9�8k�v�ӹ����QH[z���r�յ�՝�mݶX+��[R~Yޏ��:��"йF[>P��]�L�:I]Ww޹i�sj]ps�C�V5"M s�W�_vv�׈��Ov$=�	ɕ�Q �zd�S�'��W��t�A�ŏ߈��ѣ)�����a��,��̛��p���+$���i���j�O�ͅޫy��	�K�U�#�h������xrrrN���H���9��L�M��f�1��=Y�~��5oY�����Ηz�ŵ*c;.�
(7(f� r�Y��gKD���-z��(*	�Ga��o}�ޤ�6\˓�#��9lq��~�H�|m�V2����h�q��w�ui�G�HY��x�=��`�d��^PjM��m�\1Ȯ$��$V(��֙
?���c%$�}T��ewƻ^��<\���Lݴ8��Sl�T���jܸ�Bo��>ה��r��_�����������&}
"C���:�W��a��@W������- m��4աM���F�Lp�)���\l-�Z��'���F�Bq�Xd��0?�J�{�g�3�"���h�^F�)F'��r�Ɉ�4;D�����
����if���R��4����F�%U9XI�1�D�^ñfS���h��ZQM5�1qVL	҄�7�BI�k-���f`�̬��7�'�{t�˅�^��q��ցh8k|C��� ǰ���H�U��S�{�/ ������ ���F����2~�Y�+������]�2���;�e�5a���-z��Yˠ_[�%��q���TM
�>��(�c�6��n��[>Xh�d	J`.�����"J%��&��R	a;��B�,��ش�%���h聕RY&/mc�Ư��oMf�����gN��Z�o|�H�f�@��B���P���S����uaP�_^h��[�z��)l�������h�af�8��Ʃ5#��]C3Z�94c�
�ٺ�������ۺ6�U��|���[~�Z���5�_m{��/Z���G�o4&��Pj=l����M'X��5�1BC�?x����P;G�FҊ�Ďcx�$��D�e�9Wh8�U��Wf�?;�ee\M��v���+�
��Uʔo���Z�BI*�M���
Y�46�Wq�x��L��;eƓnk��V��B��>�����Nbۂ7�n�7{�ҭ.&t^OѪ�d��^2��=<��!F'蹖�ʩojo^����oU)��T6�>���1����F�ѷ���̰Z�$6XҰ��{sL��6�������)sA��4;���V���!@��2i��j��U���*	�yS�r\B�+�A&Δ	�m�^�-J����6��1kԬ����6�������<�0@}xwH�x���W��M��P4���̜�ɍy~Y�t%4�8BPC��R�?�y��&���S�I��dpn�[���TY�M���d��K���h#��*����m�cg�ZP�cn�p��dT�@�3b�����S���F�>J{�T��ZC��&�Ƙw;FH��(?�yqY�<����c�ߵv&q����9j��%���j�@�X7#.3"��W�v�C)���-B%XT����1�G��b;��4�{�16�2&l�R^��\�6J�f�n7%�d8�<o�^���#&`�`#a,���S�Z�73[��Ψ��.%4����q��  Y_���=g�x{�62A���֥�_NH�ϚJ-����a;��4�=<#��çl�$ۿA���l<��-�NH�:<O�mR��A��=O^9�ݱ���u9��E�:E«}���&��F;�]�U.%��w�m�!���B[������A��&���D�Ƥ��Q�-��kn��*�\r&
fw3|����8��SOl��uw�f�`z-Ol�N���h6>nm�0�)���#充�yc��Ʋ4pW�P�~NIY�����T1uV�V\�[i�uP�C*-��l*��+<�_���iɕ-?*�O^��Ϸ�I��q���c�����:�Tq��SȻ���UC��/����rA!�+��p�l��O�~��v��EO~�q����u)�`�k>�/p|o�o�����?��<�/��^�I'��9����+^h�s��whck��:���p�'���O��&�dG�/�;�P�t�8}���LZ�}2�~X�I܄ʆҋ�m��u���KC��{D˨���fa�0e��z�u
��q�VTQmq�PL󍼈7����(/���V;I�<}�"���Y�N����H�"�Hj�n�(���i�=;ֲ�+����C��He.������6CD�R�؄��G�s�3��@���h҅�o<�>�Þ5C�ru]���P\F��-eh-M4>(+�%�P���mM~������';�:��*[֞ �I"�#o@��Y{��f� ��,��~-�Ɩ�Y�I��b���./��)ʶ�%�l*��R�Uv`V�)���%
�A|�XK�a3���j�=Y����g *��͡أ���G#��H����hO��|�.���V���{�4*I��AD��a�dw������R��Cm�m�%ꏯ0����%}[(>M#�: ��d ]��ѵI�t�EK�c`��T�����h� �)z�I�zs�VsG��G�?����xK��E0H������@��:u��86��Eۤ䧼z�U7�v�<L@�w�*���xA&K��9��e�N�[u&]���w�Q�B#Em.XA���
�	��]�t,=��g��� ��YҨ����׽�m.���#���U��*����[p��?04}To7:9�	8W/��3dvf�y���}s֒��|�{i����Z����([sƴЂ��&WX�_����T��u���p��& ��pV��3��񨚤�X
��3���+����&�u:��4�ĩ�����:=���Cc{sEظ-ޙ��Vo�>��v]#Ǭ����G����*-�_�C�C�����>f�с`�@-��]�@v<� �e��
��hC1�C�^�DH�qb�0��7$�e��ɧ���	X��>�:���y�Q�F��;X׈�k����L���u��Pxo����l�sڅ5�F!.W�i����ao'bՌ��~��}sJ9a��F[y� T!b�\]Qe�o�2��X��nT%���,3$J�3�jSXVQZa�$���E@��/�TA@V:�#��?�C�����*"7���+�{K�fo��>�څT��q�нٶ���e�%�X���)S-|[��7޵�$˱n�4�� PB/�/utH�j��a�4b�T�:2VN�?���.�@�I����o�tku�=�wےg�%E
�냀�Lг�!#^�?����볗E�tK[_��uyg��<�{X:�r/i/���/B٢\!j�e5Hj�8Yu�"lg��9ʮ�L����Nqzp�תs_uj䷗�/`�(�r�x6����<Jf�ʤ�q��kŞ��w�/f�E/cOO�"6`�b���O1��Ef@�&.����(e��~�!��g�|'�S�1�3��j*jhX~�/g� G��Ї��?���dt�{�9�J���?�ɞc��JdjשּN���p&��V*Cȧ�)�n�c��k9�{���/�Q��0Ay�d��H��3�)�S/�S��J�5�	���z�_�_�����]$�?Su��������/a��y���P����Ic6�D|�Xk�\����4B�qim�a2X��N5�JYI��jWDV���K�}�3�!��r"f��*����Iu�!^����F�!�sl�/�I{%p�] v J�j��Քh~�1�L^�� ���\�.����!���'��> ���
��J)w�������(muфf."����[�~c-�9x����>]qC�Z��4'����:��9�T�oXcF
d%��;�K��nx��^�#�ng1��g��bh�NL�B�/�����e��������YgJ�?���"KG"������mG:���;Q�=	Bs�y�&4���"ǆ	���:;�"]��`����>���j�X�i(b�A|�����E���3?	�bv��Q�h :{wT�WMj�2��+�1�F��)Q,��/�+3dPi�-�?��ٲ��N��P��V*����w̎��ˉ�L����$��t
RM��Y �1_m�p��JD'��1�5E\�����Y��H�v�r�Da�?{-K~ΰ2�va��F �9z�t���^5�тM��Y���^�!�0�x�"�cfl��eo2�׎�����~8��Ydw�\(�~|]���I���c*��%�f#s#�u��������:������}���r�����ԡjZWv5ts�j�����;����wǠ��/�pN�x�*�i@��Ż�<'��#���)X� �2�k��%�/z�Q�JP�^�z|�b���Q�k�E��q�fj���uB�c~Sg6���>9~�
.N@Y@-&���*� v;������\�o�&̲�>�mV5X��W/I�n*�l!��2R,^T���௒�Z�f���i���3��������e(=�t������3��D��!�$S�ɣU���:���M��E�-0���P�E�<Gk��ԟ����ѿ�1`!Qd���7c;(��*p\��Re�Y8���q���2 }}iJ��ԗӎ������oGֱɻ�Ѳl71�E��v�k����U�4�%��A��zS�����*�c����6P�VA%Yz�f����Q	d7��g��׏�*������%P)�
����U����]8s��g0�!�C�'�ֻ8?�|Mu~�D���^�;?ZIRE`,)��x�8x���r�v�Z�V���ڡ�I� ��s> H�1/�^7��?����c(c�l�a�TsB�9��,i;.��A�H�$���3�ru1É�˳8�{�:e �J�S�I��S����V�e�'�׈Xm4�R�-Ʃ[�S- ���Ls�E����"u	l��utEN�Z����Y�f�n��:�'�ua�_0��c�L`�K8�ĵ�oy��6P+��]�t�X+;R,vZ��w�bTO�}�1D�1ˀ�֙�oI�!Jl��j��v�e %�ߋ.D-���
:2�-	E��X��:�b�7�p���2R�N0� )���?̊�O�̢��ca��◳�b��!B�/��gf�m�>����N:���>��S��ᱴ�O��	�K�*�20��b�3�4��ܪi�:p�E/>���:�u����w"9>��3�v��K��:?2F�D+�<׳��UL�+U��R��Wa;��a` V�A�Ir��\�xN��A�`I�
O+w߲���+g#z��pT�\)+�$�Yg�}G��!+Wm�?�Jf�U���X�7(�׭�;�z»�t�mٽ�������>�[p���Qlh�u�ݾ�{�!�Ӹ�נ9����~a(�r���p��V4撙ԑ�,��pZ㿫`�RD�4^~N�yEt��n����ª�l0�x��C�%�Umg��z��ES�tj�Ն�(���L��F!)H�O�)�K��B1B�Z�y8�ٿ!����=�;0zB�xD-��7V�/�jYT�g��u-�E˻V�J;Ȕ���?�6����[m��w�9-�IUwY��?F��n����'z�ch;��.�&IO��u�k�rd�ߔ��0