��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4d�#尭�ǕmpC��՘���z����m�0��X�fծ�+oa���}˗!i�v�:¢#��������<#}>!�K֎[�y�����,�]�glfs��y'Myh�ܧN>r�|j����'n�XZ/-<P?�Ah!LQ�ս�����]�aI�aM*�zZb-���o#��̀PZ�|P�	����ŏ�G'׼�<�-�w�.y���R�$Ei~�t�8�ix�98Oe��E���A�?�o��5cxq"XOw�at�"b?�Ԍ��'��nh"����&̆�h���q��2
�6ε��|����o&���'ě�V��G��}m�p(���Hj2�ItINB��W��&XF�O/>�?rf�dcGG�[���+��� �S㋑8Th��$��w9G�?&��9�����~1���v���u�9r#������۹��v��?����PǴ�q"6��4��}�˶�>���"��"!��;��?E<�d�zI,K��}V��|t�4����\�eM�rĽή4*.��@qɮ��&K��i���d�&f��"{:;���; �$(,�x��^a��F6'hd|�v6A�ύ�\l����Y=�Gd@N��4���D���F����ϹY��R��\�U'>:`E�9[�����1��9y�VD]��l5��V�:R9�����\��2�U>k�� )v
�י���m?���M�����@�k��B�*r��ʈM��J��&x����b�G`M�6�Jóq�h����ϗ�h0U�>�:^�8ǽn���n�y�Q������%ddg�oaRG�Ԓ&����,jj�ndD��3~��b\�÷���r�,�z}"K�����H^��_D�!$
�̘������N��;�v��AX�����\�o�lJ�e��:z�q���֖��X��Y��h1�e0҅@�?�.e�&m�L�R�թK�f"B8��5��_x��5Cg%��r�Q���
_4��q�qv�F.?[9�D�R��i�k����=�((�?K�����Hqݎ�)���W��f�G�U��+�,�)\;����!*�	�� ��!� ������	3ٹ�|��(�r3���%6�����Ӡ��n�T��]���POwq*��s'���ł�7�N��}�2�_ؽ��Y�AӪ�3]�M��E���ER�<0Pc/��4TLWd��9�v�IX�h"�%�B롿�D�)��O���/nG  ���� >�޵�+6�K�����a)@�>��Ӱ��a�ܬ���s�����h��@�w���v�ʈ�\G����9s=�-w%'�E���l� �8�}�X��zɠ1W͏���}t<��!��"M�n�z:�gp���p	h�6 �h���(��)bIeA�;nr=�(�_!�q���t�i�+X��}T�t���X��r�=}�m�?�?k��օMTe[F��T1rl�+�"?��IR����YR��ߟ>�H�&=�h�G�v�i�3�n90zn��+
䛈nQv�Φ�Z��,��^5����K��o60yF�G�d�1�Z�8紳yq���	�g��2��OgeJ���,��p��@}_���cX�G�������fR��]����"���0�Z�������i+W����@�窙��$��n�W�����Ѷ����p:�X�L@�;�}�漤��[-��8۱6����a��;��
�F5(�h�hF3�QX�}8�=�(�~ֿ�d(50u�.��)5����~�������2L��Xˏ^7������3����ӓF0��歿#8���@��p&�r�;t�y)�/�=P��SI֍�<����������_$�ߒ�%n'�TF�(,)�C�L��,��0o^"�U��e\�}��G�Z��
4�MU0wu��F��B�R�>��i��l5���n�^C�>��yz�tz�:�w	v�^qB�P���Cp��i�az���5�a�a�9�A���\_�I��|�M�ӆ��%�E����<<����2���H4����K4���r5��ތG�J�`%�6!�f�!Ч����o�0bk�|6��F6�M�>����N ��ZtRg��HF��D�lƎ ��	5dD���Q�.�x�Xוs�gA�:�K�LS��z�N�T»
WK�������Ŭ�$�é9|�>�'U�{o*�蚿ֽ�E@�l��w�K��ݖtM:�&�iȄ���'��=���������L-�
�����$6��	T:d������/w �#�gK���1�ʾ5���b�+>:Ag&GKF���_�*:u�S��~}�
@��K˧�:�%����u���v�[�@m��lK�i�{*�`i�����O�O�2���Q����s̭���#���m����]�.�n�10ȏDS��XM5p��&T���F�0�P���*9�,O���s���.�𣷬W����s����;��uwV?g8x4FnHd��x@�!�nn*����ڹxR<������^
#+��C��gK�S�y�0���{q�b(�ΛCq�H�1�np�o�$WJ����2��15/�*���i�� ��T!����_�1L�`��my�.VF�+@-����15߅�lx�-������+������JMa�Nϒo��m��%^����3V���<.��҄��㲚ex��?�O-����(0(��Fk�ݚ:����9���o�j?�Bܵ+� ��WM��z���˪ɴ��>�6������� QI)W�@|J����v�C����?凚Z���(R��Z\�}F^u�CI�V�=�����C;�c�L��UN���i�P��v]K qS� w.;�p���C�<��h�֠��Z�/W��!WO�0i9�R����;����Pe����/��0�FTX�i�	6�2�鄪�y $��Uq�Ed��J?����F�#v���U�:�a��V��_�<! ��q>Fa���śiL^x�	�H%:8�Bp�z���i���ᑴ��'����p���b�J�<�jʅ1���~?=��>�цڐuy��q�F��1OY�!�+(2_j5+N���^�HV���/�gQTkW��B.���b�%��uζ���
���wNW�����	"~x^�����ƿ{f��E�x ׃��C'(��!�b/J�C\�ᄃ�̲���ʶ�x���0^".�'�,6�[g�2W}3 ΑG��v���)a���x��è�z�Q�Jdv��?�2��B4$��=q0iF��ȴz���DQ�m��F�����0kJ/c��}�mv-	.oH
]�i��FDu`$\uHv����|ŗ�eZ������A������G7�j ϟD�wa��i(����p��,?�m)�ՄG"M3�ٰƉ�n,I7SA�c%�T�RoɿG( L��\����-��c ���19[!���A�;Wx��v:�q��,R�lGp��H�����g�N`¸w9Չ�ȽK�	tHO�Ӗ8��܄����s_n@��]�ÓqW�Z��̅6-Ek3}��/�]���׌�A��ۄ���}�.>.�Nv3_`i$ʩ'.=̘5��k ��QGl��i�hy6k*$rZ>Sw�v�4(8D��=�2PFo���H�Ky8�Imw'�wp$;���F�0�P'�7]n�z$���]cv 3mZ��f�Z����x���B���}Oxp(+�J+('�A�fd�iN@��м�y{[e���Fc�x�Ra�<�98F0�r��2XW�^�_�qf�S�{h�L�D�kB`����=��#��ؑ�	��yk���d�&�hxT���r9���b�������D�rR#���W&����;1��e&�542q����+�/�6Y��ד�.q�$
��o'"RQ�w��Y�WZ(@oͮ^.U��`]�����"��<#�U&\@6O^�֯16�!@��y5�b�D�`��4tCVE�ē��{�<)�\S'
�O8�ƄIﲫ����I��?j�J!�oؔ���3,3R����69M�Jqن�<��X�=� �!y}�8��_GA2ٸ�܇��C��0�S�
{R�J�-ݘ�O٤Ͱ�����_'$�B�jA��H�(F�jv�+�ES�uf�)x�0q�Z�gp�&��.rR:��'�M�|�v��D7�$1�Ss�[�ǯ����F!"����E�)����bX�u�W��cJ	zX�^P? mX�r}_e��>�Hi29�A �5�Ҍ����S�s������g�������-�|#* ��ڿ�zJ��
w�v�lH�HSKr�#s ����~)Q�U�
J��~������\'��,��G�`݋���~d��:�A6����'{Bll�Gtf3X<��=�i�A��]��ͧH�g-��� �u��l2ʏ=G�:��ׄ_����E���3�#T�5�7P��=��������J�&�W"�׻0�{����Ϊb7=�by�(2�n@Ű��4Y��/�����_���1!�Ԁ��ĵ�a&v��x� �Ƶ�e�-Y�q9E �xoP�01v4�����x�&a��R
i����->kx9���'��%x�8�m��Y�t�(��C�@��5�˂CP<)) �����	�I"$6w���#G����?�=��[�T�Jr����q'5����~/;���9��<��i�S���/}����'ۀ_Q8���+`�R8h3!�S�+�B����5���CMv%���&�uG�ô'��J��}@�l4p��~9Û�V��?밙AV��?��wC�a��b�^�G�r0�rə�D�S�<�1Y������8wh�t��p�������{y�.�=�]N�[��=LL�8�Ҳ�N/H������"m�	���F�}o�^�QTL�jN��^0~WSp��uF�*$\��V�#�h�Q� ^��t3|��b5�P�r�u�۪b���Ï;����� E�U����0���S�.�-�Q���Eܼ���3p2��P��l"� ��ы>�
̭�x�FBF1�f��H�=��a��Z(9kנ��u&��i��p^$�!p��y�P�?l���w��厁���]|)��z����;��*۱!�Ӝ��44nXQ��}�:��� ���<�o�lT�߂�K�8������"�����'AH6d�g�6+������p��cq�y�b+�Q.c����4��
NJ^�%:��~i_8��VV}���)�¸��q6wyH!�����Ƒ�������ϊkO�ȱ%�Ps��N�S�z�^�c�3 �ۚg�
J�~�ko�M)q9'��J_f�rm����#�C�!]�������ᥫ�A�٘	�h`��H��� � ���wߩCL���vr-b"9"V~d0��z��Mޓ?�3@\t�v�;���O�y��-,Ҋ�u3u�/�٥�����9i�!ys�-נY���5^��N=?@�^�Xc�p/�����6.�y�!�����z��Wfm����D�y#�#�RQp5*�����Ŕ9 RKt�}\8WD�������4㈹:n�B�LY�6,�Ư�e�r�:����e����%�X>�_>�jךL~��n�����"P�$OPI��0x�8A��(dR{x��|$W#،&��m{hw��_���O�R�)�P��,���lUZ9rb���3�W~��^;��$�N��/�q���Vn.R�<WzUJ�)~�R�̵�ȉ�>�y�GC�HVB[�[l��g��a.���L�/�[�tH���	��鿋��@�0�7���HCx�v�*PLy.	<��Y\�k�������T�J�3��f��vկ� #��;\l7�z{"��y��r��m��o�i�/�B&�O�	�%����\`��Bn�	�7��ke�k�(X� ƞ-�5���֝p vs�Y�&(n!�@�HH����p3/&&���+�X���A?DL�A>�-
���.����x:ݾ�����]2�^�w<z����k�w�Sd��:���J��!��s��Z�
��|��m�.h!�F�!s]Z.�9�c�+[C���e�_�w�hVS�<?2#>�Zs�?
k�M8L�:�8v�H88
�Y���U����2]g����ࡆ=��Bd� ��3�!e=��4��ޱ�s�y��\N���΍$�-x����K��c;U=)�5��t��,���� X3���Vw�W�?F��*��p<�s��ň���⍫|עF�Ҥ��W��qs�İ|�=ȅ!���g_�v��l*�F�0k��8L��<�0���D�d^嘝����hF���IYXV�Ɯ�ъ���(�K�Ԯ)���i�-����Ly��b�xvn3����t�u0��8���>���[2���G�?�v�9A���~n`I��eW��X�U�%��u���yw9֐=w&���|!�n���?����3�g���[��}�(�$��[F�1G��܀F������͑Qt�l��Ӌ� P���%E��l\�L���(l��Y+�`���"Cr�#��r��ptEA��Ҏ"�L�bO���+{�m���<L������};>ǏJ���/*r; m��5�5r9�����/�������p���4���Jl��sd�p���z�6.�o��6�O�\�we
 �ns�lZPjy�B���:�t���Z��Ά�s�¢���.�.3![.W#]�,��9��k��p��QZjQ�p`|�E��Vj}L?�O�<�)ι���I�tRB2K^��v��8a� )n���:�Kt��U	��=y���� �ȱ�<)�-3��/�k߻ȹs1a8%_��T"���
�))�XJv�"��k�,��f�r�{�����!�A$X�7l�ε�̌��{��-Dݭ*g
1���������s�B���{>x��nH�7]Yw�범�	��q��(�m�y+9K-f0��a�69X/��l�l�? ����D�:DU}M�cb�<cra҈0����E�G�^䬌 �充.�J{�:x�g�详�E ����V������p�3?���mō�� �#����V�s�w�\'�n��|p)񇰥��
���,�DO�<{x��/~�ϻ��e_�꧃����P�_�iG%���w������M�F_ס0al�67��:mbkz���j�|�R�Ua����ѥN駠h���q����]±J�d�H��`+���l!l�z�l��J]3K!��҆�����bM��	�FM�TG�.��=!f�BA�Y&rZ}k�SW(�R�ܥ`�rÆq��L���E���1j��*��x�r���n�ee�;Kf�2�ޏ��i�W'����t(�]dM��ʱ/;�����i���b;��'*�5e�{G�u��r�)���m<�2oO�!�9˲�C��/�O95,~��A������2$T�5ȏf�%R��:�ٯ�Ǎxx��O���Estu�QO�=; �\-Τ�@B\��N1����A�Z��<ǥ�u $��9�tXܲ��8��ȸ�ڴ!+De�pK��=��G�{�hJJUc2��it�q� ��}O8�<5�Q���է��`\t��#�X�ܯ굢R�(`ސ��2n1�=>�<�䲐5~��q7�,Y����]�"=��5��rzR�Zܦc㳖z�k�U�t# ���|��zj��9�s��[�4�i*u���o�:;u��Œ�Nώl}Ѿ��?��~����|Y��H��.!����*z��.�jW���ЋN�43uˉ�;��&̀d�B�g��td���틿 �;����J�[�:��_�V����ơܹ�f� �Q�K��0�'cGUq��0��0>�S*��k��W��]�D��$�,�q��}7�?<���1$T��=Nfʜr������%l��J�����O.�0Xq)=7gQ|;�@Oh\��JJfaNve�?�r����R����
��܀�JΚ��򣃖^�,�����~�y��?sy�=4uJ��v$���pżN�P �[W�qA�����]|���C&����*~2�yfۘ1j�a�8W�6R���jFMo���1\�@����j�#�V���|'d����q#E�פ��`G�K`}�t:%"�X2�Pn�� :�����A�FI�sXY��E���_	�9�g�wHCy�7�/M�g� �`-�*�/�
��A����?�\r�c���T�OT��<ŷ���$���3�|�����0�=0&��{`�f:[�-���X(�a��)�I�غCVgVV��m70+�Y*� �rR�������yOmA���>� ��U9pv���5$��p��(��'N��܉�S����w^ҷ������h�ww�&w�)��I��7�-�[��Ajp��Q���l��.{��))N.r���H�}���	��Bl��M�����L�ʽ��黎��B1�d�7�1%��>��*m�m��_ 5V�Yj!�:i���oĤImM�἗K|qS��9nT�%�f�1������
�Q4)A��֔U��/��