��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�J��"4�=�7(�T�JѺ�ő��,\��s���ӣ�F�؏tlu
��¹���>X�I:�;6���u� ���R���3I��6`��p�=g�Ń5��1��I��i-yz��.	3�$+�u^t��!BLԄ�A-��J
�q��������m҅N��8�
*0������Մ�)\�iG���i��݁�n���_H#�[�k7���a�`@�A �}s5n���3
>O)�Ξ�����{�,i�1��%J���H�/���	� ��,k������d��h`s��g<4^�sP.�KeB�^(��{�by�$��7���M�=J���hӛj�<��6�G�4�D�D�����_��XH`�Ĳ�D�3g&L���x�,��{��[�6q[<���T��_�`@�e��U��'R���gvI�T���5TUSH����0Ƹu?��%6P.��*;��ϳ�Ez���3'e�ѡ(׆�fL��N�a�q��f�aF�Ԩ�9��z="��O.�i%�jj��>�ѧr�T�`��dl����GG0�z��������J�
Rns�8�ɓYc��U�@��{Ƹ��m筩���Z����c�l5��h<��� ��?�cڕ�"g{Mzt�]l+ղ��˘�^�E���1TS��:b��t�p2�t�nG���k"o���9�vI����V�X��}t�E"*�[b;���g��V�s򾵡8��8��rؘBn�zL���+�)O&����w{�e�̘�'zg���o]Uq�����էے�g�t��n�����j�S�AN!4#bW~�֌25� ���iLQ�U4��\���,}a��4����\br(�ݰ59d��G�+�9jhfŃ��p���0�<��͡_:��B$8��n�<a<���]C#]�q��~0���.��1�Jc(�By��*ra�Y�t��)�[��?�oW�tNj�lr[���֓��J JQ�AC2��������!��J��q�ػ_L�G:��Dd=�l����N��|�`HB������x
�{�����%�=�w��%�'w�'-������3N�@}c)������5�j$=�W��#l��mĴ�q��@��L}�c%��܀�_��w��N�yJ$�.٭���\f��Cd$�9@�ĝ��@��:�#�]��ھt���P���l�u�'87�}�b<�~���?wu�,��o�0�jw�k��5Eǫg<5,��:��Pf��q���9�%�n�UH-0��_��'��9یaa�����uԱ������!�վNp��G^���m�ϒ�Te�Zv2;�^�v9Y^VV$��������C�a�K@�z\��Pc��X�
'�D]U&j�m#�3qL��Ρ�pA$��b۝��{�?��cj�e�p1rw��*r�}����{�g^�`�3��9$�,=$�\FZ����q��λ�#���
 F��!]"
�T�h�k�EY�锜ڢ�Q�2?�t+=�4�ߞ���>1xbq��x��)?EJ��J�����Nrs�k�nx�_���[�P3q�qه���թ�hEX�b�����)3V�lt�&	���T�d$����]{y��-6Ϥv�����^wɫ��F��,�sc7'e]��~3�=J=ץ]��۵('V�""�/#0l���d8�	��;K��ti
Z���G�괤���Av�0$�j�$!�2���'�#
q����Xha���s�tW��D����Uf�t8��,��[�����ݒ:~��Xhh�23�D}�ʀ����ԋ��.:��!�46&'�PVZ)��--Ҽ���NܖL����� ���vMM��$YU]a�l�%�i�'ٖX�����X�N�%B.{�A[xΟ2VC4����7sb|E�Ďą��u�R�S±��ě�� ���8���;%�l���uAm�..�&�1�
xظh��g�s�g#��>,z�V�������&_tЁ⍬�;aa�J柱�@W�SjٶhgA��Y��_S�g�-�����[�>��y�����:3G``�k�vp
����H9��"j���[ኙ��z��N?`��V�)����J��;��~��7�X��o�)���F�!YLE�P��I����n��W����v4
�ZI{l�3��U�Y���l�
n�/hJL�pT���@�/�%˧�H��Ǚh��.�����=�7r�x1<*u.9�|�ze_�`|�6��.1v��&K��kW�¨���k�}?�o���M�-�m^r�z�"&O5^�����
+9�Ӯ��c�������m,���%p�M����Y�{d߫=�Y��p�����aÝQ��#�jE���2}!�k4���ƞo�������ů��d�r7��,4�07=hU�k�����q�>)¹y$�1�!G�^�%���ShH��0�%�{���@#4<~�"�A1��m�3��%!��	
�Q�g��r{�Bڑ�w�ȴ�W|�+��&J��U .s��Ky��2��YB��5=�ޮ�9���)F[k��4��Ua�]n����Ďq�-vW�;�B�%G��I��v�|P����-�(�u�<��GS�u�v�e�LmA9���ʊə�ṭr�Q�\K����s=��-�<�Wm�
Y8�Z�����+&�+V��5��ւJ���-����O3��!��GL�[�o?��L`��?��[�;��^uJ�A�4�p�D��E��c5�fV�@�V��������c8H�^�,+!�:߰mF)�E���Oe��R��%M�2���:3�|���q��^M�(y�vɦ�K	\���BvŽ%����.W�>�����K�����)�����x�h:/+D7��V�͐}�GZ���%朩N���7��sM����MX���Wn^�7W��7�8��$�.���Q�!P�u?��Ue�OPN�{?���2��,�1:��Q�sW}Oֆ-��{�x�f�:0�����V_]ְzE� �S�'�/Y�+�2c�I��S�ī��/g���.a	$¥��l٠����H��r\�uZy���)	�f�O[W�������/#C\��cBo9P��p,N 7�nf4�{���q�#��W��n>��>��r4�E#1r�:.]��&�[�";���oF�W�e[9Y$���S��N�G����:��Ι��5�"�'{��++�Mʿ�b9M!�*6�F_Bu�i�7m���P��, �:�]h�ʇD�0a�7��Ufp*.���0����m�����6��lbN���V��P/�Al8d5���y��lDd��V�%�����/E�Tf�V���Z݇D�Б?%|�d�40f�K�����BT-*�56��ð�*	�Z�:�̱����Vi��n�X�g�`��c�S����b�"�H�=T�0x.���D{�v����N��+椞>��T'�CK�EKcS����J1�Hϩc��UP��d��./X��1"U���QBN������<�8-�b�1\_�s4���t�=�\9����P�j�����c�_�A�s�! �!�T�������JEw��@o���wb��Ѫ��"!RS��y�Y&��[3�f	՜H��4|���_�7�,�g`.���+�c5H*��A�^nftL4�	��K|\�57Wǿ�����J��k:�?�O�Z�+�	ב���Б�AuQ���-�kd"NP�i��N���J
�t��)����N��!�n� U���k����,@���z�V��:��|a����B�Z�E%N)�Ⱥ��E��;/���qA��S�q�B/8�!0N���^�P0�m�0��4�?�J�>�~iK{�� �������2���|.fdF�
Jb]�1�ع5���K*铑'�^K��@d���%�D�(Ygb4���}��Ql&�3�Τ��EN�s�<�'�����Nۺ�J����U�?�C���JdW'�}�� �Wt�rw�+��_2�3gI�ޟ�+�w#��N�H4�7�۪&ՅOH�3!ąJ�ӡ��o�X��/R�S%E���a[��=ZP	�g,}Z�5�1�|9I��<8DIB��&�	4�r�c��[����b��,>:i� �oT�,���V��.��Wpk~����|�&����?*�Z,�uu4�h����@8h[�O�ٰw��Wt*�N��ݲ}�i6�YQ�ϙMʤ �͝���eÃ�:�Xp>���/=K�5Ԁ{6f[͚Z����W��*}1aͻ�)�!U/�\�]}��%�]�:6�ȕ�9�����Q�� �gl���6����c=�<�Y��._F��fxF��=ҴT�f�۫�ur��U�f���X��T=��V�W#�*U�ˆ��H�FA�g܆׭���������s���s#�^��7{u�r [������d�,�-�����=�y�a�7E�,���l���$γ��!zF�:o[Q��&��b'za����+�eb�'6*1�.�BO�eNM�*��lq��̐��I�	�Jq�1�rN���`�0� ��W�4=�	$?��J�ܡ�9�%� .?eJ�+F�çC���}Ŷao�D��6e���ē�Yc{R���P��j�N�YfT�.����� ����pF\���weX��u_��+�O��yR�_P����rꋓ���K�L�ܬ��ߜ<Bw]a�O��vj0Q%J��}��+�xH�Ⱦ�Q��؊�\����a���r B{��m�����4�h�t)��1~0��z�#�vqت��w'�yUE��S�*p��8^V	$�:������md��
y�j&�����H����fo��HC��2����nv�A=����|�2���?G�gL?_�t�ho���s�H���	8�XV��R��)ڍՀ���P�"(僀����)a��'+�ʿ��K�m2�j���?�� ���XM������{�%�.��*�/�I[b��9� D����2���ܠ��hUs`��6i��Rn3�f[Joh�0(O�����۽�F�Ks/0��-ӑ?�U�-ZLn7��Tw�X韮��|5��-(A��s��cu���[�\T����J��mп~#Q<�e�NP�=��܉���R̜	�%'{���
�i�U@r���6�$��,��[�ο��YJ��[�}gE�~���Z�(�}�ڤ��(-�b�ǲ2�݊�s���d�V��?(��a������M�n�t�2c{�����-O��e�{�^K��{+���P7J����R�H�ժ�޷�eѸ�5eb�d>�����N�2\�t_��,WY�H|r���n�j	�������}��g�n��fsJE<EԷ<�7Ə�Ʉg�����Y,ED����Vxޚ7�	�ti^B�CS�2g�<��T�1C⃭33D����L���P���3�ᥴ$��y��N�=���St�ݠ�q"� ��W��G@]��3��=,�c.�c� ��=g�}ѣ�v4�g�-h�ឆ����m7j�Z��;rT�A�p��C�5 [F�KGk3/I>Y�(uDAS[�a�D���ygac��Fz��H�:�j�|�����%?	�~���3^���ʨ��w�8�><a�S�f�SՕ��C�8��8��-��=��N�;d?,�������]��ƽ=�LMB��;��a���^�����p��Y��r߂~�胾/��t�)���7KxZX��v��FD�(!D���ý��;>W���/�6 q%�N���Y��f����T�j�Ht�D�� �f4`��UE/.6V�әq/�z�	�Iۍl)j	�=��ϊ���*�㽃
o���F�2�����e�A��v7d��_���7,�q0�nI�pe�����è#Q��)"�4U�5�ȬP
-W�i�]/s�:�R�Yv؎!}x6��G�/�V����!h�iJpԊ�P�{�]9�5��"�B���Ռ����T"sEtnm�Fi�+�g��F�]�~�^�E7Oܧ9��>l��!G��HO�~$M��E���F�g����^hD�������:5@<�p�K�)����m�~���D�Q��W�z OCU�:0S�+�*�P��B�!���M`�8��\��x�樉��p��ʨ�e�C7	���F)$�->�g�M�I�Z��Rq�]�����FD^�GD�nP��o髶lp��H�^V9��*\����Oc4���'����ս �u��`�w�K�u~XC�1\�:�ȑ�3���{�""�Tjk�\zg����/$QÈ	��Y�ޚ@��Tq���%}���ys
LM� 'k��xF�-����۩J�!���
^
��U����l8�L��u3.����;��jYiS
S����g�����ބ�<U�'~͸&j���q�/��3e��7ci�[�7Xt7���Y����`��z��i�>}�4��чf�`��Q���z X��ZÉ�o�zJS�F��|*����Uk���Ʀk{kAf�_囧�	:��
g�F��1�,Xkcd]�]�]�L�`��h�[x�~ �F���ݏ�!��^������F��v!?�r�UJ���;O&I2}��:Q��h�q|��$�Ixr�a*-�x$��4��N��ς�sd��rėߕ��U�K��͙���������M@�"o�&�f�`>4j�N_T?F��#������,�э�m)W���4��0TW�Z��C��(yK�Ԥ���|
hV�Kt�f@Y��s�w�l%�D�0��n�<Z�{ha��0�!;��S����n�j7�6D�j��3��������x�r�.�0j?6��IC�_�����U�Wn�ᖱft�|Z/���>2մG�t|�}3	��h*NR���Q9j�������4})Ґ�baL�B�P�b��h�Tۚ�nFNVKVq	+5�+��=?�7��	�͏��7YBo�{�Nw������aזu��3��b�^�K^����w9��>s����x�#	�>��h<d���j�9bP�g�A'��T1^,�8-H�zVHΏuE0ЧJ�>��7���4?%��E�{�uk��+͗���2�W{�/k��Z���H�L�����o֏����w�_���:����}iԆځ�]�O�r��81��M��:�JCn��(�Zs�h%|*:�>�%����,��i�~/��.}q�(�X�YQ������B��Q�!4��^8��Ē7��m������+��j��*�\�#U�)m��,CM"��  }��l!`ɱ��4�2�~9�Sd���\#Pc�J�.O���u��S�37��6���:H~���/>�\9B�V!Sm���^���y;9-}˺� ��I�J�I�J�+�V�v(S�t�İ��y�;�рl�J�D��F�F;�o�p�-B~�����eDѰ[\]>{�#�**j���b�� F�
��V���N�$wԅ\�|�@��[�o�&lU��K��X���8���ޱ�(O����u��fqEf�"8A�KyZ�'�4�T�ȼԚ�Q�b{����0��-q�w� �,}v�/��3��t}�t)Z��ov!W[���>��m=� [�!2?Y(�nDS�N)��1�e�-�ngL<WQY��\
Fj)/�޹���b\+���ž<5�}�o){��Q�0u/����,�ˑ�¢Jf��'j4�d��]cA�.�	��H�ߖQF��~�5�3����O7o�*G�P���z��@oQ���Q\��ak�}�� �P4�1�������/��ac=Nv�X�o,��� �����ct����q]ű:����*�|m�۩�TJ��7"SD҄�*7rڸ�w]�^�p�w��ϞU�鯯V�� k` ��O��
ef�Čҹ�5��<�=�s�`�:얂���i.B�1yA'�Y����9Q��bW�v�iYV<x�°9�W��9�I5YS]�ru93���̵��=ӿ��[bB����>����5NO�,��PE^��M�+m�B���c�ˌz�do3!6&��� ]Ȁ���k�����G	=ϔ/��+�wV
#�Gҳ�X��m��bp(%�1Xw`���zU����b�I��.�*w��A� ���xW�����J��_,�H��8@K��-����^�6��L�VH���Y a�ΌE<�f��4� \[�w��}�'��X��#s
�8��HZ�C�tz�d�����7�H��㟼�Yޭ�1��q2�n�g^k'�S��tG�59�����_aT@5��՗���������r�:<]ʋ͞���p|;�L����,����~�}!/���7�sFɁ
�}�s��i�3�+I���e�X��9��2��ߠf(��n��:#��� Ѻ@Pc|�(t���Q����h��
�U���D�k����Y�siX�m.;�W���Ӡ��T��]�(H��h Z��E��Ѐr�����l0�<�ie�a�����|n��		�*�%�yՍC��
F�mώ׷"�F��f�	���\9�X���s�@Dw��Cyλ�$��$b�F	��Ks')��j�(��\7�ěX��+L�������1�O_����'���(F�\�l�I=�"z��ߕ�|��M@K����,t��R1�ȴ�����G}�5��S3�z�sq0R	��VѾ�-"�VK����6�EWg>�������\��K�(Dƶ�^�C�ڇv������@��(�}!�6� �H�AA�;��� ��f��եGG�!iԮ�m)r;�PB�n#�������g�J� )-
@H��������N4O_��m�K)�^�W��8V�c��R��,�C'O�1�ć+��ŗ���9�W��b�g����!h����nX�;Tm�sx���r�q�go��rJt\��ub��Y�!&����g =�� N�n���ՇQ�*��v��!Qb��)q��d���3ֽyn���ݑ#0���Y����\�}�Д�H`�#)�V��m�X&���	��p�r�1�e�_ߜд����D!.y�9n�oF�t�"󂼽DȢԂh�� Y�4�B�z�Ġ�x�5��8�\�^=RZ�݁�|�6�lEQ�q�a�F��R�M��j"D8����Tչ��ڇA�"`��Y��S҇3v�eǚ�!j��2>r<� �?%/B�e�g���<�4s�]{x)U��͠�Fd~OiW�'����n#O8��9סU!S�.�8�h��@/Bv.ӌ-xK����N��0�ܕ҄��@i
���#����jRؠ��>�l�F��SEę-k�в��>����:��A���;�/�d{��a�哄��X��� eͬ�O��c�!��:(�	|�h��Lm��:�f�#�ꬲ��z~ ��)�ɧw���_&y�%Y~��ѮHD��4k�\�`_XW���h������ڐć�� d�x�	I�~�k�&_���Y��7��@z���L��i��o0I�i���Tr�32̿$2쬵M�ڞ>����l/*RU�51�~YE1,Imf֍!�#�9U�}n~��f	�`�]D��&���~��hCkʂ���gDG}H	B#M^��|��KP�;��7z~�t��n�&D�X��VL��w���G/��Uw�=0�����]���_k��Rv�E&#�5&�� pg��*G�gGucr2D-�� $��U9�C���MZ��3T��6��%���G���I�C۱E\�~G\�1S3�Ko��G��U�P�na$���E3�a0S6�﯈�E瀙��:�{�x����]1�0
��|�cB���0��udZ%�2<�e3��U �bv��� xSќb�\Vd�����(��3�^��4���h�,E�]_<�����QcHge��zwVv�]��{��{��ƾC���Z�3Q��P��ѹ����sË@/`��"���
��S<X�E��UHz�����j��������!綋э��|�2{l�d�}�F9�W#���|��l
��w�������7���a��a�f!���+$v��6�E3�O�V�-�
�͖ͼ$�_#��SKw�S?���a�$V�D���YT�e�44O��*�Lt�<��!_�Yy��F�-KB��]҃��=������`�mq�t��<ri3Y�1����t�q�76ȃ?>CB�'�)k��`�B�`���L�p'�1g�3�R�2a�ށT�~�۝<�I��a͸B��MAo��W��	�8�[q(�*�=�M��@3f�8����e�[�>}��X��b�⠄*��U����E�Glo���B[SjȞ<ddLά� Q
�=�8�y\"� �S���jh>mw�+!��o.��E�S��,M�,�Ax��˔����~"q@_ .m;e4	�Ml����Dh���%�&�)��ׅ1i��K���;"��uذClyx����N~c�1�O�e�ɠ~��i�)u `%������@c��i�uZ`�Q��R����$Ħl�)tr]�1�7�^ �.�B��w�x���:/�lIO�� �=�ch<��/�`sy��Sl��؁�����%��>�-R�U&�l��~-"���<܀3Al��8a�xr,P�>�P����cL`� J��.F�P3�Pk�����v(���h'��yۇYE���C�n�"�JD-	��P��P����T�8`�X�*N���ǎ��"�L���(w��E�8���a�+�n����-�򫟖��[w)䨎
7§����2�C�"�w@�B�u�BT0;�q�f�@J=�5�S�|hW[#��Bn=O����I�ݯ�S@zn��~����f����f�f-ꌶ�*���#Hx���YsQL3�^�1%�v1!Z�$t�`�4��RG[�P�eeO�i?�~�.�YD�`�j���u閆��sx�:e1�Q�����F�����@.�.k�����3��V��m�d��\��3]���w錀з�����ũO��|���3�-ڃ�t%�gUؙ�z�8BM.�iI���ey�o6ɖ��=��0�,ԅn�����y�<B_��l\_�fM�#��w e�ۙ/M�0�t��������o�fn��w2���h��&�0;0Ő�epv O���	�����Ֆ�D��,��ta�9Ê!����k��J֎���z�ŝZy:~} �(��W�Z���}x&�ѓ����w�+|阐|ܐ�-�M����Ё=�G�P?�~>����M&^(6���GVW@�8�bA����<-�6fuKb�X�!�@k��	2A�"�	ց�$��_aGJ=��+pVl\2:2��E����a�.�Je�%�&҅���В;1y��k��.����{�I��%���.οB,�V��F�~+ƃ�o����K3�)��y���J"#�/k3��ҥ��v�G�ƽ�d��/�qX�5���(� �]h�xvA��z�~|Rp�]�X�. gi���TF��9�~�ʥ��hk��:ɽ��r�C؇p,j�	fXh�UH$��*��A��+h{�7Fs���{кZA|�;������h�|����b<��p�����W,�?Nh�7����8�r��{o�`���s. Uo�?h��"5������@�B\�j�`:��wt�կ�9�F.�.�
�9�<]<G��a���g�M==E/^��ۥ�iD���0�C�������Ilx�����Vm�����c#a`��}J@cb.B,o55��ɦN.pe��5��O�oBь����wj<�)N����yIO
q�j���	��n�;4��-@�)_@�o���\���&&aD��Ru��)��m����?M�‎*h��G��	7�W^t ����r�l��r�ܙ���%(\���	�fo�FE&�Sǋ��؂�i���k�{ڵC
-�n���7(�h>�!�'/�	Cģ�p ���4�����`:#5�z���k���i����Ӂ��И�,_o��4��| ���g��
��aA13�#á(���k/U���a5s���$o��>-��NL�L�T�����G�;=vm����k�rr\t�@�V V�^.�teW���V���U(�{�}�?�5
`�ܫ��|!��S�EF
�d��+�r���HG�v�&��C� 5M��X�j2���4R>S$�E~z8��>3+��눁�Ī��p?�u�#�X{��lKXio�B�7C���羭 ȃ:0������̿`S���2J7�$"��jH+�[wDش]}V"d��2�R�zvBu��峋`}�+e�[��ᙊq�?�=dV�$�^�j�Eh�P���ч-��j�AN��+p�K��R�����DuH�A�:���*�b5����U����z����e��?����BRU�>!�(�T�=V:Rɂ`�aXn�i�V\�$#�M`��˟�͗���O��8R���*)�PjJlj@O
����m��!W�A�w��A��ks�K�b�p�QҴ��������8�C�S��S��~�wj	����,���S��LJz�UZ�YBu
�D��4#hd�5
a�ˆ'�:v�/+n�����2�w��%��O�<���R�����W�*JtOp|�!�J�l��y�>��x�a�>�����n� V�.q�D>����*�FP��a����s�:	�J�}���j���IQY!ŕMU ώ���F�:鳷>��7��Q�O�E�[����\����D:�g���A�v`�=���64�Nlx��
�ZO-��9�MP�9��U���w��EM���3�S{��/���@��Ξ���!O�,D���)lk�	E�����B�U���K �ΡJ`J��;_GM���Z���L?mu�+��&^��i��i�?"��U��8z��?�6�ˁj����x�zF��LN��M���8��M��rI�i\9N����d�W�\�^ /:N>.9}��$L~-��8�ah�ձ0�F�m�'��ӛ5�8���P�6L�nNJȅK���ώ��]�:|xpO�����[2�T�S��2�����K�Qk�o�� ����@ľ�A8�>��iG�5�#C�6)��_���y���=ie��JŎ��X��^�"���◌]u��^,(����]��� ,'Ʉv NIe�����#��-��6����.���Svk3dCXF6XD��eN}�8DZ:��S
������#3cdQ�2��~=ne2�sWY��%xC(`L�֧��0�	�&��%�8Nt75R���g�e__h(��
��ۃڷ�?&P3�	[�TbH-Ϋ�aC%'�:W������'8.��Hz$}�Q�U�C��#R͉J�ȭ(�F�l�?Lk��+=	�w�����S�R��!�M�lDl$x��\�U�� (V�-�!�.mL���8�1��Xޤ�P ��	U.�<�z��Q�̻��
q��{���##C\u��3�P��ZZ����X'{+ .�Xk,�ŗk���7��n�I)�E�G����BT�b�څ��Y^V������X��*���hl^�/�	���?�EЧ���i��� g�T��هFK��B���0.D]��-��C�s����"8F7�֌�G` I�2F
Gm��V����)���^'�-�O�W��m{���8H�"�rT�.QYOT;j���nIp^[��}P ��D̪FDX;Z�ZpW��;V$_T\���~�Qe��S�'L:>�rG����{A��g��IG����}�U��!�C�J���M��G���u/����qA������������oe�	K 0�1�*�̲֗YҹR"|}BB M�t>�Cr7�t��lAqvړ�!Lm�p�W�ٲ�"V�8<��GH���>������K�{sݬZ�	]�(�T�����N��4�^VUo�)_U^}s6�ڛ/E��)��j�w����,ٝ�����ͧ`g�_�̢ez���B�� $:�v]S�M,��+��a��'�1:������}VY-*TS�Q��G�b�L9��� Q*7}�n/ImH�� ��lR�i"+�412�!�	�Â< �h�$�ɘ5�q l9�D�ր��i8cZ�ɚ��) �s%��	�R����|�A��㝳��lc&Zb�@1`�V���k!S�?�)r�I�:W�K���T�iN�j�fS����ŭ�A�7�Y,I�����.l���	?���j�Ģ��D�c�� V~pd�y�����_�d���9]�"����*e����\Z��G��w���/��V�%IK6v�MI�]�wp��=��Lpю8���>M,��;[�J�Pgb%v;U�x��(2����-'����WmF���K<[j�Wp��I�t��aP .�Di�Q=i������d%�N|�.S&�U� �s��>����)�C�޻�&Tfz¸��p˧v��¦kG?E�c(�:۽��5}�dr�U��)2j�_V���:�o��䜺>��5Ce��=�Cf��i�w-'���-/�-����Y��<mFp�d�j�݌�� �V�hIO�1d(Ʉ�����$�:�Nq�즄��'eE+���>r��jO)��k���sY!gqo�6@�'����ek�$�6�:�G��`�ϥ�����d5O�A髥K]�9N�pt�,Ҽ����b
�G 5�
'��V�
{�Kƚ���͐(9�b� 	����0�-��0���L����陃�ы�x���$��v��Ѻ<L:�I巟�H�m�`[�[{CF~���؏ǫ�d�2���Juf�)v]\C��p~���mi��0A����0�F�;�Z� �N#Χf�Mk��T�5�S��f8�j�#�2O���h�Pw4ӂ�Iv��i�rG��q�7*�8 �m��5&�s	������뀽��lZ뵴��ʆLܰB�-��>��s(��^pDv�OH �nV���C4_���%N��g�����Y��H�edlh%�N�L���'�=�U�f���e?�h��4�k  2ʑ��XF��Q�u�:@����c��i����܀I
g�K�������t ��"�q校l�1\��7Zdl�gk����E����U]��^H����f�\�{'�R�LOw3D"�������� �@�``�9���O��ҹ��mT`w��a�=�67������z(=���d'?�[و��A�����M�y#hMH�MWbb�doz�ۘ��5������*C�Mw~�}��1+��?��)ۀ=^b�jO�5�����YH�������G�����wG���\҅uyPeg7=��r�Vu}F'�4D\B�i�)AWP0����Jw�h�>���%��o>�/�eH>��}�׼�d�\=�[�d��jw}D�#^pi�hy62N���7����{�{H�
��@ɊчI��h	��
5�u�!*8o&������h��' ��M�L��-�J�0v�,Q�^�O�p���X�3��k	��"q�VO�mue8�A�`2��Mq�-�g&�ӫ���*:ढQ�.?b�)��{�In�2�">���W��$����dӿƠm�확|�]���E�m�`Z���K���GL'-2�&��:~�x&���e��(�Z���|��ŋ�J�K�\��B��|�^�l��IÈ������]5i7hk]& ��Ii�:d�i�oT[�VW��9�XT��;y�ϻVj��=9*��G�!�ވ0���F��F䷊��3~�6�����_41b]#�{�����⠩� �C�9T,�,�܋�h�(u���3Ì1��K*�I4��pb�I�Җ�$��r�z��|�C��4�%�vG�}��Պ�'
�O3|���r!����B�D�t��֚�D�PsiЊ�ߤN��SP �#���z���ߜ�)f3_ȯ�T�IaB;��;��lD���4���~� ����/��M�xL\L�z	��F� ����S�"PeH�^�m�Zm�a����8�	Kp4�����dM��S���d	�9���b��	�^����B��:[���^9é	Q��j��̛:a�	�ؽ�U��7�����h�J9�u�f��6�&%�_���h��P&ұ�fH��q�Z*d�)J�A���,�6���h�q�k��6b$�o�:%Zĥ��Ö��hZޝW2����Ϻf��A�E!��r֐
1�)�y��x�tKt9�42k���?�?����M���f"y��/�@&�}��̞&�=0����v�]mA^��.Yl��QFo�O��[�N�1�e��ڹ�D����,��({I��eZz6�J���J��è�bh��'���:0giV+� cj:Zf��� �A'�,�ֈS�ͨ��ŴA)�+���|�h�Ҍ�N�����k�w�[�#�X�M�N���k QiS�&���*��� [�e�-M�w�5���2���J����b�}*�i꾿�D��|���V���؎����㒢��
��]��A��;`[�/��<�]��x�(� Y�)����?w�`�b�(!���z�GJ��\��Ϭ�r=x:��XD7f(�����`��	r�O����J�se�݌o�䊣��:�u����wVN��E�q��G<�Ո'�}4�1e�y,��Ư�d�+Вĺ���E"{I�$����S㥈B_�*���[&�%�"�0���,��~Dq����=�ib��1Z�^���ݒ���V�7�+Op�PH�k�l����⛍lh/��l�t�SdG���yυrMa>�F��a�cZ���)2nw��=�Xw#�#�	�T_w��v���O|�$��Ϥ���,.���]����}�1���Bj��������R�t۞�Wu22�wE3�f�.f*��Z�[? �����;h�;�e�8����$I�`�%�t$u��݂�aԡo�A%;i�¸2�W���-pB��G��XFG-?��!/N��oZUV��*!{4)H���S�\�?,�,�����7p�j��R�kB%F(O�I���Z�ҤD��ؓ�g���f%���4ɥ���(=l>�k�Y�^���r�T*Ej�@H���`\$��pA��U�MݡQ�Q�G��}��,���,5)��ܹi���[y1Ӌ��-���D��|�ʤ�a[�^vH���^z�C��������IO�ZPc��#H��sU����PZ1H�+�|[�1�\!���M�۽��`u�8 ���B��#j΀��?ҥ{�vm�xe�C��$����J{85oF�Ƶ_�:��O�,C��c���/�5���Xދ����f��k*�|�2��ϖ��1A��wka�k�F�@N��D�%Sv�w=Q��iM�/~]�����u!�.ȝ ߓG;+��o["O�6��Їn���,E�B�L3ST����ܑ�kΕ>j`�>6R�hKVyx}�4)��k�
1U<�Z"��Y�hGP��,�ۿF��,J$eϹn&��h>͉�?��nښ�ff���@�9&�Փ���:��D�_��̏k�[�?�}	���2�cK0�ϔ���`�h�f�Ϡ�̑� <e��d�t�k)��QUb�x�����|L߽1�9(�}�JcT� ���w��i����[8X���E�N�Aw�ʷ��Z��Η�~J�$�G�J��'�hG���ϖ[.�7L����Q�N��P����i������
n�tYG�$�*˵���wC�T��Vo��E}V�BG=��v�}�
�@v�/ M��?�$�jw�������Q���t��sm�D�]�@�T]�m)�(�i�92�� ��Fe_|0!�5K��v��7�7�չ��5{�Me$�_�6 ���?xd4�7c�ʶ�1���C-X���VI�׊7aE�����W���X��P=6��QE�^,_�@�.�Wb���
�3�i�u�_�R�/k*�o��!�i���/�궉C��G5`�3&�d������~�|��F]N5�J?�E������q��s+'������ $
)Pf<��nw�.� P�Cη����>�/.Ijc����%)��?�����Y��xr49lo٣Eb�O�R�K[�+ ��?\J��H\��/�႙�ɨ7��U��	�V2P���_�����$y�3���1U%���l�a�'t(mz���N}$Q�8���cj���>`,�o:O$�C|�3*{jV^;v�A|A�%�� A9��t��,�5j��,v~`�sM����:]*�'�:H1 ���
x�Et��q򂞏�tc|�e:�\ �T����kK�й����D
���P���-L���,�+��_����rGWgiZ0Y=qya�/祊�ԕ�
��޴��UB/���uX]f^�-l��K3 Dg �S�r��A��g�n踴e��o��F�5=���������jY�p+E�s��ҫ��駖�~E+w�V�Д���T4^S)��e72 ���ZB�b�x,)ҁ{�:2~&έof�F�����fxkv�q{�.�A9=z��v�yvS>$L�*��A�.���I�BS���4�j��K����C�Ͳw+~g%��\a9osAb��-��I�[��QJ��|�&g)!+)�Ao�g�|���>r��ꅭ�2L.q�:��#S��q�A�gǀ�s{�Y*�Cgt����MX����#«`���CQU���*si�G[;�q\�^Lp�}�/3��U8��J����!�3x�Xt�&��b����N��������;���N������R&%�Mp���UZJ=�T46qR��� ��K�5=�$�:UN�L�Q���g1��֣S|��4���ޔ��m��S4#z2���K��3|�z���+�W<{���N�?)GS��B#&&���Ef�;�.'5�R6���+ae�ZP����K��L)�Ը/����x�a/|bp����Dڼ��/������n������ �_���;�8.�q+>r�_�=1�H�`-���{�ή 6-Ǜv�K��2�|�?����谖+Z�18�p���P������h�eN$:�*eKΤ_8��W���J;�EUS�����Y�1��u��S���/����F�c�ǾF��`�)�̒aZ z����m}A�!�FW���1x���U��0�6+���I�n���	��K�Dov�.�j���]'55�z�e;���zs�u�3`_���WQ=&���)�����S�2�'H��W���!��R��x�Iŵb��A�������R�eL�O���j���-�u�
̄����d	/�s�Z� ��.!7iư�!'�ZѪ(�����`󑬿(XH^���L"Ҙ4�w-Er ��nd��Pm��5�?�`�S����]&,1��=��'�)����1����.aђ���Q�>S����~+T�>�Â?SMڸ!�hՆQ�l���z6li��&?'֕P��e���e�Q�ۊ;� ���d��� �u�}_��t��Ӹ�v�Ȏ<��%e����d���S;�A^���PA3��5%��N�]V�+�zc��?3P�!C�u3._Q׻G�9����͹�[+�k���X� �'J��+ዖ!8nT2�w<^7ۃ�x	��D��>��_O��$q���>.p u#;̓��x"_��A���,��
�erK�>������;&gZ�j��I�Ll�q;�K���з��+�ߺ��9[ϩAp��E�ҵ:�}Zy��E?r�Pm?������Ѐc��l`w$ � TMܮ��"��a����!=��+c�����/�жg@D�(�B�P,^(.�v�g���L��� ���z�h{�I-�6�П�Xa�`�oG�h=�"=�N���5T�#Bs��7�ӕ�R��})�׽�ZwO��KS�s2y9��1������Z{�^V,MQ"."�]�{ʑŪ�S�7�������F0z�{ݯs���+�������F*�k=n-��CZ
2rQ	�V�▫}�g����ݹXY���y_�p�g ��M:o������gs����ʽX?���23�Y�Q���4������0*;e�'?���H� !������.����XyzyT��c��J�R�<�PS�'V��9�;B���ϜW�F_���.�$de@�B\�R�po�s�ڶ9M8c����Jϳ< �b:�Q�_�Y�au�Ն�|SG���YD���|��͏�'�E�͐�F��d��1�/��#�&6mHi!N�2�_�+*�tB�Wmkviq�]9�o�$��s�9:��#�Z�XP�T�%
X&���ZW���{b{�a?��z����{3fw��o|x��t�C�w8\_�<J�1t�N4���	�����Kbm�%�f3}/0O�Q��.�rS?�}��K�_z������G��_X�+<�<H+�Gq���yLp�z=�'Du�!� (z�IM��x���5B�!�E ?(�0I�"I,[6��2��~�4� Ə����������t9"�$��c���:�E�wb[�0�"~Y�+����1�^9�r7�q���U�xu��>�҄����\ɦ	3��,�l���zl���4 Z*�D%�A�J�Dkr����9��ʏ{������r؈!V��_q��<�1��BS�؄)|�#^����6rO̢�ay.Tl�)�?��큙ء���U��-y9�`V��X�KE��I�K�v��5Π�g���E���Ů�璬�O꼄u����.zD΁0���t�%!%���Z2B��2�HQ>>n��@u�]�K���܅�(���՛���pi���jLn��PZ;,̛aX�U/5�1�|%��m�������>���!{@���̈�@BԿQ���S8�lQ��$��*Ha��mI���y��V���v��j�i�S?i?1W�j�@���	��T���7c��M����l��<����$���x������3${'�ZL�щ�B*���r������&d��q��<��R-��r<��g��/9B.���6${����/���|�H\d����EU���xȽmu�����O�r;�cx�6F̍K�b�1
K�����2�h�*�;��ld/r��W-N �C��*���@b�	U�j��t.߶+�},3)s���<��x�C�q�0��l�sy��+���r+�O�*E�(�u��~�oK�Z�-P��dE�Ғ�l:ݽS���4��Y"#Uj�p</��d�Ec�#S��>B�����v5M;o�p����[��)����dY���V�����ծ����\܈��hBh�G/�?�A��72�{�{����6��kz>���/<����P0͔, �d�ـ�	��'1����$P���^�7}p6�X�`��m�t!x�o���|�H�=��*��_��}��qig��Ch�Y��%a+��w�H;ݮ8Rf����i.Siߨq���aT�M�f��kU�9�z4��j�<��gg1	�����6(
��똄���;N��/G��x)M�08,���i&O4��;��$��f)Z�guj{Io?w��=|�����]����8�?�	�L}�;���p�5��R�5S3���M[Q���^D3���NѴ��0���k�#�!�e��;F�S���C^�q�E)J�>}�{��hc��I��4�U�Ь-N\I�������?%d�e��wg�U}3E��3@���a��Mq��� ��㟊L,1��~Y� ��ܤT�R��EQ��v�ؽ]w*�����A""�V݊��ߛ����oa��0�	�w�
��-%�!>�r�/��Ѳ2�KMˡA����4Q8�ʡ]m�STw<N�:j� ����zb������
�<����P�ݵ �	�ײC�ܫ�����g�\ͤ|���J��T2��Q���g��7n�����Ai!e=9�\�$�;D\��T�K���1�գ*[�
���?��K�|����1()�3?�����m�MXڔ�8�C/h{-�c�"=�܂ٌ��L/�7U���`��\�^_g���
zYI�_�sL��P��l@�&�E
4�'�����n���G=tH6�o<i���u��]�W��k��OO��* �yJ(�P{���G�4�FL�O5�M�G#MJAqZ�j��0�⻣9��!�*�}\7QX��ws� j2:�+ᩬ{0|���%�e����ȃ�O$s�f�,h><Q���vC;���<JвBW[�t�"�W����m��ey�; $ҳ!{��I����-V}*�_�O���j-�q�L�V�J]T�B�����eOz��_N���#��D�K�8��pP!�)c�<��^['�I�d��=�H_}���^�QF�f�?�v��q� �Ѭ���|6f��D��:N�y��������E�Ձ��[�y�Lm|���9�Y��)����FS����N�H��б�举��FŲ�l�:�R��vO�A*CD���S��&�cXL�E
Q�vq@fI1� ��r�f�G�zÿ)��=�*r��u��@I��&ޠw�җ��1�[��k����dW���qg;{d�g�L��]`���a����K�����t�%�gE%�蕞A[��T�>ڡ�b���@˜�QM�Y�P �`�F*$���^��e-��r�q���aҮ�a	����n?B�d�]Uo���ViGr�#w����$2$�X*B;2�!~2�6��lҬ�K����[�ިKQ����B�Ay3���ٶ���o�R9��ȝ4�˄�B��3>-�5��BN~|�7�1'�6IC4�f�'7����xU�Š�#�8�:�ҕ��v�_W������<�pX&C�����W�ׅ��:�����Y�߲�K�Q.���C�g�Dܪ�51�^h���X1n��UHX���- ���b�4e�� A��(b���w�Đ&�8V��z�h�I���\��g��U�@k�����.\ĢL�w�f2�ĸ-i�����3h?���#-lՖE�̫�[(��λ�Ȫ�*M9���0���}����i׍͞ou�3Xx(���G�}|�Ë*QE��O�����^��i3�7���w��W+����%���� -O�\x7:���o�An=���jaɿ���rs�j�O#�|�bo�������5�Hk*�YGsK��Xq��<��3��3�٬R�L
y5�Ps
���b�3�&4���T�.nI~�io�D=�s�K�̡;�B�v�p(z�丟����;@W�eF���b�I�d�K�Bǉ�(^�4W��ӊ�����F�c��_J���@�+��\��t��'�e�p}���~m`N���TkNV�\}Զ|d��7��w+��oG��=�� �;��Dr�*�`{���y;���]y�!��ɟ)/�m�6��X4ɽ����}���}���5>J[L�)Eɢ�1gN�Є���=�q��")���+!Bp`U�]�U^�t��\�E��~W<Q�e�"7�Ou���Cc`&��}�˾7�O�"q��w������j%Z�K#̈`a�ۯ��,m����yvn�Ak�j�K�.C�^�ȸ���a���~��$3P�MB�(��-����Ί]9�JkvkR�[CM����S�6O�b�Ǵ�gw�m���C���!\�S՘�7��Yi��l��UW�������Q�'�����h����CS���'�r���J��c�U��&o�3�T�֪��;�5Jr�-jf']sΙ~�^x���Xlh��j���X3II�.&fk���j͈U2si{�-f��К%ԮJj4�m�pD��FF�+�M�G���8��'d>fz6߻������t·%��'>Odc$8�Q^A�Қ��l��D6j���O�a�ڂ������$R��$�nU��5S���.�Fو1c�2�9�j>�ȵ�hЭ��yq�\���!�ҷ�j���y$��.ȸ��h��sD-�m�*NbAx��=���B�	��C�M��.��E�$sN��%����0��w;3��d�u��F�Qng%���y}(��Bm"ci)Gĉ�w.�,t%t�& �s��P�H^�B���4��f��<�#���S��������6/�M�xL�ƿ��_$������$�(��aو�������H:�>��#�R�th�XS؂Z�zJ)6��6�2�*��s7�\�.ڍ�Z.���^�:!�>��8u*}}��Aũ ��q~��=���yVCM�Ƌ�N�4l�{a푨@�?ZkZ��>r��_U��a���7���IL�����Y����L�x��Hǖ����\�0 ��o�y�"�ZohW�c����b!Y��$a�����,H��m��Q�a31C�'y ��B�^�*�����[}ť�r�,�򗸆���=UVVq^���FB?э�V�S1tlÆl��N$����n-��a�wU/�1֡H�*U�{//D�#�WF�?Y�x��B��63�W��_Y�= ��@�!���Y.y��#�k.��(N��C3������`�n����X���,�\Z�s���a�s;��f�4�pu�� ���EC�Y�� �f*�W-���>_F �����z$�yAw����c�-X����Ѡ�Q��J��Jm�搝�����䩟K]�Eo�
5{�Jz��N���8�O6��7<�Zc���!]r�>��Awx��Z���4B=����i>��ze��;;p�s�t���IwLx�����5ߤ���bѼ?3�ι��ELүV{E��S�޷Ѕ�?�3�	�C��Ɛo�`�z�n,�/�qU�g8�n��qc����� ڠ�� �xǠrFD���V���st����5��4����oɪ����<�uX��~�on�@�џom�*���5�.�Aok�]�Gj0%��k�Ep%CJ7���,���*�������ZZ4��0�Qh�I��Lu���� �=�(�
����j]�CE�t���������fk�u���tjaV�|�e���ӝ��L�o�)%Ľ)�	Y6�(���ȵ0�Mt�v�2̅����r?���qW�=��7p�1�LtT��g/�����.�&^T�"D�bM�����ўw������{��:�>·0��EVM��ť�r��
G`�����8��Z������E��n{%eKNXZm.N�-R܎J�OD{j֦j��B��2��즼%���c��T(�����f؅�1��6��!֗TB�h��~/z��p����>:�Y�:���-8�*S��ܫ*E�'N�Gr�x���;�ơ��bJO�Z^@L'�e��<����\O���ƚQ��n�d�?o��X 5���W�#u[gl�a��ݴ��d0����W�����jq�b^8��iC��d�$	j�HU�.����+����j!��]�Z$e��˘n�;?`�S$6�UGYz�a�3$�DhUL~t	iE��Ԕco�.���W�*��n��8�d4e������KbfC��r}�WD<�������8ֹ��nRB��W�~	��¥���V��$�Y�����NX�NR�띋��p"�A�gt���̫�����#V��A!��z�o�BتYz(N�����S�\��Wn�_0)�Qx�l�c�:K�i������4V~*�idULnA6�+�	�Y�3T�6x���� A��ya�T&P��O}��f1�����w��7";��e����F�!J��T�l4�������>����lU�@��
��j�j	֜r�����{ې9�ƍ17��Ӱ�ĂB�l��c�;>K���!.Q���>*c�Z�YP��!��QJ�m�xEI���sU'�a���÷@��55I?���<�#ޖ�tXRU���YtD�J3��26�>���;<���,''�zq�� �~��'^F��g�ׄ���z�UVy^ô���7�)��2+`J6	M��'�����R3
B��nߵu�M��l̐����xN;ի�ġ�c�vp	�x�_���8�fme�k�`ʟ*�%4x�c�$���H*FǗ�Ù���6�smu�ƹ�H �l���|��]�����~맙��*(����~�c���(6a�����,7�,X
y��:�>[��ͽN�Z(�V�H&J�:�)_k:B#�Z6�t{����7���A�l�7�*ͣ�������k������~���-A
l�h�l�[�Y+Z9!ܴk��}��,)c;�t�`.V���S7~���Чp�R����J����!@��o�ɑ>Xr��b�/��=�D3l?���Ǘ�'r��h�� �(�t���z����T@�cj���l4�2�����K!�F���A�7	��ޝ���틘���6F�zH��A���"^�������FA��CO���Ц�'5���O�sqvV�M�O�v�����P&�Řጟ�vL�R,zrD5E�vy�S� ���,����؊�w���(� Ixr�;�]������;�@���do4���֪�I�똍&ڔ8\�.�CTR�����?ɔ/ױ�=5<r�v�:=*xE�?/���;f&/����]�"���짗��+%��د�7I���á�� K5ϟ`��/�]��F<�'mP�g�Be�2�\dU�Eˉg��0���� � B��5`��㿲�b� Y���ؒ^��}/�O�e���!H�U��ف&1���`�\��#_M���Ⱦ˦C?���^��Zs����#g�=��GIx�T_�0�O���ap�^���hmEy�&j�D�!\Ta��@^j�6<�`�HŶX^��}�SF0�:ˆ)ž{riH3 �G�N}��n�4)H^�Wq���Hy-��M|T�enғ�M�ټi:d� �ѝJ�#�0�~�B$b	��{��<�6��F �I���
�����Q~نp,�l����.h�#�" �����R�i����xya����8��OQ�_lW8�IP�П��As=�%��)���"�I�˕�JP�$���M�h�\s_\}|L������&�@�ny�j���GO:�E�_�Z��������%yi��?ү]?�m��ħ2���n�4A�w�Oxl���t�����[S��6I�M�!Q��go��Њbv�㘱��T��M�а�@p�!�	���ѝw��+��}<�eI@�W����<���]���T��m�Vɤ��֗�7�e�qW)�/�d?A�����	(��2%3������k��j<�a�wp�@��G�����v�%aT�5�����d�]2*a�B�W%ٴ3.��v|b&�(P��j� @bz�Ó�:��*�$h-����udB�<�����="�XDrc�\}�}@�3��uV�M���(�=�M��"���<B�0��,���"��� ��&^�,�,�jʂ�񤟅�E͠B�� Ť8�Xjn6���j��ɿ+�g�"��w8��Q��f���s�x�XiFO�٨���r�yDr#;Az���I��i?����{��t�H�h���� �����/�Si�m$��DwK�4KT�4\貸س��~q��X�\�0�̀�I�Hv���D������9�c�<�oO%`�6x�l���4��]�����"5�Ѷ-ĝ���*> B�{k��SS��B�V��ϡ�O���+d���-B�$?־��lS�O4��Fp�J7�o����GG.i�vr�xh�͒�A�a6�jg��&��z�O�|%�޾�T�X�#t�,]�#�
�@����q4���X�z��<6�����V�@ɲNK*��_��5��x�-���������L�T��y���C�͚���Z*a�U#��:�k�K�#U�u�;��L(�:�X���jG�`�;�
Z`��������b�n�\���*��p�Y *��B��>����vB,ψ.��Tkw�'n�#ܢB�١������j��c��8�� ��cT��J#��k�V:1S5G�x_�Y�%�ܝU�/�4�ٮ�nK�W�*k��>�cB[tX�,xu��v�%�i�4��yT��U�QZj��� �دh4,�M�˦�N�S
�$��v�;�a)g�c���-�
C�Q��Qu��'�������2ئ��-� �n]8�5���j������l�t\kI��zC�j����,��:G�aj�=��)���7��GV=��4Z�O9����}
���;f�!�מ³�zV�giܡ7s���5��j��5�\��P.��W))�i�ʘV"=���t�D�X����tf1��Yp={B?.�{5�t�2�8��l����>	t!�/���*���
\��/�ۺ����g�.T6\5Yu@��/�y�E�YG��:�.��
=gd�������i)ސt�	@�hO�{�<ͧQ�;�� h�z��Pp��K�(ֺ��J����/��d�!q)]5�����NKnT�Q�՛��8���&fvR�5�I�/!�([�@i�UZI�~�j�n!�%)*�G��@Oq�I��*�/ȓt�E���4��V��qԊY�ʐ��x>m�Wc:&gE�^)���]&�z��S���1��
�e�]�ch�n!�Id%1��-�J��&�`�D�#����:we��{@I)0�܁��'7��L�~��������Y�Tռ۰�T8&�UA1$�VfL�	!�u�<��ʔ�sܧ�I�Ե��6��X(t�Et(��<�""^Y���ea?�3��qCI������g�
�s���/d��࠵�°DW�!�M, ���DU��}{FJ��7\A)�`~��Or�6ʯo,iZ6�C!ˆJ�\y��?������A��8e�$���@״�?��1z�����#�T�p����Z��Y��
���5�I�)�=���Eta���naa�4����\��f�Q zc�R�fE�/K#+�ٿ5��,V>�Z�����2�v7�5�����γ�AwpT���.IR�8a���h��$��̇�����	E�ʬ�-�雲���'��}c��RV7���-�vV��x���K."���u���@���%c����p-��Uotg�,i��Yծd���-~m[Pa8�b�Ga����x&X"�b�X�Rc�p��ع�R��d�Ur���M&�<Y\,J�!�aw�Z�����:���r����_ �j�Ԕ	��'vF�%S8�h�������6SRj
�Dd�κ���[�����J�r��\Uѿ��Q,�Ō�~�;�������Ĩx�����Iv�0�����EiHhM��Ę�千�Z�ڸ�	4?Z�Q(&�%#��T6?U_~����	�$�v��tM�&~O����<�"Lv_���$	'�z���%��/ހ�MqWk�Ǖ0��$����E@��:;E����1A/����m3
ii~����35y���� ��Z
�獛֯���:D�Y��/�l�d�7MN��P[Ո6���L�J���l�Aj�CkOC�@ϝC�G�zKnc��)�֫#p='|H�����n%
T�~�Կ�Q��K�pͳ��=��`����I��9���RE���j�2�m<�e��?�AC��(�,�^:UkK�����D��>R)�g݀w�o�0u��O��o;����+&�].��HH���T��(�kTqp�ȬCPJ�)L��,�J!���	0m_�%�&!�C�J=&
�`1���F�O8�{�"�M}�����|:�aF9���	��U�>����>nܟ�5�_#ސ���@wRT/�[� $��đ�
i�9)��qbI&�F�TF�h0y8�U����b��i���l��ÕPe�O���dA����`9�q?]�S#Oԭ� �Pe`�H�~��c_#4RVkH��d�g7�4�|�v��PYs��+=�g�9���Ό��<
H���`Qm�܋�e~{[�
$�L�2��_�rgՔ������Mk���q��a$�Ik�2���V�~n �]�]]"���zC��%?� �9�i**�q/D�-W)��ʳ.��h�:S^�r\I�.!"A��{:��A'��\"��3��4M<Ȭ�l��s�Ą��<�ToԘʑ�\����/*8V� ֝�R�v��X����# ;����I����a4a�m3��ƾR�2L��7��)X���_"��6-h{�%��d8/�7
8S�yL��Xf�^�z�?�8�_���������^/��^�N		f�q��e���/�M�L��w���98b档1!=j�����������Ѱ�z��lŋ�ܾrנ�-��}�T+�2σ]��7:$��?��*��C36��<�x�������pD]��'�M� ,�%�SR�|��ʃ�>�Bf$yk�����$�d����Xw�<