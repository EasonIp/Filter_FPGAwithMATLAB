��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjfm~���*9&ʋ}�T������%[��Уt�'�}��������l�J:��	�gO�p�?�LkR{lmj$��H�����ey���t�@��cg�/�\�����>��`��0/ⱳ$���R�� �K�� *���g�Q�J2'�	�=d�E���ϠN)G99׷���(���Þ����n��8��Ÿ��� Hk��OU���v��'�� ��)��JINMg�<���8)	����j�.|�q�5A:�g0ƭ�7L8�
�hf�t�W���|��Ng�Fn�}G�_I�I��[�#`!ˌt��{1��/��'q@:O�qG�K2�a��,��S��ǆ.�&ٖq�X^�6#c�
��|/LY�/u~��]�6D7�ۥ�n����PN��7bQ"�g-����*��� l��x����H�Mj��n�L��|��J���9i�q	�l��m�O<��
���#���x�4m?�A��[&Aql��f�ܜ�y�h��X�[��[��BK�p�ۍ�O�W��zg	Y���a��<՛æQ<*�wvo�/X��*���5f�x��X��*"l��@*�*c��F�\cf3�t�p�Q�P/o�.���^էc|7�t"������}��mg�ࠡ���zy���������u�g�S��͘٠7���J7�ܪ���)7#G�/p������>Z%i��N���<�u�kE���T	�,�Q��+�b`�JH�`r�A�RM;@j����t>�[0��&����r��z���\F�w���H'Zĝ�|�8�7 +��ޫW[C9��=S�ρH	�� ^m��(�����(�(>��u�Q-���m��[�������!zh�`{τ�"Nݦ�)`�;��5?��e -x�x͜�V�H�l��H9]+*v(���p%͜�����Մe�N���Ѫmp�	�/��Ą���t�{��;c�����6��r���|-`�(�z���W?	#�tA�H����Q�
n��P�zϧ̦�Ȉ�9��]��7u/<ˤHSI���I#�BD�d�,�H2�Z��(�1_d9TY~�6��- �.�ЭYW�d��k�n���]hI)�9%��B�l�r�.$?I5�����v��A'X��>�t��[,��M ?��!�Yr?�
�r~&�,�*t��0L�k]�e���6���S��G�En��OT� ��B��yߒW�Y��N����X.�d�à�gB%z����ۦ��hNZ���Q�昊t^sa��ju���>3VN��;;��ˎh�]}�i<d��v���ƋA�S:K
B�����?,㽌����@��F̙7�v��?�F ����+`
t0M'��u�����[�B�o���7�.���,�	X��s�v��=�[9@�f��툡Wb���h�$u�A�"�qG�!��~ɳ��q����l�HN������w*5ܪT��'��A���%W�o�MK4��ORJ�#~D�A������PI�ٚ�n��M*;�x�Фn�Ax�L�B|��w0T�����?�?n��< �h� T��Wj�G�e8��c�#:�	u0�	�� �f��W�������J�W�om����(�|K�P4�K�,�f劷�ü�ɣ4Wp�}gM�/rI"-��[�^��M�C��hP��)O�30PF�%3T�+�~rs{��t �U���%��=����	����T��"����!Į�I>����;��g�Xj3<���<j�����}��~��?@����u�fDO~�P��F�N�E���|%Am�z吕�݆JJl;a"�zQB~*��j�����)|�<W��.��cPd�'�v�	�y漣yk�QB�{ d��ѿD�D�2��;-�+K�8̓�j����w4�]�:&�=��k]Gjў�,_���}��|Z�I�į^;s��߁�s#��{^�'�u����Q�(�����-h����|������s�aܕ:��*�j,_8�U������\������ʥ���D��@h�$�Kŧtg=;��=�Dr���#@K������w%Z��i��7��N�@�
�9ކ@Zߜ�d��ϐ1���y���b���F-3�=������EW��q7���z�]�KN��Pbϥ���rN�)�*�;N'F��ی��/L���ċ�2��A������l��AB�?Vae/x�Z�;��d�j��=���7;SK�+�.��N�����鷋�'�S��Tj�0��a�gs��N�p�\ӷ��pS0OY��/#�I�=�Y�΋tۘn�AG\���~n�x����%	��#��n�e�/.+�]0=];�R��a
=^H���W��kw��dkF��E�7>|����b倄gY�I���Oupdn���F�&+=@H�����K����[}��ښ&�z���>�[�J�aE��)�{E���bM��.`Y.��F�@k�����ß�MP:l���-+�0c��Qz�����3�x�S���71�z�˯��̿��^��G�@�r��K�\<�~;��E�<�aQovˁ�\�J8E�wˎW޶9�R�����D&��5��@!W�av\J�!kU�ܡt���$-8����Y ��B�
��g�LA����m�-X��1u��-�=�N�7_r�C)ˑ�e~���?�h�d�W1��Y�]�2BH���d+CEQm&�#� i�E��F�"0n�"�аg���kT�R�y��`����k�xVc�wLw� �L�"5(%�QhR���Oq���E�ǡ��Օq���-�����7�J�*��{��_d͟0���Խ�z98�#b��l�3��fk��f�kU� V�F�����LLw2��,`�/�X#��/l���T~��|多�j��͏8g�.D�CA��4̫����TAVjc�K���h	�>UL �����1�l҃��i���>�g��s��;�q�a-�P��[�1y�9����sRt�v��o*!���8�6�Ο1��m�}Jß]��;ٻ�R�r�B?���>��
�l��a!��/���������D�,�$�F�ߝ��'�6h�w>m���x�G8���`����v{	���^�����0+�(]}�`���뼿� obtюq��d$�O=&�\���'
1��a(ֲޕg&�%�>�ěk�C�;8eON�xD�<���X��.�]CԒ4���tf}��0���L���8�p���F��ig��Ӑ<�)���͢l8��?4<#��T��N,��k�M�QT��a��ւ]�u9�y�+�0P���|�)G�ԝ�ky�-�`���*m1���[��2h����4x���<�hl��t5�C�szN�P��4�x�;�ك@tY.��0��[�K�
߉­3�ܴ�8���d aׄ$T����]�e4ѫ-ZBb2�w�4&��vN
,r����
PS�^��&�)�\��	ͭ������v#<�4n��L�M���=�+��b�$�.����ݱ��iU,x�.p�����}}�d�;�r���"z����(�I\��ǐ�K0�m���/`�IW�S1J1@̵\�T
�7��+S�	�*H�R����0���*ݹu����P���	���Q!a�ѷT��_œiZX�Z���-�x][|&���ߥ�� �I]�h{�rV�d�|_�� E&U럣�X��61 �J���������c�`t�9�L�x�'��b7bf���vO�fpS`�-�.��\�D�D�Tu;^�MH�ܗDh=����=��Է��{�Rk��fy��;%1����X��j��G��Z>�@L�Dd�Y<�)	���������Z-��_1�/>(�tt�>)\�@]�'� #�W�K�G�%ls/Td3�!�p.����Ww�2f-E�D���9rDە�j ���� �?"�D �,cUt58��Uט��4yz�U���;!�J=�(���I�E�
_���i�S����v��v3W��S�m|��I�b��9Fɿ�a����$	�w��G��۰�f�}]��\?\t$pv��H}ާ�y����,�׉�4яMA���e�^�lv����Ê�H�\�!���0��̦	�^(��FV�kH�^��	���a=��~��P����q"�aX�Qu��K9�����p�-���?�-��&����s�S�3��c��� �a>��G��G]�_�\o�y	YA��.�s����#����F�*~�St��t�'-[��zU�s�ld�_5~���l���������[�W���%�Bj٧k���8N]�]&rZ^2)���;Q9d��W��;�j��T��(Kw�}R����q�?�;d�{�+:��
pC�ݬMR�dzd坕��+�c] �}~�TH~�r�+�����ѥ�1ù�c��5O|����<�q���O�v��2���-&T��Zc���܈��As�^�~��?�ɏ��lv�"�����v��m��3�s[&{w����s܇cC8$��F�H��1TrC��2��RD��69�S].s��2g@���;��J�I�o�q���N ;��:~S)Xi�p�<b�n�rCj�=;��#���&V��r�
P��_����F\����@E8㘶�Kȹ�򶼜;I�-��j�gp�z��jGZ��b���\��U*_ͳR.[B�W�&� и�tL;��]���-^��K$�9L�=@�o�"�
�8	�O�]*��7
������f$'v霪6@]7:�W�Ox��<Z���H�R�����~5�_�T5.}����{\���W#i�dZ*y�B��`e�R��0��x.�vwo�28��S`���Q&aT�K��5��g(w5ܹ���N�-�Q�5(:KP�}r�l���IP�}�v'!M���<�m�9��Tȫ-c�k����<��>�v8m���za���C,%�Ө�3�Sn�{�We
�������}�dls
y�/6$�\n%�C_]�ajGV���mw
�Û�(58�(~������^���ω�3��R�ߘM}���w7�c>8bO%�Q��I�'4��v�г{���J@��Nim�x��I�cR���x�b���%`i��
ۗ7U��ms1JSqc"�hѸ�,�����6��i��w󋣊,�`���3L�pVJ��
Y)Dh}�o�֤+<b�l�;�V��m�#B���YHy*�~�2&eOăU���BY�nP�Q�.~4��p�s��B �أ
������$r���rT�(*��ѽq����FC]��6�c�ZXp^��-Ja5��r����ک�6��Ђ(��s����i��5F� 
5pL�\+����j�R�{�*�?�'�6{��e���e�n�5�{�7V�(v�U�e>��Npі�E�#++"�g�*�[p�
��V	�e�6@���+�=�0S�mW��xX�
������E�ߡ
Ȑ���
o�,<;_Ma%�z�4���z�`$����+8ı�.M��j}2'g�8�a��B�-��	S|�O`��4A����F���.��,����D�3.�trW�4Uxa0Df
j��h��8�z E��%Ic:�p������Y��"��9@4wH���픱H�DE:=%8$):0	e<8�����u	��Է����1��em)�hRiB�3 8��\a_mFi��y4䮣�-:����������o�`"�J[�T�:E�Z8�ލH�?'a�N�)yc��v7��t���z�,+��b�����57�}Ә���H��"�r�b�tR�������L��x����$Z�Or�7\ڐOA��H{n��46�4�	EQ�,<�W�=)#[�û������]�>�d��y�Z�qEw��I���M�}B�z�<�� ���G��p�{�@����)����},j�׶".��7����S��9N �\0��׎�J꧰ơt�^r��{�܎AT������޵!t����ءS��2�0��O�;�6���k%-��Ё=?�6ǁ�q��ĺ  ������������)�7�@j�p�Y���v�eș@`�Ԩ�',�~��u��C��s�z9L�y�Wc#��&;�3�dX�����*��!W-D_����%��� 2����3���^@���Q�F�B����+tWƋ&C
&�~J��Y��xM�c�����]~'����ut@9j"�<��W�0�o(��&iDɛ3�3.묋h�s��A�8e���q9�
< }��n������H.�+ר�6�����0_���A^Mun�M�J�hF�	����I�{Nڇ���U@�U㺮<� ,F&�̂�`�^P/4�ޅx^@n��j�?�g�����T4������I׌s��Ȳx6�e(%H-��V\���x�B�%�����d�z깓���P[���"W�0�pwx��w��ɨÚx�M���d����� �4���E[zI�Z�ɫ�.X���o@ m�BSk�y��R+c�~b�8�;/(+�a�aE:����6� ¶�F\T�M4V��E8����F�p��F­w~�RG���)��U0���K��VGCv���/<�O��+�b0^;���r���S�Ge���V#1p)��|{��!�z�����0E����2R��W%0�P������:Z�%�]z%��D?qH�F�ō/�4ڮ9�O`��S��mM��K���k�z��;�Xj�!<,�UX��8Z�l�Ǹ���GL���:
����F,��n��̑d����~}���4�'�p��"���"��TI��6��W�w��%��h���d�	����{G��V���{^/V�Sn6m�љʮ+�96�U��4��!����]�^:���W5��=
�H�!�C*�8�S�6ՌG���nFI���Ԅ`��5�g+��Z���b�iy&��	k��K«���vJvVV��2�����3�9Q
� z+;�Y��MTc8qʤ���6��=��t�> Tq�(����{-�h�Ùl�47�f��o���²���p*�l��;����[�����	�|ǵ!$d0�P��>b�\�u뼲g=��\_T�	F��
�!��iQB&�ꊧ�r����GN3�;r���gtTyx��e^6���<���#�$2�������ߢ�u�)Yl\���r��WMIb�d�oen	n+�|��Þ�p�9�m�;����Y�9���q9��/�����}�db��[��6*�0K�[����<8Z�%��}��'���.�����1�&oB!-*�&TFrֈ���u�R���{xHL���&T���W7����'1�.�gv�:�;��H��>�����BF��{۶e�j*��Y���3��e�4��&)*O���ԂK��]�yb\�s(Z���H�����Ex�����Sr�y9�5�P��sk&7���w������w*��~x(�k)����2n�G���hΗ���6tf�6ۚux�`�<o)�	� ^b%i��ᖪ�1�uE�6$6��C��1u����<�܏۔S��1mj�'~^ok��G�v�2�pI�U�^Aj�TE	�������'r�7��3��)���%[��׃��L�������������Ҙj����S��������I��4ҥ�я�Vݸ����/W���$?�:�-9ө�:��(6B��t��zi�|4���7��8M8��Y�`O(��}3� bP0��d=ɠ�.ý^�n�u}�
4�\�y%�|S,�+��d��W�!�� aP�T����A�v:���bh@���!L������/! �U�������wW�qbK?�7��*�]SdA��T,gt�1�@����ߩ�̬�CeL4��*2�|r
�a�%�����Ƴ{Xbo�$X�J�a�n���?�7�)��ɟ�c��x�dλ-�|��Ǜ�}���Qn������I㟇�T L��Ǥ(ud��?�a���T�X�R�8%]��L����~h��bw�.����r�Q�O�d�k�i���\�"�?����p��h���"|<���Pm"�L��^�������O�PJ�4Q�]�	kδ��������?��f��hw�}��ѳ�5K�:�j���2���AR[�=u(���W�e���s]�W�&�IP�����mpV6����`?u�k��:'tHM�r��̓ʁ��z��[��@e^����s���v�#�P ��Ri���nٓ���!M� ���ao7b�i�N�b��� ����(��<�P����� -���G^�G72&������F[ݹ
m�������ּ��9��VY��/_�h6���ը$���bYS��s�s����� =:S�?�X.c��M�m�,ťׅ�(�v]�Aj�؋g��?T;��?�Q��Wo\_p���ZTcT�v����<n��<����tN�W�6�!ANw��2��=!����e��ɟ��b1��
Q��X�)�N!�O�f����W�E����jF�))%I����I7k�N���%�1�R�2��C�kk�]�@�Dj��Y��_�G%��t��f
�Yo�7�xx��5���~?���?#Hy�c�N�ZAu�,e�6�8�;��%�X)b>�UQ�c��)hClrxȕ*I#�F"�nj�4u�N+H̬0;��f��@�8��@j�����+UA(��j�D��=��Q\�����+��m/��ٗ�,6!�J���qz,���{z�rD"x�� �
�����9��ijN��\
�b�����A�/Lmv+�i��Y�#R��t��������j�J�o3X&�ԤD��z�S��t�_�k��A��E�7��� �i�i����>��]�Rj	q)I��4�R���z��d����(#�OY���Z3�/�?���]j�Nt�A�ڀ��z��)+I��+:!�"���z���T���U��?n&*�����y}e�/W��-dV��i�/y~�#�.��;q�=2�t&"Kb?漌h�:�,.��[ќ%̚&y���X��vt6{�?,�G}���.jB-�f���$��9A��@��
�=�w�O7���n>!����b�(8��%G�������)S�����\��H�$�/iO2!���h���W�f!	n.g$k���V�J��{Em��	+"]K�m�s/�ܶ��Fd�,��.�Ǣ^���L�P-�3><�ydB�G�xne�@t�{o���q8Y/�_@S�kjȿ�A��Œ^)�7��Z<X��>:\Xqi�M���i��L���٘����Y�^	���^��v��O��4�4c-��F\g���,b�#����e�8Q�ߨ0�ި���?+WZo��G��Y���-�!q^�&m�"I,w��u�5�3��0�����f�,B�R֒9d�|~��kL�([4Cz�o�4�)w���}��(��>�/�z�Qos�c&�+h =�l��Ֆ
Ѣ��,�# C"��� i.I��K�p�h\3i��W�\*��j����K��'�1�/A䊫+��z�Ɔ  �S/S2��a���~=%ȎC�!]hƥ�J8,�eh(#�������x-G=	GX��r��7��P*�l�%AŔw[��A31K��v76��t�<c"�a�:�ʽDC��GN%3s$�@1#��"���7�]�^-�s�ث�O,�!P%�wy����P���W/�����K�C��3@@�g��g�8�,#`S�^�[�N�����D�O2�;�� ��?�Q�8�"J,?�3���Iˁ.��⃑v������Ҋ��~~O��ہt�	*��ă{�O��Z%C)�΢�?���45_�tӣ{ Hy6;�>��K�9���w<o�*W�5B��hP�r�+�[��z�9����-\��x�[���s�P׏�9���Ҽ	{�uv��@d���$<��9���Ŕ�:�m��*)0���p�w1d����k3g�>3ʏ4Ո�� XOS�ыπa�����.�ѝ+"����,��x��a8U�O
|�ԝ�A���rWoxS�}�f����o��k�i ��?[�5PۅQXzm��-�a��y��Bf=�+]�JȂ2xծ�G�q48@��qD�!ȋ��K;������4~��ɓ~��*���5{!� ��o��ڠ���GA,��в��>��^v���7fS��2�|�Wջ	Z�������8ʛ ����i�h����u�3x�wk,�P,Y� �]�F���N][���P��5��ݘ�嘠>Z��������,��w�j�[>�|~�
O ü1����&$�;ܬ�9��|�w�)qr��6��˙X�)�m�;�2�8ff�.����E���ˇ��;l��e��0RЁ6�̻2��6�k�z���H�1�Ye�s���ll-?a].�����x����a�~�(0<��L���<�������� 5�PpvX�+�3�##6��kDѴ������Iq�EUo�ˇ��\�!/!�m�����1�i"BD��M;�(f9��W�)���[t鍓�[��	��	=�k/[�;eQ.�?;�Et�N�'����7�mz)�W��M6N[���؃�`otR��Ra,Hs:*b�>������,���<�xJf�A�p(%J�Fh��4ٲ���[?>w��$���u���'��JnBG��e �(O�9b�F�-��mi��&i@la�#�,�2E�Az]&��l�u��7�S�������i#Ȏ�y��5^L���Q�×��<�=d.��e/N0J��r��#x��::x�$�G�Lo���.H�xɪM�.Bۿ��^�
a;I$���5��*�2j�$�g%I�GǪB��@*���Kn��S�')��Qm8,\�(�.�]q��zdW�q��G��/e�D�j}�0�A����Z��3|<�ŔSC���z�f7|41F��%��)-�Q��2���]
���*� m������鹿w����Lض�[��Ƒ�w��wW��#Ǐ�!B�i9=�\f<��ǁ[L�3b߀j4��U������:�����$dI`�`�&���	��Z�ޱ�~a�oaњ�����^y�q$�1��=�B�������2�� g�n�� �s�X
������G'm>�9�:̻��1��^Q�Vʁ'�
�a��h����H���P�L�4�	r
�ܽ��J\�#�\=�ڊ���8f;>�a3��|}KO']���X%�zf�9�B�� J _��!�
�^�!Ri�Tg|�_���^e��Dє�x7#��Rn:X�އs�1L૳��\��x?��o��՗�[��R$����6
����7�D~���*���"�O�s�ސ����W�87�&u&����� 6욞%�h��}>o���֏P]��}[q��QX���a��0c�{(*��4��ͼX���)Δ�A��pF]�-sw�Қۥ�P#sf>@�;&��{v�sY�ƪ1�h�2_�"�����X�����z��X�\$!{?�W��F�$�!+,�<Nw��K(/�I�
�[�5I�����&`R�,�i�O�����Un��,�]2�.��;�{�$]�O��{���/�g�Gp3քfpO#�GdQ�C;��8	�U��W�)��-R\�������Q��16��?H� ��XFw��!_3��|W<dt==+�����M�ơ,��pRӿC8pS���h
��Z����,5��V��Af��͘61�8�x�a6�}��6�+Q��GO|X�݀KF���Q8����Fژk$e��"�#wik=���Z���dv�U�^m��KJ[��D&;��x�#rց�J�� u�����v�y]5/�]��Bv�vꈶ��B�kX��E g�%Q@�w�L�H-n�}��7����@��2���K�V�E�"�7a2У���g��']|��]�)��\cd$r ����S�{jq��f���Y`TMv�e�`����v���%���	�����סfR��e>�p��s��M� `�U��g�5q�c����+������{S_Q5,��:���c[c�&9S�(͂(�t;"Qw�?%�d���ݨi��-�����ۤ�vi����UhY���p��r͇� r��lANnS�{��R.��'�i��J�S���1�h�h��<�yE3M0����$������阅<�(�/����I�Ἧ�o��~$���n�CTϽs�B��C�M?߉:L�rЅ���󂣝�T ���a����V�S�(�i�)���ڵ�h�b�c�Uj�yv�K�b*�6*��Vf���W�Fb��l:��m��^�e���J���Q&E��ZE:S�.���Y&p��)˴�B���MjD��81�pt����^�&��
�y0��T�Y�La�}�K���Lh%^F��?`3S:����X�6�qr���|��=���k�ݽ��}Op�=ra����A���>`?��\�d���(*kkH�i�9���Mb�d���9���+;�|��Ȳ1氕�"_;��P%�x�g���?�X����F1�� ~��oq��n'	1�?�e}q����`~g��:����ӡ��yZ/ѴP�A�S��N@�Y�H���!ۃ��^�}X�|�����o��*O3y��L,k���m�[��I-�5 Ză�ڲa��%'br�Jl�Ȃ�N�� K����u����猷��D}sڶ���Y���g��G�qԤ/Z�E+�y�(.�.P��7�N:��&�y��1�j��qc6�T/J�7�C���� L/��>>X��eŀa�ng���v}�V�GJf��+�]IZF���ˊ�7]�;��.�vmPJT�������O����A�vug]B�]�����S$a��pb��@鬧��s���K�j��3��3[�{�N-���{q�da�:Oq�!�L󇤏 �Ek�N���Ns�z[�vnT�-c�jV�Yp���m��0���"2h��)b`��]W[��*E�Ϊ����*��ʬ_Ѯ-�=��jx���3U5���Σn,��dp�~�L/�g�]ɳ(s}hϼ��?(T�ˬ	�˺~#��%^;PG	��N��d�ݥ|�˙\��5��/�w�l���غ��̡��d�u9ڢ��]�b�7�q463Ye,�Vӳ8��e�{��X��J�9"»�%s�^į �摌��/��h'R�u@���x�$�zY��H�y=�ٯL����:�/+ֿ���#�c�}� \̮�Wī� A����8�ڊWk�?��DE�e����{j�Ly�D�&����M����q�\�� F˾�G�Δ�(�9,.�����j���1U��_��l	� 8ډʣ��Z4�)؈�]�5�}�'œ����Vs��/��!	������:�]�<9��.h���+L�REd|,Qq���)�������~q�R�@n�=�<�f,w
�zP��'�HmHC��].O!6k��UL9,�Sԁ}�?�!ZO"e	
[��6��ʧ �VH<$���x�-��1Y8�|�
�.;�6a`��W�a��Z|�Y��*z�S�>Qe����h���.ܴ3mtuYt��t�R���L?����!\��?��Y��1H�d�c"Mt�����(s��,8j#�kY�l#�q.��?� �y�h�l�{�#\���'��[�CקE�:(���퐥Ch�����~���huأ��VTX�]�_�����i�b�G���<T]��L���B��n<(x���-a�b#~Kܠ�j6�w+c*�գ��|ހ{!�H�<$�j���'/o��/�!R��,�Xz���w��vfG˶)��7e�����Cɟ���T����x���每ҩ ��_�:���B�f.�b!�J����1  {�Q�)����] �Ӭ���`T�*N%!�)C�K�7�7��ճD�U�����v*}�m|gc�x
v0)�$���^{g.=?��^�l�q8눓.���$��bm>�6\����Z����$6=X�߈#f������R���f�������y�q�Ԥ�z/	裂w��ϵ�tH�;��Σ2�\2�l��[�3��,ޅt�zwx�t&�D\��o�v��o�;y-���+wr���41#]��t��ex��M=���&`���q�a+��R鬩η�r��H�P,�b��c^M����aW�Y���ހ��
e;;�'�:EіB�,?&}Ý�BZ"̸W��V%�:�Z }��]�:	�&�,t.p?-^UH�v
6����A��2.��@�\,���V�fx�ć���Y'��t�����:�Iig3.CS1��ԺX]r���H:%��� �:vy>�G�@�񩸸R_zz��w�hy'9d���*
�<e��+O��}�Bb�
�� �<Hr�7����T-�;����#�i�Ng�L���Va<^7 ăf�j����;Wu�3C -�����c��;���u��[&ݝ��"�������P5� Hԙ�=����8�p'�:щ(=Zz`�U�'9�ίU�����d�(�������P�Ԭh�;�=���N��4�� f._
{�*�.��̻[`1��v�����'%���/ڶ��%��OWn�3�8G���8�T��	u�ʥ`�y��. ��$:Q������p��^��
�q��&oS2UA�Z�X.:��`��W���{��N��0�^�~�E�Z�ɡ�6��u��NXw%m)�%N�.�c���^�5�����"�F��o �`΃�w�d��L��_�~�]�B�ɭШv�xZ��1��@�ϙ�*��ءX�6>�!
&ɯP�� �l6������ݙ�4 9� ��L��ծ���w|��,�X�m�K��e�Ԍ���}]b���Z�j�gU�챋Ly�|��$p(����S4�r������T��:�['�R�c���� �"�����T��~��C|� ��ӎ��Qa�Y@����D��(��D�A���V/N4�����-��T3ׁ���RR�)�̀B!
xQ��������蓨~�����{i��5N��z�<V��LNtw���Q�PD��T����wuȊ����O����|�l�`�0�셔�������H6�]��ˬO��u�C��60�%����@�%V�y��z
6�g'3�X�kƶZu��.���U*�\�/�TU�O��Ѫo��`m��5��V��+�L�dl��kڑBc��U ���=�q�O��x�{[h�� O��CJ|� ��ܟm��B�;�,�N���g|�C
�;��f��|\"�Q�w������+;��·����,Y*-rm���
D���D_�π/��`Y\���i���y>c
zq�h��ِ��R�j�&��@^�q`��\�/��d�*�$l�RiL��8w㩄�8��ns
\O��4�F���UfG�<R���g�gj��@��K�C�yY�9�y���:iF[��?�k���~�M���#ı��v��6qLP���NT��r#~%2�Yn��+�~�r�e��#5i���}r
o�O~�,S��VG�ֳ{�/��.
��˶�%�����%�F������-6�w�id"\97��N�d�feJ%�����Qk73�,|��c��c�o�Ը�ՅV����*p橯�3�XSF��-���Hr���n�ڟ6���ͪ�s�!�vpa�H�؀����ixzo����e�����`.!�yma(� ��$+�F�w�'P����#eKw�����j*ۿ�|���@�/���`0����G �jz���m�=͑ܯ?��^���U��Z�0����Bl0���w�Qan�H�F; '��Kl:xc��y���p,�,�.���:���K�]��`jlO%`Õ�J�����7�<��Ŧ���?��%��	�k!u��y�XR'kX�?��� l�E_��/��ƙJק��s��:��m~n/�'p�4�W�gOy� �hx}�oVCS�@�X�J��'�+P����=�^&�.��Y������A�s��W����C[�R3��/l7 -4��u�Jft�e@1�G�q���?��l���8[חJEuO��i��s��.��������r�-y�����Db��m�cy�p~��-)�mG*���Ny)<p�<d/]�\�?�H����;�7Z�)�D����#�����+��� r�=��K�C �Z`dY8"�� 3���a�	�]j(q}@�C��=�zb������_.8�[�ˬU�.Wd~��OG���@�0�{.^�R�e���$8D`��}�%�Xx�5���*�v��g��q.�w-:A/~����9��tL�wxn�����LG�i����I�Y�Y�ƕ_�@{�^
��Uٹ�vYxW�s�m����~��=�[�!m���@�f��dp��#i�6��5t����ᥛ�D��s\�^P�qd\�F�﵈�2��e�����u�ϒ�eܦj'iry�_ҁd�����!�f����X�$\�g���%{����R9�5 !��y�܊��P����μ뎺�/x���hu½�IDX�*�AA��*��>l-1*Q�質�1���i�`����Ǡ`(qX'�둩l��rt��3r�&�#H���j"S�/F�Y\�d����O ��J���$����X��̅N����s����%>a�fU����ͧ*���A���^o�f.:<T��`������@���횂��1��q<.�9̕IY\b�������$.�b��I�c^��U�j�����FG�W��|�a���5��Ӆ��yuɈ�.��F];z1��9n,�h}�CL��&w_8]��?���h�߯:�r4���*^wL'bH�ʛ�����5:�!�m�/qB�|j�(cl�	�� YE½��M^�bo6�{�,�����L�~O�S�U���񪘥��j�m7#~c��q��]'��_����T��Ci}�q�����'X�L������w��_q���]�/f�
|B(w4T2 P4�AH�P3D*��2q��UODM�0�
,�O뭤�|�Rň���(.D�X�0��h��|�e����(N2>���Ġ���*���E�h<��M�A���ls��M[�> O�&��/B�,b��g���x��&ߒNu�(/�0@�8B:x{��ҧj|�4�O���d�d���IV6I�3�TT��J���%�_��я�u8�/��2W8�!Gp�I����3��|"䜬2/˃+^ Ҏ��>�1Ƨ=�ͫ�Ej��xz�G*�95m�Q�JCto����u|�ʾ@K��;n�N}��l�����F$����p )�))ZiZ7jw<��6�]$y,�K�"�Kd��1nd� {�6�J���Ɵ��1�vw��^�����
O����}��sϜ�q�@97Њ��*V�~�kv�P��S�v������H
��U�#�;M '��t�Ka�Oqʺ��9riѳ���N��sd$��Pd$�`K�lu�>Q��/���Q���q9Rd���+^'�4�����/'� F��xᨷ�� ���hL�ĺ�<a(m�;k|0�(ЎJ�f��5�C����=���M �H߈�zn����$��͂��D�?���xk�՜Hl�t�#�pr���h�KgFĻ��fI���`p���#g����)n�[kJh���;�߁�s$&z!��4]�)vd�k�fqy���Dw
��_�o�H���%����k��0v�L݊�3��gS0b���_��8{צU��'
�Rx!�D�T"]�j�I����
/,�-�D�e�;�n��c��pJ}���Qp�T����N�����s��jV�F���Ǹ�����7���ԏ�n�h�{���H�;��9!n���)n�<o�O�����v� u��]TӍ�k
�[���oV��N�x��^{��'���zM�i$�S<���
�Q�?���3u����kV�ɸ�l��g&����\"��Wp��تj�p�˕��#�E�;%?A�C��7����b�Ҥh�?*uk�n/b��� �-ֲ��ӂH2�9��ڨ�z�7�!97	��A��@lK	��
�3[���������C���=	в�����o4 �d��L� ��k���	�7:����d^s�����vȳ��j���Ij����t�:O�b�1�w��LE�}����'��1a��ƍ�u�X�P�<����C��l,U8�	�Wa6JR���P'b��(`I��:�k�g��(p�;��k������k_�櫰�Y}����:d�� Om�/�,>�'���;���ƪ9���:���75|ѡ�P)A�)�)��5���&F��t�6
27�5�	-:�(���c���p�F7��~kAieEm"O����ۛ���ɸQ��t��&�{�qR@}5��,$RSqQ��,U��5@6)]��K����	�_�{�PqaU_���9DV6�F=P��'�����J���rEs=(CIZXƹ�\��N��c}ˍ�5�G�BGQ�W���<�Y�Q�?N�o�μ�Xhi$-��@��Vi#%F�!^�E8��S�τ+�cMS���;�Ms�B���.r����K��m�����h���fd2�l�|5%[\�@��ƽ���hu�P���_�$8jv�D+=�Ħ�a�ĳzu�b{j�Ey}b��,W�2z�>HC�X�A�����K��Z�1��HJ��=g:;L(�b��h�ڔ��6[�e�z�!t��qF�
�����[-�MRm �rϳ�0�xOyY���E\���	��D���Bu�m���;��*2 	�����O ,AG�Ih*�x[Wʦ#v�M�i5��/y�Jؠ��űh�E%>nO���a�'�bJ�s֔��	��]f���J�Q��҇W��Ņ����r[��>;�����%	�CzPK�q�MG�kD�j��}�D�?�˭X+����c���n�k��}_�Q��1#�O���x�j��TD<��?vO!���JϜ}a��3��|����؛�UC�����'w4XCbG	|���G��94�X�^<����0Z�p!uVb)Ƚ ��#r죖 F�*�x@2����a2-f�xr�	�S�|� ��B���XflDH��ݎv[4Қ��t�ؚ`�DV0��6�L>��'G����F8��t`��������I���Q�Ҩ��)L����
��rzb`�-z�=�w!���̎�������20�Ә��������kC:���	�ZX��"���3�.n�c@,+���0�9�wbw����}E��6�w�b���J�N��\x�7�����R�Ɠ�*5I=����R'��Mpe~D�����	���wl��	A�s��i�r(ӓX��㙛�Z����$3L���Ttx��Qm�ż��7e�Kh�jb�P�:�\��Z�<��f�L��:�&��T���MF[����m c�ɋ����)v2�g9#m[+K}	3�o�&��J�M��8�����,D�l�<���*�t�4���Z�����c!�d	X���^i_�p`�`��
�~m�Z�m]x��[�Ĉ"���XC7��$y���G���Bگ�׳Pj)6����bȚGF�O�f&��|q��Y����l�&�r3��Lf�rE�4��+�j�MJ��ĊCq�H��Nӳ
Ǳ]�7�D��wɵ!$`N�N	5��;��ئ����
7��X�1�A���r��E��@���N��)_��y�x��]VO�G��D5�<0�s�\�ZO匃��(�T�~��i��	�"�s�Ӊ6�0>��<� L�ܩ:��o��T�C�e�F;�/��{ڏ�Z��4A*=�I:�	����Y*��iH��	a)Q�b4�t]����8����Cx� ��a �A���^�]SZ,�}1~���Kxf�?f��D&�RP��Q��ՠ���'*�]p�g�rO@�ǹ��`h���S���q��rd�����4S���݈3T���"V3�*"0�����} Q2�`+,�@i��ܒ�<��sm� 9��=(z���f��#�K�r�4*����D3���ߔX���gO�)�����E�]� A /I+ρ�C�9�hN�BEE\��rh��/�|�=ty��2i��_�-��2�s�2�b��sU���%��ɗt-�|hZزy��P�3bH��I�p��91�_��6�kԩؼ�~�<���K*_N1�����F�x��k���>`��ܴ��_�P�"�qy3�9EÐ=o�m�/��n�i�/	i���'H��:3Q�&��_ B4�s����Z`�;�X��ʚ�o�He[77��[�4�)��^�H	���T��S�u2�k�:�R\s��3;}��'[���:�./*0������vW�f	��G�g>mӬH'v�`�������v7g���\��lӪ�1;�x)	���y�xX�������+�˹�>rDT�����46�����1�\����������V�c�f�_vKZ����b�C�f�,��x���h�$^������Ѽ�;ax�?D*���h��(�8֯V��y|��ApC����	5��}�� �C�Go�XC`�O��C�*Ѡ�yn?��D~���Q��I0���&�J��*&+#���C�s��\��7eJ��
��>�L!�����Cu�r���i��J\�,�a]Z�M�Q";�W7�=�ސ�*�
�B�X?�zN�;�l��'[56�߁��p��`��>��CH%ƾ�<'�B����N�W_X�j�rF}�q���~�W�H6;��\�(ծ�C}�JZM�7k~�_�ďN�"X���	�a�9��;�����<vYM,;���ˆ�v8�-�~�%x?w����Q���!7j���!�el8͞[䆦�b#&�T��W�Vc�v��C�1��:������i��F�4�9��`���?CNE숸�X�S������Y�i�8�9:���Tn(���$��q9m���]�>�~�tݟ�ZY���΄�w��=ą��M�M�j�|r����oG���K��ϐ�L�,���[d����V-U��뼁��r�#�����@�B��/�c�!^ИI��������J�eR����*�Q)w5������h
D��9˫}:h�ߍ�[�X�i@=��P�j��,ui9��eȺ�͈�!�N�a������`cQk��?�d���z��^Ո�1�Ӆc��ҭ��J�r�������C�s�ҭ2*�c0@$N��~R.�ȊK���ܩ�&�Ư�!���C�t��0j�<�2��eU�L�ə�Ph�{Tn�)[�+� ��}i�4'F2E������D�Y��mo����WJ��ļq,d�W���r���=)ʁ)���X�/S:�<��
�2�ϭ\���A�����4"N��0���}�O��ԧ���v����@T�+��u��t�t��F%�S�[�s��X���?/���q{��γ�*���'j2��B�����[|���}��N״W��=��Y�f7��ϣ>�R�U[ �Z�n�U%z�5�Ig5�0@:��!!�W��_%<�a�rP�/lǷ���|7�s�@��,��� &+���.�dk����Z�9L�v4�OE�;Ci�~QbO�6p���͗br!�i��σ�Q�l5G -�k�E���[�z�o}�����l?�������,Z��d`�KS�)l�����DW�L͸Ng�X��E�S4H��3P�ez�����C�/����x���|�C�p�!��=%�`A������Hb���H��o� pcab�>	l���]b�8Gr�I꒔(�D�m��5�޵�9cPT�2Dێ�2�.��)�Xc^Y�S� ���w}�fS�Qs��k�I{��
�J�1�UK����f{(4c2�U��U�L�|�����k2��l�M7���z�mb���j��>�=P�G�Q@�}�b�D%_p¶x�i��<���ѾP�TY�E�Mi�5�I����ɺHZ�L��ȶ�\�L��K�T\-�9���B��2�����Зd��(]n��Ԥ!�)oW�>�/����C7Uձ�d0V�K���N"&���H��0�g��������a`�|�D������ɨ���l���rU������~��L��M��)Y	 �be� Zݾ���KRł�F��ꚫ^/y�i��*W���*�����-����.���	�F��{,�lf9!����8\VdɄ�+E�r��L��A�	u���Ȩ��b}���x���dXmPMH�ѩ�.=��w߫������k��f��	����Y_�z-���.ޚ�95K��*���q�6*����%�v���~��X�J�.8������m����pd"pz�noS)}������wD��>��3>C Oj�_H��k垨��Eߙ?H�t���CI��_�.��4ѠQ�k H��{Y��55�:pG�E�A$W�l�?c�~̜k�U����7'����h��X�������d�����
V�/�P��Ǉz�5�ւ���O�t�xf�d�)g��6�1�2�_A�D.���v���1蠌OQ���>�����Y!x$�$�hj��(0�Mu��8�:$�fV軘z����p��`��U��2G��u�Tj	����h�qcP��?v-�u���i`qŸe�N5J��,8����C!~�d^�(ٳ��yhr J��� 	������bBQ�tM+ĺ"����pm+!�	�'���T�t/����i5.�4]�67KfK~�p�Y�� <dHEo6��t딻���%�����ωӷ�h{#��N��{�2/X[���b�S�3Q\٠V;�%�	��'�p_S�hK�{;�X�N���7!t2�l[�6�p2@?����"�� ��>��*� $��q��^s�30�T�V�y
�*V�`�lc�0�i�R�H���Y�S���s:ȴ5�����8�=�41����.b6x�u��Ep�2BI"������F~x9X��M�3s>f����~*���%Y�_m�ރ�5e��ko>�.`�=��eJ�-�ߢ�]�/�1�63������!/�������o���F�.��r;�CX|�uGwW��g`~@�h�U�䝌=7%=��$����k�<@�P�;<�r���{ϧJR�ιH�\�r���8���7��0r����|E����[�;v��9����L��Q�I�?GN"٧VU;PH��
�*�A�A��ɦ(Y-3ۈ) Ԍ�7O�\������g�
���]����m{¬	�.��J��h�3���X F��Q
,��[�������~c�-;�I5�k�#�V�ۉ�A#��&��4wqʕ�J5/y#R2��x���a���+��5w�/{��U���_]��[0��Z�+C�4���=��qfI3��,��('E�]jL0I��#�\��4�t:e�Ą��">P�O�&�?�R�8˳�m�҉>)���ԙ􌴟���ɻZ��5���g�gѼB8��.�R��9 �,�����<
ru���D7��;��]��^��'m�p˫�?�1��c�͍����8���,��ST5]L��{�w?{c�#g�����'��l��!3)����2�
$"����H̴N�4`��˯���cW���c��7�:��3�D�k%Q���>�'�S�lrB�m�Y�@K��	}0��9튕w [i�-�_8�M�>U�A�iZ3-�67�$��Tj��V0�ݖ^R�v�n`G|xt�igQ�uio����ƗR���he�N���B�����an�ţ�N���91�E;�.R����`��&�{�i��&�dGo�����ⷳ@kz��O|�lJ�s&�/���8������7"b3z�,� }e�}�X�Q2�y�� ��hg{BaSL��*Dz���@�ҽ���:����Y��2��>E�$��:t�K������n�r���U�����#o`v�cf\�r1g�ng��+��3���k�g�u���0(Z��2�f�&��:���~�y4���4d�l �
m^�}_�M��9�.�T���B 7%� oe��h����M|��G���R�z���VE�}�L-b�g-�Grkn�:%E?�D@�芝@��¯�"��ħ?�s�@*r�|ŐPJ�m��<�ΗC��gtqO+�$��
�c��ǅ���C�����95l�C��7y���,Ȏ�N>�\>"��35�f8�nYV��|�5Y�T~"Kz�Mea�B�8���s
�9��9	�]Xn�~F5H͎F�(y+'qd��N
�]C�uP��������3��Vu��ŞD�~\���fc<�QK�V�~���)V�#F� :�����h)�U�}(CU>+ա�U�"w�P��Ӷ�c�8l�|�����-A}���o�����u�Ҋa����W����33�Z��S�+�f�sH���L&�@a�C�����(�#.D���7���x8�e-7�$�b�������,��!�s�1M��h$�l�y2��!��|�����ٜpY�^\���p�w�Vo�fc�|���6"d,x�WOT2�}�Z��<Z$�3�*=���Gv-��%{�@9���l�i�k�Ϧ���j(N�&�v�q�@
�VX�A)�܏a�;(O�0҂'ٯ�|.�:ߚ�z/�Z�K���<m���d�p�$������Db�{=�6��(I���)�&k1�={8E��1�VѢ�m4��'�^�J"d���v�E��W۱R*ǜ'�Q���&���䘓���u�c�4O���n���@V��ϔx�`v���/�^<J���l֢<�\�a��z��Kg�5¨�!��Gc��C����"��*�YV��d&jq���[��n1u%��ƃ�exp�o�.�K�3���zxq>�ʸno�8"|��k�
Cl%��g�ES���
U�I�o�tb�
G��@'qA(��W����P���ݕ8"�{b��7k}��(�hNq��]:�
�x�I5��}��@9\E+Z�"��꥟�N�{���E�V���=�_U�`ǔ��H1o�n�D�����f����p��f�-�>�䥺���Qg$�:m��p���m��\U�(�go7��Qۚ�@1��]�A��k|zP��w��%
nw��4�^Fb3�1�pcpVw)��#��r���x=�.n����Q�m�Ys��2����N@�iݶ�T�� �%<�e|O�%�����cV�&��`��ГlV���}����%\ �*����Ȃ{D�Nv|�b;�߃�L9�V���7C|����S�-\_ 6����ܨ}p��;~pU5��_�?�b���I���ԑv����{Cߨ��T�ldh8ئ^���B"��Hu�6�z����ԍeW��7�F�HN�"̝G�x��W%��@��zi�֫^2Ƶ���k�V=[�a9�;GH0ԡ�#�[�3�/����쑺��NQ��$������9����ޢRB1��(i��)��dR�KIsJz��[�h+4Swd��*�o�+M��X~�<��2��\>b_�pc�_	p=	s&�VT�1�6�����p=�˕���Su3,)X�2X?,bZқ��Y�Y�0�5�*��1�h�'
�V
�J#�i�0nsa�����M�7܅���gd�.@0A�њ�s�h��j�ۘ�FE.M��[���%���]�����K9�t��]u�p�͆�.�7��zYm��C�V;=�_��&K^�y�PJ��^�tCܱ�XŠx�M[��7Y��<
r1����b�Ң��Y��h62ӗ��n����R�SA ؞���A��о]L8�%m#;��(�
�}�S�ט�����3MP��%!\����g|m ��[�c���#X��
�g��xC�-P���8����n�%�l�X.���L#�Ԏ���ǅ���N��ozzl��P9^���Ie�v}��^�ZN��#Z�ʂ�^��7����W a]q����i5n ��_�����YW.������$M!~�"a~<C��(����h� ��Z����'�'Oh}5�6�/�!h�+�R�-��SS%5a:)�r��r�hGt-�ez+�����H��ٯ���=쇅����$�Xϥ�TYy�euD��|*�-�vb�J��AfoB��2v-�QU�shA9�p�|������H�h<�i�@�%&��-�����w�U&蒌Ho�����+|�W�8���q	�Mp�a�lL �&Y)<��Uew�nSĉm@���{hl_�a�xAK���� �q)#�yǶ�m��Lz�c癶�he6eҰ��uM������z��v�VE2أ w���m�R��t@3�Ҿc���&(�}�@�0�qKf%��9��%cY�T�7U�b�4p�(pG=���9(�2K��8�8�6�-ފ8�ͬ�������4y/��̢-c�E$�ȯ#�z�/ؿ�|'�m]p��^���P�:MR��@L7!�קZ'�%�1u�9d��#��WuDo)�s�����#3}�O�2\E���g%�=�_d9{�2F��+>`+cM��w�4����<�����V4�;�LWG8
VN}E$���ԉ�`�:����?-_�E�豁��t@M�RS�	�N2"������g�9�t� M�:��UT��b���@�A����t<�6
Ƶ���N����A[�ye��̹=��mO���������Dh��,c��Y�D�� �;�n?՗'׫) g0���{?��OJ�Ⓘ,7w�A�fE�tv,��5W��'	R�i�3�U�Xp���b3T���c�巪�G�������M3�� ��T�ӍA��Ea�.f��V&X	�[���")D�϶��Sq�t��x������#8�.�b�^�s\�D���5V�^L�W�F���!5�e}k�s�w��'�oزc����7@��9�B`�=|��AJ13��b�X��	�,&_xyOҁf�w
/�6�@h��3�A=̃����/�_s����W;�2�±�O�ۡ����kN�q���R�^�W��Z2yYO��k�Ǖ9_��پ=�\�9f�fϫU|��I���;[�E�k���#:�����|�9�8?2g}B�h�Vq��P'�-��'�2,��+蓯d��cz���=4Mie4�ɜ��@1kEy
���3��T24@&4���.%Y��;|���e���p�Py3N�(��3J���J��D��w��`�x��c�x�RQ=���XDR�����w�:֖��O$Ӵ��zl�:@�Cw��P���b�
�G�"���:��s������Z~�}��:L)�i�ѭ��n�R�3���%��B-վsC�A>Iz�w?]7�5�P�d@H�/��=�Gݎ'��]�p$$4�$�8xmBaW,'����'�>��[ QĶS8聻`_����`U�����Ah oB5R��7Ⱥ�|³���y�`� ����\�~-x�{����.�ۄ��X���ه	pĬ