��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α��wԊ�6�a�3� G��λ�:~7 !�v sh��~��P�'|#��x�C�[�~���{-چ��!�:���)�#aE�C�;� ���&�'��c�w|�:�)��$��Sއ�Y�K��N�4uFLN��6n���)G�Kh\��V�5�Hro�\��M)r����ԙ�r%�
�߱����5�����W=� p��yo�����!��˂1��)8Dױ*gC*M:3]n���_����ȕ��bJ�j��P*$7����T����ԦR�rBae�ܠe[�G��v]9�DIpq�Q�R��!�m.2�b�*����,\�>�ǂ�pѦ�P��\��q 7F׽k�w��A�X�5�������߾Ч4h3Y�]�P:���I�83���f�ڀT*�������ۏ�$�����y����z%SV���9��1���H��f�Tw���(��z��-G�k��*�=|4"8�$f���{�a��E����D����z�p΅��~�����TF�!�6:= �ab�s�F�@y�t����1XZXs�5�od��.�K�K_(�mb�g:���K�;��g?5G�x�*�tp��]s����of7*����0suQ���"Tz���� {)��/Ѐ�M���:�Ft���6��к�vw�q��N-+B��t=��A&�r���>�s�:<�.tC{ؒUi&9������ɟ�KR���m!��
��{l}x�����E�����qz}��t?���G���q1$�X摒&yU����꫖,�k=
���y�v(6*��1i�s�1�O�1�� �Ƣ~B]�#D�!<8�v'w�2�>q6fBGCǐxU�28���!H3��?��`�YF�beL�U�D��B���,i�g
i0Rl�'�3���z>"kj�0� \8愁H�z�E��R��z��L�Nz]o�O����:+�_25��y�fЋ�_�q�9�FD��WZ�w��"����+[,%"�f܃^K��o��a��4�y�������r��ZC4��J�.���C"����)8Xԉ�~Z3���I�i���f.�\�\�㰕��TJkr9�'i�ly_�ء�����$Ȣy-M�I�5���+a�E������O��C7�/E¶���	S��<�k1���>��/?2>��ǎ�$�B�B{Ls@)�pkBt��՟Et��{HB�HՂ㘁�ؠ����̤x���߂����r�J�e�%�:f�D��vcpj��2�$Ou���}��� } ����k����ֱ�"�/�k�UFM��Y8�j4�e�:���<oQ�����.���dw�}]�AJf�m:��\�mI����X�Y����j|����ձ�a|���ψ��|�F�(Ddr��:A09N9Tn�a"�ZГ�k"��Cn?��ס�;��\1�m���n *��Y��š4�	P��=��}U�I(�ˣ��s�@���՚`J[=@�ܞS�Aܶ$;2/��V���p����3����
_Qo�Bi���2�.��)KyPV �(���l�����C���U9 (r��,�ο�,&�
/�j$ߘ R����6���S�^������~�ǚ� iA���k�2�*�P�P����|��1*��Y�x�D�p��r�,�ƒ췜�'bqV��um�Ѧ�v¦^t���7&�RjR7o��֪��;���P큞.���Cg�B|s�W����n���{�h
8_ہ;�=�Cfh�߈r,�9�'b�=��R-�1EW�y��Α"����M�c�>��$l῜m�=@�_*��Z�	�
����3��9�,��C�^η�M���W8�4a�')	4S\hٺ���B�o9�����H�U�u��쯊+���B��c��^�����(>}�y+q���l�jR�b�l^/wE�O˶l@�O��A��*t�^�>�6l[X~	�98j���ula'v��q��N���Ȅ�%!mt �GY9i 	5��`� �R�b:Rׁ�<��?"�����%4*�,HqKO��ɟ�>��ѵ�#�ȏ��Ǜ��Z@��\9̑U�����H�4�g�o�i�Z
>�W�����y.IO�]{���57�a8�q-G��$�r�O�U���HH��."����V�q�:0;L����

����"�g˂���<6���IX�Ǫr7� ��p�gƹ'�tD5v���%�FCZ�6�`�r;(�}��+!.�y &�y��F;x�hD�Z���{���O���<���w�r^f��z@I��|���sȒ"�����	C]��F6s]�F��qjx����� p�
�3t9h�s��ȂL���Hy�=X� tl�����Y;[��ޕ��f����*!u(
q}lG��~��%��4��t��I��d�Z2�1���}�b�0������F���j]���g\&n;��=�o�L�L!)5�i�#���b�k$�P��;��-�;3�J��3 ޽���ʽ�T��U������UY%��&��"[~�n%���BA�G���Q�509+;�ڽ7�� �5b�*v�x��}ܘ'���.Y�*�G-� �����B�D��@�J���2�s���0I��9�t҃����.P?(a�Ʒ|TX���|���rϖ9C������|�[^�MZ�iy�O�o��6L��	H�e���J�i5�a�US�Q�cZK��O5�m��y#=!����� ���
�����]ŋ���/��܍L��KAҔ�Bc���J�mZrN7L�I�Z�pE�rVQ���b�YV�5���n��m��m�Ѻr�"���������h4�iY� ��B��ܨ�op��
� �
��~�C��v���S�xĸy2}B���=���瀡� �(�r7|2+}WD5"#i^�5�<���F�_�{kg�Gf.xA.mn/r�ؼ���x`�
���$��s�oTB H!b�Lig6���'V(*oۄ���I둇g��[W����֜�W%3��\�^�{��m�eR�_z��R&� ��U vv[Sv
��+��.{��<|Rc1%�2	�'�!J�u
��<���ϊ