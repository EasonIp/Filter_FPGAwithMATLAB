��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ��nͳ�R[�ظ�_����Qq���G�]~��\�^�W.Z��ke��X�?�I\�zA@���Y"���a`MBl��$���X���/~%�cg��OU#,��;o�w�F�~�wy�0�Sa��qC�$�_됲��ݗ� ���D��.����v��C��k���<�$J��3��I
����<[�P�}&ʁ_m3�P{�
A���-X'�H4Eml�}-���i���[�f�c�:Z��� �Bq��Ƴ��v��g�e�ӳD*�~^��v����$�>�,e�0Dt��:�VlY=As�UPR{q�U١��'�5-ᯄ!Z��=�o�h�W����v�y�%x����� G�|ӑ����}�(^��ڊ�(mKa�/>*�����b��e8�U ;�>Q�e�`N!i�ߒ�O�/魭�|�lF�����ӣ��ϲ��Y���8�qA=A����d�����Z�AqFo?=ʨS�F�;��T�$�ڊ��?����3�E^����(��:_���s�}���
�w�i�����|D&5�ȗ'^�&P婄���ď9��
f�р���0~���p���{e�<��M��AG�Q�?���sf�9�����hT}[�ؼ�,<8�`a�������ױcΖ��_�������ּ,�]M�qB��>TWG�A
m�'Xjs'z����e`��=&>��g
y7MC	���� O�� 6AX��E��DG�LK���=��)E�P�KVX��=�Ccұ�VE%��Ⱦ�ɮ:J��`�7���F�<����hk֛}?o��~�N�Za�*؅M� vm��q�aPm�40�$����y�X��K�f"�Ĳ�7q?�K(J8��r���k>�ʿ��>$�zr���u���MD�-
��^����p�d��ͻ�@��r�"_M�u����P@������4�P��BQ��s����|F�c�
�L�r8���)�\��G�n��,�n�.h�LcWZ.Et{���b*6���ư~�0F��"��HU�U��#���Zjx�(��3�SZ�٧�>�A���V�&&_���mt�a06�TN��~��')�LL���Ѫ�N�����t�;�f7<�Ps��F�7��!;��H+�(9I��&���*�{G�>���4�j}>�S�n����H2[�pX����˞{
�0�T�UQjS��Ye��F#�U3��Vb�:>������$�ioPK||�@�7�2ݔ�9����=di�!��l9Nr2�vB���4a|6S'݃�B�:'�F\�{|}Vepa�}x�q�:zJ�Ը�<mQ#��/��.�b_�86I����n��I�_���(���N,cj�I<"�d�B'&7l(��Q�x	�9��0�Q%|s[�[_)d�0Bl��
F^�����qe[�1��P�d�)X�vbUO����C�����.���iC�ԁ;G���?����E"�%�J뻰�$�Vf|B@����[*O0�{w�k#�o�9
�6�����[T�z*���	)��k/+Z�L�Jp��	Ǔ�s�a���\$zvp�j����s/ή;�BN9`^�'���'��^���y�9�"6����dM�T(��Ȯ��DI4�y2	�_S��I�eia�E���H�y
�:��-mE4��E���Y��$jP���#p�#-�y[M� u`����y��	�u���~�ȊЁZ����zX!�IZ-�8G�R����^�u3��sU0ch�wE
���k��@�4fk�/��O v!L��G0��n�Q8eͥ`~�,vmTF�S���&���G��,��A����@�o�2_ք���]�-!���" @���.�9� ��~l���NG*G׷�@��p�'��h�|鰃D��D�C��
�&b0�{���Q�Y(	@��Ui� c�jp���W$6�'�0kl*&f,U����I�L��R-; G��Zm*z'a���sUe ��r.D��K�y�oE���]�v ��e��7� {�4ue�{1ʗi�~����$i�p�8h��u�"��hR�vY@��ڈ�����'��+�M��MߥH���0Ǌ �8Kʆ���)d�9/-��>�=�S-U��%Ƣn�-���I5rUA��*��'�<�q��-w��[@��S�Z���qi�ZPܔ6?�/���u���>��QR��.��3-��%><o���(������2��Ư@��]�t2� EH���g8@g��ʡ��o��^>R�QG����
*2d��C�]���SR�(l��r�q�5y�-��O���a��
	5~�CT26 R����� Q��]��I �n�G�sl������ˣZ"@bH�m��2���v?��W�
<�֡D#y����k�8m��[�FFGh;Q��i�_�J�l�mǵ_��s��\�:Ōl��b�Y�ԩ�P�}@!|qv3Z��lS�u�m��x깫���w���i3��Pۀ]�)��ь��j�V�8����v��3G@\��D<����H1y��qE�܎�JQM�I��N��.���ܙ^}+{N�sdp���&-��yZ�V�Z��C�U��q+Ü߄�|��r����ߙ��V)@�� ���{���(@�L�rޱ(�� `�.c�6��9	����J�C	��F7m�g�#*��_��E�W=���x���0?��m��ߤ�}Y=���fY��EJ�:G�t���Db�!<���H�Ai!��Ħ$�+?�^�e�A-�dN�mx1tH�,o@W�	��_��D�<�@�	��Ikd�)�J��(t�����F!]*>{�	��T�֘PGC��k���4����J�t��_��b���'X�p�����PA��ӖSpo.��m��\�`�N�eR=	��C���S�q��t���ޡ2E�	DfٟE�VO}��q���VZ��j}C���j]� 0/l�f�]�� 	Oӕ����!_7�=�mu~� k��$8e�MT�]��s!���@�= �!�辡�Pσ�e�Vm.+�V��$�IO�D��A@ᘾ%!+V�����v��9�f���׸�<M\M���`�G��d����Q���ڽC��_:٠��M�҅a\�;�����y�ey2BHQ1�v�:���C1�j�0���
 �и
}�`�4�|��ʈ���vRH;ۉr�z���:��^�ޞ�=�N��#^O�(��b�N� ��.>��(�
�M!ɜi�o��89ndӐLQ�h�#���+d��8�?�(�\�?h����F�T��>>��;� �8��$�r���}W(����J~A���_Ͽ�<8���BX:�
i�:O��Gs%��_[��@H*|���S�l�v�����E *���f�	 zb��J�tÊ|��VK��MT>��黚R�g��7W�"�I���;�Ri�t��^��M��X(�6A"N-Y�&�C�Z��\?�%*r�zD�6�/v������UK�\�΃|)�a�]ŧ�h�.��Zͺ��VԷ^2���P���֧�.-<��0DO��|-��j=r��F��,�9�5�lN/�c�I�7�$�ܜ'��o�.�(I�� ��`�l����1�y�y�8�o8[��ًw�����釙��Ͱ� �
�d��s�>E�J�t�K�G���l
 |��.4�
�8w;��tG��.@�K�(I�����rDMV�#�S/Z<�;W �����tgt����Y�ܤ���'�gz
`�&�cq�7��t@.o��3�J�]Ű���(Í'� �i)���<�~��qEg�1uQ��8 I�|;��)&>}wWi���ތ�Lq��l��V�8*��Q+yO��>����Y���a&�x�
��I����"%��(�������g5�@
�ᮻ��
�4��7�GyN��	� ?��to:�ͺ�B��_J,��t�]��M��Z_��l9�y�y�v��X���6�$3z�TvF�N�'�Tk���n����Z�~;7��4��G�ZOU2!v�;	l�{������g�ͬ't0�AC�6�U��kW�Qr���0MY����9�+J�᜗�k����	u�r�/��K���e'/��H�Aq:o��<g*����v`��;sR<un�џFg�C�:��ӭK��k6�$c����k���0�`8�1���Pѧ��wlF�zQ�8��Q��1k2*��8��sC��{�P�zА��Iyo��6�k-V�tB6�Fy� \�)