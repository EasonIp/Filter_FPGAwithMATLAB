��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4d��oc���_LG����*k����۾�T>x�/>:��e�=�C5!)f���86�$����ԤE���oZ�&�x���� ]1����V'���Hci������I���-�;����{�gr�HR�l�q����~�n�2�����̴S�c�6�'o����f�?L�2���r�����uq/�Z��a['R�)9"+",��:�l/
����#���U\3�$π��`3��J�,�;K��=.�ʄ1���c��ą�&Y+[&��z{��/j��?|��~:�%��?�!M1�3?ߤ�	d���j"VlVg8��j&84)�|K�\�Y��m���TU-�^V <h�Τ�4XU�/6�����X�_A����W!��i��o��>��B��.��9C��iżׇ�2�%>+o��q�(t�
�%�\����·�*,U��y�oxmX S�`���;�F�S7�
�(���!�e�5�I��Ey·���e�`
&NTv��n�������Րae�m�d�9�<]����kw/��׼3`����ǧ=��ό����d%;�4�����"?E����R�m%���<�:F�Z�䕼jp�j7���P�U����AX�����:;��}1I>�[Z�洽��J�(T��(A���ik�sO����al�	�y�7�Ady�3� Ck�ѐ�9���#O�XM��@ŏ��X@���6�-i�� �*D�ӆZ-sa)K�7�
�3�`8�"\��u������Axw|*�>�y�Z��eDJ��rs�?���P�ι��Q \�f�Q)hQ�&��c�'��n.l�.'I�X	�D)!���s_��@U[%�Q�A���"��L��֢��۾����KJϽ�U ��T�/�f�MYA�����������=��D����e��|E��T��_%�����̸;�[�T�J������i���~��9׾$T�r�j?źR�o��*��C.�������uׇ<V�6�ĳ��Č�z<\�^?�����h�%X7�mp�Y^}Oa�V���_�L��������|fMX���M�T�B>�W�~l�}zvLW��8XQ?���|/�U�<3J3�����  J��m���%N	,�>v"$����d��p��s�/������&1���v���+�~h�q�&�_�HPϜ���r��!���PJ03"���q;�QP����3C�|�Y���H��^�>� T�jYU50�ME[��t���QDt���Fg�" �I_�#!P�� ���7���[��chV\���/�I�bS�H��A�^��.r=s���3��	���5���1�5�ͼ�۷x���*X�E��N%���a���(�%��瀶�E�29�~h!|HHz����
�z�1m����\���l�x�K	�f�X§,�}����ӳ���,�h,��w���_�П2��C�ҍ�ow�E�;9�)0/�E���������+�h�Nc����5JUo^d����e��fF:���y�,[�݋b�>90��O�f\Y�"�s�q�����!�4�b�	�0�g̈́&�~4X��f�l�<�uao*��K$镪#/|\�6?�j��졆�����]�o����6P��_�Р@�Ow�X�DlT"n�!��WL;�r��}$�}V�������艦s~暸�6�3
D��;E�K��כ�C8]yXV\5(V�~/�>�B��3<6�Ӗ�X�\��Ay��ֹ6�hXR1��{��
����
�>�ĩ�l�!N���yɾ��!"�ĩ�F�F�����v�f��̓)�A�P�Uǖ]]�C���`B��jx2�a/R��|;�Lr+ʋ
���G9vt�ц)2�v'��.���4Գ�ev�D0n�Z�]-�`�@����:}s�h³!���S&��6����_���Р6-��>n\~�8�Ɂ¸�V�z��W�.���)ȗ�cIE%G�S�{)���~-��,9�U��:.+0��s�����o|�W��ah��I]=-9ȡR|�(IL�?(~��-�卿��s��c���:�gW�fW���J��kH]�c���A�/��HF��r941V?D\Sr�5u0j�m��[��z �NI�TPw��_R,���n;>6�`�e 5��Qz�$���{�����S4�l�������^�Q�z���O��U���o���G�9Of��2$wh���.6�ʟ���TV��~��?�z?���S�%G��7���9�zOsg3�4�Qr�X��'D�	z��9���ҋ�Q��%��X����q=�>�f^�����OM���`�d���|�4Y���X}������z
� +yB
��Q]�� !�A��H~����Ca}lu
ߊ>x/5�l{)��i`���D:DR�K�C��*�&1�e+�8�^��=@���t�i�A��e�EGg;n�^}£h��~��Ы��=nsk&��%��|f-(=C�pf�v_#FSO�C��������Cu��f����|R���$Ҡ|�<uGO�D�Q}EJ$��}�UX�"u�����{��W^�6����C;��u�����'$��[��K7Q&{`e�|�%8���A묤�\3Gj�!��]��7����#g:�}�`��v����~�����\�m�±x��Ӯ��x�����t����k�y�בo �J�gV��S*1�۲i��I�Z�O<)�g����Bq����A�v�ךz�hS��gB
c����p��Ɓ}����re�Xz
���NkǨ]����a-��m�?Pl�E�Z���'^��D#��јְ沃�D�w�$mq��dy���o��ƒ�V�)�S۝A�Ly#����:�p�p,���[ɷ�f�`��sP��ʿ:��>ĂV��[Q�w]$J&�JE������)�*!i�So��#��~j𝨑^$m�$R�r�����YB2��V�"�k��.X&n>����="i�nn)N���p&ڙ(/�R	�7�7�o������D��'V��6�e���k���GO��}qW�k��}6��5��
D"� ��u�j+̭߽o灖��:e@�g�������p�w ���~ǰ��������e��-֜�q�؉�b�0m{�y��H�
�%���p�#�Hc2��l̠�)S�_��l܃Q��tu$�^f�[�#BN��W��T��,�������|�21��7�Z��j����Eo"�}�A4e#����
��%�b��%'F���+j���E��?}B���PnN��GW3���k��C��jN����x*�AR!�I��%�k��z�e���_f�B��|\bJ�� �h�#��=�t��%�P �*t!����{�q�ސ���{��k��
��c���z,57��%��U~�"���V�1�JJ8qg���G"r8>![��w�x�A@�6t�� �"�{�$`t�1��Wޝ$��m~�,,�̅;<�	�wC�e�IL*�=8xW�Z��,cw��ˆ~�SA�,3�%	���,�������3���qN	y��`�<'��ݚDuv6�WϋV�pZ�����Ӭ=	�����W�%|��kz�0�<��MS��߶�:84R�A�;�į�[�S����^J����ȳą�m��u�����m����/��8�B<�U�[����+���k�`_��8kcF�����ޒ��,8�p�T8ݎ�֖��p�BW��VsE;��S=���@�c��	�]OF$4�C���5h�W�x.����R4��HJY�����Ԫ�6�����e�Xn�(i��}�Z��-��d
s��Ɍ��u��9DA$Z��?���T�*��w|@h�����ڠળ��`x���p���]�![�`�0�NŚ�� �GM���������]s�Eˑq���,]��Gz�
q'��}�Q�qg_�z��f�j~c�J-�1�%P�}� Ơ�~�K�3n��,��*�N��O%I(~��%}w!�U�U���|�IO�a�1Qt�#�D^�����-�ϠJ�1z��Xy�9����D���2��S�n��R��[�_�Kewg >@�Wwy'᠙�~0|q�*��M3�'�V���(��2�F�of��v3=��cj��eA.�a� �a��ݐ�QFǝ�d%��2 LZ>\���μ�2��\Mm�L�x��;���l/�T���!�4#|u?�~�'�{�\���?7��2���܁qfy0�0��M��c���M�z������su��z��V��S)��t�T>&��P�DM����XT����+���?R�L�r+�6�Bvw(�,�ľ,m.1��؝C�y-����Pٲ���C���tk[~���d���ɳ��["�\�j�=i <�"j�ξo�C��j�}�B�=Vg?�T��P�[ϩ>�P����uP�:�{8�=��ʈ��u�a��s3��A�n`�cc�qJO���h��gۢf�g�o7�N�\&��A����WB*�C�ܰ7�ޙ ����k�Sn�ZbV�&����
]�6WҌ��i���17�D��D�*��F�y�T��$�4s�ĈϤ���ԃ�@MO���<Y�,R����;R�X�A��gw��"�yHl��g����I?½6��B7�������5#�䫜���QǤ_J^�oD�p�6�t����S3!l}��d��NfE�Qh&k�2[`;3TaL�%lI������AZ%�%��֯<�_�-4ԴZ������M�Y��� �����:m�)v�pI,6���' pVV���C�	�|�rX���T�AX���GFƨe�e%'/�@�R4���*�޲O��m?���b
2�})�DT�{`D,��2�栩ZK<��-�\�Cݚm����
zzY��ܴ�ޥ����J���HH_#Bq�a����-�Vz��)a	��>��~�F7���ΐi/����Q����Z��^���K�����=��������ȍ�I��n	g����6EZ����FAjes=�<M��O��f���xº5^\D��}S�d;�	�(�~�b�~�g+zHO��X������Ұ6D	��"�ĥ�2�`��2�p�\T
�LpuR�4<#�ٟ���F�Q^�Fd0�����Uz>wi��N�o;��+u�]t?�\�w�~�gv�B�@�fC�E�����Y|�R�=-��K[��Q%vp�@eH�P嘵�V&��Ѐ��X.�c(�ߔ��e2\Ӡo���	w��	���!K!伱��qhJ0�y�ɜ�:(��k���e�����V��Q�E2�i�DrOǤ���D���1���/��ެ��y�>��P ~����w?x�I�ܖ��
w�إ��q�}��q����Ƭ���W?M�<�L(�V�d�D��D��y�:����=LĬ��5�����3�/=��z ץԨ	�WX�&}��9�������;�{{D�a�[�Kyq�[Kt��̞r�mm݉�sA����ò�0�FF�G>u�ѕ�\,#0�o7K<v�+��B�HRc�y	x���ZA��"��)���LB�uw�]%�8s��+z8?����^̙xo�"�r�a��z#0a|�p���X����=-���!�:7 7<���O��C�ET��\�� �:��G�^ܩ�#���%n��v埓�J� �h=�#�>5&jQ�j|�����"0�r�wV ��GC�ѓ��0�F������B�t���HΖ�?)��!���6�i]������8 ~�l�i��0�?rHih��$�),ҮMj���q�q�P�S���n�Z�掌��Y�suu@�,,ţ�0�1�(�>�W"M"V'U}��)Ճ�ż���ÂË���u��� ;B�3���B�L���<s��:8�7�й�8 �Q�P�{C�pO��+���D�X��OR