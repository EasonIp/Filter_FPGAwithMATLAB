��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M��*����g#φ'����T��6%.^f��8{�^v�wK�T��fAN(.�oC�Yt���Ao�>���� �h�*��9礩[s�Tj˧��Y���oG� �'!�D!�#S��E3@b����}��doB۳��P����F�.r�Z8Bg��������K~�g\�l1�i����r`0���Sw����X՛m�ɒ��Fq{�GT���܉Ub��o#���;��V���
��ħ�u#ĳY���Ei�Տ�#4�P!���	j�c0G�'�(t�g�5g�O�U���H�x�{ؽ%�qT�ˡ���٫^�)�׶�rn�.c����Z] p�ֆ����s��b'��qw�3�Շ�O��)b;6��!dg~ȁ������U��mD����a}>���<&��HA󧩩Ͽ�[�Jϲ���4B�JޟǴ�J�$��$�*? �$O�fhq�Eds�ӥ�r�-�b4���y�Y�hG����Pqȫ����" f�$��p�:ЬT	��c(����qo�?V�"v9��	e���+b�H���g�MGaNJ�|��!b�Ggȴ�Okg�y�K�2�lS����Dȓ"��
�s�TN���Y ���ZxM���?Z7R�\��������޾�	�d;�J����gc9�	�E�}tg��Az� �	?1�k<ID|(�Ce|N�y�VՇN�FY�_�G�X��$��!3� D�����g����9�m���t���H.4�s=e?C�ᜊ�Ct��v����m	>75oP�nu�8��W�;�۠�V��8ho�ZZ4���*��8B��R@/��}7�E��R�5�bb����E�K��7���W���6�e&w�ȹBPk��B�cNyǆk_�t>�w��8:5�|�՝�a1b�N>o@f�����!�fD�o���Ztնe�p���e�AD�62�����g���t���|��cM�锘�[��8�i�-^�j��x}=��)[e"U�%$�G���d���&�#�wx��	���y[�$W{�?4�MO���#��WD� 跔�v�w��W7Ca/���������\8�[��AI*��1�b���!�H�t��9�4�8���^"bXh�p�͎��dw>�ބQ�O��ۉ]B�/(�fI�1��R$h�����P}�}�r�>R^�9�Tr��M;�	ٔ��Q2���V|����I+)�Ce�߇�as�m��;�l�Xv6A�#�b� ��
Fp@�Q~��dU������*T� �[��rx��Xv��مF"�v_���Ё��E�����[���W���82T��^
�<}�u���%��*\���f��t�r7����W^����;��9+�υA{v��E�|�{|A)0�U�������䝛�=˒u:�(��co���(h\��|[�ý�!�ƢX��I��{�>���p��(�=�f*�o�y@jzS�&-���*z�_aX��,x:�-�HRH���3z��{7qx�nǀQ�|�竣#S���io�@N��� [�]�Q���G�F��	�
~E�]��s�,��z�����<Č��,�"�T��1�`N��!�|e�`i?��V$�mX����'u�������m_?خ�v&�v���T����D�e��=f�?\n����QO,�#3s�rټ�3wU`E;���<����u�]'����;b��3�P1Vq2Uۡ��8vd��IԪ�;���S>Ref�>
������Px]է�T��}��WjF|��XDj����*�]�yC'���6Y#��Ҙ�-����;^p�ހ#�z��2�ʭ�t�$�;�Ż�Cԍ�P��B:���8�GhЈ��l�k%������oãk�I�1uFl�ZZ�f��Sc-K�Φ���;�� ���iqLU���!��
�w�r�T��
P���͔l����aO�),����e>�$���IA�&��U�b\f��Ċ����]4RO��'m�a?�j���Z>�傤�����t��G�<j ��p<MM�����;�_m�D�2�����sg?�d#���R�{�a$�E~x��[W?d>�����џ�{m	w��g��P}zq�4d��^�D�T~�S8"���|#,m��]8J��w�uiEK�:�ft�?�{��@.�wC�MC���m���O��du��F��A� �޽$E(�������9���F�Ǣ�d���������
�V��ڇ�DR'�kd`cc�V�ExR�Bf����y{�J^�/�rm���;�\]p�Z*!�k��:�G�T�^%�t�q����݇�Tr?�k�ء�}�U���e��ODχ�2���a ��)���u+�=�P�[d����k��ECO��^<���|%k�K�����&���x\�np=_s�mϧ �p��A{�-�,�Kc�3 c�+dK.�sWb]��ҹ����`��2���zO��}�ƕ~lT͠����ymj\��dY�dE���E%W�\�0�/��K�B��K���i���R
� �(�J�5{!�*K0�� ��noĄ���N���b{��%�b���K�sıt���qE[�H�_:��V��4x෴N�(p�A-��T!sB-��ؼ~%�A���9|������K�i�N�5J��r8�  �Cn$�!m3�]�zV7���OC _��ۋi�S�w�ņ� Q����'�O�|C9E�ܹ۟y��¶�ݽ�ڭ��l�a�븽w�\oN��iUo��3b��t���` F�>]�T��Hѻ�Y%� *��|fj�}~�!������jFu���!([7�i���!�{1�9�䃝��S^=�����yÞ�ߴ��g<�u؋Ζף���\�բ��L��"w�?��A�{)��j6����{���}�dܘU�w1?�K�x�{��[�v5��*�B{�h���h��NGN��Ȗ�ʳ@n۶�0�u!����7"n��3�+���=�{�5�!?���b�q(����Pc)N�m�<:�3���Wn��n���i�sF�~��RH�ru��>���U��b������z�w�:�aOS__�3N�7g�M���I;��:H��3 x�椦Uy�����]�U�f��6�dVz����)sR�к�^�@"p�����}�("�LBD�<�~���qr�$OQ$���/��[7圆}GϞU*}�i��Z��pxx.R��W˩��.-[��ﶗ�����5�Aۍ���V�7����ܞ�S\Z-O��*gȬ�Q�V�ȶ��Y�	ǫ�X�a�Y��Ӿ#ca�E]�J��$���D��	�;�G.`j3�*���JՄ���حj�VYgfZ8�1f�?��^��R�qt�g�Q��K� :��] W��?�a�4���~����J ,�"�iRS� ���E\��)��'�9)��5�9_�nH�r#��$���,M�)�ԭ�^t>��{q��%qn:q�T�Z=Kȿ�W��a���j��j�}ʢ|?�s#֑��Q�?�=��]7r�<��j�S��d�~���f���'_TL�斜����h��:�*y��Y�#��0Zq�~ҏ����1I �1"�^�d� <��:����G��'�i�d8�MpK�LB�WOƊ���ߺ�Rɕ�@���I���䣫i��[���,�@���6�C�7)�+�xj�׋���g���Y�q�.@�Z`�X���\����~�6�������8U�NGrR׀�f�4���|qD�LԖ���~��A�.~���E�(�?*!$���'��7�6j*�#W�C�L�����8����F�X&��X3�tgK{v�lD�O�L����Nj9ފ����[j�R�b�4��y�e��>�gq�~���@��h ��~3�?\�ȴ�]\V�Ό&o <� �"���cF	
m2��Q0�ɜ�@�
v_�F~��)ͻz$x��$PL�h��&��U�/�w���̃UZ�fKU��*�����f�[�N�!n;/����s�-���X���8t�Zf�Bѣ�B;a�^�����AO�J_ٗk�V��Q���}��`oPnHa�0����� �T�+����"�x�����~Z����9�F'.��w���(^Fpe��0����u��冘Dg�hvf�P�C.�3u���}��x�8s���&�����N�w7����+%DX]DRߍ��%�J���#�[�����u��c�,5Fⓔt՚���!�����3<㌚����6'�0`	��j$�j��v�W��ޖ8C��\��%�J+�z�'t�ɖm�HT�8����'�J�o��6�΀@��O�&��/���rD�&~�����1�8��E�p?��aU7�$�i��@��.��u��}31�k���>��ܒ_{/򖐽`&,�Idc�؏��\�mހT6`�����$,�R��$�JDuPPZ+��!�.S_[����<�o`W�(�ػjg����Q;@�I�˔�@,�~�p�ֻ�ӱ���Ս���'Kb���~?�<��6��ޫ�Z��!(��]A�J� ��x��9TfPL�|C�8��f4g�RD`_���A��5�#�rʭ�#9c�4�����󩰞��˾��ĔFE�N^�뺌}`>OE1�>��Tt$�WqRG|����Q����q�?T��r�y��˸������  ��r�+Zk����À�-uw��t��oq*��s��ӊ�/��L�Ӭpu?�V����sa�>{S�f*��%�Է�*�\8�5����R�)��yX"��~�^�ڙ�nvsM��9����(���g���	d��{���*xΥ\/��O�[�=ڎM���;�w�^�="Q�U�=(�(��*A�x6�D��	��x�k�~��,Z"��<�e��d� �A�S=�`�Z_J#\u~�V���y��SN�Ч��]p�;,���Eٮ�`���T<�ȍI��t��TD���O�y��(M5�r��-k�~0/n�#^����mr=��m���lYF�+�4�*a	5��\���?�o��v�|kC�5�2����wR<��0J"��V�9�P���4�����c_����[�0rt�sBA|�½{�ؘ�aov�k{�N~�>�f��b{l���M��X�s|��G�I�m�wf]h= ��4��Rӫ�/�%��au�p'��9K�����N�HZ#Ȋ�X����+��]�q'��ɽ拿�^tL�	H��*�G��z��5�J���J�O��������Ikz>��@؆ջ�TY4��T>�� n���]�зsX����vJ�Bn^�6HA�-@G'�����t���Z�F�;?_7�x$Eо��Z
���S�_��=�n������h?�����LyfP'~�ip���=���e.4���I�l���;��C��l�:q��ɘ>����1�/uQ�LP>�j�M�pg�����ba3������i�5b�	�8���
��EY��Ÿ$s~�G�������۵��a׳�ZM~}A�ɣ<��#��,�!��r�)�0$(�Tүي�e��,����$�s���~��m��W��;-�#��}�*%%�X8n��f��(��RM#?f��_
��4o�&�8(b4Ĕ!T�᳊�9�Asǩ���'�u_��t���C�˒�aG�֭�)F��藨�&�߆��0q�RK�>���x��5��b��}��W"���Q��"L]�,����̩ �'�u���K���t��[Rw>4�}6� "l&�g'��Nuy��o�Y"3��\�\\�e6���xP�4ϑ��ED���O$�p��C&�U�{�ԉ�dvGjBb'w7�OMC;�G6��j�9B�EHX(n��5ji;��53�)�p�4��q�&��x8��A0��{�u�L�6-E��0�^�����UP��h��A� �c���]�=�����ͥ�G��6b��͚ݯ�|���W�-�L�P	1��,S�Y^r:q�����92���h���ݍȋt� �<��9rX_��Q��wl_���	��|�W_���sh�X_���z^�|�#�o��33Q�v�+�2�ն-�3"���KX��CV*s#�����,c%?�����z��^p�2�!�V%5�*���I@�x5��?*7������m��U�^��E�	%(�}�\�u�9�����S�t$J�_"�4��,ݣ��YA��~�N��gH�A���ة��@9��
F!4"�v�3��Z+҅����.I7ű��x1���\~Q�h?���L*��S�47T�Yg73$��Í`78fp%���x�0Z��o��X����3�,���T��t���m^���;*�DU���ԉ�< 5ґ���U�ݛD���h����k�����F �C��u����^���{�h�<��"@�OJ}�~`6;��5��6t�I^Z�[�DK�i�'��LI��ư�u �2ؚ�!w��SlL-m_�
]BlN}_�/x���_��I��u�o&q�폰ho��K0N�L5�,;��#@���)��Ys��2��!�$��Ǫ��ﬤ�2�*+��3h�f�K�扒b�$e�cƂ^���ɣ	���(��12~:c���Nf�ޠ"e�{�������#�E���[�9�����yRb���_dh�¼5r�+��ɋ��o�`7N��!����ի��R��#� �HO����t�EE��F��^oM%�K� ���nsΑ���b��a�!���~�e9���.̬�}o�v��?%J�p�7n�C����k'�������LI/�~�R��nzN)�p
���l"�O�p�MJ���������A�;f�v���[�0�;.�p�[��e�x���s8YgQa��Y*�w�VF�sD������+�l��>���`(�v�n�Q:����P uv�~D�k��I�a�Pc4t d^:7k'��Tw��R��l�ćgN���(��2�����2DsH��v�dӡ��v9:��8�AS�=T� ��q��u'B�ʮ��с/<�r���"=l��%&\з�5B)+.7M	�s�k��E���lMd�m�r�."�Yo����2���
��nD�l�h���{sq���_�2ٜ�ZY�~^��{�������R���O��̗��8�9{����yH���K�դ����ke�͙���q��W/-](S�\��N�;�������Y�2!»�)������"N��s���:HO���A����P�4)��e��$v���:W0d̹�Iuq`�ZDs�JhH8��i]�������":�)����6�d��CS�.�}(�P* �'V��KJ��T7���Zu�wNž�;*�yt�x�j� �f��cM�;��Z�XtF�X�H>�8��2��:S�2t�ao$�>E�^�L�݋�I%'q}ל!O9+:?%���ؖE��ɍ:q㦍�y��4�l�K�6Q(�G=KEIKZj��RΤ��z���jU�y�I��M�6��-Y�Բ��ҿ�c��i��w��E-�ِ	��C.������t�M1^�gV��e�z���;���<�	��t$�k�K�g+p��"��׊h�!6�Vm꠪�C��)(��B��?��C�~�]ӆ��vv(`٣�!D�2B��N%��ŧЉ�/;�~Y�bqߧ���\2(�%ņ�����g��?�u��Тp8�|��]��m��S��/J�Յlrĳ�m���̈�qe �	�B%s����Y�b(�܁懴Tܠ�P�P;��Ϫ:v ���2�M"���$�c�$��>W�T��I�GVRn��ţ1=qSGe��\�eF���
Tq=Z��e���[/�P��8�Xщ�������$A�oW8��ϣ�y-��䦠��.�E�@�F�-êU,D~|�}�~�Z��������!�&���3Y��R^���J��z���B�ZK6T��ĭ��v�I�kj6�+�Ƙ*-��
�a!����e���w�Ю�p�^%ɲ�[4Ŏ��T�sah�q�߃�8/��͛�v����u���n�J���v���S�02��\�־+`���]���k�r��|�Dm=��Y�O
j�	��H:`j��1h&u�F���n+#�ס�������MB	�2���.��ԫ��fO�`��*���k��Bx
z��&�.��6��5��������v>L��@v݁#�̐ٰ��b��{sZ<�� �'��㷾�t1�V��,�O��?��{���<���_³:�9*v����h�e�%7`,�ѕu�&�G��S��r������
��_�A�6ئ�|��*ǂq~ʭ%����b+2X��!��d���#^W���Wx"�8U_�T�/},&�����	���{�ע�%-�um �����Q\�U��مoV��q_/�!Z���%'�X�����ɇ*X��_�[L]D=���J�76¬�>[x��é	^S���{d�� ��`�Mg����$)Bp��������w�����:�Y����h�>��{���s����(M���e �xR�0ʅl� 3I���sĬ�'[�B�~F�J��glvp�_�4��\=	�SW�/\9�Si�x�� HeԷ�l�y]�2-Ƭ|j��K�(AA�Bn����;�<
�,�M�dy@��F��#�Nn�nϟQ��)��9���;�iGY@��M97��(>@G3ާ`,��S�;Jە��2��uy��ʁU�R�~�x:�?X�1$bFo�;Ե�ϙ���iPFY\Q�7H#�j�S,b!_Ǵ�|���=� j��0�?9TtPvه_(�S/ɘ���!��8�^�i�l'm�l��:J��f��c�nx�]�Q=�@u��N�f��ޅJ(�v&Xtl����v`��^���\�j��_2H] ������lx����}֪1���gG��#^;^-ĭ	�NX+�G$.��Ǘ𥿯�?p�r�#L(N�.%A�G��&$A-���w04Z#�Z#�+N	"���{No���9A �[V�PB�e�Y���4�&BqCM����9�.�V�L5�(g�T�n��bw�X��B�Q��i���뼠ָ2�z�������q�H���RGF���c_m��eΊ�;�yD���`�Qf�"�.(r&P��v!.t�_�%�+\���U�l�7/����0��$v>7&�;xvJ���X�������`�Zz��q34M�F���=r�r� D�����K�ck���|#J��ʤ�E���ϱ�wxC���48��D�͗\U�g��	)=$��(�j�d�,_��J9f�S"���TVR>�OO�w�M������"�wãm�lː����Whyg�!�E��<�9k����"��6�\�,��x�j�7G�6a����';_u"�F�OH���\��9�̚p����ԝRځ��X��xu�̴�x�4x<8J�#-�rK��P{_L�M�o�Ş����B�o;��NhO�\�_1�h�!@�Җp:��bhE�����@�S��]37u���bR�􉴹T�	��{'���$&��f:�<O����Ê 1��c���D�p�3$�'pu��T�ۑ�/i�W�9��g���3:^��F�6�w���!���_p &��V��[�q^�-k��}]F%�!Vm��:�w��/M�[�Ak�R�K)�K�7�ʣED����+yaju�F�m�sRz����j��[@�NۻDH-0�fj��/�L���w�.Z;*L˓�wt�mS������P�L�Z��t'�%a�{0�ڣ���V鸼'���uN�'�T�#���� (C�O�t9�N��<����%��Yf5�r;�u���-�X��z{�8�qc�oE ��x��2-<��!�	��S��2�	��ّ���pӒ�iC�N>B0�3U���I+�=s� L��a.��%ꮘNɏ_�)`�l�u����4��l��g���ܣ'�OQZ�[)��Y����q!��F5�˷{���1eb�~�G��0�2�X��<(`���	�S�	�����A�ƬQ;��+{��:�Z�9���{FMP��P�����)�N]�����pq>��u�DU�V5y֒g������7w�F�$��{������'�K� ܆�c�b`�v"�3,{��������9�j��$s��x��O^�j�����m�p�F��F��Q�ˤZ� %����I�C�#m^S�r�žS���rQ�-���+�4��K!�dz�H�٠hR/RUieE���%�f82��_����Z�A�nE�,�	���V@�]�u�l�u�����D/K
|[� L��]�[|�V{�����/GE���Q�V�ϑ��g��#�T=�$K)]�
�����_�J�A�����b��ȷ ����Q�J.S��0&�gM��,���E���P�~�	�QA`���r AY9nԴ�PQ��${h�"�j96�E��QsjE0`*�3��̿I��A�#�KWp���Y3��}�/Ã�;�C�Q��x�Vy�,])L���ѓ��9d���b����Yr��&�!B[]�TWb`��M�E������GE�ER�b����X��;�s�W���rE�� ��B$T#U���'J+���
�Ȃ&,��Z=������<�4�̯G��L���/5LP�FZt���6��L��pE��~*6ng��yGug>Js8)%"�骲�͆���ᜯ�F��H�{)�$3��"[m�sY܅꯸��U�WV����m\�(f�F�!�����ױ;�ZR=�۲��IS!8�t�*��n�ƭn�N[�K�wW��A�f,��(gK3VpD�:�!G�.�s��6Y
r��ƶR�{��[��	01�.�\
����Q3[jsqu���"Վ^��R@�T/�����	��`�υz~���طpE��}ڸޥ���GJw���ܱ="?�mSu�QW�sŭ���\��.�m��Z�W�v^�A_^�Ϡ��2�f�H�S	ȍn������ܹ��� ��)�5�?�L����D3��?�1����_I�j�A`ʪ��AMx������`���̭{�K�%�0�Aձ�؟F|ٌ�{U�ۖ���5TM�6�_���o3��t�*Pb��=�H�N� � O��7�Q��刻X
�����IY>�$2=����(��m�'�y`=�$�ZTf~
_��\�O��b�	�ER]�J�c`�8��:�sW�B?U/�O�7-ڶ��!k��W9� Q��D�<m��Ilɋ��u�1ޫ�W�u��S<W1)��Ȣ��#O��۳B�d�P�ΖEt��a-e�k@
�EM8Ӟ��w:�}���xD]#�ޫ?�8��ǠZd�V�QPT��Đ���Y#η�0�1O]=�/��S	�(���VO~�6���&��4M[6X�2L�ҖB+��}�M�o`��hA�������5�����m�7{��eu��ۄuq�L�t�b[{�\�6���u!�32��$@)U��7=����Ts*Om��`���>�8> �����
_*gQfr͔���V���or�nP�V_�6�}������A�/7!�`�I���0MZ�v=J��ͼI״9ԘS�~N�Қ�''�����}e��O�ŀ/˛	��&=�Q@c��Ķ)��Z�CW
ܓ�H��i����ϓȟ`r���1 x�q��z_�rxL~Z��1�r�\X���r{�/�!Zn��Ђ����n)�y&2E3wDq��~�"*B�U� ^���$�>�M"�>����z�8��eЦ.]��l��A��l��[��*��^jWX��E6�^��%�4����i�F�M����2�#J�xe~����dN�E�˄+BR����/�7)�c�2��	?����O�J��=)��lRH#��x�x}�u�˭�$�JNϐ
�m�g����J��{ڛq�
�)X���Sl��r�&7�K��=!
M�_5?ҩ��1		�H(}����rH�o�Q��e������R��]K����5�*-ο��X�-����qu���z���F��p��J�U���%�pw/?1׌����g� PJdM�c7EF�z�I�N�j,��c��3Z]�7i0�~�}PRSL�8��W�@�tf��+�R	��J��$j�y��VyNߌ�4~c��?��=Ғ�|1r[�Ha��t��-��}5�<���O�WDN�Q�tf�9|��^��;Zv˿<=:u��zNN����7 p�l�d�N.�L��?2�����OWG�3oX�a �3��]@j�ߙ�� ��
�����\��x̐:��L��^<V--��&%2�iyP���q%}�°�����B�����G8G* � 9ν��ʈP���O�k
�����Fߊ�i?�9�+�>!]�%��q,5��Wэr���!w��xفW
�=뷛�3*1|s$�;*%Q�{e�>��G���~�0� +uS��7imI�b?&`�J2�w�[�����23?�	a�z��?���|r8��?i>aG�e%�ןP��E8K�ǈ�V �)B�sW$�i��0L���@wq #��7��S�"�Pˊ8/0�m��h��k,����3c�:61��Zph���q����'>H�C�z9�fR���R8oQ����ݎװ�-X}��iד��$)`g�>*��ǳ��=�Sr�a����ie��U�.^@��y�䘵�a�@�K�?�c�7� ����Χvd�]�Y��{ SLj���x,@Js�.��(5��{_f.���6���	��~�1#<!��0�Sz:��z�7�`�������VE�`��ک9�,���ѼV�༦�d���@�	/�������
� �b��yF<Gp�Rz�6mr�&���Ÿ�{��8���>Ak�K��eS�/��"���۴ ����j���b�ZTZ��6�22��q����M	zIǩÜzy|�,:���߃�Ǩ^n?`Mc�+�C'�R,�h�� ���&�2�l� f���-xO!���@ͣm���[�?��sZ�����2jWb0W�x�j�4���3��S�~�C��v�C͎D��<�"����N]��M6j�ѝx��M������:D�U��a����9��+�\�j�

�NevyUJ����	��̈��#�5g�{��jִ�(��2Y+.\.ۊ����~��ٚ�'�K��c\�k2[���W��|].�՘�N��W�d�ï'���t���s�TB�;O��d�7�hٷ���4!�7MJ�C�z������e}N
��m��I���)�vC��=�D��?C�#����Zf��FO�䩭��/Yao@��q�3_�]���%\��f ��ca��n�1�:�-7�i3M�%��)�Ƣ�z 	�솙fE8t��P�,x6�������	R�=�If֓��L�y�V�u��X��9%JQ7��+������V�q���g`RK'��^l�'�T3)א��u!%3���\���
6N�

`Y0�D�I�U4;پB�F������`3�i�Z�2�$㣓J��~�p1Z��ysD��KOǇ'^f�6��O?�,�I��!�9u����=��k��n�
�U�����C�h$���E��i�*X.�p�ʢ�ŉ)u_��c����ڙ�@��ٰ�GM��ܔ�|t�;�&��]�l'_� r��w9Vf�yK���@�%Y�N>�R�t��|�z�*�^�u���$�Cͮe�����Oz֌!��}�Ux�k1�fG�r<���p�EБ��]���� tvx4J�}�y������M��,3_pY����5ኣ��4�/;`}/b����疿ī�E�����~�J�:{L��j7���ě���k%�a��E�N�X�:��N��D�7Pp�$�u�D "��|{�c�魘;:8OܙL�zl�ٙ���7��;)�.������@5tҽ�1{���U���0M��r����{OD�T�����ޗ�ݐ�Q!>:��Ec��IT��Ϛ��j�1�����%��+� �wﹼN۶�ր�S� ;7�-��6��J��"��*��G����G��m؎8R_�~�xp�����2:+��g<��,v�L/�`)�RO/}��}zĠC�oɈ���M����T�W��Ҏ�5T�C�T����y�KiiO��,ہ�;�xt�2@�Т���*�`F����[C=jLs?��'�ql��UܭP�=й���#b�|�8��?"��d�aޱ�n`@H�ƼEsQ.EY$��Z=q N��?�1D�O�����kC��.A�$E��ưd��k�m5��}Ǝ�f�_k;xO^ر�����5-7�u>9��Xޕ��,gdg��掀 [6�v�匬��⑜�.�&21>YR)��v�q>I�~ֱ�}�J���`�q�l�8R��mw.���&Q�չX�[�#:#��[�K��O�Q�.:�y4�z��f�?��W&e��$���"��k=�s8����m��w`�t�kH�K���o�˘�U�3�J3-85Y�5�OD��SܚK�T�$���R�
��^�J��2����2 �0Di���z�ƕ��'v�3R7� ��@���g49Iv��$?�~��"4��v�P��6�d'��H���7�ØffrH<xϿ1�d$�W/v!�X���m���F��D>8�+��|^)�:�I�|�,d#�����٩o�!�=��b)\y2���Lԣym�Ak�X�-�ؕ/�$�}�B!+�\�#NA �b�Խlh�3�ӌ"�:�N��_�{*q]�1E�2<?:��4��DNrk���[�ȍ6�w���fJ�2_�E$�G����@� O���`�*�^_��Y0��L%�m��Ud�ͭ�hZ�T�N�q}��*��uZO��g�����q��2U۞n��.%c��K�J[�ӜuF8��.:�=�9�D@0��5�x)�������l�[����eY��U���%�*��4�3RT���0o H�%.x�\��l=�.�0�Q�rS���y������i�L���)TYw<�2s�C�!�P�e����A�+B�ȶ:(��;O�6��^� ���ܾ�b&�8$1�[�qE
�������gA 1��A!0���rB�Kp������M6�s2�E���/NiE�o~{L�t߄�
���Qg ���!b��.Q,3������ʮG[�P��3m��7
U�A�����<K{�g����k�+YU]��f@<����o��O�FVj_�$��@g[f��(��<����2a�DLfP$���!Z&�!~4;eʝ�{�|~��������"d]��m��Ǎ��<��F񼪜X)(�~3����(�������
�{�<F�Ba��xd�蟀��-g}������%�ȵ�iV�t�'� �hR�5Y�Z�����]�����4� f�m�:Gꪫ{4�������]��+��|��Z������S�c�>�s#��v�{�8���H�y��$t�:Q��)˩�x~'�V#�zxw����=㑗y�w̏�52�$i��H�Ă·�(�o%�~�u�1��Ȅ�w�����s�$��`b��Œެ-�.:��������r�������3ao��f�^�Y<��ٞ&�����1݉��!|r蘸���B�0�\>��%x��!:�&��0�4�ۦ�6�����Ǭ�F-`�d�R�A�\:m��8�������[�^�k��ptga���r���Y��*}z[�����(�ʙ�;#/:�Pa�0�?k�����G�:���Ϣ����PpX��є���./��0"��h}�R:m��,��'���$�ޛ�����`�S�&��y�"� �݈��[ ��u+
 ЈǌC��Ap��������=K����T07��R1�?7��$�=Oް�q P�v��B�^���+��U�&�ee�\�\��r� ʼ\���$49�ꆮ`�>��d�VѷwRj��ߠL8(���Imo��R�-X��B	��$�'������,���x���](ʍQ���dY�����W�+ x�`' r���4�}��� �?�c�=c�/�Î����Q�@�� �k;�t��:Z�+�������k��\S�
���_�d�-:R�d� ��F�4E��l�`���upd����JN]G��c��$�"�>j�kN���ע*���3.m�z 7�����U"��ꖏ�д6�aV��[j#�m�����0 @�C���ʅN�*��q������Y��(�kĖ��da��z�����.�~��O	���;�sA��sFSؗ��*S�o�)�7@��E���8���`;��`_$N�Ȃ��+�@�qݹ�*�Y�h��cjҘF<|�qk���]��� �˖�m#�����"\.BV�H#1�W�'O����p:�aѸJ��rт- zAQ�҄�	$�O��&�W���Ǽ���FxrH#� �j�Ƈ���sF�W��ܓY,��K��aV(����7u��H.����%cMUѕ��^���Y���m�@m#��u�RC�����n���̧�K�����6��D-�Z��:�0up�u�vO"��̵=��)ra?!㥾�_E�L�?V�ؘ��U�^� �A�oQ���&"a��řZG��Ԯ����#��VQ�Z���%V�0Ԓ�d��\$��Ի���U�Z����u�ݳl�U���8���:���Z�s�d�k�V��d�2�7�*��ý�[�Q0�mn\�*E	�6U/�Hq�'�;E��0��u�L;1JQ
p��y��b�RT�{"��Y���Qg7\UT�U2@Z՘ �P\|�9k&��q0:=��'1̛r5����R`j�E9�E@ ��
�������L���5ݿ��~�o,�hC8�sz
���b.���o��7����͇O�T���v1*�eWN�p�p��P�����ez�CLî�o0o���?�y���U�(E1v@=�,pf)p0�O�C��fR'u3N3I3[��<� �ߨ�茀�&*� �j"�����N?���ϡ	��q��Z	�����<����sC��cР��K�~�߆��{� ����?|w��}Q�*����5��-�pe�9P��i�O��Z$+]����E�m���@����7�s;>xn�9?{�x2)� oT����e�3 �W�tE�p)�SN�*S�%�mb3�+��s*�������ko*k�#7]l�����r�~=�>f�S��xb����JZN�5>��۞�q�ﶉiJ�?�3���o\�u}�ڹ��]q��b�D�)������+ğ�b���C1�3���0KaS�9���n*$�o ����̈́�ꁉ�V��B��a�{@}]�ů-�/�v�|���JCJ�r��{��`B�Uv�_��R��˜I�%M;��7��i�~
����`:�-�1�f�6�ˤA�THB�g��S��Hp�!L�fR��u�u�b��a�/�{x����lıy#�'hG"�\�ۉ�;��J�T���*K����b��ǋq!����O�5���8��a�Y�kA���^1�G@+�8O�����xF�m������Q�\h3P�_a��p֘� T��˘�I�o�DUZ�����"+�[;U�7/yr`0��S�^�j�\�
�R���X���؃R_�-g�/pp�F�s�l��`sEU�,�����v϶h�M�:U�PM��so(��A��|cd,w�
�	*7c�b�n�j
1h�< o�����;n�/��T:ߑvͧ���ܶɁ�9��a�����t�wxV��DMt7�~t
���a�p�B(���s.jc}�zs��#H3sV���c,&ň�\e`��~�Z1�1�-�&<�*�����*�����R'�92/A���޽�ԗ31���}E�[��P$�Ʃ��d���'��p�;���#�ҲXJ�;�6ģX�ǝ�2-�%ye�4�ՠRw��e�d�vʊ���7��a~Ro�녨(R.y��"9��M�t��ܟ�oh�T���j�%s`��i��(��]�X#��6xk�t�c�pqSێ��)SC=:|��;�3=TgE�q�$(Ȳ;�i����ϰyB&��@_��<Ʋ�p��||�n=�>�[-��$U-�ܢn��+:�G!�PR�No���)��/zV}v���5v,����9Տ�A�;��*��Z~��&]Nͼ�c�Z�}E+N4v#��+�0{D������Y�$u�
��]�nʫPhi��'R�+o3S���O���Jp�fwt���M�!�h���cDɟB�-��LD�nK�Q����^Ά)�V������,���)IC��b�(N
U1��2�p=�s�+��	��6��[���Xi�:m�Ju��D��t� �����ށ��:Ķ76v��r�̏{ϔ��1��u�gF�c�_ի�e ��<WId63���#a�aM���ř���'��w���Z�Cz��=h�Q�%�g	rqܜ3��Suvݐ�c�����j��"�QAJ��<M={][�o�{��:���ݢfG틬Z2����C��PNɻ�����#�G%��G>>��LK��d�fb`sR�	�Gj7+���e����d�p�)a{V���
{=��8����@���>��qT��|XHP M�����8t4GE�HC��>˗ǳ��X��n@,/�8A2���CG8쎥;���'i�"�ܐ�B��53�Cм`����Q9슭�d�t�-�����R�Mۄ�N?8c�َn��@��\�F�8\�dkn�)ZԱ�5��j/��o3��)�D�F"�u��sAo�}�MI��{�t�'+ʸ2,'���eFL^�a�"��ܺ�����XX�9t`�ߖ�󣎑e�Z�4R�W	�'+����&ݍ��3Xy��վ���}ݎ��wD�Ǐ�����9�fmL}T���7(�FC&4��b�h��?�,�
�O���~�o�h�����`��p(`�j�J����fֶtɬ�����3�X�`��cz8�W�4�ʪ��#�	q�%fpA�{���8q��,�z������e��JЙ�2O��V��X��3�;aG�~ҁLY�L���T%L���5��"�+u����4� �1{����]#Y������2Gkΰ��t��D���d���.Ǧ'����ji3��V���P�yJZj#矀�C��w���\,5R�}�#9w� ��dgi���wԪ���u���z��g���M�LBo�#qTZ$�+K(��Hw
Pә�9ҋ� �3<�E���.0'�ł��6JMU���w�0r������-��Eò	N9�I�2J�Կm�y��5٘y;��`��;}4d||�����)�`���I�/К�&i!���=�<{\���K;M�/x���D���T�(�W*���c��ƞ�h)?P���QW�Q;S4���`��r��#f-F��zU ;r�P�0��S�Ґ�q<:��C���˜	�躬x)������bP��PE�A��?���V�Pn�����^���>�7{�-NHEz'gE�XCِ����|�oL�]��h� (J�(p<�P"��S"D���:��-l�wh��hqI.���Lz�o��W��7M=�]�m�C�o��W�Z��E��s޴t'L��e��;���.-uJ@���l�G��|S�����~2�%���yx�Ƈ��}�3��\�n�+6+�ɝ�>{�'�a��c��͹hvDalt]/m��*x�r�8��@׸�Ʌ.!���n���=6�[����a���f����V5&D��{/c(w��&�V��n�Jx%j��T��0nJ!��#�K;O�.B�X9Oش�ֳ��h��޼j����Ā��2��E�����s��)S���@�w��b?8+�����6�a�� ��P����������M���[��5���'��q� ���N�~�XZ�� �zB�׌�,��έ��#�H�(����}bh�W��D�w&���{���QB��p1u���SG�J/��S��;62�3�Y!������Qc\�v�/�)v��B�'�J��x%�� miu�"H�h���Q��[礞�g�dcV��`I�?j8��e�'$���J��
�b��h�qm&F���<N)?��˂���-�ChgYa����ޠ��T�jd^�"���߂��]�ڳ�,��uG(<jltFeҜ�Q�5C��|�}э��@>����y9�'�o�+�B(�҉TD�%�- �F9좌�0�m�x���MɎ�ȳ�b��-g;���㇟e��X�ՃV(<q�ou
	yo�&��A��V̅��),u�P��Zڧ%�ԞC��xN��\=DUY!6��R���JBK/��	~��_Pm9���~[{�2��B��S/0[NHU:�̠�3��pO�}G��`���쑸4Ԝ����C�Ċ��M��3��k�d2[[�}tϛ��U�5$����$x(ؖfSXQ׷�Kdb}Φ ;�y���/�=��1mכ������`��Cvb<׿;��0�����
�*�:}4��*:�mZ��np��2�dߣ�AvT@�ZdKȀ8O���	����Z:����N6�� �^G�_�0���e��+T��J�h���t��!V�ݻ|�^�M�����+*ոi��v�d�5���v	WA��_��g6�T�E�ִ��fi8�
[E��Ԡ��|�y"�E새��� �ro7Tw0$�i)��-9�'HOQ� ����&�Fݡ����]��m�۠K%���w��-c��4�^�ܷ��c��iO!kT�ZAh|j�̂
���g�%���l�+��$�?�7>`/w)�U�2��Mv�f��.֚/v�2A�� R����h�|_cr��� �zȵ�x���O�jBl�����?&�Y��w��[b�!U�]l�	-0x��yՊ�_q�*�7��9����
ږ@�	cu�r�����c�D8�T�-ǱSR��a��_EX�"tjw�)3�YU�jBC10J�I!�\D��������Dc���|v���i�M��=���5w��T)C@�C��KN3��v �D��|U�tW�r��=&�����	;��W�W+��1wYG�l�;F�׺ĬQ+��2�S�4�P�7���c��,Y���_v��t֊$`2#%���̯�c&��j z���.���,Mnȹ#T�Z},7�ĝ^�W�?D���OX9;�*	yp9|B+��'���3�K?4$�ā�F��;���5�Jɘ(m�@��s�'���)qF��,G�����W��r19�u��-mE��b�a����q���8m�b�*@�5����]t���"%Lz��ہ�QN�4d�B����PbB��:�3��X������r]����^KRë�'���f�&��l���?��)	4�#|�<�K�5��E���q������IS��A������t�+���֦\��s���p?�SK� ^�\��,& ��g5B����93%�=���X)��^�y��)=v���I^��ٷ
��*8���w�k�Z�E��c�Dfwz�l��� �`��쑨C,�o��9S����d��Zn��:�t�t�A��q�l��#�p=��~䞙R�b@�Ʉa�~B~%u>W^<������C�6&��R^��#]|�Ky�_,��'�Lf����@�ܭ���4�$����AV��ك�ȥ����bE�(�l���+<����V��Wz�H��Cp^�p'[�Ҟ2�T��~�!�\�E<�rs��G��y
�����|ب��\�h���eF�e�����g��z����0���=����xz�n��v��ˇt6���:���Ѧ5��p��x�U�[(�{Z
���g�/d�
\cմr� �?f�*�ck��"}����_� �w�G��-���Ǘ\�&�ԇEvZ�s��UӞ���|�����Co.@�Ťw�SU���"=�s6C2�w����[��ST�<#}��-�� ,�Io�S�����4k�:��m�������	Z�U�I�F��ŪB1%�w^@`�z�Gˎ�,����	���OW�����}�c�D/vp���_��M+$D�So����Z����3�M��g4hkڒ�i���qd��:%"@�`�^��ܒTY_1%�1*���`�M桚��e�X=�j�Zb�4�/S�{0[,�$G^����ȇ��hF��'i�>��\ҙ#9�6��.�q$ۮ����Xy�{���<�g?jP�ɇSq45@��R���|�2D��lݿCK�j�(�-t~�(���퇥Ξ��,�
�sp�V:�,�9p����&c�mJ���Vnh�� &q�{���AN�Rw�bUƵ�#���?Z@O,�;�8�,�	��F���Ӽ��"�7404�<�U��2"�Ve�?}��'|TPVɭDƙ��\��1.����8Tb��+��5����֌&g�J��>�U�5���\�5d�=�B�@(1݅E��Y�pc6-�}��l��poX��q_ӯaZ�U��� _��1���f玗	W�rΏn:�Mq��_4�ɕ^:1���,5��m�.E]���� �p+�8�D�z�K̭� ���,�Q�Y���9
��t��qa�-AO�uqP�75e2O�T�
��x.��7�u�{��H���p�# ���g�t�f� ��(]��u
�rͬ���p���~x��1n�R�W]˳J�����~��0�2���NY���n�ٞ5��P<�kV�U�mI'������q��:t������F}:mT`�[uXPYY���G�$�8��Nga�<ǥj��,����'��[��>�mO�2̈́!r萁n�Ԅ{�e3�A���.IA)����o�G�����)�޳�"1����}Ǿ��XL����3��<���{�X+V%{���jz(u�SР���d�]�{ђ�\�����sI�ڒ��E���L:d9<�4�P�MM��\���.:�{1&k9|�L��y�z�}�P�wтeuC��п����h��e2N�	�C�@ߵ}:T1]�����D�.�����no�L@��u���Tr˄\jO/J+W ������'�
�7ע+)� �J����9376[�wU�؞u�ƣd\����yف؜P�a9���,�%�o�a��\����ocJ�,@5�^L7�:l�j��^S��̨j0�+s�r>�-��aq��z۩t�2����8�|�3��39,Bo�q�w��%�@�Q��b�J`�v"Q3�͙k��&|������0�}{��;)1XBZ�j\�gyu0c�8j$��|)���)��QG_��Ca��V��-��mE�Xi生`=�̆�R�b�B����I��0ٞ8�������4�?�U�����[�U^#6�����OdX_vUg8��=f�	")SI5� �s>��� Q��@��o75����T�k����+I Y�%��m)û���%HI�u��7�&�^�˲���(,"��_1���}IVq�]�#�k]|+5˷S�6�Z�IzKco�Y?�`x����=�����JjAΨ�ȋu1�]�I���^�秐�nQ� �Dc�]�6r�n���%O���l%S�t�C·I�h+�V�>�a�NƠ���ra�m�ֹ
�7)y��7�]L�6W��m����PI�C�~��貴�
��e���}`+�ɶ����0[� �cX�5�C	5��$���