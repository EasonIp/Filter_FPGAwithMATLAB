��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~���"WYj����i� �N�7A!�@<e�]N��?�jj�����W���a�q���#����MP�F�pdoF.8��+:���h1�ԭL��L��[j�1���߀/AP�0,r�F��x�N��>�RziB�M�\�P�ua��B�MɥBe�U�����v��+�R��|BC�:6u��8�B�����趟���*���I�lklry�.T����b��`��qe*@]({�Zc/��:r&�}��E�#h���c\iH+�,��-Ď[��Z�&����̧h1����{IE.a�]����C�;"ur���9���m�W߫��H@<Vh�/������х:79����g�{��)���[*B ��?v��,�k�g�)?c���:�C���Kq�����L�`�3���FԹ����B�tY���4��;�*�U����hL{����]0L?��	|�G7�y���J��nT#�@���~͛��j0�U�	�RF��s�K������D���X�_�+�Fy@�C�5۲,%�z?�Q\ ýZQ�s<�;��‹�q0�X�u�1Of��{w:���]��SuF�O�{�_��Ž}q��m6<�H5Fm��G���M	g���U��{���xz3Eqjj �E��%hV��{v[�9�"����Kk�:�AԎ��iI�Yb�}G�C�1r��,������3�5�4j�zs�y��E��\���eX�k��9�4���?�嚖�0c'��L�Z��'(��z��la�A�	ɍ�	a�}��zd�g� ��+QS�r����mǊb�cܔw�NvA�Ց	4&G��;�hw4S/�z/<-��I��$di��a���YO癦	�������o�].�#MN��Sg
0o�����*�%�N�
�VG��U���m����^mh����ܬ�`�|[uH2>����"Fdr^co�.�:ꦍ>2�ˣ�GVs�gV��a(V���@|�ȼc35���Ʉ}2���}���%SRZ�|�˅p�r�o�h"P����.���b��]F�[��� P�%������n�dtv�bW��`���_�į4CrX�H��RW�����ī�OH	m�r��M]D�[��)��\������soAML����at�d�����ZG����UX����t�L5�@������_J*�bJաW�p���S�7��cq�盧`�r���9y|�:�N��==����R��D���u3>T��Q�뿬0�:���.�vkꕿ|U��-綪aT *jT;��*,#9��1����Ƿ���#~�F0��|�iÍ�[}:�/�u�>e��>v���q{��Е��(�)~���x=!�NL�N������#�A���mH���s��0M*'�sL����ͮ���#U��ȋ1�z)R������7]w�n��e�nH����$,g��K֘�@�-D�ŕ���Rŵ8���*���^z���o�^)�J�^;���m�ϴ�h
*ˮ$]T��h����(rSL�`��R�s�Î�����iJ�_Ǥ����|���Xx��Wu|��>�v�y%e��;Ȳ�� )�q��,�Xن����CJ�d4p�b��@*t��2I(D7�YL���5��͊�8��VΚ�R������-�<CǨ/��5b��/"w�ɯ��ɇoDӏt�q����f$i�ql~1�/�VS46��د�A4x�@��!>�h��˷?Wߞ�_#{��3[��Ŝnn2D�/���o�輶�#K��W��Ї�1Y`:��J�~�#ˁ����oB��<�*^|��7ń���JH����&1"��@�L	�h�]o�J̻�g+ܲ}Ŗ*��ǧ7`�m�#����S�����4q�]S�";'�ҳ,��D>Oz����}.՚[��]�)�=�+�����e����)��Im	JwK��G#�kF����ʶ|[ēĿ�tQ��޴Y9S�L9���,嘒�.74�}@�z��Q�
�<0�[\yt�\?�����0pFy)l�6��ǭ#F���z?A+����[l&&��wR��Sq����Z�\������"�$Z{�%�ę�O���twꎗD���'���t�l �Ze���,�xk)�y<h�-��BT��䗱�T6�����}�"�a���)��0'�ӈ�Hw�HRqq�IV؟��~����fp����L�IO��t�����p��P>���c��S�º�J.M�ˑ�8_B5���������3���5�{�Ҕ�8�vB���o��z*ƚv�����M��uu5I�nyf\IS]��jl�1�-��d�QvT��|:	?�[<Hm�J��:�1�s8�,]Z�<S�M-9��Q�zʚ�g��Z<����2�~@*�uH&�����3�WA�Ϝ��h[O�O��)¡<>�����z� ���R�<�*��M]Z��}���`$flQ���(L�#}��<���Ac0���H5�Y�~)�l5,{-�.�b?N껽��J�a���X��LR�����!m8|asc]�1����R�	����}~A1�rە���kQ-��j졼�P�|��)F��Zyjt�M�j�P����B��V�Xt��C1���;/����Q���T��
�\W%V�����F1j�dXM�KK��c��5�%����KP�$J��u��k@~�1�K�
C:'�nn�Ex��p	�vS�2�'�=�,:<��D����W�_��q��[�j�u��˼Իt�M"��|sj\?;��^6��(�eq�ۜ�P02�Yr�U��ﭪr�/#O��;L��,L�� 2�^�~�.d��+��P+R�Q���yڛ_��̀	�7��߳;d�#�/��Ճ ���>Mw�f�3%�<���9\˳�Y3J�~�u��6rH¾Y��re�����ꉥ�*%�m^�^C���T���.�M������,ѧ������f�u�j	��E
�4NT��M0���Z �EՊ8qebv5<�XY~o4��!�ZX�;J)�������w�4z�a�lG�V#��=�gu�;*��c�b��/�p134+5��ߜ8F��&����� �L��*�b#��w(؏����j�w�C�b��#(���E�x�<ny���Z�T���
�r�F�911�v�p�a����(�a���Vm��&V bML�+�V��WoϞ��8N��9�j�Ī����q�,�Ck�7����sCO�w�Zx[��O��Z�8IԼ��L�m��O��YW��2U���WAأXm;I��W)�������B�yydk,��'f�J �[��z*X�!�nuP]v!P���
^�HM�r��h}��{Z�'j?5�� ���1ֿ�H�Fy�%��5y�竕�e��'l�}X�+ �n�-dw�!C�=wZ�+�J��TNc�$�	a����t�M�"���4쬃��՛%�y��7�b1F%=��p��Ke�H��B�g-�x�	j�JgqQ��IL��c7''�$�D���v�gU���x�٩�P!#���	N�����j�GKrX���������&�W��g�*��Ck�.�~O�7�'qM��6�|�|�/�
Sc���E�y���\a3;P"�fymk�g����d�7Y�idQ�ĕx�*�
���ː�ܿ׾���u��;�g#�T~��*63�b_��Ͷa/ ���-Ug�y�Fl��߶�(�*��q���rbzyZ>��V�{7�-iq�h�*��6�?>7Ԥm�Y�wm�������z,��p�L�&:��2�Oj&�ZAH�oK���� �\+��*��O�U�G�t�K���@GШƆK�x גS�Yґ�d^t���:�	=�qiޠJjH0=��	:���XV�E��kW�e��<֮�?���C�*��rb�uIgAbdDl�� ��� t,fG��I�7`��frQ\tÕ�E��գ\�R��s�?rAu�;~�29��-�<�W�X"�Ff��SW�Xɰ-���[�C�<�k[�1� s��U��d  �K�ƾGߠNHw�ÃvDҍ��$N�`�+�WT+$r����}��<�R<�t��deH�0.N¢B�Ʋt0}�����M��gU< ��lb�͵�v!fc�&`��9m�g<A�A���Y��D#�I�n��<���$Gޗ�;zjd�
��,�5��RM�%����L�I����u�mqۤ���jx,0b��*��2����ͭ!�p�-9�[[(0�a�]7`��"I.3���h������p.cp�,����HG�G?�3w��|%5W�[*����8����t��\�6Z�gi����TĨ�'Pm�=�����0!�B�Z S_<���jO��fSי0A��c�t�O�]
Ś�1�������TB2c��+��c)n�c��Nm@WV�
v����
Eh@#�>�[��j$!MJ?v
��\�xB	�G��Vt�,�냃�r `��~~��_՜�� ��|�w�d�q�hu�5������Q��k.l)��ȇy�<�i�h�1�͎�}7c+��M�<�e�8��MEF
zL5��!4�b��"Í��Η5�w �]�pgD���eD|�fɖ�����X���]|�$k�.Ӏ�2�����7�����3�B�B��_s���3��o���I���!T��P�^}#m4���=G,"T~҂j(�p�M��}i�{P��:�7J�vV3l~���B�>uL�;z�)��B�o�c|�'fVɲ�Tlb���K0r�i���
@�MH���[���В�N݀�D��^���\>�E�9� ��vvP�M�K� {Mf�/��âK�q�,��(���Ƞ��gk�c�̆fē��8k������Z	MI��:��ᐶ}U�kj�\р*�}7�Kv�ZO<�����uf�0$�O�E��Yͅ�	�	Y8�#IBp�Ƽ����]�m=��%x��x��9-��:ס���o+���H<i�9mPw�7|o�c%9��m���̈.>a��_��D�����%��+m��f��Y)%�_:SΆW���x�
t�>~F7��ȓ��Q ��a���T�^��.n���3T�3�r�����N(�C�� H��Jņ�0NH���a��ˤ3�F֢}�RӋ�=Uh5�O�4|���S�h�4��8�.��) �����q�:2Ld�����c���b����n�f��I��%�\����I��G\J�Vʡ���U$q�G��Plګf�K����	Ȝ�ق�nY��f�!�W�>X��������`�淬Nk���ޥ���$�r�(���6����U�ɯpP���H(�Byƚ����]b���X�i�hj���0�j�-������i�S�ZJ�7���)}t}� ����i��'Qc3�I��k�j�n�=����[�K����\Xgk!6����{�Cg L���k@�0�y�ͥs�K�� 0�g�GvM���s�ߤ�	�q9^K��,���0w���zH������Z����2ɘ�i3�`g�����S;���#F1<�:��#생�e��Kv&�����s�ޟ��)���9�'zX:��e8��F%Ʀ|L<�9μ1H5��6/R��vrYxۋ���~㙾���r�Gq���>K��>|�-���̇"�(R��楷)a�D��it%�`��*B�!�L�Q���0Ԉ�z	����A�<=�~�4�2_��%�}ß��8+Q��y�f�GA(�@bHa%x�V���Wؚ��=q?aIԁ�P!����ὂMy�p!�=���Z���1�k�s��NW��̞��4 ��ǎ�P~��<�	BHR勰nfzqCi�`�^e`:��_�>��B�
~���?��)�OzRh�%�°bT��a72�,*?`��&A�P��[2`�Gw7[J�S��M>��1!֩oZ��2����pDݾ���_<ÿ�wWr'7������ M�w3:Drɞw�����)'�"vU��!VxP�}���H9r7�iU���W�3�|��!*^�z��]6�b&xP;<��~FR���
��¤��
Y���{��kDcQ�T/l�Ν6<`���ێ�����I�Q�r*�~ⵄ����沥�AT����4��H��3:��p��dJ�I���$H�����IoS�rn4o7y����>}�Ƌ��I-�W��Un__~�y�3�UP� �'�z^�N�����T%�Tძ�&���w�B]����׭�@1r[%�Iw�R���.ǝ���F�t�*uUǞѼ��	�w��y���6~jh=���˒�mM�	(mQ�Tr�2�p�y�����
u�`kۚ0q2Bhm���H�٤|�P��R�ڲy�j�����h�5�b��Xt,��,3�ё�w�=V��Jd/�=�<�?\��<��JS���}��$o/�;���\���@h���\��\J�����B.5��Lt%�RD�ޔR������k����Y�����; 	��y(R��tr�K�^e4cΑ�ފ%f�ef��ݬ��8�IZDq���2��s\��-(�E�r��6��inN[�tN*���nWx�'�Ѫ�<��o�,��!���j�����t�{������pđ!Q�EO	���
����ɒ�;϶�k<�7�|�Vi���I.�Ր�;�������>J��vw�b��A B�K�4�o%}�6Bg'���ھ�&��(t)raG��v;*��Raڜ,~�N~��Ƣa
�4xo������N 2�|��T����L1Ӧ6c�C�fnp~��}M���bL]�z�Q�uK�Q�i�ā���W����k	ocD�&Α�:ᄒ>�+�%z�(�J�!v뢺5I���g��L2���,�E���~1�W�-��������ę�w��T�_c	n�]ʅ�[R��'�_��MJ;IP-��bn� V$| ��8�ӛ�k���|
���xϖ�D�X�����妎�L�F�8L|<�L���ݓfD�+�wOOpY��.��8zԀ)��`jg�/Eغu\����&��=M���{(m0PZ�����y'g'B��0;��}��1�V�߱�䇆���k&����q@�1�o� a�Y�/�L�J`�B��eN���C���eʽ=�5Ne�b�[P�/o���B�풻�#���>Y�I�'̫}	��{��{UXi�H{rќ��>�%��¯�$/+�G�wSz�>{�S�M	�_�1����D:b]ʳɬ��뇦(ʐ�f�AwE�CM�&��fe��_�Z�˅�c����JMU�}l����<\����a�Π���G�o�mB��b$9�01�3m��/Q�O^�hw{�|Ĝ���X>Ԏ}��\��)�A,n�\D摢�y�hݜ6�K�X�l��Pxdrl^�. �y.�k�L!�Xy������v�h�+�Q�.Y��0y
��{���y�:I�1<�)��*��ea_ё�V���jد^?�jE8#���:7��!+*G~��@��{��@�)�.-��ɤX,��?�xQL4"�0�Tu��gE���������Qmcy/�0�cXx9�E�q?�Q�������@2�������: T�ݫ�b�8?�~:��>��c"C�� M7��/���'ǖ����,�P�ۊ�/kb���_�#��L5C�q�(�.��9̢��XC��X���A՘�˜���� �g��Z�����mܥB��Z.�1��?m}!�<�¥��dAv�hf�G�e��5�'ֳb�z~�k�4)l�ʹ�H�{t���&��p��P_���+����<��)@v#��Ҁ^�̎�-��ns�����Ӯ��_�H��͜_�o!�t�OGI���6v7`�T�j%*�{�TD(�M����0��I����6��xu����9X����Z�ց<d�}���u=���9��l�X���af�+)�`��7��jvZ��gy���4S�P��j������4G:C�T]l�C��s����ݞ+�￣��OmąP��Ì��M�I��J�����$E1(X�b+�.-�����7���}2	]�J%��xD�:/�B�s^��	AO���ϭ��J�,�O�0��[ԙf�@��\-�V<�Ǯ�a���P�E�㢆�N~h^�p�b��B߭T�#u���=�GѻhU�:���ìݧŌiF.�� ����.�o��x.��O��=�K��ݜiz��*�/Ա|�xM�9o���2��v*�d,��531|��"*Z�U�J���ƋS�/�4`\�[��@t8?Ǫ%�Tu�֏�X��<)�E �wAgn�.SL�\�׿��5W��sIa�����ɀw���3�`d_:،�zϚ����J-��ʌ�W�*�Z�QԞ��>����|ۨ�ڰ� Dҿ&*�B9�Nw3bj�P��2��4�:U�������� Q�<.��w���m��3}	�WH�Ɩ����`.�D��v�
$'\`��n�h�g��r� �,wk�� D��<��y�O�$4�;���=C".<CS�̍�< 8�r]2>��D��5z]>\^����̼�gi�������c������Lq�PʾND�1�2�|�0/PNψȭ�ܼ'P�S48�I>G�|"陉F����k������2��
$`ȇ��f@!o~s��<ě�LÚ,SdLd����/���E���4����!�YM�b�� �%U-3�h��{��c�I$�q�Ŀt 5~��#�G�5�@�ĵ`v�@�#�B�$x)��p�~J:����ܢeM(W��C�}4z����s)a�C�ʜ/�A���;:ߕ�[�ut]�p�&��nw[�Cq����_^��E�b;�7�X絥a_��LĜ�Ǫ}n0>��:�v)������)�m�\Rt�s��F������O7,Ą#�j)��0�0)A��	��NCK��R��Ac�:sTO��\}���ε\���#���ȳ�i���԰#e��X���4�y����L;�2��3������&E�Z/Xp��:9�$�r����2�H�ZXh�-2�M�yX�1�A1л��Zlfm�T�6ֆ�����LeW���f=����憵Tp�S�5k��G��]���L�X�4V����/���K�ܛ�?�Ε�yB��hB�x�)�_��~ic����.�9Ǜ����M���B 3=��"���A�7[l�i�g ���,��4�{� ��h��	B��l~�}OG!N�)A���6հ���3�ՕO=�6IW�R���4!װ:ЊgmVnY3Ϲ�Y �̢�I�A�}h31G�nђ+�����?��7U�тA�JJRp��9]����kyʸ�q1��?T�k9��w�!���lq�hf�^AX�/E3��Q����ܤ~G C"d���{���fw��ȫk�@a��~�����?�]��&�Y�t#T�2&�I��g��5A[����5��z�X�h�j[��խ�s\�oN��Zb��H�.���y��"s��A7*
 P��5j=W��׳��FH!<�n��"C^����?l~���.%��$��L"���v�i��/p�R=v?�Z
1��}�оw<������o�`��� ���-B�ҿ��M��G!��W������7�钇FA��%j?~�Jz���C�7�{��0��pe)9���R@�H�����B c%�����n���pqb���X��/��f�%,ܒ�d]�c�T��|�ݫ�v$��CrM�ehl�h鴱�c��o�"y���꠽|F�OmN0}��z���q������Ps#�-�2�#����Ҍ�8���ǲAͭ>U��Agç�8͘�Bk���kEj�7��YQ�S��q��\ړG�ۼ���g:�pk�KQ��;i��$�l]��0dt'��HM���-˸�-����+�xc��\}u���;{柠���3sș��`�P��x.=x ���T2�ͫᎉA!�A�*��oA*�	��>g�3[��>轡�Ed�ԽE��Fe�3q0L�TpAQ�{q
Fв���sA^g��! ��8�T�>W��ɗ�RH�lK�=�����pH[F�Da㙹w��h=O�=T*U�I���'-,}��Q7�����T���I��o1z���q��&h{����I��q5�6�G?��[肚��"�c�y�̵�:��CV ����-<j��ݑ6�9��C���<����(;��ؒ�Y)?y�`t ��聇�/
���b=�\�Ϡ�mb0������ �g������KSR�&p���@ם# g�'�i��V�'Ɇ$�סV���S�7g=�>���{і��eQ�n|0^��&�sxTv��e��
�A�i#��m��8�L37ۻB�d4���j.{�Z\�J���z�����s5�VU�����	$��9�6WHa}1����T�*羱C� dG��w�[/��������Q���{�����I�6q�4����ʭ�f�n�8��Ǟ�=�niB?N.vyf����]X6PI
�:
MN8�#ȓ�A�.Ke�ܰ���κ�����M�rI�r*V�ag�~�ظ҇�>.�əx���~��G�	������	<���EHޥ�� ����0>�^���(��F돩�����5�:�6+�M��U	�n I*������@z�G���W����8�M鎣(ʖ�Α�h�a���8���j�2L��|KQ�͒�G#R*��g�$����jmv�pT�gz%V����JD�@�-:Pb̶rFK|��Ϻ�	>����:0�O�t��q}�,�O���T
0|W{����B�9s��χe6�� g�(^K}"I;�Q�\ϥ\����H��eJ ���|�<o�?���>WgZ�+��,�Pozܞ�>7�d�M"4��$	Z�a���)��]	�/*O��n�T�+ �s���~�nO�1�\6����y�d�� �|���
7S�|�.|�1���ã�>�'��z����ğ�����7y��^�\~��^�c��YaI})�J�#ά�hJ�;���}��ϴ�aC����Jpq"�)	������� &x��S�p�ZM��?$�p���6{�J1�{��\�ow ��������<��>Н��h�+����*0m��U�n�����4�g���:�]���?�HCT���?�y�-�`�T!��/�þ�19�R#�T_��ǌ���^��~����>��	ξJ��Uva`���VdPRI�zֲ��[-�� r�22�ޛ
M
-��_��m����a�ɇ��h1?xT�����l�Lz�)��I����k�.�
��*����҄�,}��;�g48�t�jG���}�5'�2��\�V@�L��!,o�)��!�e�n���pO�w�N�3zX�x�[�Բ���GgzD�����{�"�,x���7�@.[��%4e�u%�/A����'�w@>C�9Ka+��dv�;��i�>�+�2���9��*ۼ�<qO߷)i,��,E��=��B���1I�@��!QJs w1���j��]vޕ{�l�)�.Q4[0��L��@r�es�&�N9��Ug��dܘz�,�Gk��V��u��n�T�䙤�;���L�+����+�C~)�������b��ֆ�=�5�	I��J=� 0�j��j%���z�m[D���k8��c'�sS�ϭ[UK� �V?Jc��⛬ʲe����2)�r��Ag��2r�� �њ�ʀk<�T�H�1�^��7;ޕ�|P�$z�Mw�vh��C������
�W���Ѷ@�k'(,)�Ujs��i���f]��G�Q��(r����>��d*c10RM�aal���{���¤���cE�Ql�3�~+�@��S&!*����0)�h� #u��u��Xj_c��� �I�xo,&�3YOW���F+ ���6�^v����P��T�;4�os���59���v�h�4��-�S�u���&bZ
j��*y#%�u8&a9�D2o�6<�`��/?�<1м��|�岼S��V��l>e��������o� �V?T�o��?��K;��{�:��Y�㢅��N���͸��]��/ߡ2u�>� �,������X�x���d����r��Q<�A�@&�߃�^�7�e��-���� ����й����:v�o(�jG/��-0-�N�Jd��G*�K]Q(��a�L��S�%>��x�>l� 損|B��T�h6KL8��=��ne>������c��o�����$�E���gȀ������x�G���J�=�kL��P`ʅ>y?w�|��c�ѻx��;r�/�=��o��J�?�1C�#���
�����?�|��	|��h�����jBJ2*B��:}fwp��b/èJ���f�s�$���W篒��kQ1�\��! �����L$v��Z�����Y��;۰��)�R�X��lQ8lt,
��l�,@p*�+R���,}5��8���T��-�	X�|T�v��9����l4;�%B��jGS��%	��󇺋dk�,��;p���ڸ�>�[l���.�s8М��۾��6nD�~��G��r���{c�B*-1�,��y~�"�
��"K��_�J�� �G������e6#N}�5����W1�b</��H���|I����>�Dj�{���n������J0����
E��������n����gFuHENzݒf�_z8�{/y�?S�`��8��{$c:���V�F�z�����1r%�H�(�����GI�ck�50J�\?C�V1C"� �p����R� ��+�80ݠѯ0&�Qܤ��\ �����r���ľ��� M�α#e�����z��S�{F׆����U�6����5�3��*�`L�Ə��<��ⷿ��a��0�wk����Dm����9�� Z���&�����?ܥjbX�VR�:a��������k[nu��i�J{�郢}���4-�٣�����T��R�C�i�+�}�)w����I%�$d#�F�Y�����cz���ʺ�y�O)� � O����{!�_ ��i�E��^��� ? ��?���td,ae��� �_j����������/� �_dd9<�g�j�Z�Ȕ�]��-	[%XL|�����ꑛy,a/�ǵ=k�U���O���Ж}�����h\�T�1P�u�(�ݲx��6��Bɏ�x�U�N�$-�9"�BK7\w��߶�l��#;R��`��}���Q�M���]����ֳU�Ft�f�x�~I�n"��l�$�5E�%�������l~]4o<�����������=e?�E�����vh	�y���Y��/��.�<tR���v��>f�RIW���j��&�ΰ�_S͢��)��1�]��#����;�^�#'�O�;�Db��X�����g�R�/+_��N[8���P�}�N��pF1j��Zm]�ӹ�bz�")H+ҋ��[gJ"����`��,fT�����o	S���^K�ElC�p�_N�'T��jNX^2�����۾p�B"Aw����h$o(���Gp:�z�����/�}����<�lk��&�G�]nG�Ο����U�Q�|��W�ۤ�-v,zM���[��8��Ϊs�_l��9�ʳC ����DxrBZΞ�p�x��;?�'��D�I���Y�IA~���Q�$�V�t'=D�T������DT��)u�q�&�'��<M��t	D�(C�2�Z:RVK��J�����>�ʨ.}$��Z��q��P�\8�ˏTfd2{�NS��Ciz�@kh�eV��|�aL�����"v�pp�o��²�iӖe�-kA�9+�\����|G�ׯH�!.O��P��:aA�I3�֞��O�v�x�ο-���K,fhg�(~n�<�d��`���j M�,S����r�ٖ�)L�B���5�Amq���	�*u����0�-
�K���1�QV�7�x�y�<�-lyD�f�������ֲ�������Pͣ�b�����5�qv�>��_�tp�I��Bh}ypP�io���ܚL,|s(TI��w6�s��h�!t���Z�U?�O���VU�Rb�qt�09[�>:_^�O�qC4�C�凿�&[�k����NGE˺@�t��I�iʔɲH&�*�q(Rp6�����|H�up
ʃA}���y�$􄁏M	2��(�x�WZSL��Mq�Ԛ4&r�r~�:?Uhc{��)�l"E 8�tq����r�j1ٶq"��wʛ�y��n�;MW2JÂ���馏�Yޛy}���b�/"\�������5��Ѯ`z��6ZX�'�U�AiI��Q+� � Ûk]�At�$3刻���?7��o.�MT����e9I�~�������F&5K�;B�b��	����As�o��w_;�vR��#�#<�ռ\�WS��݇�����}`�ڴ:���Jl� �tM��j���K|m�P�V(�� @��G�s+.�#��p��Ҥs�y�}�����#�J�?���6;��E��I^v�+1��I��^��B	���P%�K��iq
���+U��5 ��;���&X�)7��0��]�����{�O��V�/��C��xr��+��D���4���r�|,��	 �9���ދ�����x�<f�%J�.y>��2�5� ��3�l���9��{��5�X�%��7XG���aU���FM��*���^A43Ӟ}�J ���ل/��X�m�������3�gsv�IC�L(����l'�A����̟5G%B�G� ��Gw�7s�`�p^��D�Ro�MX�vm�H���k���!���%��ٜ�k�箉)O ����'"������;�W��,^q������i� ;���u����"�D�_�F�3x� Z�_-9=�UEi�do�79 �������`.��\�5��rmfa���@� � ��x�>1ѳ���
.x�u��i,�2`LG�����Rh\�E�g~h���	(G�� z���c��)���yy�����>��Qv�'�U�.��U�ρO�Q�	�[�56�E���0d�ް�����QS�Ѵ�K���~p�g\�e�uI��0�]��]�L�>ɧ�w/�d.N�q�8�qORmB�	�ҭ7��fp�호��z�*���8^��'6��_[�����$�[k�9W��	lh�;�].�x��q�=|��;h��_ĔE�a�[R~Ȼe:/Ph#%s���>��BmW�7�k$�DX�MA��=j�fs<��YR��������������(Nw��h[�9�Z�}��ճZ�N���j.Z�j�ǇZ�C&���.�o�q��`$E9d��[."�[ ���c�r��
H�I�g�r�m;Ւ �ƀ�<��g���i�N�Q=3R°�u���Du��c(u�f����rz�6���6���3��h�e��0��z�6�q��:�#0�;�ߝ�%>��攻W��V��"�.y=��J�1��y��[��(�凁��r�3T�1��8}c����︘�F$�t {9�$|v(R� dT������m0%{~�� ͻHɘ�k��	�bOLR�ٔ��C�a����K1���)�a���p��'�ۦw{� �w���|Hu�� ��t�v*y(@ Ew��rُ����Ih$��I���fv���&쥓t�H�m��u0��ۿ爢)�D�皢��.�87��8e�b�s�_:��
@ӓ֤|��2b��^#å
]'_B��B�4�泯m�{�(7p>��	��m�U _�꘺)xxN�Y~LZQd�8w,��p��۶��{�:�͋\_���rz���=�-���*�����002�%Wɒ�j�"(��sz~�V�	��wr1����i�6EW� �Q�r
��k�!�x��Bn�z�Χ�<��9\��ۣ������^��j�8�b�,�"r��ic�+��;\�BxQ� J�voTn�b�lW�eۦ<^��|V
p�/�E�s8�X�w��˞��;t.�z|E����y"A4����j��Vk)���B6�`�`��aR�S�˽+H�!�ƽ)�<ےr ׾�RR!_s�A�g4��;�Ov�9����3���dg�Ӌ�a�_�O�@�?}>�]r$��������\� Q���IZP�kSF,�r�l�_햨'������d{��b��6W�>��#Bh�p#It'��-���S���{�C��-�lʯ�cn+81X���gh�U$�P�2�p��n��$�S��\�_.�wcʃ!��M��*�$�8Gc_��9	����-�N�k#k˥1��Of^�����	�����]֫�h�c��-�dL�1����ڀF5Ϲ�J�<.�j|�TJ��@{�@��K�W:)��eR�,lfE[<�8�ʐ!��m�z�2w\�>���eI�w�5���u��[+���O��X%@+LZC���2�����o3s<�9H��Ҫs��5ڕ�� x��!
M���`���Y��!�
(�Qa�6��v]緐5�Z�#̞���� I�?(�~�|ƻH���b%v�n�{}υm��b����B�q��߁5=��J����?�F�$5Hv��IHYj�'&D�Vhm���Gjm����ӤP-�L�cȥ��im����Tu�װ7����Ym�)���H���a*�T� ��Nt��"���ݒk������*�>�5��/)��<p�_�pf���/a+ÿv<N�M�U�-�/u��v��rJ3%�L�7[�B�?	4�1���R����Z���8�~���k5T�G�~֚��ۣ�hS㗁s��H&�R�ˑ9F�?���_�%��ƿ���n^y=��/7Ʋ���iˇ�Z���סY,���i�t�an���x�7-��ku+��n�;�K��l�ځ��-t�����mط7��P�<�k���;e�S���fB8�o�@g[���#�B��#[��Xz2,"z���?�Ҵ��Γf	m�/�������yx���F�8�W�`ʹ��K��~-�w�*_u�G���	'.��	/(����u��`�>�B�<�X�D,Q��7�ߨ4����9U������Q�fm��\�_�bz�wi.�5����1������n�
��Q�����dKAio�2�T���ޟ�xf5mX�O��߼~��U��gp�(�:���mY�^��?ƃS04}G�a�]	�ۖ�3,�`;�ЊZ.����F4�x��$ޣ�)�2d���p%=��F��苏������R�,Y,c��}�@Kl�yr�w��׃Fzd�·eiУ��� ���:���'q�a�|��B��Y�C��Aex��G��]��ep�4��l����t32�cW3��9�[�4:�"��)�[�=��N�$6�s�VUfB�\�R�Y5l�T#�ie�g���8Hь���R����zw1�G#�8���|}���
�[f�4�_S�8{
+r���:������8Ǖ���g�~N�A��� ��/��po�{�7&0����--�2g)�g�$�l ��5���}���ӈdݱ���'
�A
}v#'��j3P��&��J�	^�?A�&�!+�kRjg��:m������˽��$HA���˴E�w6!������ߡ�-�5�?m�-�B�X��+e�hȏg��8f�m�%��W_��_��	�A3�t�3��*���-9q1�cd��]X����"�7�aѸ.�dA)�
��e� r�e76QC �3��O%m9��L뛠�S��ݟ�2�/ɿa@���N���� �h�%C��'�#��~�co��(��C�x8����4"��U$	D���Sf��0r�י�U�rYP��LpRA]��M^�~!��Q�x�m���Y����t�]~�\�5������-d��Wc�rψh|���� Pw�uY��kZ1�)J퐘g%iD�/��<+���y���T}���ӈ.�_��UUh@09C����D,��8�����A���e��I@爎�D�)0q�>qUs�'�j����%m���1�Y�j��w} ���TTč^-�@�nw���(�v��ӥ�&��B��N:�̾����j+%��i}{w٠�������ec�Ј؁匍�%�V�*,ATg��*��I����#�.�&����	 ��!ϟ�Q,Du+&����G�N&�%��':�>���m΃\W�!��x�OO1���"�ӹ �$F�L:d�6e�h�� ���7���`a�P�B)�uG?l���%e�)P�]�2�c6�!o&b)�>���@��j["K#�a�	�>R�2�C�;�����?ј YCk�c��;�/�����_
���3�)��Ӣ� &�@߭���U�[r���}��
���QvCPp������)��l���<�%
F�����\�hG7رĢ	+�������}�M̩3�`T2���#	�@�B�H�9���d���3�xE���T�ez;��!P����� L�*�vX��1+�j��ꍧ��F� ���6��iߦ��DC��Iu]�M��]BR�Lh���5*H6��u#"#�u2�2��kbքO��&����5�ܰ'�)�?���gT���!�l	��4�����D<=9L�����0�O <���FJ��Q������X.���	�O���-�'ױ*����y�n����F�-sl��<g�U��'f�?�\ss[���b��:�����e�#�T)R�G��{�Q��i���.B�~���fa�	�����y؋.U���'Q+t<!�bp"YG�a_���f�uy��r���i��G�K���{��������q�"��.���ST�2f�.�VϿf5e=���-��P�����L�f̺����ՙ�~�,&}��x!��	�Z��Q��%��	�� �I���6����sK�#��b��~r<QM�������_Pb�k7��m����_�U��/<I���a�Uݻ�z��Uʯ�'F�W�A�4Y��	��H-{��&�s-�F��9�#S���ņ�����\'�$���t��d�L���xY����G;w�_�Kd�b��^H�?8n���7��߃�Y.���>�.�ْ}����`�P�&�$&�C����3"���}�9L�s��M���V�?|�F7��[%l"�A�{�,=��6���7���F��9a���R,��z���s/��:��/RI�	y*0Z�ÔuM8w )M6��}w�[z�ܿt��Ε�C��` ��� UJ����Ѵ���_�6�'wp��(i�:L.W���Q�e{�cX[c��]�ָV��\�$1��!$��o�f'g8���P���&�Xu$���kW�`O�v�?=����{ fi�*a�m���=�]v���Fn�A=�yl�aWG)��·��~J����Wh���f���w���b����Q���Yqh�!��~���SPo�Ğ�Mh��绿�r�.6��H�w=��fU�����)�1v^�&�v�j�Ӗ�p-�9��Z�4��_��C�L��?���-�&y���^���9�"��AЇ���@tg��%)D��C1���?�l%o`E�8鏤�ݏ7!6�>��@	l�׹��^�A�����9�Y�Áނ�/��_\[􎥗~��J���"S{�[���s8�z�7Zk��Fv�]��H�jp���ș���+�s��� �:�����H������E	!/�D9q��XI�r:�YT`�s�p����V�~r_��n{�ì�B�*�k�+��y":���/�o-B%��Z���Ўs�Y/|���jW���h)�6ވJH�		G�wR��5�)@o]�i۠js0d���і4����{m�z욍i�x3�ߩ(<��C���'���#/|�a�2���A�z}�u��eP&��-�Z(���h��\B1~F���4��%�k�P��(F�?��@�.�XX]Z�噜��<�9��hճ�����E��e+"I-A�O��"���v�A���$*��E0 ��b%�)Ё�tG	��a�G8�6<H��͎�\h`���!5v�;�@�c��t�$�}���� �L�Qk�f����(��*��:�yv!7{k�p��T/���cXH�>����B�A�d],��1Rj�N�,azD������WN�7"��r��)�*�^x���-���Wb��Z��"��T2nd��<-�u!�.L�ة<�/�Qʴ���6��+5;�W��
{�5z��*�<xb��a%^���R5��ؚѓ� ґC�6��
�a^��%���cq
j�k�-Z�}`'[�Ê&tO��k|2�\���3sJ���������d��[�wnԒ�VR�5LDo���?����c��1����_�c�k���K���^�� �m囦��bȘ��)�%��.͔�����W:f��	XK�YQ�("M�pfmH�|I�ϓ_o/j������w@f=w�ǓDpk!�)�ޞ`�\�}ods��˵���D}��N��.�-����o{x��S>��Y�6Ǝ��Ӹ\
��pj�^[jK�&[���֔'w L&d�u�_�3�L����߬<]a�3�dR��嚨������d$n�������`�6�����3r���/�L��J.-j���5�"zL.��W4���cH;H$��M<�9+_s�Ͼ�b�8������Mn�f��
��,|9���?/:Q�`n[ӏ�Dݧ�6BN]2�|��ƽ�d�R�x���t�ӕ?3�����t�sI�U�;�â�d���<>?+��
5(�ּ;��~%-n̥<��pM(k,I5/n�[Uᶹ��$v��$��:�/�<-���6,\*�Ѽ8w���"	'������cu��*����sB�����!��C�q3/�Q�e	�~ܪgԮhd��<����7��],����]�h��9�>-hRK��1�>�a̻�[r"��%�u���2u��Ryo2��ױ�u{J�R疲�4���8T�QHEv����n&�Q[�ikK��W
���ѕX��BKu9���W�d4O���Kxt*�g��s>B��t��L�l��
��lЪh��
p�GLc.��=�	��>Ǎ���Hȓ�j1��� ��~�6�0T�^$��¯\���F�c�3��q�Q��")U����:_�o����AEfn;n�0J^U�[" �[Ts{�nWEKő=O�_Q l�Z�myZ��0<{W٠�4x6B�C�\�����~�iG�I�;IY�5_:.^�/��	�&��fJ�:KS��w�3D�"Or��v����)$}����<K���^\�K]k��>G��UZ�{_���E�r���^Upy&�@)!)Z v�O6��9Ԡ;�k/g��,sBZm�����c�Ph�_��z�S��V�-��uk���H?���\D��J[ɏ�8E� ���K�a��՟���d��ܻ@El�������%�<U�ւZ�u��p���I2� ��^���V<wCA7�>Ԍ�[
���R���< ��y���@.���pdrV����w��~;�>u�5e�~���:"�4=dPtH��4q~��>��F�(�2w���g�����~�k;�Q[��WMy���4lq�E�Lc˱�C��͹V-��-�m��K�?�e���l�j�-�KT4�"2�Q���Z��*x?'�+����� �ϱ�B���,+��(���36�����8&j��c�6�&K�m
��9���fՈ?w�\ac���S�SC��R1��z�v1����?@BG��d�dL�I�i^X:w�����xI����a01%�@߮��Q�����r#e�bۅ,�j+/�vOv��UR�YM,@�+��㫸��L*wu���Ss�:~=�q���u�Z�qL�������x<B�z��ҥ>�1����LY�MD�*�l�\�-6u�^4!�:�̅��'��%}3 ��+���-d�*
��n��T��|u�O0P>�fE~�ޢ��7S�mM��4u4�l�?�><)���F�p�]'0*����y*v�_<���,�m6���4�A�Ȑ[2���e"FK��B���;���!���zOH����K�׷������2�t��u'��+���I�	����Rw��77K%%�҄��m�o5%0
�_su�Xu#,J ���h=�aE]1�*
�:PU��������M�����yr�-c}Ҙ,�k��A��cłq�3�X�a�ySZ�10�9��^��`��{>����T�0x`3�!�wEr������K�=�'��·�R&�K�O���M,E�0��o�9-�:�kY.�$��0����18�**;oh�8����т�]�� M�ݓ�ך�T����`(��O��<��ψʓ�zW�븅3�o_ę�L3^��Q3��Y��%�o_���r[�B� wi�Q� ��/cz;�˫��%֭�;Gd�.�;���!\���B�#���P��&JfO�"���� 7�/&���Y�%�hqX.��0I��-��4�Y�3�f���	�E�5�逴r����M���j%��v�W�%��-~�ѶԱ܌#�����q�Z�	�j'R-��ȯ1�.�8\!�����%qZJh�Ӆ����b0�N����s$o�'�Df�\[؈N#��]+� �f�2�]�����䃵���T��e�톗�P��ϩ�)����I_Q��u��cj�ܟ]W�gm���yy��L�v � �&��a�*�7	�?�f�&_�%�v`��9G��gC����y�����.�Y����.L��k�2�~@������EϪ	�b�uAjZ
�RF���9K0ȷ1z2��a~e��L7�v�玥�@ѥQ�����u����q�%+��q�b��y���^j�h::�5S03�b>�7�L�K�������������]%;%�H!���+�E���0!��y�So�R����q�iF��?��=�N��qEKlG����=1,�
��{dA]�	�D�-o��C�d`L�E�xj�{XH��l��ҳ̙c3|E�S֚��U}��:pD�6f�'�l���c� �[���ŮsKaM�u��#Թ\�E�7���E">z�>����������P��kmv.$�]��BN����m&5�QO~_nuY����Q�XU���E(���� B>�E��4�X�A�C[��ZV�O��\ F}�V���;&{������IX�+�-X]����+�7l�n��������J��:8�מ,:t?�V�iNcy���@���H����B7+�w@���B����A����dٹ��������J!x��g�L����
�1�~A�ba�E2��$�Ji�<�-0E�/n$HP�mme���RȰ��B�9X,���ܦ��I�[L�gi$�$�+>�x?[8�}&�^fxf]��8x�g�����#�}�e���82�����PwT|�z�2��k@h��RX��wܐO����csU,9Y�GX���ca������|_��}?ڟ��"�\9�WN=�[��s��U\�l���-���%��p_���������z��ٔr��?	�Z�*�:GO��� ������������ٽz��-� �ڜ�J�2@�oG�j�	���#H^?0]�Ԇ)�GEX��,:�`87���Ӑql�r���� M��j4\'<97�Y��Fc�����P
5܀&P�,g����IR��o�.2�j�KC�vφ9���X�<X6�ǳ��Bb/�M�(-�m&ʖ�B�G^��D�e��CD���kٖP�)w�M�(�s�N�}|�J�!������B�y~ћ��/><�E1��t�՝�j������i���$ %�,/	�pt�؄�H!�iS-�S��I�� ���ފj�'(�s��6������ �Y�J�9ZQbI�}Y��K �'/Qn�ѹ_s�A��M��Eaʪ�M�${������S֟�ϯM�?��q9�n�{��\�=费y{hZ��r�Qie��_O7X��c!نs��;���s�4�P�_u���/�?�U��l<���,)��h�(� a��na�n�tE�;ʝ�����#e���j	ֈ��^_(���#5s�4�|�����^���|�!\�8cx�,:͜.2C�Z�o��X���[.Iʅ*��&��X'�d��I�D變Y{�S� �YZ���ғ�MF���1������;'zB�(Z�y��'%1�|�cN_mB�o;�MXs"YV� t�����.�)H&�#2PQN3���5��j5)���C�*�9f,�[���Kٟ�u?^&��Q��]?��Q��d������J
��ڎ����gG��pّ|j��C����>1����L;4�W���@��ꏁ���7?]{�B11s�%a��JX��8���;��?��3רY�"��,R��|�
҆��+a+�M"�m��*B� �{%^s��@�D3�1�rjGEY6��F��v#���AgZ{o�c!d5<�_�iw15G�����Uyߋ:���������O���E_7�T��hj��1��ˮ��1=�(#�E�|-Z�Tc���	�M��>̢[T��Ƴ�6�����~e���B(!
(����i�Bְ]:Fp��Jx�������NǗr��)k�������*7���lɦT������
ߣk��`��靦br�$��*y���j�IV!��3%�n$>�l�}��cA�Q�A��<��k�q�Z��d��0�3o���A1>�t�3$D����m:J<����O}1G;�F#���tN�r&8��D��Zv�9PmY1Z��un���;�l
θ�����My�����P����a��� ��z-�gnun�� Y�1,��O��p��[�n ���
PH�b��veػ]�@���>m��Sw?�ɍ�v+�X����&DA:`����AaW~���?��u���lxdsc�s�+%4d R�v�x=/�w� ���౅�E+�`�fR�J���4qק���F���=�c5dU�=��`�=uQ��|&���&\����R<�&�N�TEW�>�$�bT�)=K��,_r�p���.�.��8�ۨ7��Y��:ʛE���qMX�?�Ț����*��R�,F���B���|���/�^�qg�4�i
��,*��F�tE�M�r�)�S5��Q%�vCM��n��M^byo���s�n%w���S �� l��DP����C�=c3�;Y�����p�)B <z`I�j�|���
�����̂�zU��쯡�[NL�cb'O�#J�KU�����YΧ�o��1���r�n��+�i;�2,��:�3wXu�����h�l��1v�}�L6]���ujC��M�/������	���>@`��k�mAQ���|���pvn�
�`<���k�w5Ek2�����s ]?Ȑ �k��Bý�sУ� �`Ib�:�G�>ܨ����(�D�cf<7�n]�~>�Fy\�t�;w[�|*6��R���R4y���s9y����7q���BN!��U�n5\��E�������f�迵'�֖h��X&Üz�?(n���1�[
ֿGV'��E%�$��P���Bӌ ~fuNA�;�s�,T�����#��h@�\�U$ـ}���÷�A��䤀&�,�
iF$��z �HZ׊t��G�}��JM�v!$�Ia��I[����t+��ګKu���j�:��d�����.�����Y�o/�FI�9�p;I�pc�
�:��� /6��^^r)"�xJ��2�# .���6b�i1��,�ʠ3sb�E�9��-��Ds̽`+*V�y�[��z�tX����B��$�-�߆Y���՝��ݒ��G��	'tL�����B�t�3��I��8!n��� �q�ږ�+R���� H�u?�6tD��R��h��)�.���N�~o�N~�M_Eg`�L]ۆJ����x�/�}o����uPl� �K����S@hoj�?$�M���/܂̼�B��6�z�a�h�������`��z|�!�j�N}��X�^�ʿ~Ml��*|�����SJ�v�X���,�d}b�����L��5�r���$�"+׸]��t����BQ�����o��W�un �}Ǝ�H��.���a�/�bl��;��C>,�A�I��Kׯe1�v�Q��[�@Ns.0�Ac0NK��m��\�L/��\s?�A�e����c��*Y4�~
?��i](����w�|Ⱥq�G?�A���-��Q����+���su�7N /vh �;KG&�0L}k��2 �Rz�7����-;OH��Y�D���o=0;�P�5�Cݜ	\��_�e��(3�=߾�u��F���C��
�)���x9}8�y�:��������DS2v1�:�g	�;�cݖu����cZ�8-�3�Io�2|����Z��Z�?��'���&Aw�G(*"[��e���'3Jn��/FSd�~$'���t�Z�Yr۾��n���%��; ��ʜ��r�ڻ�6�.ҜV��ED� &҇��	��Al.1�zS#�M���]o��gI��Q���\���us�V��~=����|�Q
�����eө#>�������7k��}���Y��	B�|�4kV(s�w�"��[d�Kd* �ӹv\���(�b{4��7�s��{�N(m!��/�y�q}'`���F0�!��1DF��5���	�wU#A��Zu>:�����(-h���)��N��9�tnU�d�O]��ՙ� ����پ(�s֮	d�U�`�0#g�
�Х6�Y�M���|o�d��p��,+S<`�~���s.��B�gZX�S�5�,ѧ��tY [�E�c��^��iֈ�a��c�=T/�%���=�w׍Ղ`D ��f�[T���0�i0b��,�2���>|�;r���3�>�j��`�?A�`����{�+�6~���R2���0���T�m��P�iq��m�T�F�4@�v��n����U����Uo���&i)� !�NU��v���p�ݍ�ۜa爛D1^���KZ���JWvP+��o����̓�(���z����ɿ��Փ�K�_���m���a��)T@�X9�2s���ˮ.,���ߵ���[��4���0�zcu`u���h_ek9n( �<�۰���e��,㠯T�M#��.^F߳��{ v�BE4��z�5�����J$�l?��v9�����ǛP@� ���%��1��_�T���>׆9�R߆���+'9��Gd���v���S��ޑ��Ȫ�mo7��ehΈ>�cd�����7�P�`a�l�ZQ��+H@S���C>T�f��#���C���x��(��2�P}��?u�\�\���[�xb�q�]JX�ZK	t6�H�{���9��R�e�T����v���x4l*f�k���	���� G�ON6�
��$.�7d�S����E�R�Fb0*�)P��Y���Y�䙹8�7-*⏲���˴T��=E^�1�
\!(�&!*~9��F%f�
?&��(�U�	(k��{
�h*�^� �MOg4��so陓4�=J��ɳ�}���뼁<�}��"�"�>S�WQ6ټ2hCy:F�\���BX>�{��pǏc��J�_O@����|���<�M��G��372�������;�4g5�%���1���Q�Ny�R]_��@IK��iG��X��}_1�|�����*e��Rö��?��.�ԣ2.�Ȳ�����e �������`l�ïK�=Tj�Az�m�~�����uR1O�v�眰�gd=W�O���ʜ!���trE�X8%"��ңE�5x�d�{�O���Uet��2B����N.л�V�G2^��=�Z<���)ZI��'�	-�e8�J�gҏiJͺ�l��&��<$R��ú�-���
�!Y}�C�כ�?��ݺ���O��i���/�
��t��������	��Ȉ2�@Vv�Pi\���[�x6ůQ'N �����|<g�ˬ�!DX�NGëQ��A��L��J�LlI��6\Ǐ��/C��)������LA�L|�xV��rN+��ڠ�Xj_��d>���+�eh�N���U(Qj��y��@0ݬ��/��	4P�u��� ��|��z0N.)�2�P*>�C�'7ë��ζQt܄��6.�����(O:�S��Clm�^��XCo��iF���@�W��Bk�}�Kލg�]1��y��Vv?i�dwc�����l�(բ��?��% 6�[��>�c<rG%�r�c�ՐuƦC��)K��cA�Z��h���s�'��c��V4y9�Y�I'�}��Y��2��'�V�L���p�Ys�N�S"�r�ϗH��{�8���v����S�~8mO+�Odw_d����6�
�'W�2^�p\���G�fXe�1�"l(�ȧ�J��絶���
����`��]x��c$]��%�oA96���#�)i-@x/"wk9~�L{�=c9�s��3���#a�� ����a�������Z"f��x�ٓ�׬��TǵcW!��yo}\��D)��E�nB4[!W<{�