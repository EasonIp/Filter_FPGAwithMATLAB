��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$������N�r��� ��Lj�cj�3	0�s�7��DM5�ڗ���Ƕw_��w����1����5i=r����$VfEp��5�y/�䰉t�R�b��=�T�F� ����i�+��E3�-����mWp=���T�+�ǒ����gy��\�>/z�Xr8�j�S��G��rˏ>��7��,�E���.�3�b{(�.�t��-�c?����x�uġ�9O�]mb��O����ݨ_��;��`����%�}���+J� (9H�M���.9<g<R��������Vu��!�&�2�e"?~T;�+��UyP�ݢ�#�&�t`����ͭ&Z�'{�n�hO����wT)�i����i�_\J /�p�;߀%O���^����� ��6?~��A���6��?�0r�K��Fg����A�s�DeS���KZ����o��j��v��=��ğ�{�C-pL�����)Ꮄs��R#Cc���n�Һ����Ȟ�ƅ��9�
Ti�U�2ꪨ-J�����n�:K��\��Lq�@,�!�rI�fmz�k��6�w�[u$��3�b��yz�b�)�I�+c�Q�����_�`n�	�~w�Ɯ�z{��i���5�`}�(N5�~�Y��*?<�Hy�秞��zi��q/j$�D��W>����՘Q���&�Ma�9�!�C�a�������FA�h �y�R]����n����g�H�jy��m_���k��}���&�F.&�:3���Q�%��. q�m�1\pj��ٓ��w�*�z���PGwz�׬�>d�.!�~P�Hdr��yW��1�v�ѹ�4��
Am6��j����27�]=�[q�������(�l���Z���⁽�϶���}Ⱦ���$;U�����
O�`)f	eK����D.r�z�ל������t@�6�$p15@iNL|j�5(y(k佻��� kg�%~����0�^��o�e�P���cy�RK+��R!�?U�x',�I��cV��ɠ��1ę���~9+����}�j~��s�csO���o��z@��;ֆ���=�c�L�t;�b���0�vl
v(�2^��}��vu*����/���t��S�P�)0%z8P�@�T1�I�Z�m2hإ��eu�_k�F�u\E�W�q�iO���F
�AN�ω�o-���K���;�f����{9�r^�{���7�E��� �yP,k1o���hEL���rȚ,\�J���O�2����D�m�����X���U[��eʁ-|����>#���mG��@Y�<�K��j{�)�t�'wuS��`6e�G0Z`ip�:�̒��	��Hi�����R��2�YhT!Q1��`�u�I�:�zl�c��׾/��^�6�,DZ/�sp����j?�9�������6J�=��.z��� I[�r�i܀=UEV���e!��IC:�i�mk^"�M��)I|�#O���}f��6����І��9�n
����R[np�5�蜸������D�u�c���N�í�Q7<?i��W�~�o�J���?y��=�<[�VV#��T;O&g�U׌S!￨hcO�>�h�ӻ�X�6�&CJ�ރ�-5�0�Z͂���dH�7�BÑ(�<��)�s�|�Յ��(p(�`�w�{��Ҽ�Pަo�T/���1`o�O����Z�䂞��N;z�4�M�h[���$�\�gCr3G\Y�Z�0x%	���%�X������؛�^o�[R}��s���;;/>��&�
Ln9�T��sq�IQ�}B���?ߵ8�&�E��&���ËϾWj�B�f��Qݡ�O�)/��y��	x�n��2ܦ�s���,~�3�d@�g�˰��lPh# qd/���/�>8uֶ���L��Nuw��:T�'*�{;��9�������M��N�`N�`�x����^�߸'�XdwcGd�/�OvM!�%.�a�I�.�}<��"�.1O�Rs�.�I=��q�5r���JG��L@s���>�%�tN_KE�Q�i���Y �Dy���;V�d��#l�ٚ�����A�ۗp�Ca���Y�0���t��h2�1 c!�h}<$��7��[�X��3����/}���Y��Pa��.x���h���`jb����DI��(Ƨ¢LI�vس<���x[�'��ٵ&��z2����ʹ��*O�ɦ��<s��W�v��t��1��$EjeD�Ҩ���k�'RN�y�e�"��r���6����#�_�vך��P�lLԧ�z�(�v�#�����(b
"A?i�qj�r�<�b�SA�T��J�t[rщ�'K.Ȏ�r�~�����q���׳kY��GA�lp��?S����C�Wq"��{�5�y�c;��>���>^M�m�=X�sS�E�_�s���I���K���Ɓ�pCŸ�U���bP�bDOg�Ҳ�����8�b��t P��{"��Y,��v�%I�hw!�6x�M��j�H��>�}+v�z�������'_j�e8�ў��d�xz�xl���{������[�[�>Z̀دbn�U&km��,0Vi�n�B��P�������z،��`�"R�E�Աgq`n~-N��Ec���f_�����gר׹p��.}�doᇶzH�&j�[��Y초i����l��G�г���ZV"|_met ����d}E?n�+���W��	8CK>�tG8�V.�n��W����O�"�,��J?!{=ےD�U ��Y	����>|8���E ���c&J�3rO6�U	���m�P������&�g�)��&��l�A����q�#�S��z;�]�°�n\2m%����­��'7bvIA?UR������n(3���m�E�t�f��#,/|�����ɋ��ZSP���61�ƈk�4�C#T�Y��$J���Gbj�*6�ю���]���d_;Q�������.���d+�@֯�{��S>�������~��[���>,�_V��C���4E��F6���9'��&M��$BQ��<��%�>��ԛ)q��G +X�
�w�d0:y!O;sg����3W/�ÈQR��LH�ZB(K[$���ƭ���MZ����0����ab~�d���t����R~(��ę�,�Yr� xfj�� �~Om��==�%�JS�tRQ�2��?�f��w^��%N�B�W5�%�^�{�P�
��5�]�� Osd��� �:b�F��^u���VJo�qsJ1Y�T�4��6s�EK�M�Ph�?H��:�.�����TKFM���ǒr�Z���cۖ���1yW:0&�7�x5����v�:6J���� l_��HA#g�d���0JV��媜�j*1ԇ�"w矪	���?�!q{�)7<��m3-lf��4�NGS�$XڴbF�NCH\.��gQ���TYP �n������SI��Os��7&�/I9Q��hb�f�sr�g���u�.s��
�㞜 �tZ���/��=S����	�M�L�,�iw�6]���ڈ" ʘ�	�S|�ob�`�jlj˚W���r1WYyF	k;��P!��x����@>>��^�@bR}���`�!���5D|�͜�3��m 6u�*����s�ok>�<}�Gy�������%0zE1+#�&��+Gb�Sl�OMH�)oK�%���:���aʐ� U2?�/e%*�Xc�gi���N��J-�{b��h_ �m��X������<䢶E�Z�� <������s�%���\<�f����)<w�Y�ak�X��r+�b�j�a����N�L6
�r��֞E&K�9��O�J_\�+OI��0��n��Uh=MC��k^l|��כ
��>��ʊ�c���6��W?�4�a���g_�����d��
	�����ǰ&Z%�y��N�i!���S��MF�JV�G�>\2h!R��1��g+Y ��d����-��0��(*�j��Ԡ�d�A�_��J2Q��#�����8ĽG���l�ݥʱ����l�,w���8=�o�ӣKwh����US�ݭ����Ԙ�m�⋘��R��<U�Ǳ���(����E��y����4��H�x�+�[A�h�T(������'f�g�^��}����W�&S���	f��&R	L�`i��:�:�"mx�Y�/�w��]Bz_ϱ�����W�k�%c�t�o%I,��g/?���EN��A>��Ў�q0<��Xn��M�6��u6�Eޔ}�ϵ�c%r�N�������%�T�yk�<�R�����V�H�O�%���ڍ����+h^I�i���73=��K�����BV[#�j9���n��\�Nڴw�j�ؗae$lE/��
ʴf#�0kSZ�k������ib=�̋,$gG	Mr�<��"4ʕ�(5��7�� ��}nr�u2�h��*�8 �����m%��*W��QC�1N�`�5���r ���ޟ����Q�Kh)`�iOx��%'S�i*�H�����w�͋�{1��[9��K��x�q�����q��^��]��k����(���>L�Κ�؁�F)���M������Q�)Izd-4�mR��;�/�:!-��<Y����|QrDǁ�h����$�iO�5��6.�(����?}���@�w��8��j ���Z��}�S4�@�q2����[�Z��+u�iS�5���+����Oi�O|
����� ��=:���q�`���P���������/���+�G*�M�Q]�������<���	qUP2l�N'z�������Q�9�@�E;�֍z܄2a���k�Is�oVh#���{�n��M�����Y�
"�Π��)Ӧ�_%����1���P���!�C7�C��D�g����Ƒ��;��os-�.a�odc�P�.�S��I Jy���h�HX�l�G��{1;��9��o3��لcJ�zEچ-�~Ifu+!I��^]�&�v��t���9�(��8�N�,C��ɭ[�����ujJZP��Ei�*d�0.|�MC�2z	����;1����ΛƬ���m2��s��Ŏ�o�䮃��k�v��ߖ�0B��*�p!�]���i��u���dņ��t�����fӛ���~�~*��g`�pCT2�U��5W���
�ɺ�t{�~|qX�i�	��J�+�K$\P��]�Z:���{�E��X+�($� aa��۔�bcdb~�ك�g��w���5�ud�����g%��Vt�^�E�B�[W�=�un_��'��)\�b�C��*�R���h2w��+a>9n��� n�P�
E�Ƒ������ݬ 0�uȅ�W%��I��+��N��[�+�C�<�j�^jZ�P�(�a���p 8]�m��R.�>��1�z��'Q��U�V�3�u�C����IO�R�;����k)��'9^T[�?2Өc0%�B^0dx�~�$��\�\v����۾R~b����V+�����0b�G�R}�F
�^]����¹����]��N4��J�(m����&K��x[�(�-^�S󱝸-H�|XT7N�/�v�R�^�9���`-�j*HQ��^g>�D�D/�V�@Wt�5�����*��|)��x7�,�ڄ�/�����
zzZ�Fa����~ȳӐ��O.�������	�Q8ۡ��b&KXǛuvK���v>7"���	�bx�����,+�.�\�o�WB�d^�-�)��� 0f ���X�$�;�.q�],���g��]P�H`��5Rbu�.R�磉C$���9�r-2������p*�:FgTn�ӛacҵ{�%��nO�� �1�v��V�SS ���w���-�4Ė�����2)�{X���yb̂;���xz'���� ϲ��ה�(1�"F��g��@�j���GӒ�V�	���,y�
zS����)p�ʟ��_d`q�vD��ͩȓ�,MO�]�npʦ�Pdʚ!�,�-6 ,%����U��h��y
�xL���bzR*|��Y����1���b�SA���p/U��II4�?��Ewv�<8[�n��;�����a�Z��?o	�ն���9f�pW�QD�+���Ɛ��R�z	�:m��4a�/b�@�2�Z�GJj�M_���s`�Lrv��Yط&����#����ؽ��d��$Ys\0D��d��_�{��6@��4^�
�_�_tNR��Ⱥ�1b���w0`
�e���ā^o�'�+A͈�-�W�|"�q��+f˟���1P�_\��4�cQ��"�Ǡ������֨���N!��Wϭ);3Ŭӊ�{P	�n�;_��+��)��3�_ۑw�L�V��cԝ�Ia�7Q��e���~�E�O$�� �U@��ZG�Z��e6�}���g�� �t����z0�*���:/������&ek����~���KY�+Q"f�ܴ.�Ʉcԝ�� �[�����C,iGN����mӊXQ3` �[��t��8k��,�<��/�Uه�z�ҝET����1#v��Y�9�N����]��Cgr�iD������}�-�aV�=�{�JOn�-w~���I��YB�}Y����8YPq����۾V�EB�OːB\C/<n����R�7䬵MGvT�V�;^|���O	s��\���La��%[���l����U��iH(/�ZTNcV\�*�-�h�e�������Rũ��	�g� 4�P/W$��͌I��M�-~��b}�����bE#*���	r �OՒ��������8|x�`!�ܷ�~u���>p����R�3�ݤ�3-\R��=	�T�4�❛/����c��K,ָ�`#EO�a����h@�}.���9hl34�iA��r����?������@싩��v�&���i�RԿsNI)*��z����'v���=�����7��w�Ԙ����}��ԾУ��L��l��<̘|��%6Qٍa��|��G;�y�AX^q�wz�d�^�cˆ��i�W���_��I�!�p��{�{��`g~��B�0
���r������`6K�#@ދd��E XP�.�KU�˯0wQpO~F��h v����k�d���y-�}��A�h��z��R�ǜ�o�!u��C�!t�Esv���a�l�L�/n��fNᕳ���_p��_�����`<
�Y���tg��!����Q�^�zu�8��ts6F��E-��}+�+��a��[fç��]"���~�&ÓIZ�`ZFF��'�cȈ|-��m1T�f�(��ӺwE���տ\�Wo��|��o��a�Q-Ƙ�ៀM�֗�E0�T}�+eW�m��Pk��Ƭ�����Z\w�i�њ[��F�/)��_UZ��M�"E-�/�]eX�(/�
�S?|��X���O���9��A`�#χι۟��A��`�C��?�0@5j�ϾC,%���ܓ�{VA����=C���Dz;b*(�����"�޺�U���P䕆���)Lb�M�W �g���H1�L��b1�L�]�#�-<J�]H.�`�@v�V�v��-���2������-A��L�7��P��Eb$�ܡm��e�U��_J�1�o�7��|�nʭ�?����c�u<7F6E��,ݢ�����R����`w4�j�p�<����b�*��i+�3�d���?����|=��J�&��Cu�LQ�4)֒����a�<�@+�`���n�ojXr�w�/�ټ�����1��蜽C�5T�N�do�̑p�ϖ�5��q� ��ǽ��	\o��[�c��c`��lD�~SGx[�й_�(�޻���wQ���΅R�;-���-�Aw��U��ݞӾ%Y��iɛwU]/_s��5*����|�+�1&����Jѭv�o��]�B^�4�����ή�i]�Ia@6����Ꮷ��D��*ԇ��_���QK�q!�k1�C&6�/(�{_�'� ���