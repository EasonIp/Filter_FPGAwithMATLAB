��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|p�n�U�_�e أ�w�T�)Ѡ$M��_�ES�3�� �����æ��c�5c��cc��N5��d��L\�b���{
��v�0	�ݫ�*��HgZ���B޿B��������X*�;3����Tsʠ���`�ߞ)X�d�O� -q�%	Ѓq،��#�0�$ˤF�Ԃ
�����!;��)O6ǻ���ā*�S��Wo�HD"K���(�x�֜0�N*)�L��
�4��b�����iW�*w_�ƣ=���r�ɦ;�tLcű�2(uS�Jm������m���ѿ�k��fv����.���ͯ�
o�i�j
�0C�:��/E��[�3��	�m��:�&w�ń�GXЛn��&P��j������Cש��R^>��I�Z)
)�j���6�o`��J7���J�����0�,"9��(�A6��̪l�u�8�J��ܻB�&����%��c3������nՉLH
�._�:�� i]�F�eVujL�hb_��M�zf<F�P��G9�;/ c1bV"�m�c
7��U�;ُ��r�顐�D��ۼn.�k��¥��nF�x2�W���1Wy'���SF�8.���T����O�Z�2^��M���(y���/�7�l8=��z��~�F���:1��\R�v��6o1�0�@?=���>̰���G�`\�;ո���3K<�E~d�n���5m-�{�߄HA����`�I%����G�^9�#Z��f� �o�Ie�`���ȿ_�����mj�.Z�ywd��챷����5l"��niZ3S��t��1]�\��".5�	`H隙\�t�y���� '��_b�y�q��`=��׎R�^�Yb��b��E�B5�������31�[y�+�2���l�Y^������S�����vg�� ���I92�M�b��0��-�J���?,��f��, "�-��tk$�A��d��2/�uLلVie�q��J���H\Q��,�ҟ[q��#�[�`؝��؄�Yd�����a�^�i�
���'�"#��v:/8�� gz���mIn��Dǫ�n�Ѳ$[T�.\��|dO��MmH5^��6����	��0eT�d�F����o<��a����U��NNc0���jB5��s��C�~�=6���Ȏ��MX��se���*RH�ڭ��f�u���UȪ��e����=B���n��g~����_'+0�1��@{Ql_-&BZ�6�l�ݠ�R;_�%1V.��m���N�����͆�P��&�s�55r=��<����9��D�֩��^Uv�.�����`V�h��֌g�{3��博��J�I�#)�����.���g���/��/i���|m"��W��8�Q܏� ��t�-����B�QӘBޞ̔D`�pq�Y���羼�me����P��0�y��P�H<!�o<��)7�'us̥V��z�q����>���	C鵥���U���=��Y�e0?Y���u#4��1�~�İl)0�X��o!�6�+�ԵP�Jr{�be��rA7#'M����y�x�)-j<b�BkO���K/6��Dn<�E��
�àœ�T+�}X?-��.$��)��PfteO*~� ���]��]c��U��:�=�g���/TƩ_�����:�u�	�@����&�W`+x �=����;k;��w����u�b��S �%�o~����68p�� �+��>g����'��/�V��F�%W~(:�V��'���V����tuV%M-�S(X��@II&tb�ݞ��^.�÷�դWd���#��j��R�?s�]�/UT4���]��F0ty�����'��o̴Wog����lq��v�C�P(����G�{ɚ�X3L�Zօ'��5������\�.>����٬�JҴ�.h�s������R	1�%��0���*���AQ���ɀ�0j^*`(a����p1��D%;�����Vaެ>VXϼ"�����V�zO~���!�7�<�k�e�co��❄�'�4�(2��A�#�DbmKCc��o�|C9=�U>Z�n���?����%㥬�;�*N����99�cؕ9h;��a�)��H��?�R��/*8:�:%��a���ai��I���ǭ7��^�Z%�&Eh���!���t�5�b� 5���
��L��u�d���Te��:f,�n6��a&{����Z��
�~Td�ˡ��A�א��N�?��hm�P�2�B _0�X�U{uF�HD�rS��7vn���=����K��@���V�����E�j��O�[v[�Eh�4����	'�5qȟ.�z�GSqp&<��S�>b�t�����i�����#H�9v�����v=�&�/�.��U���b���qU?�������[}�u�d��Q�P���b�ޒp��/B/!̥�����7��.�������U]�LK��ߔDŢI*/���H�ظ�	�s
w���
�L�yUP��6�������[�5Y��"eԨ��Bk�m$_�2"�*�y�_n�q^O1n�<#����w֢�/'�z{g0���X[)�0�y��cӉ;�3�Z����/�٢�:��(uJ���N4?��\�D�e�7�M�Q�̚����fv�n��!~%�o�P�Zɍ����,��a���f<:_32(���jcl����8�Y���	(q#���6��ׄ���,E*�U5Y����|�{�����<| "��"�g-)?�j��6�c�Ye4���(]�-F��)9]Ř�p�|��􈾵M��2�:=�g�Ҽ�'�������&�N��y�FG]kM�f��-���x�.����â��\2i�o~��ƬBk\��l�9 �7���VN�W;�``nc�@�4X!�q%�i�Xc�/t�Y��z�J�#rx��K͉��L�N�)!m�c`�dli%�/J)ց���k�Hj%d˰F? p!p�S�v5<ާ�	`�����o~t�L4����6��e_��gv��-�jb��?7	���m�jۙf�qM����
��no��C��aμ�հ�?����O�n_�ܾ���=���K�d>N�WQ�KYN����+A�5��K�w��Nݑe�H�oC�L<h�Er�[{�c�������2
+�[�0�5�K0��5���xD���2/.Q@6�Q�9c���IV\�i�'y�����n����`?���N$
����_�rU��� �˴]I>w�U��^��,�e��)~�J�|v�4� �|�����[���3��FW��*d5�6JW�����A������8���8vB����x���G��\��Mc!L0��(��6^@-��������L��+�,��������:._�(W��Յ����t����!�K�x��j�D���ݹ�]6�vC@j��c���G���z��j�g��r�Y�u8l?N����]��My�����~ۏ�VH#%�ؠ���ft-�W8��2�x�{X�8R!l�R������5I�߶��ɵh�S�=˴�OI�+��ƥ̮+��Yd�C�!jvޥ/��Y̢7�n/cU�p��ʀ�#T�v���v�܏���?a�
����AD�g��i^o����R?�V�x�G\�:񮯦��Qm�QFGX@.�謉g�G2��(�U��}k������^�`U��u�e�j{�	�e����-/ܲ&7��Co�6���������L`*�	Z���?Wb�9�pY�������vF\�������z�e�{�*s���%1��ȿLb+L�3�mF����
 ���:1RoJ�E��J�[���$r8e)ms]5ቿ�#����U�t�4�	����Ғ &W�qL�̾��zG�M����IU}n)L�h:�D���/�p-P#?$e�	iJ �濵鮥Vl�� ��vExW����t�uK��"S�Ź�����F��E2}�`�*b�(V`���u���Y:�p�ސ�o&���󓎳�я�N6�]3y�m����X��$&�(�b���(����=a������1rBB�b�+��P���a�aeN�^U�p"vJ��޽C��l��N��"���r����ڧ��]i�Y:Fz����{Ut�a�x��w�����ps��+����[�MS(��)���,aL�����Y����U��4���=L;~M���L�����Á7�R�'6�)Zj�����U�_����d��I�y�B��1��H{�Z�o ��|�gU�i/!��7�1�+�͍��KS��0��2S\����Y�m�S#���������,�NY3����`Qx*sW�D$��H"WwU!Ǘ���3�o4^�^f��9�_�Hd��T�ҹ�����^��*č����l��R��=��	��C7����}�؏f��Y��z#X��5�E������@R�r��mE�$4��ٗJ%VؔrS�w"V�,�{>�焕4T�}h\�P3�&�6��9le9߸�gt���Ü௖�=t` �E
5Ó����V�� ��P��J�2I�;[�Fs�Hp��ڊ�|f��U�pi0��H�H{d@{!�ݶ���숚Uds�C<z�[Э5�mf��*����gOZ4�k��͓N�5&d�3c�:�wj^��9���8 �p3���+�r��#��龴Eh7��
;���8�K�A�;�3I��|ɿ�z��|�:�KDeBs�G8�}~�$�8�FF/�a"��L"�@	7�:�����3��3	�Q�����Z�2z��ţ�ӮC�{�~fs%CAp3�o@۷,�s�{T��a3d��rp���=���ƣ���z���Bg��Z�?jCx|��F8���m��/F�8��=��z]蕘م�T�x�h�(�A2���c�EPX�F� ��Y�#Ϛ0�g�s6Lu}k�ܼ%T]� � k���n#��1���>�@�	[�� }���}�_�^,R�Z\����~h3I�{Rџ=�-l�L؉�}pN�fOW ;:�o��^a^�l���K��׿C�6W֌"�[:�U}؆�N���݋�o��!��p��.��B����(@��tt�-�?$��R\�*ߐɌ�!� åq��7!U�x��,%P���J�m���]�:�y;�aJ������E� 5��Yq~<���;�M�XF7B���py?XD��[�YU��'�E{��vs��ڧPgF)UFg�9L;���ł�Tv�ld&��GG�g.�P�g��a�������1�#Pջ��`�՟u� .K/"����-=�)y����7tx��tz�"i����{̭ԙ[Ə?*�<嗤\L���NI<x���������-	�Ej�,P�_XOc�8J�c�@�QT|t�4��R��a��>���D�
���m9k�xM��R62�~��nX�V!O���Jdx��&�qF"�cb�&�T={(*]��v���3e���g��/7�}|�8س�?����H��"!�L��H���#��˯�9�>���Λ[���'*b�tG'y��?9ӳ�i���C�y�s��ߒ���04H ˅.YXée�����q{r<B���H��7x����֢���}ڇ�}� �B��R�i�&Y7B9�_.�����l�=a ��4����:<>M�؅���ߓ��_��}�W�I�n޳GI]Z��q�����I[�*Y�����N\u�����qh����9�I��2�>����CI�lN�Z�ް�vhؔg���Wc/�E�� }w�K-�B𝲻Ors�
�@.r���I�,��a�����G�0Nv�FJv���E�.^n;�� ��¶o��*s��sx���µƋ+^T� ф��5�Y�e5S�"�v�
 �A�_�$Z�DEwF20�z�C�;��,�Db�S�q����&A_n�݅�%T(he���Uan�@��p\A4R���ȋ�,�#羵�K9$g�5�J:���3��v=02��L"l���-�#)m�-���?��eu��B��yA�l���s����խK�L&�_B�GO>�	�������@!�z�$͕�i�eD��@}�;��Fz㴣��!�}*K�pe4�C�i��=�:\X=�������c��R#Q�3��6X�Ys6�y)�|!$�|��x����$���&V��dtb?�w�CDo�P��1h�
� @i"����xGJ��v6�u����~6o���1�5"����	�����P�ʌZ�g���r�E,$�}��>�9�������������@=�K�g���#�C^���SL�xQ���t�Hw�������%�`� .�~]H4�5��4h_̠��6� o��1Ʈ	�`�W0���y{��D�+80�A�#��MƑ<Þ���HB�fd�.�I:A����XZ�_�Ʉ�r�e��$D����o�c����L���
�W�{�矁1�@3=��F�}1�g(�2ٴ�Y�A�S�8>:��,�}���ń)=	&~)�m�b�ڂ�Hf���S�߰�rqx�b�/I�G��	ˇ���I��'Op�� u�n���Z�1��t9�S�w9�՚,��־���ȉ���������"�1kbm�R�Y�}�Kҥ��U�W4=z;�>�L�S[���Mg�[��U)��cE��2���{3�K���j��-�@/���lgj�Q���L"ؽ���!m�����>'�g���B���by���`[�RW��`QeYM�H�[kk'r��'�'�V�6�����iu[�V�Ca:dv\���a-m�݌,$KC��z̬�{l���hM�\��*��o/�;x]�c�W�n�iA��|cP��(bW���ṙ<�������X��-�M����["	��Y沨⠙ʷ),ڟ�N�c��i\2�"��`�E��U���tx�c\�����f���d+KGqzxe�߿�<��M�i���θ%��bD�<;P;?sJ��7�}�A����gfT*{�}���ivH񐄦�+�@�qc��E,���l{���4.)����ݽ�����
��λe8*K�ѣ�j8�nO���E�������
�� ƹ�k���Rb ��	��2��R��D6֎��5���W���H����!�mM#�W>Y_����J��g?/��K�ܒw�-c��`�v��윤-M�!Հa���.���u��'��q�K�G95�XS��@yy�ӊd��!��q���$��e����:�H8����7\��q�/3��7�7��}��bm����,�����/8l�ɖ�HQ?G�Eۉ���P���r\0R�q�IX�a��DQ5�������IF|���K&�m������ӵ���ި�F���$r�Z�K�8A���x����>ƀ�F�ǈ(�뗜rMLIM'Ă�pį�2K&�G^�gi���W0{��y1j� ϼ�&��k�}�L��c�<c��W`��a*�Q1����'Ip���w�bn~�
�{�5O��@]�hP�)v��ϺIU-Ř<�䭄��ڏ���"B����_T@��0�����j��{|������a��z	�Y/[���O�-D'�$Ӿ��*4��;�*V�9Gxc���jE�rU	�y+=�X���s�2�u�ش��>�hF���Բs!�S+��Tz��w��9��54V�p ��ý�2f�����)S�JB��ĲK���#[_�=����� v?4%�j�=�I��k���~z���Y�hЛ�r�ć����N��s�����`�#\Y��BGZN�{�#ڬ,I(4Mn����I�5�����Fc��u\��s�l:ܖ���&v"A�"ms�>��G�����"�[w�AEF�y+S�����=�;?�����cl�)�_��!�{\+���E����γ��<xv�{��%��V����.i<��A��ųX�r��2-ؿ|9�E4�Z֢1>�tj(_ίz��fi#�9�{����>��0L<J�W����,d�9�Ӧ�N��$��*�ؖ���n�3Tۋ�2�g_Z��H���[��#��������~W�
���!���X�æV���^([ħs�]�땘��Nj6�N��ʕ\3��?B��:e�sr-��>8>L�
N����"��N1�~8͝�nHD@\�L[�/�a���|>��~w(�:J��~)H��`�a�ED|�#Lj$��'�}3���h��Vf����H�6G�,�[W�6��"^������2�&���`�eŒ�0(�E;�)	�❺���<u��; @��nioj�����Plz+C9R|Qy�q����\d�/���wݗq��a�3�Ҹ��}QG�M��D��ʑ[w���0M+�2�8��6�=���\��m�r0�a�]*��{��޾:��y)�͠�G�����ҵ����L�GXHH���u�P��gi�&&�5�mY2U�W�MQ�$���5�|аM��J*	��ݲ�!�s�Nd� �����eq���<ᢾҪg��Y�@t�W�O4��1��n���rg���淸���v�f
U�"r�Vu�? ̈́�Nl��ak�çt�M���{E����s�����-�d5ۨ�~VLۄ`�=�SO�ce3�ᾋw�X�,��5���<��OM=�u��}�إ$��LٌԖ���|<Fb�t@D�����6f3��z���5��NtE �, *FL�,��6E6����e;���=�4�N��ٙt?@��"�Ԭz��H��XS4e�L��I�ͩ��6z؅<t���&(��W��ff���
�5��!���~к1�Ҩj�+���<F*(�;��� ��/ =4�����Al�g�?�����Z^���鋖�֖0�F!Iai��ug�Iߚ�����D���XF/�0;�=���(le�wh׶w�k��h��W���UI���#�&�\_aj��D�q yȲ�V#i�D��Ȝ�1T#��P����3/�^�9���h��Tp��$ѧi|��%�>m=�)G�chj�W��o����\Y�^Rj�{ږ¤�%~,�X��T�+ۘ����%�N;>t�ZL�RLԬ޷+M�*�:+�Ql^p��:*E�b��K��z*1/�?�s�����>Z��E�lr[���CE4]d�cp��Q�j5���>�v��	)���_p�=IH^_��;U�`�y�;�.0�% 2 r�:��jm�u(Wk�	�������s����r���Z��lTb��ĩysv4pƳ`i�=n��:=qT�S��K���ī������BQ���6�0X��͍	%(N}
]�8������1��q:Z���lH2Oz]��]w��,�l�t2@�-��H���;G����4C�������}�H+�K*_�t%s�d�9$=dpZ�^�5�E�l,]�sJ=��g��_��<Ӡ�U -M�[?�V�xB��LMF����4_����"NN#�Uu����D�uO�7=!�|G�3�ae�*ni]O��=i;	K�<�ǉ#�����p�M���bQ���g3s/?�Vj+��u��r)Y|Y����%=F��r/���4���q����� �+}*��\a��K	����4���Y��q�b=\�Ҵ��U	<����b�^+w��]�sU�Hn�G�����w��P:W��_��	��U@�P˰փ����q�d���^N�������{;��*� }�ȝ �K��0vx�X��N%�rh̗̍�V���ԋw�Q��6�s�y�ɭǧ���4^�'I f:�A |oqi�'I����e��� p���`˸�'yǷF�2�+���jE�ܚ�^˛h7���T F0EVs�"a��G����1Q��"0�9F����������6qP�K� 
4���a���X�����/C1�b�a��yr���G�Ҁɋ���"��?%���%sX�B�K����3j`��-���p��".���_���;5BwP|f��l/�\Kb�F6O�ìh�{O$���a�����}�x1���}4rB[�I�),�2mB ��`='ȫ�*�J2י���4|-�ڤ!aӾ��ʠ�e�4"�&�.~��eE��PK5]��]�k2;V��a'� kHOA�0[�w��ɒ,z�R��EC��s�CmE���|f�TPӶ}�0��$Wn���g;ٺ�d�T�ж��o�!�ۥe�{�m���ۊ�{���17�������n�'B��^��:��D�HT͖�=g��G���"聼�p���c9�4dTJ�����td��ч��js��(p�7�WP��?��<	����~���Qؤ�7=5��[�h~���f$��G(��j܃r{�����{B%���� |�7M_��}�����JIͭ>����׹�>Ʃ��x=s�4��K�7��&�ͤm��>��8X뵠���)��Z����IX���/�ĖĽ��j˒�"w����������._��L�� ���V�DMtE�`.k��偺�p��f�v�(_�aS����A/�lx��,�`km�s�Ѫ�@�F��W�6�Tm�a*�+k�9P��2���t��6@��8����&�QS_���Nt�g��]��s$��9���Wּ����	����˸P�.w$��}Uj�۰�� LjI��J��>�L��x_�_m}N$t�Rs�;��K͘oUЛ���n6�'�������Jd����mcx�	H){&��(���w'�p�����	V�;�{�p9@�4�ټ�~/���-/�ϞYO�"�� ��2�2ۦ�;+�SԩO��X�-��Ѡ�S���E3Y��]�+=o�[r��18KV���	��*�;��HJ��e��C�����,��B�fL����?�̄�U0��G� ��S���������d����PLĒ�-��uP�`SQ>��4፦�p�+q��=s�߲WI�ê3ǃ&�l���X�H�T���-������F�z'�dGN8��h�5�/�p�q�p2�.&"*�#"���-o��diÈ�]����{�����mW-�t��:���>8|C�'��HZ(ZD������[Ӣ7�т?�zM�0G�b�FBI�E@�e^g׹���e��:�H4gj��������,z2ѩ*��af<.�A6�$ʖǍ�q<�4OTEE�h���p��ثx{�oJ
������Pͦ]٣ٌ�T|�i4�w�+��3��z��S(����w��Jy�%��/d=`$Ūrwh�Aw�B���#��ʳui,�x�W���� �l=����_ƙ���dc'�O<�h�4�r�s%�Zq�a����p�GrWj�b{��c��5nU'+t������Qј��k K(ؚ�N����-�����6jvrEN��v��f*�o�	�'x�6#��Z�F?�,H���I54B�Hf���cf�F�K��:�6�}�]�I���L4�n��mslmy(����T�N�9�PG�qe����k�+%�'���N�C��ǯ��<}I�}3�DQx���^v5���i)ٚ(}A�?�/���g��fq)��� >^t=�a5R�t��87b_3=:h��!��9�I֩��D�=(�Z��C�='�gm�٬��)�Ru�V4g��S������Kڔ�a��=F��`ʀ��c�K(�R�J�;5C|�O�ٝ�d\^J�b���:�T���$3�(
��}�oi^5@��논�[j?MA-�����R��w��� ����庄�����co�;��������U��|c+`��1�[e��t?C���PWĤ��wW#�EC�>c�E&� �@����4�= +��!ׄk��ɗ�z��s�w��<�`�!uW�(���b��ȯ*=�frX_���7�Ŝ�U�:-�������?R�&B��O�$/�-������B�&��1��qw�R��Ō��-�T���1��h�Mt��E�Hx��#�_�^�A�寎�� �5ۜ�HJT�T��՗uR�����qF��r-�={��C�Y��rwg�+m�g^��d`���閘˷:x?�id�[G�:暖d���O'L�v_r�[D����xٚE�¢Ñ������p�]ﯦj�gD������vXg�
�Z��P��6{�M]�"��ѿT�_IM_�W�3�6�J�ןn��kѼ��(��*�Y��0��Wେ��--���R�Fj��s}E��w���Y2���_�D��[E��*��]�t�1�n�^Ϡ[n���_/!&Cb�c�z�CxaN^�{��5M	s>�Yg>!�UxS��>��cJ��(�<�&k^_��ظP�
iD48��k�������BJh�ۘ"h��{a�p=��wZ�4\7�ͣ�kJ��k��'WnO �I��9]'a��k���#QT�Śx��};w�o�k/��mm�8��{�ĊjV�Kd�μ׋o7mvw�#�ؓ�L��t�;�P��A�]����'*�F���NO!LR��Ok9����p��Y4��b�^�'a���~�nB!�E���E#�9�A�?�:��Do֕{�*�r���� ٫7Q����o9��t��&=�i~ң0^ZWU����>>��;��8�*t�%@+�mJ�����P���1ǋ�n�N�g�9�_�m��ve��C}+�����7!����#��q�ƀs�������Ӑ����ÐitdR>a�)#FJ��e���q�3LsA�t�.�r6Z��ɟɑ����cOH;�5츩в����WNpNZa��c�h�i>�f��"�@L��W�'v�$�i?TV?� ~Xkt7���S�/O�X�f�f�Z9}� �a\�H�NW��y�	ɱ�P�|0�J3[��������t��v)���I��r� i9�ӑ�iw�x|j^�!�' �i�%˫ؓ:5�3�����|z~A_r��m���� \��m��q���D�u�?��6l��|a����K������He��
Ѧ-91�k���w���ۊ��N� ��,���D��J/���V�i�.����eOx��uv^ �����J��I�Hػw0+O��]�wg�@�
U� u�G�Hdd�Ԟg@�"�e�G�{��gD��g��l=��?�0���<����M���J�^�.�j�G�6�;�]��k�yg�._�LA�Z��F�N���`g��6��J����m�����p6'�c`X	f-�0�/���r<�g�m���_$����5������hPZ��4���ɈSPI�:H(� ��z߇#B!_G�Ql���u	�ko��E)L�,h���e���-�7����u��������r���.,Ä.�C!�����ig�C���$R��^�G�h�t�L�-��ANj�nY�|��;��LU&�s��ԯ�HȞ6b������ydY��S����b%K+���y�uf�R�P�1���q%����B��j���*��e�s�6(k��ѭ�7m9F?�Vs�\R�ـ�u˹�C@՝��,���ǖ�� _&HJܒ:�X?B�'���8/l18�^��9�Ԓ�J��$���+���W@C]˿X���.�f�>�ն�R�$���4O�M;��n�?��*��~YW�����k�Zw9K,}q�c�������^,>Dz�U:�m٪V�xU�ᶓ��i�;\�6��G�jOy&T��#�/���M��y<FP�W'���&���ϛ !�wT������p!Lg�H3o%�_m�O+���dOoF�l�ً�~Ɉ-pפ��b�,&��/4�/r�/���-��\��6,c�%@T!5s���k�̤����=R�$*�2�����)�^�07
�O/
���1���x�(���BD~Q��5o��m� +�h:���N�۠G�xA	��\wP��4U��om&&�ҏ���e3��=_�J4�H+�B�-u�4��" �����+���uAY��Ȑ�h�=Pgc5�aV��|���]t��� ������Y�}�<:���'=��b�:�r�V� ͊����)��~�� /�j��@䗾��3:��sO���������������d�M�,��	�!!@���+�-5&U��22���,��`l�CW�����1��L�Lst�i�9ț�{������eʯ1o�n9 ����L�s�{��I@�_��E6zℛyXS{#�h���I�#1Z�hs�N����3j=������`��v�?Q}\+ƌ�N��<6����H0���#�L��ӳ���N�b���MQ�6������/r�Y9Ok�(���}�k��֭M�`~"ç�}:&4r�� 3|$�)�q(AZZ�T���(B���(��U�hg�,j������;��^9�W��n�w~��:8��؄\�*��<UM� =Wp�LYg�qyL�k���lr�4�G��IoGk*���A��t�i0�ǭ�i��|Ҳ���\��`}n���a
gz��ht�AϮ ��
Ꮷ�={��Zŋ?�g�9�����ѩF<����%{���)��@U�V�w��E.!�_�Lh\�w�`�.���d�℡��*t�5�F���[�U��mH9�א�v��2� փ�G����<�<��~��%n�L��}|p���ks��[y���u�
O������;��VN��B]�˚y�o�4��'oHMz�pl��)B��kiD�φ�Ǳr��������RߥTV�[R���]f�̨��,�L�Bcr����>�����6�W?����C�:CDǽ����a�:e����l<SuXĉ�W.KfNM�$�����&u��V|,m�(��N	�輟�x�5���h�R�J������K��ؐ�Rj�e������=܍� ����j&��c��C��	Np�e)@bX��-����	��}�9��s�;��$��E�t�^�O5�Jg��H��7�͖�]hA��ɭ�F5zZ����O���ߌM�;aPr�� T��]�k������ƻ�u�����C��س0��-%��5	��"W�����|�-H�����O�.��ї I����ô�j��1K��z��@v0������N5H���F���9����SU:�I>��%�К�p�;砶�m
�Rb�ť����+-=��eC��`����R�7h��"Tn� �N[h��~����8��U��.ŉ�KSXD���kw
3A�*�,�*�=g~p����7E#�Yr�f�5ޞr��E
��"���Q&X$�G�\�=Gӧ�^+�E�w�4�<�K�f�|v�L����b�xF�eybͣ^��p��tas��tK���� ��S?mJm)
=%�"��{7�+�0Q��@���̷�va��w���M�1i��fW�:���g0}�k�we�Ҵٜ�ｘMG����,�^��h̔�Ken�����ňt4���-�~|k�泸���X���W8��a�i�'n��A�b+
���|�����|�B�MUK^����Φvd�q�Шt�r���6�Y���)-Jc��� 8'�ۇ>���A�G��g�Wy��i��|�;��1p$��Spq�,�1(m2�B�T~����ĆD�
[�EU�;�t͎�@�ZJa��xN騚.�	�:�!sV\�`��ɦ�y��))�]��F˯,^z9	�6!�������3�U�-5u�YC	1���8ĵ���#��Ŵ햯F
��T$?��)��3t>:�$w���B������)&�x�&�#��&���=4�F�x�@^�)�&v4�7H�K��K��!��a����]u_�D4W��1��PUd����f��]=�h
r�y|Sj���BKpoe�R�%N]＿�6q�:΁�Ӈ"�����3���BAR;��?�y|U��*i��s�X�Qb��[C+�����O�Q��M�u
p�����|�mVz�>)35D����E��/�͎�ff�;������ z?�?�r��&�
�U?���y@�ƫk��2��ٲ���/C'.��K�F$(��xE�F��U ^��|��{�O]�8`:N���7w@S��u�h��U籞@r�����o�&೵���>����f��Z������f�Sz4���T��I�1�ZZf��L���O� \ "��5���h������.>uԕ��?E^��ؙ�.��(^Q��N2�X�b���V�iXނ�`����)~���w>3}��k�H�6����5&[z#����D����Z�c��"�c=��ee�#pנQ�
)H�ySOᕭ)����w�f�$����_����M1)�|����zǱ��57\�T���+
XN|R|[enz�*^��	ޭ���F|���Qx'Th| ����P�6���y��ĕ�K�a�o���i��E̛8�y.�_��녺u}��
9LJi!��Ɨ������e��.ZI�!UDV+s���\Q���e�ʜ>n����J��m��!����|�M"�@p�qy�ɰ���IN�I!%HH�'�`�I�\�l��w-!����,yCq��!O��HwЦ78�qP;�pnm]���^$/��m��=�8`	$|$RxH�A������80�P!��K���A�錳E����X���m���'��+u���-����rǰp3����cxj/�g����x��rYN�1�	&��j����Do�e���}J'cP��Y���s�P(:��]"�� r�wf��V8:��������r"�w��:ge(��Ld[����=T*�s�V�O&���Q�wlbd9�X�����$~��(g���H�~^�����c������]��Nk�}A�+t̩.\�~�MQ+���Qr��U��hɥx�~����)W�p��N�*�LS���jT���l�nu��������'�ѐ��p����ₖ ���Mݛ�%%��?`i�Zb�q�#���ω�F�� 3����3f9�	<t��֯aUc���
��H��僼a��e��\?`0��}p|j�r��j�A[R�o�5�>-�k���dF�pQ*]*��:�v�syy/ЅM�����!�^e�;�� \ά����]�Yj~-"�I��hA+��RV�TlAbo�.qLUH�TMD�Y쒄u ��Y���K�Ϳ�yc�O�\�B7+,)ѽ�ѰA?�QVX��v�+}��|�@���"��xĈjr��:��3i2����'Gc����6��F!;w�35�q�L8��Q�v�hJ<w.�_Q�&|����0�w@����� {r�|��F�o��:�v@ ��4���辐��0��+���#�p�/��'|��������	�!n���55$����-�4��[�v^|$�^�Yd�j�"�8i��D���'��htQM��|��w�aza]8@Oi���(��/�H�7�Y-�L`����>�7��"��E%���ƞ�g����JN���)S5�E����g������\ěH�۸�7otm�8x����J��5T�)-BmxD�V�	�F�T�}%ŭB���
e%廊ɘd��J�y_X<?.�uy��i'G�{e�R!�;1lEK�J!�>���F���NӠ�r��g�uw|{�nXE�Gk�A��E#�<k@��������ͅ�l�1���:Z`6�D�:�nF[��Ֆ� ݼ�$�X�^�zT\�-�ֹȁ��i�Q;�ˆ^Ʀ2�7�g��u�0-�wG�!�J���RN7�P�{��!r��t=�~7ʤ�9�Ԃ���}br��lDS����	�7;���B˒�t��s���\	>��r��7i�k��~��f҈;��N��J��.E�V��OW��2�|�8����C�<�#YU)z����~��sr2�q�d��
�\�Z0��PUvml���h���(7Y�n]��Ix�-)F85�s����[=�W��I2'҇��q��+�V2����r5�^�=%R�Μ�����6���e�ŋJ���/�JM�S�f|i�7��C�Q9��N��vr?6)�� �U���I�+H*��g�CT�e8�����7oU��_J������R��_��Ɨ1���&�֟㽫ɇ�gH�۹P����u��K�hW�r����x?��Ġ�}�&�"'I�H+��4��H����"k#t;��M�'��5@d�d*0�"lX>� ˆl�dp>("�]��[��a��4�Ej�+��%��Q�_�E]OE��o���>��\�X{�@<����}IK�h���t�I���vݴ�~�G����'"����d\������_�9Ij�O�0�\ �]uy��F��fE���g =!�Jĭ^�7�PP�=���8:f{�^�����F��]��9D�]<\�L��J���%�f{���H¥~ ��G���I07xNV2/�Y����A��غ2�A��ϕ"��Y�UE'�Z��0�qs��  O���p��`�U-Tn�=�I�s�q<�߱)���=���Ӵ<	S��t:D�1>�(���+�������cb,���f\N�u�F�cĸ@/�eZ�ը�A��I��
�Ġ��{�>��$S�I]jC���	��,W��b͆�x�u,E�m��'�;�gˉO���4�K��w�q/��#���uůA붧��Ņ�ܽ�H��mؽ�z�
�bl�D>G�"���z�ۺ��A���G\6F:^���dx���u�(��9)K5Æ;��	U3�]g�Ig��q��˙>��/�J9����U5�*�)1��[:�4�dC��>$�b�vmfއ��xu��v��0n����Kv��y����o��)�9�ۺL�yU�M�m	�Ȏ%���"Sf��=�gI�*UU8��Ԡ�WZˀĔ���2���� �Y��݈�ނB��������Ydу�tms�Y���+<�5��v��b��뽕����6���/��V��m�$��#W'c>�Lub��x�Cm�X���z���Ld����RC����C�����o����1qL-<wrm-v��{�YЖt�w���Ԛ^?_���M���R��E=�} �$�<��ܪHŨI����/uG��G==�i>S
*�HY�xXP�͚�	*��	&�������a����53���4�0���^��N� G%�7���M�P:��O���G�ۓ������p��~X#��eڍ/tJ�����gO�4Qi�r�m35=�'3o G�����ެ�2  %rd�d�İbGe�6��j�� #�/�9[�7��a�1�p�V� �ͮ����>l&&w1��߭	�[YuZ|�bM��d}���+�=�?@Ոh��v��2�U3��������+�AwhH��R�e�c+9��Q����RP���erϿ�3���Ʃ��ɇA�O�ax�U�sCBc��&V$Q�[ڬ�M\�m�+8r" ���	9���x��j4k_�gB��C�� ����*�r,jhX�W���@�]pZ��'��pe���g�q���P#���-ɲ��Ev��f="����ɋ���F�_��7C��� �A�R�u`�mx7��Z�Zb�x�$1Gčオt�I���
(����<�W�@��H({h흜�ыJc��_2̖��q!�{��*)�V6�ث�a��흟�Jݾ���Wotȓ�� e��0I�ǂ�KH��i�tf��E�i�7���o;	�C���V?7X�k{�[��vV�ˆ����+�iS����#�*-@��CU޴.�;�X�E�7���hW�LX��u���gu�m�'��壉���םfn��ɯz洓�Bn����V���J"�h�?͛U��点�GC�t�0O؀&Ѩ�r��O�6���c�g B<'��v���H��X|�:��8��p�}�,���O�ӐFVKxK�sN�K��s�K�0'�(#��뾳S)�b�Iƈ5|��|�j�R���&-X�D�Y�a��(�v��GD۩��'@��g�0�ַ�����&Y�X����Ԯ����R*V��&�[Ry�n�4�uDaԛ宮��p���9�n8�!ҘMo��[��H�M��G�L�|ko� �	d�&��#E�=֌?I8b��ֺZ�|+*��9p4��`տI�?J�ɳ�{��o^h�9�����*��b�3g�&sb��i��_b��Pe��[�̂A�!�E��糮��G��}� ��dn���l�7�>8�}�M�g�.���u3D��Ju(�j$4E�J�@��U�U������f׵D����C.�١��K��O��5�$��h&�3E��-G7x YǛ(N�a2*G��0���2�j�/��V���nx(*�o���8�f��!ى-��m۹��!�H���Y�\��'/�v��ЩYk�|\��̳��p��\��˻���o��ꬄ�>=~�p�o9T9b�m%`�&� �	;Ʌ�p���V�z-������ F���4������
�a\�I��̏�S���x��َv�=�s����?�,��{{壸!���j�j�G��{MptT��iN��W�u�娳�<�����Ʊj{BFR�����\Ӊ��F&d���|���F�����Օ����M��ƽ���=n�(���֠�|R�dV���i�:S~B,�O-��������)ٝ��D_�@Ҏ���I`�y^�_�t	^��}
r�ŭr�'U�EC��8�����%��X�6B�sH�-��A�p��D��<�b�w�ٺ#�w�B�	M��D�IQz��A<��Q���|��C`�P��
vK��$�h��\��W*!.���\��y��k^p���,F�>ݶ�,� xd";�Z=��Q���y$m�p!�?@��l����B��_)A4����	cX��w �4��������Y�޼ ��:ʣ�$:&���qQ�k�oQ�I������?��y�gt����B�;�#���:z�^6"�u���d4>�������O���p9,5�DW�����.
z젟*�kЧ�u&˹�W\��~򳥇+���Զ�a�4��()��Y�MB�]�i, xߨ3\��1�-��ý%bb�;�cv�-ʣ�ђc7s���T���b���]��"��zL���N�Ru���}ͼ�K4˽Q�w�I�˓��+K����\P'��i��=�nV���l��r�m5��������5���?1���7�E]�uӱ��O��d���W�~�d�+$q��s>%4ؔ��s�B������!��𓱫HW{6F'�R���eD���t�	����<�OcGԓ���<�2�I�rq����P�L��-�qT_1��ֆ$���AzVv\l7�ƸA ��Bn]m�97�m����ߕ��B��^vࣿU��ޭk�N�M�~�?`����%0�AZG.��i?N�T�,*�G"��AuX�C��#�Kˠ��շp��q��X7XS�UH�bB�m��7ψ��n��d�O�n���g>3�W?�ciY�ú���T�k+o>���)KE /	9~3����G��d�[9v��=z�D�{�z��9Ҥ|p������L�3p���P�"�[Ӄ\����p��#R[TW0��9�5�d�|��\�T~�E��c[)�	�*`^#]�q��Z嫮�wa��@4�4�i�[��`��E��U���(
�����q(:;���C8������.�5710�ML�!�<��i��W�����9*i��g?���es-?���UNXWj�ק�|
kT1[hs��+�������%��������V��_��0�+���������3,EUqġ���7'��M�h3>���>%2�2û��U ^�7����^�k����ӷ���_V`W���20��;�F�����%|
1 �Y��Qpѳ�ݔ�6A�r�ِ_G_!o���:��x�dƋ���Tdv%��Z�J-*��\���iU���`� ��<;@�[X�C�F��6�\��T�q�E�����Gx�5fH.Sp�k+�ޜ$
+V3�����w7�s�~�w5���Hk)jx�@��(�+S�r|��b�^�oa�?���d�e	���T����g����3���3*`o�vJ�*��L#�-�q��`�6��+��k�dN@�q�Fi`�2���+����Z���sR~�:H\��[k��.���$&����������Kј�wZ;ɏ�lG*Q�����z5�_lx�X�  }z���r�^�7PE��S~÷����k��fq��S~����yCl\Z����p����v���ڢ��f�nm�y4���,҆��v;�4�ʩS}�A���S���0��=��_og�f��J�K����X$�w{B*��?�[ͽoT4H�jhN�Dk�U.���5����]w��9heV%v>���]����L�fd)�Hl��H�����G��w�Y�o�,��qK�+��yM\`�:P�P���/�%Od�B붶��~��.��졅_�I�҉xc�� �� ���u�Қ�V��:ek ߌyb�o[v���e�r�	W����I�e�s'���jӌ�B�=K�: ��b{O�ٰ��Yal��N�	��ܖ����ij��hއ��ʛz/��	y���~�s�^YU�l�6���V�q��tۃt�j^Du?�+D!q~$��ƎҊ�6������9tzĠ�Qd΢�'�[�.!����9�^��oU^*�,[�&l�>�lɵ�rJ���*����ȷ[�wM?W���=hW�U ��q�.ݰ��������1�%�g0��_#��	���@����3�&��у����~��^E�|B:�!�g���~�D�H40Ϸ���������B����EȈ��e�܍��&/���H<�@� ����o��;��;fG�ջ6 ����ka�M��S����*)�Zy��j��7<C��S�մ�]󺣒`u�~��hE�m���e��^HA�X�����e1����mf���IL)Y�j�6�i@[�"�dy�5nS�|*�Z!�n�$��c=P7����5Rgx�%�c/����*̒��r?*RXb�_�7��a�^�>��Jl�e���r4�ʘ(����	���n33�Q˰R�x��R�<;�[?ps��j��[}z�']�7Ke͈S��@�p��u���KW=��
��&�4�U:�7|L�}m\��}eۈV�S*�S�b�������h���e!�|�pw_WM�l?�/֜�ۏ�N�>q~�yZ�؝"�e��nfDf(��V�q����I:����C �vU�2n���h��	���P��a����+n�L! N�u� ��������l��Q�3�?'=Î벧We>E&��V�O$�Ȣ-Hn
u<p�5�i��rˀ���!��2I]���#qY�NXZ�?�l��
v�W ���%��OV���ʸ���4�o�ga�p��3�е�P"7x�'�X�L�hS����hK���)_��}�?y��V�B�9vٞ��|�_�f����j\��&Ps<�Z� tᖎ�ɹܤ�g�=���pz�����fw8�f)�f���p�sR0�B�B��