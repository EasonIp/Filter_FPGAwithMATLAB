��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|۶��-�E�8@|Jq�^����`څ)h�(��Թ`�4!�s̆d���GR`���"b#	�ޯ�2�������_'/|~� ��� ���^����{h/f��Z0#��G�=Ǹ�k���M:��i��a������bH�C��q}fX���o����*.@�NV��x���x%��\���I3�Q����J[�<,I���yM�D��څ�Yo4lu%�[WJ�<��_5!��@p��Ȕ��ˀ��y��_�D<x��uo*C��|Iv��JB�v7'|M"#Lw��rCV������/M��7���W�la*�%��q͋^`_��(Q��K�Lz�]͌�?��ګ.%�h����ѳ�N<�N���w>m�"�Ɖ\[��د�u���̋�%����4��'H�пO�f��݄h��Ym,=��֡,�8���t���gޠˠ �frr�!Y�u� �>囑"Y)�5U�a��J2�����1l�"ٲ�p�?����Xw����t(ߺ6��c��g[��X
����@T4��{��sf�Il��f��n |؏i��9&Iv`��n�+=5B3��q�p}]�o:�J�|�$�7�B����*A��ڊ^� � T_�H\XYH�����'ш|�/�8ZU���w)�G�7�>�ޥ������L:sA���`�r�8�a���3	�|��K��}}u�0߱6�%������� ���ti<����Y�A�q�{d��6�
\N���X�B�t���7y~HhIJ�	A:5��[s0W�ϑܷ&�<.U@��4Vh���?��\o\��7�p��hfG�1W�֡��wK�)0�*�"X]eCv��{F���n��p�&����U�.�K�2 L[p����$8���+�'�U��Qg�=��,6��Dp���_�Q�H�z��J�r۽��F��/ȅ�,�>V���1������A��HͬǕwq���\j�1HK���KK�Ə�� �da�u��y�sZ'B���i�챛NzP����/��}����8���=���3�)�38�\������Y������r��̮�]�x~6�`L�e�_U6�Ѳ#Q09_�銃��46���Hw(HvD�ͻ\!�e|���ܵ!Њ��n��>�a��IU�Jv��v�Y,����p���:�X61۪�Sڳ�A��h��s%~�X��ü�����.*�D��\!N �aLŹd�7.:c�F���-p�\u�/rԝ�Έ���|�T2�*P�EMW�u=]�o�Հ���(+�\ׁ��3���7�=/A·6Ж*u�ӂ��{t�4L� +���C�Ϝ����彽����وԊ��4�N��Z������Ռ���O�n��REK���\�X=A!)oDH��t���+=�*�����B�g�����m����T��$L`7�'�W�{��(�=h����#;OQ�a�e�:*{S�vR��>�pִĻ z��V2~�Iơm���jt(x/S�/�����Ǐ����y�����"���};�}pXEsh�#�x���L:���b<q�+�nթ��h���OܗV}��*�gb~�(�%?��^Ɖ@>^إ�[�l6my�㨋9_�B&q�����M9��O�}"�e�D\c�{����n�G�f{)����̖�'	j5�ep��a�
��)�������/JP>�K~3ҝƂ��N� 4_R��q�9e�0,y6@Dh�e���JUЂǄv����(V�><}�B]a�I���zw�t�tK:�z&�S��w�#�y��K�U��X��	�}k���1���)�������H�§���y��N�S�%�R4�U���ٽ�yXg����p��y�^�����&B��jzl�5��q�����x���L��{���ي��.�1���	��|S���VjZo_>�8�<T�Y=�opq��f9{Y��ُ�!Pё��o�y�4P��^�^��Md����<J��m#|�E3��h�z��� 9e 'I����b]/N�H(7�x$<��k6�zx�4毤�k^��e����J���Y��P�PЮ�aGzx���������Q�[e�A@�̪��۳���0*�[��m�_�Xy�w���1	?U�GԦv��~ٵ���#F@-��)�U��&�2�Љ�Q������O��^i%��G�(3���+�k
u]=��l/�0L��S�N#}28�`9�\��}k�R�̼��Bg�J\�=<��{�f=��̈́���d����Δ����	P��+�Jp� )�����/�=ŵ��|��s��A�^�0?���5�p�l�1_W'+͹��|U�mﭑ~��0�zd���Q\P�euUzɚM���J2���z�[��44,�H��,&�r�l�g�����PW,د���`Xw?��K�2�a)]!#]I.[}�_=rP�*׋�n�|l�QR�9�A(O�NcL���H���|j�)R��9ܳ�m4-�?1	P��~��7����V8;JFUN֕SiQ�YZ*RIn���k���º�U6�%ُ������N�MZ��QU�;}�-#�� ��T7����ov����l�R���b^�H��/�w�������������l��$m�9s�&�9-J�r#��y0�ah~.�:T~�&����C�5︅w��FYӻ�ۄ�
\�����s=T[�%^���吼�o�c̢���etPVS"��LQH�5"47ʻ���Y��@.E��t �0	V�i��-uz>ˁ'�������!������]��/r#_��ej�zB£�<P�q���9�_#��_��N�|F:�n���uܫ��"��a/��)��2�p� 	XNsߗ\Ahz�@���e��<�u�
�%2�i�mdL8�v�;K!v����ڛ�k<!U�����ÿuZ�����B���
�ػ����@	�X��9"�(a�,�ߜ�p��O�6��٥:�?"�'��)cܻ�c.g�����Õ{s�E$�\`ޗcB����"�-p�'�	FE�"� ;Z8�T�aa@R�ݴ6�Vd\>�� +uȤ>-�/���땊�������h���gm�a�����L��H���~Xt����cq�d`j�J���z�T�dwꙟ&7e�=�׼�!�V�si�k{��:B���}����_�ŏN��zԕps.�F�s�Pf�z�������1P�������c��oLu�mE\w��!�P!�V��� �w`?shk�]¼�u�/���C�

s�B�a�$�
N��둒{f_��Ґ�?ޅ���e�
Ć^R�,�!<w6$��Ӵl����E�)�,$K�씋0��S��⩕�ʰ����E�6@{I(��
礏� ����)ݔ�)H� ���9}/�G����ݘ]nT�qk)�y�
��]"T��~��z�V�k�~ʿ. �uԿ��8;�_��
���	��-��/Qn������Z,*ת,��@��-e8�s����~V���N%煿� Iy����/��.UA�� �z����|<�4AiŲ����8i'�2�^��O�e��ִ�ȹ����xC �[{̜��w �G�?epy����jv��h���4,k2ig?�*��E�π6'�� ��7�x�m�g��6����%��on]/��I���|���#�,%gI5*���6�ó�,9��_	�>E�KT����3�u\��������@��N�=����&9�sS��y�W��+�șЀ���P8?��&�E��nj�������i�p��>��G�	S�T?��>AR�y��ܶz��)U[]��C߷J+���ٹ��P�-ba�"�'x�{tp��v�>hjE�FKs�)ڑ�Q^���n��S�6HiF���A��Q����`�c!s�1.�d/*���G�^̞-���Ğ�GfSỠqދ��%E����g{�WdY��d(2�ؔ~z0t0���ONZ�)B�]������͖��[�C����w��/�)h�0�K�BӾWqn�)Ov4��0���A״O�lq��B&Łe��0c P=Xt`�% �v@N7��	���,�#
��y6�!�-��a��g�VT+�K~����k\�7�2�L�P}�Gd��vjs0�4{5K�vm���X���qw���R.4:�����vK��N�II��%�묒<�1|���j�*�2H��ƅ�K=��,��9��ˈ����w�Xq���B�6�uu7�8K1���,�H�vO���Ư�DW5�OcO�TsQ��Vm6�P*���=f�&�@2\V����}E��:�w���1�b[:��hi���i���@�}�al�_�Ї(��2�S�*�������o;����Ò�!+l���d�)�ؗ��`�������.%����h�s�c��v,�ի��J�~4_O�⨄=)��8p*	p�Q��/K}��=��
z	�.��W(�/u��Rڷ��WZ�E���!��CV,�A1eb�0�Otl�^8�L�x��]��cA̚�-�ZUI"���:~65:iWSt^΅�\�xc�$�,�TQ�|��?'�@��'������Q8�����8ꤓ���}�
|:��f�!Eo�i�|��S<2o��hOv�����m��vԠ�I;ND��ͤ�w�ejK��_�l�����>�:���k\_H�}������t��癑I9�����:> �O�����K�)�	-�}��6~�]*V��O*(=dʺ�����2��?lF�-����27�/?s��y;ySr\���C�P"A��t�F߸�4��>������h�`~��,�:L��e)J��M�ANR���?p����MqSy;���(�f�~)-��`"qVϼW�#�b8�O7���E��q�R'=VN�CÁ_M�~��k�=a���[h�w:ɫ���lHRA�)����� 1qQQ��b�p|�p�Ig¦�_�JZÁ+i�K �
��>ѕX0�i��]%��BJ?;9��`��9��F�%������\4���a5ŇC����g?�r��Q����dy�
aj<��G����MUOZ��8ؠ�_�����=]�}�>-��"�#R�.�>!�>k{�f��tM1j��M5�:g7�p�y���i�Kk�
^�'tQ���_u�����z���>��p5](#\�d�R%)L�T���O�G���͇�L��������.7��P]�{����"�{[��n8ñ"g�R�%�S#��<AZ��l>������a�M�>�?[R�8RI1i`Y
���%�\d���P����%y0���!Y,5�<r_�	o^59�1����}��Pأ�_rþr�>���1��\Z�&{�8�� �i+�UZa̼�!
�C�[~���O#x�#s�([�o�=W?���)��đ�򫫣���i�d���:E<C΀t�K��y�ĉ�nĢ��m͘��^ۘ�^r-��R����4M�叕��<�%���D
O�Հ�-VJ+)K���[
%��"F��b�ޞV�ُ�摛�Q
��C�b\[m'�/��p� z=�Yb��r�������� ~u��T�77\�I�@�ќu�
�+�F7O9�f�ţ{��<O���h��Z�s8�t��N~qc�}��	��ol��h�\Sg.HN�)�ڷp�SUR+|(��`¸ZHv��eh_��� � 0��	�m�eˉ�b�~��Y�N%^�Я/޻aJ6u�@8u��mj�;���aa�JѪ��˖��iC4������mf�l�jy�V9�������L��Fֱ��,A0!*},Fz��z~`�x���svaz�C��9_�g%b�:MG����Ֆ���㑷w��U���~�q) ���n�s�d�F��������k!�=��u!c�fN���6�Q,Y�ǫ�BX�4�	p��̌%�r���D�[�֧�ꗐ�`�I���-f;�v'E�-�&�@���8�d8�1�
~e�C���W �O<x�2��S�*����h����:�Gc�.x��?1�|zc̦0��IOBhТ�� �hf�*ʇ�ܭ��`���w�4�ܺ���oJ�n�%�ct������3b2���yag3Sl�E�"���4�rU}��9�;�5n<[X����S/B;�o�S�6���G��.��� "��߮�`zaD8������uQ��Dk�U�X�5�� ��0�6UU[�d�O����h�7~����&왯p.�Gf݋)\����:Boa��b��8���V �o[��&A��sW#&ѷ��R��k�	��3��Ƽȇ�~)݁'4.&�("�;G�ڬ�5j�1@ar���R���2�婂��,�������&X�gmBSN�M��a���#hۀ�ߎ'��ݽ���0�	?]c�S�T�T{�V�����/����8/��n���'��v6��پA����W�
m�_�-�o�� ����yȜ	:8��m��l+ ���d���9V��-Ss�ltǑ0�ma�&i�W ��c�p�K�R�-�(_VeΥ��>��3��Z*|����3A^Oq5I����4�+�������v!����r���(>\��Z����|+\`�['I�p_\M����Z�^KT��%�Lf�e�1��S���֯��7P]���Yy����t���z\5��X8�&�t/8\!6ʛf�P�E4��1���y_9/��C93Vh���h����D��d�$���e;��hS`��2�&��M覢��<(#oڻ:%T���l��
x�kK.0�q� _��G[k�����JH�u��a/�E�U'>}��8�k� ���z��y�|���-"w���>�`{�!Td��#LFȹ�ޕb5�)\�f�]S[{�:gzŸ�n�ȣn,�F�%��K8&�M/o�G� (�E�N��)/S�Aw��P#�;��ַ !�P�s/1f��{0��H&�7U����
���w��_�;�z�5�1����HA�U��Dq �A��(ˁ�k��QM�g��# ��:�k�0�T��D/�]���ZJ4
�w�ԱS�`C��_]AGc�2 �g��z�8R�����tZ���m��Z�m|��H��������?؊ʎ)������Z냦bF�oCq"�)t����D>�R��m�~�o�y��J	�Ay������1uF����ܵ��gL*Z{��JR�4���UQV��>�e|�y�p~���ٱ>&�I�������,t9�ϟ1����F�w8��x�4
|�K�c�p��F�*�D���eI���a�v��3hٰ��7�{<���TLY�#W�_�X�FB�u$��"��n��Q�m��q?ݘ�3t���N�׻B2cw؈H*���n*T�3��q���.%�%T{L��S068�ט7�Rl0$���K�5=I|i9䂨mU��)˷��A)|M���ƿ�`��]�SEk�B�Z�����QSc��ؽ����3U����{ρx�#*(lE���[;ҳ
��%cP���,޲�Td�f��c��g��+��͹G%ܨ�Q)9b��/rV�W�9�d�0�y��/p�\;R��H꛴^L��P
��Up��aq�,�wa�J�El�vUs-&-?�k�!�*�NBV�/H�kC���;L	 u���i(S�Q1�Q��y��Ƕ3�7�:{�I�/�=�ptڣg��Q�|�A˶U��xoa։G�N���J�2�R6�9�􂐃��k�����;a�U�.?p�BPh�	�t�/	��9G�9�0�RbS`�_�_)�Y	���a8�_����$$~����9�O,+P��sg��{=
ݬu���c�,�� �%��J�Z�T%�/���_fvC�ge���z:�~�nѪ�s�D|:����):i�ͰoeC�D�Վӥ����)����N�,v�zrk2�TXOw8+�Vy?y�n\}&�}5X�+PV�vH�]k��/�z?笰O��b���}"��sn�f����٫\2]�s4{�J�3T��������I�7N"[e_�.e���!��H�%�)��P��8���g��g�6����m����rm�b%H�ؖ�qK{���U�L�3��!���c�1����wt�.�#P�{]��.�(����v�$cuY���X�FxF�`�
n:u��@hurT��hm��r<��;���T*R.����*GHXLտ@:�̝cڨO!�b��[��#�l*��"铺�K��S��c�c�_��Q�{}$�''૯�Nd餣�� �l1�Ή55�J�%�>��& ��) �aO���R�S�D�{ǖ�#�p$�To��G�3@�a���I�9?H�8�en������S�6�����i�� }��Y��u���O�H/!k����ci�u^�0��/��t�>4}Ϋ`r�U*{��Y�X�3b���ī��c။�Ѭ� ���T��9y%���QZ��vn�����%~�x�u�\e�7�u�r�Uvf�#�6�E�'P:wV��}:�D�1-��)3	��H�@r@�'_DX�y8�E( ?��	�Y���:j\���9�u�Vh��QyV��2v�I̎31
/Veh�˗�%6.�7sk���U�tWp�aI��:����}U�
���tbGcd����)@���Ji�E,�׬�G\�#�2�٘����Ej���%U@׶u��@Kz�0ɳE��P��Pr��E:���p+Xi6��lfI�����9������](��O�ɉ�-E��#Q�F�����$�L�Ӊ���|��?��c�6
��:���w^�6I�V_U�vٳGG�9��9ۥ3$�M�m}������D�V�(�kGx�L~R�8!Y
5G�K�����Gq~v�Dg$���!i�_��J�A^0:�J\Px/�u� b�z��L�7c��,'�}��H���4����1)R�
�ʒ~�T��R�]�o���<���堣Lb�jzu�@jו�1�����9L���|,\�%�px�j��W�\�}�E�!-�����y;��
qcm��"������r��T1�	���]묭��#��'i�: �40`�Cĉة� �K�e��'%3�v�LʉW��`�wQ+v�Ra������m��D���w,��w�L���0��L����
~�����%�N�xQPx���*w+χR j� w?��⧲H7j>s4EL0��k��l�
�QE�6c�dS�i�\  �H�����r��N~���@���ޅ:��]wMduqû����v���+���ԝ�p�{�>�@��ꝙ*�R�gO�! U�U�	9��'��ޏ@wY�3^��7��.��T:フ�{�#��x@Y�AW������|��S��>,
�/3�����?�Ɏ�@-��[d���|\<~�cK��dV]�t`�=h�Y��K�yg��*��ܰ1���7��8WDP7`X�)�f�KK�0v b���L�) �8ʒQB��S\�L-�q�[�Q�F�)$)c��!��etт����Q�ʯ0�q�� wP��W+ �;L�����bF�a�u?O"ȓ�.��c�T�p:����l��Q��%7�};=��e�\&ly7-�D�n'�mq.FfE�P�p��2��2�|�󔋤57+��S��,֚%M_P��Ƒ����0���m��fb1!�~4��?�R�!t���L�Oz�ˠŷ~ d9�}�GnT�:�|U��i��"L�L�C���۽
:��v�=��2���
�@֠j��q�.��l��#�Zzז�D9�?�>*�d�u��8]2?}� :9&w��C�V��j��-'�y��M��+ �R��s�Z�ξ0�����3c@V�Vv��^bC��z����"��G�7��e D�L�e���O���[c�4����9��J�|�~,��*(�u��F�(3�&���{�O�b6�rk��-�N�=FN����;A�J��-$�`����j|ƄO&�T��x�sl"Q�܉s����m ��N��]�!n���҉D2Y�U��gɾ����F�x]�ғ�G��}���	�(�w�~��@ݚ�ZJ8V0�x7R�5��^�I� �<ԡم�ř|�����2D���M%5M8Ϳ�ā�V�UP��c_�<����nlm��H�!xۿdP1Bȴ��S���i��ZZw����?a��}���PqW�^�����x�`C�vU¨��Z�7O҆/C�T�HU�n�SN.�eȉ7��g"c9׉J�Z����^�ř
���wA�ӨjC��o��J0i�6�Y��7��Υ��f^�O�{,�h=�h^a��^�1�1��<.c��X{��&�T���$D	G�$/h5	|h� �`G:?S��L����*ፃ��7_M�߷�h�mN�+���k�^�ϗm]0�s:�l6Jd)�����⼪�dՏ���z�����4z�D�_�*�z�-��\k7a4��A+v���T�Qo�^����ų���ӊi��F{UE����(��K��f1�<��v�@����T�8s�z���/�79r�x� �OM)A~��5������pA������8�qXv$ǥR�tHuk�=�h�l�-(9�g}b�`���Ӝ��Ϩ�vґL��>�$l���G=���Զj������fq ��O+�yc����~��#Ŏ�CC _Ǘ���T~ǖ��ƪsn�v��^߅���i{`�=�b��~`p -��*<$Dr���?-���L�����_��b?]�A+*[rX����Us��E5(��D���&?xyLK'0C��^#�@-	�����P��<��N�d�\痪2�FY�i��/��][Zٷ�T�C��x�R���B�޳u��II;l�n���8k�hm;#�iB�|"��s԰=4Y�KC�f�W�X>�X␕.�����q�'�J@PMثH����2Ҿ�o�(��� ��|�+y�P�g�Nh�z����
�[p�L��eSc~}t~���הD��슴�H,�Y.�M���[���i�h��q��w�� ˠ��[�V��ņJۧY{�EpO�5��ʉs_K5lu��c=��X�3��t���3BA�x�`��u�nn�<CB���WB�1�B��.�tǗ���*�8��9�^-鶷"�>	F��kN|�V2Gu�')sdv̀νB�N��~��f|�o���&n�֧ڪE�p}���h�-C�S���z���v�8���w���Gf#���+�bGe'�{����\�{���6��(V��� +���B����^0D'��> (mw$�A�7������ƾ\Ȅ��$�*��p�0>���D1�PN�$��x���FZGx�|& ��˶P��z�|Q�=�8��M@�կ��@ �	���$ȫ�$�P�R�Uvu�ІK��v��=(��g$���C}qq�cK�70G,!��R�C�%���#
�wY���,i�T���?,�.U��3�뺥w��ߑ̈�|t�`�O�"{��"Wi�?{?���_#l� 0��,�Lwq�|�	��e_`������0��Ñ���u ��;}]ZoMN��)G�7�x2��I��=��ƕ�_�Έ�M#}�=�٪
�S�bO��Q1! ���9�7`TK�<$z|6�}��۪����M�CiڧYԃ��Kzi�7͸o<mCi���B� �<�>�7�e;=Q�M��P�
�Y^��0d��&��^����$y��H)Lp�V걌�������h%_!̇pB���J�t�|�}�C�~(xs���{A���Z��P7#�\���H	�c*�Ek{o��ۡ�y�9��ej�/#�8�"Of����+��;�D�9{�"`�G���M\�b�zD����\;6�&W�������%5�t�����+a��(l%.�	���j� ��	�AI��w\{��B����%�s�_-P��>RO�T���l2&�~:�@��G2q����Mx.~�8Ň�U���TJ"S�H �{Ips���}N���g��$LAcP����t?p�`������2�����+\��W���,)Y�|h<���+II�҉v��?ؗ��s6:�@^[���2����P�*�
��>(���0+]�Lv��!"&����F��I�c��������'2���8n?��\�e{������]�;�	pJ!�i�y����~�8t�s�x:ݤ�jFM_�t����ey���3Xˆ�Z�<~��Ra!�T�wb~��!�=�n�u�H�Ĳ�����/II������1��M:=�����#j�џ�s�bZ���'�����`�k8����$���p���u���oDL㗗$��?2&��W�`̟�t�H=}E��\"�o�+<O�H�
�t��jP~	�j�]�ak㩴K��w�c����uk$��.��m��
b�2K��5�|��O�l?}a.�PW�C�>sY�7�܎,�3�`ǟ#ߔ�ʶ��a�;6`��u��0����3�!��&d]:�h(�n�.*�<B��Jx�X
	I��>X�@[������o.f�Qo#zt����JF"����_��9_�gn:�����fZ���r|#I��l��w۽��ib�G�G���̷�ӧ��h�l�%Y� jK��5��� �����n���|m<��oZ�Us�����@�9!@W�^��I���I
S��O�k����J�?�˂��'QkV\ǆ�K`�>4���=��S�w�=�ף�`���<ĒWR�����0�?g�dd|+���Q��D�m�Ɩ_*�ۄ��Z5Uo�i*pz�|EV���^�)$��w��o4�[�w�{`�Q�@b>H����%(�4��;�@�d�6c���Gޣp�4�:;�������)DkܠE�dĕg�@���7zN��u�.|Ԗ�����o����h�;]��6�p;قS�
c�VRB��,`�f�W�������w�)\2$~+c�*x���e=*�����^8�m��?�ÂQ(�3��g�&�|D���꠱(n��uՖDdx��­H����W�1�sj � ��a������A ށq "��8���c��Sy�6��|��U�����<]tFj��p2H�d(`H��췊?��(�V�ޫQ?vo{l�(,�(4Ro�A �t�3a�B����'DO���v�f.⡋31��-�8���r=kt�f�K�����U5�4�x��ZQ�;D7��n!��-e$�*�h���������jbk{0�H�`���<�=��}�4�U���v3��|����s��Ҫ�,�(��~) me^�:���(=zm�n�y���T�>�x;�*ɞ�^���~ȳ�@
ru��(�qD8u����wՒ�j����"��+,���ʫA��u���a���J��7j�B�K'� h�'c�lg�}@��S�H(� �.Z�y���"%r�a��rI_�/�(Q���8�"�/�"M�?�j�M��cڳ�u��l�Y�\���y^'�|Z8l����R&��@N��N\Lw@x@���MH�Wė*�C�-��;F��K3u���{�'/Ll7��K��
.1�V�7s�PT����eW>y��|j�Oy��OB����"�<",ɛ-bu/_�����>4�m��qx���%�[�P��t*�������M_r�8}jm,S�؆�8���ܕ2/�ۿY����� ��Q�_d����_M`�n��,I��)�31Y��8���pzI��U�Ɨ��	�Tl�ؾI��ɜ�p�a��dW.�:���e,�3�[u��ɣ����y	�hꀑ�H� ����ʎs��Sͣ~�6�C}[A7�{6��F�*ze���H�z
�m�w0�;cW2����H��d������?�&�ߑ��Ī�Q��Vr�n�vi$�=��^�e��c7�
Ac�����"3�,|��o�[r����i���dv3��O��&���}�O㞷!z�]�$�Ug�V..ܔ٬����J��U���S���s�I�6�����3��6��r�}.���>��$�d��sj��\�LU��N}]�i�����op��Z�����vlP݋ � 2��e"��i�_���pA���)u��eLJ��Se��������Τ���h�9��]�\a��+��@*��Q��`���['H/�Yzg�-�)9�Il�F:9-D7�f<k����|�T$pR}2�vp�N��B�_��7r���2���-�X�S
��h����*�kʆ������b��)81sd5A����UpR�}�d��V�T��'m]
���tؿĶ����l4��Q6
������{�����KE������m"���j>�V��^�� p�,y�|	�*R������1 ݒ��A�զ[��C-��i��#��Iã��`|1h���a��b��U�uU`��g��cc�w>E:����xW"W���h5o�Oit,z�;�ݟ�=�h1��H��7�(ǸG�Lf�������*B�^I����s��X;u��V��k/Uh�[���d? ��O����6�Ӻ��D��|�|-�N=��ʖ`�+��+��T����!d�ބ[���E�r7"!�a���b4_楤�r`�OI�<��O`����Q׿�Q�4�d*�/�ɶm%���DH�ҖN��]2�͒�/W�f-7���%̻�������V�|�6�Gl������]�i��nU�؄�-,qg/�S��"N춍ГWژ��F��е�09��#N�&�\k//�Oy��GJ~6���R���5[��d+_� 4�@ݟ�S��nS��X٠�zf�2�٣}��90E���"� �/B^T�K�;��L=�3d��T��I�q�@D�J��X���[ζU�%��z��H��N�v��.It������G�KR�/_G2�͢����2��C|��}&K�xG�h��S�����B�s���lf�q��)	n����+��g�p�"� ƨAV�N
�o�t {���Z����pI�Ń��A�
�,�N�!�9�Kt��#d�ܰ�̯#섲�K'\;z���5G�
�~��!�s�kW��&4P*ҁ��}��_y�1�B�Gu���0�
��6��_d�Ο�&� ��;5R�>O㲌M�mh��
�‰�̦uHs'���GMV��*
U��[+5�4Q��GT';���ܤ�o3��b�4���3�Vl����T�e�X{k^B-�P��B�P�/�fD�2�J�OۂUȰ��7���&B�I]�^�2&s����B�	-��y
�N&�9����4��/>���I�}��z�wU�=�+�T���g��T���!�Υa�EOE��߉�[-I���O��dY�2E��F��!�	Vx�0
q�|h���Aꨇvn@�g��?��v�t�;,�5�/�r]�>;��te� �A%O�����xg������%�aS��-����S�&��缝�,B��Q�AP����SS5䍶�"b�{�ﱯ�$!l���ia����L7 �n�D��FM��I�݌���#m׿*��jp@9�pϐ�B��w�7o�� ���dt�>v�s������e�ޯ�7)��0̓ҵ�I���;g1 x>���%s�친���q�'ɘ�}W�W��tΛ3��F�z�+=���T.a�&!1�*�o�=��!���l��ں�Y�@G�d�C��Y�l~2x!+lM�C�'��W늙����Ӷ��~Yk(�Q/�̘~|�ub�'(�6���C�>�@ �@(ؙ��Ie%Dt�H'����Ա��ފ�[6���XΩ3��*�g��
�5V���
a�D�/j�p�@"��n�Z�q�*P��poA}�k3��ă�{�w!֑�=��EKA��?0�?_��g�YʪX��p���08��%����|]��s�� T����u##��M�A���+M�ȝ}1�o�Z�)F�N�smA�d���D��Ђ��i� /�h���#�B ���2����3�۾��9�PBy��Y�Ͱn�������z{�uD˅U�B"�+�<g��FU��wb׵�q$�xSS�V�f�!�7�$Ԋ%R�D5g�)̹)���If�팝����!B�\�#�H�����&�?�]/<��霨��H���WHΠ�.�ނn|4ye�-��FWT�>Z �1ŧƘB��ި��$�L�1P84��߻�svsz�Wk��r/���blL��S�k� ��h��������N��h�՚sӠ�k�ol�<�q,o�!H�@�T{���f�� ���ţA
"�*�_���N�T�ፍ���Fc���L�sq�SϚ�������.��_S�s/nnK�Ѷ����H�}6u����[鶞.�6'7�q����#@i� ��Z���:x���ZιZ�B�9:�z���g���1�Dx���$��7���G�L���	�b^�~����c��c�gX��{x��ް��$~N�|�v�H��)���1B�f��|h�t�e��W�+K,��\����T,ͧ7��zO��5 3��-������n�h����L�]?y��	�^z��l@j]t5��Q��v�����8=�ihB�����:��_���I�c2�W�T/���C/����df��|�W�N�"��{h]0~�.��ӡWK78LwB�7�Ku��֡��)\F�G�-��T��[%��!��_ {�/
V]��yѵ*��nq���+O�M�]�LdG��:��v-�J��F{3i��t��j��=9�\*��K�%�E_���\�m��z�(�֙"6!y���J�$�(ځ��o�x|i�q����{�yl�d��y�Y|��>���5� �~��?Wt�9�S�,І�����%���#Ӎ^JfS���U�8��=W�BX��u҂]��u�����@�ip�GIC�λ-�U�൵�?�}�o�c0z�%�*�g5�O޹���il��ERTq���v��3��K˘��j�_f���WOΎ�3F��l��}��K�bbG�-�'_����@��'��M'[Yc|�'-�����d�:_>�iUI�F�f-x[��s"M�86����p=̈́/�;@A�-�p����)$��<š�eU�Dn�Y�j�{�=bD�>)�B`9H�I�q�@s�\��c��擠Y{7Ln}:x�xgE�9���9��� �S=_Q����_�;�z�N�Gd�~�g��4��L���O�&�m
�˸~\B`�bV��?�����z�!�S5 C�yV�������n��
�6c8=�����j~�z�Įx@ñ�P��&�s�̇S������[�/��2�U�sx��v`�ldʿ�a]Zٜ&LA oM�Y�_�;����.S�|7��$���Mh�ài����i:��_�I��%
��/��y�|r`X#����E[F��sŶg�SKkOp��Np��wI��,tZx�cP�����4��æ�P(s*�����7������&z�U-
"E���q�sz�Kx��q�Q߁1�'
�@��uo�2ds��)}w��lrް����OK&�T������ɦ�g�_
��9$x��������S�^A�~5�\�F>O'N��5_@�Tkh9�>��>����j8t��-Y�
	��e���t"�~��r�#��M]�9�c��(\y�����(T8�|%5����<N��� ��J��~�������Z"�����SX�[� l"+�A����,1��J�7ݯƭG]ʭt�"n=�r�*���P}�2M��=Ţ_HN]�#�q
j��l(��ɶ���᤬J�­��L'���}ACLbO��4�
����Y����~��v��^I���.�l�ǃ��<Ej;����$ �Ƒ�S����HyB���8���t�*�F��F?d+��$�tY�8r�jt�2*�4HP���֜���*#��v��;�:�:���Y;-���:�n�)��ϔ�ga7���0����J��\���WX��	�E����Bv� �Է�%�3)��=�v$�a����x������J%�҇|��3��am� �?�7���?)�9�P�%�@wUǎ.v�2!Y�EmU��Rr~m�,�e)��u27}ȔҮQ�s���:oL�4�.i�u`�ۊ����OРӿH�3�2':��mo �;��{�P�`A�+=ڄd�4hg�:��2�ZTj�vl�Mh*���R[-����i����JZ���^<�S;Ķ�G��tt9�H����i��� ��mqȡ���mn��������C���_;Y�����7`��;��T�ڍ�:O:��!����
�� �F�P��v��Ɓ�e稜��-:��F:�$n�"'����C��U˿�	#M�J4e:�� �m�
�(�V`��q������%�Va���<=F��'5��Ϡ�~��"X�| ��G�&��:i�Q�j~���)(ͻ�c�B[P+����z�'b��2�K�\�^L�R��/aK� �h�-�����A�>�;Qr!K�o�mϻ�;��k������  &�z�U��_�j�.�t-�͌�*8�"G��8/���`[!厛V8f���<��%nk��/�6M���(<�ıZy��[��)sA�����P[ѡt��F�V��3�.�;���;�M����s�;=2���=E�v(���=6ɢ.$��ߗd��.�߭᳾�Y3~�N/�T���zuU�p�����~)�P	LpNU]�YD�k|I����M��
����ȴ}���7��k�Q�u�AO�ur�9�Cd�X;�� ���j�@u���'�&g<{��kp\�)?��tڦwݏ�*���8�h�3�i?s�/�XJ)����=���~+��tK��i~N�Ė�g�x��o��qS��5gU��,T��o�Ss@�Q�?��t>���d��L��É���d�������B��YF��ix�+`~q�3�~���_�#��̻�7��|��1���{J-��e(�]�@b���V���G_��r���黥��l�]%D��}�y,P8B�v��ܲ�`�� P%�/�-H����7�<�{<����iU�sK��xeVNZٴHj�#�O���+K"}(&�V"jg�vbG�p���:}��n�9���R�v��Hj�!�<�2I����
��gҍ1������MW�G�'`B&2ښ��'ӎ ��Tu�v���������u6�Q�!'�3���fg����p"��<���E��0v���У;��bV��։NN�]�D�����dnTp<�⪋�:��`[�Z���7��_1=���	��a�d�6S��>���Fx(�sQ�A�5�/���#K�xcwE�.����H� I��D� ̃�@�K\t`;,4��H�r&���ni��v�D%L�P')=oIg_����H�M	[���F���N9��V[�_?��5@�>��ӽ�>�Z��j�=P�c��L����6���k�����kQ���h�`C��3��������Km��ƃ�U����*��FK�<26����F��dTs���ˬ	���6��o���� <�b�:�43�q�!�"����J������o>�oط�X-�}�w��R���ʶ�듓�:���o�ҶM�Kw
!h��/�Q���?��q�Ԙ'���q����>�%X ��ǿ��i�9q}p�3��QVT�G߃^�-�sʡ�4�cLO��P�B��U���1.=v�[�N�o3�$��7�,b�3, ��K�3��2X��bmP��B!^JM�~^6�/������dh	%�z;��ߖN^е�����e��e�vD��)���\��\d�y��:\k��*�H?�^�1H�콆mi=I�vs�Q����e�NU ��Є}��G�)m�E`9v�<�A)�
�g�
V����	���uQ��W� b-}6���0>����!6��xI�"6����JP�����)}j�����p>3QbV�jQl��{0ۈ���0O�r���p��"�W�������y�e=ɓ0���Kc7�*��"��!k�2�E~�Yb´�X޼�ǿ�bD�B�C�J��)n�E�e��AK��~�4�/�(~w�;UbO%���C͢�����2���%Ǐ��|�Ŕ��pv���lI�m�6��"�R���G`����Ի�X�O��
W�Q��yT�J9/,R�0����#O;޿�����d]*�Y��� �@DYx-AFhib�R>�C"��7*�=��AW���w��ZCü1.�t�l���%��푟�7�����̊AMF�R�u�P�S�����B���Iq������E�����Okk_���G/�&z���Y8d��j@��05�o8߷���O�b{׾{�B�ʐ*�W�e�PsA{*�6d�ۻ!{��^=y�t�x)�oR�$�r�	�h��I�E�Y��2�$~���T�&�;]g��5�a�w' Y?�_�`�z9��~v_���Ѝ��z���C�.��U�-Д�\ ����vx�2	���
��jB�fږ�s���V���~��<4�v��.kV��N��~p6����He�<(�����ϰ4{P�>�]"~���S��[����}WJhs)	�׭lY���K���i��p�G���l��|N��@��
�]w2_��F�ec��n��Q���Q���QJ7��g����ΐ��l�L����o��6�'x�m(��#O�;@G��s�|��6���~���Yu��Kt�hG}"���I�����}��0"�g��D���d]�KɝD=w��2�5�rW����(��PbI�0�~� �u�Y�8f�J�O^�J�&�,͙�7uě ��S)���O�������m1y˔��o����L�;1��[�VE��*y3.��/l���{�7+G�1L�fk*A {�4�&��
�Q�r������_[�-�*
�G{Z93�7m	���LqFdO" s�>ذ�h��Iݻl{ң<V~�Zz.�u5>M[p��
�7�3�!IT�I�[�5sf��H���*�".�S0|����1���'�����hL������C''8�D���g�,G�Z7l��?��_t��LCq��k�Y|��>��mo�
�泶���pS������c� 2��T��?�O"��>��=�cv������F�.�3��p�~���|�G�sK/���U|��5�M��}�8�hݽ&ؠ�w����ޕr�\ߦ� �-����K�ó�r���*zុd��?UN)��|��������Za��,JQ���-���*K����9+Ϸ*O��F`��m����k.�c�_x���$�_�D4�������+�g)�!߲QTL;[�$��õ·F`f]�u8բ^��#ϝpg[��=���)��EJ��@H�9]"��]-F�G���`��P��`�.q^71Ȋ�����wv��י��iL̈*���LD���CG����o�L�ϋ�N�&����\���w E�a�7d�p�	���
��*�W��^��pO���x���� ��:� �F �O8�)�c]�!?��mD�����{�=��!�`ޠ*�_Z��F��p���V�B-sA�?�|�����{$lA�*�<2���f��[���_��#%�����:�RR}7�*�YXe�n_f$�*�0�y���ȿ�K��d�m��đ	���T��b�|
-R65�bWi'���h��B�D�zWrש���b�EƮ��&+t��J�E��s��G�#;�lO��%KY�����Ձ��ٲ�R�1��b���գ�d�c�蓚�B"p�r�H�?���o֧A��<�s�ٶ��!�H*��ooC֟zb�	 ��5+(۬�O+_ �&\�5�%ISfG2��ρ�B������$��Cy��V��d��<��Ȗu_Wx����j�O�vf��w�7m���Ԛ!�|���&C��> v��6�P#�|EL� �d�z6��hY��f8T��Qm�}�&�q���K>~S$��?A�I�bQ�@��eV�q�^���`oX�pn��1[�q��ɤ�l���b�|v&w��r<.5ν�P/bv�A�Y���V+��q���=��'��̛c�9`�E�Ƒ�~�����J�I^S)V^�fҍ�r'������]4�Lu�oG#8=��T��J<� �z Y+����V��Z\x ]�V��z��쬟��ɟ�ǅ�ab�v�����K|U��^���ec�)bB�B��g��Z���z2��ã�n'2�-w<��:IT�2�3l���Pb4�Q��+N �?Xr�6~>��[MjF|;j/č����?5x�njP?�;c�p������ˋQ�ٳ�Zx�ݝ����j�j#ʴ����{�a�I��z��&��O��2��CB|�����{,]���:D6���L�m0Ѫ�x��Ӑ잆}��z$7�=���I�G��`���1V���Q����Ѕb����̙֬Mx/ן2Ew��BJ��{�(�`�?��� Ԋ��^L���N%��uY ϒSv�-��/�B�,����xoVE.ȗ�E�0IV�?M!c�c ,�}{x�s�,��A6�)�e~\�%@��
#��:�p��T��l��r���g7���~s%��rQ\f7�v<�������=I�1��N�ϓ_�c�r-�vVP#DP1��Tv_���3���Izowgߍ������o��6���u,��LٷUD�	?ǌ�זgӘ�\V����hzBF,RA$�W{`��ƞ^P.�m$cN��Z'<}C��r���Ψ:[�՘����S�J�7	�be�U�Ic�ŴɧVl!M�p���w��L��R��e�6�%&Cl��N"#��4��6��K��+��O�FY���koz�Pc[1��X��|�q6��G�����a�cg��W�N
cKL<�:GU���F^ɗr�mV�b8�*���5��"
j���2it��
zQ�h��683!8"~��L�䄓�\�G���3�\>@�ʔ�bF��Nq�U�	5��d��F�ag��q��NF��z��ȣ٢UPȺ&���ڮ�؜�N�����W|FsS��^�Y�Ћ�^h�`g�.���8��D@VF����>V��zE$�Tw^:kR��"x�[�8�O���C�n�	��'4qX�j�;�Ğt#��dnz��V#uD�JS2������7���Ԏ��tF���h��G��B�cn08���IX>Kж��ڞ�[��q���1��F�))sD�q�Ԭ���~��<j	�V�O�{_}L;M� kcR�!�E��"J[���D�1$�#�g�����[R&���l��N�+���}��ծ�:�����,����ڋA5t�;	�^�ss�6�Z��@�vB��'��C߇��F��H(WS~���(��,G5L�y�շ�2�ʾ�k��@��k��w��W".�I|��Buk�1���+���i��?PT%09k$!�<�ÿI�gp�Mn�KT�訓�A��H���h��R����V���Z�F� �(�m��#c�Q���p����*c]Z�����	�K`#��3�LHlb��>�g�rlA�C�k3J���AX�K�{@��M!`_����]�<��;�:�����
L@kL0ٞ8�k{�{w"w�	aA����AO	cz=�@V&0Bp�︛#Wx+�2�wޯc��d�k��Xj|^@�ksqXn�
�.G�ίf�}c�۔Č��� �,��Q� ���p���H7����QY�}#���u�ӆ:iE��şJO(�'��-����n�ɾ��`��ln�)Ò�)e6(�~Ӿ��,� ��^*U=6�W�ᑖ�2�o���ڴ,�Ib[���3M�8���6�ʪw43�B�셬�C�n���K=rgMRjת@�K5]J����] �nWBe~�[�j�2y�t��Ε{6:���<
��*,�x�i�8�Q��ä*xM�= Dz@l�X���'�Y@��$��2i/B��9�,E�v�&{2k �қ��G�ʝB�n� "_C=�j}�=�4Jxk�W6a�f��W��Y^�P���k��[r�نO4� ��[9F���x�\:sdI�4��wއӾ�d�c�/�ߧo�/��4��B��u�p������Ys^�b��%%�d1�X�u����B?�Y��Z�����B�EB���{������F�mD�i���镝��:�sh󯏠�U�=N�N��>�AZA����H�n^39F�K�urUo��7����)@��B*R�
�g�+��#?6���H���jR�"7H:��
����xd��;�Q!��@��d���o�����N���]�L������	�a �R��/:3�c4q�O5o�mA�Gg���~�肎/�D�i�ǂ�1�U���\`��d�5ƅRdt�������&mC{�/=���m���y̆�u\�.�0���b�f���dM�#�1j& �ï��ߔ�������L ��eu�Ϫ����U>�&��c�h~m�A[=0�)UK)�?�����຋�W[���X��b�I�n�d$E_\e��'o�>$$�	�U��S�1�[Sޣ���/�ڡ��Wքb�Ӥ\3�7�����w��(l���֔wz2�R�h��d��6ew�)8PJ��	H�EY��l{���p;�N񍛏�;D���5~pT�\�jι 
���)o��%�Zk1A�
�o��R���fJ7�C�T�)���f�u%�İ)���p�5!�qj���D毺BLy�6eEv�L�v��:���h#�K?�0�*2��^N��b�	�8�n}�i{�\m�e>悵<�&7"J�o�N��vpm��`S�$5�T������f��Hm��;�V-����^W6��%��;�c3L4c�d�W/�<t�W'�Rl�Ԟ�\�'��N��� l��CJ]ނ4�P�)��Ͼ��|Be�g�����ŚfǴY9T�yɭ@I�>�H�Q��/i\`�f-�.� _�c��<�>Jߛ���P]�8�b:�����x:^�Y͹^&<2�V�w�X��R�n�W�ʿߕ�	���k�8f�v�T"~������Qkhk�$�3�b|/B�k͗��'��A"@�U�N_��Zk����f���r�&P�v=O��
�����sT
��?�q� �e�%��R�n-�DB�+,\�8Ek�A}l���z�ZG[�̚��������>����_	d����:�D��Ի5"��ɃS��Z3M���r���5e����L?�s̪��^1�6�;����r� d��'��������-^T"�'�zǔ+�p]��Sm��7�����d�Yea�y���<�R�m�3ϣ�l����S�[�߼%&������"^k�HlIm�ذ��֯����[, o�<�h�����ї�P��oPnB��t���u7����x��hjZ�o��y}ey{��/��ā�"��!��,�� ��lmm�y�	���;�麥�3Y��|�OBN濭�eF�To��k[w8����Yr�\�N�HO��|��<%\=>�fP�8(U�c�p�P�0f�G�6m�	�_�H��j���:�G����w���K���M4��M�(��S:�)ҙ ߦ��&p��L�AA,�Q�5�?43XQA�gv��Ǐ�W�����@���~`����z��⯴Cڰ?�cvЌM�2���l#A�xs����ǋ��6���U�j�/�m�Z����08��oddH� �t�� ˢľ*$�2JU��P������ïpt�En�+�.�E���->ѝ��1<�y�}����1���:�U~�NI��,�faLe�)��(Tu����&�Y/���>��N4���g���"����nIg,�����K�Ű��~ܟs�FR�ST��#B�� ռ��7�ﳅ��9�-9
I��"�������� �'~W��>M��������H3�CVX �|R�4X�	'�sP�F�U���L話v�1�3j޲E�P?�����`*��3f��?	�,F^i!4�/kto�z(���JHX���Ǻ��ܕ�`sQ��}��l�e�k��%���0�����\_ްU���cv�|la$��QDC��M���d˜@<�+،F����w��";�\�d���X�ԩ9Ѻi:��md���Sp�=��.���dkV���w3 hS��!lF%(>�@����X�Vr�פ�� ~��T4��^.޳-d+Xvy$��&��6�8�@#Mf!�Ȓ4�)<|S�I���M8��z�z�����p�5Í���'���m2L�c!���6�ԏ�Ϟ:Z��_Y8C���e����8��&_�r���	;c�U����lS\��MXST}�:����b�qs��t�!Oڨ�}l�gb����<p0���߆a$��p����3$f�F���ٮ}L�IlD�K��0yw��o���K��ÿ �:���1ڗ�5bf��M�u�uH���C�H�Dw����$�� m�K�u��=$�J�zXB���u��_�C�6� �2��[�t����zSp�^K�	���W��Vx��+���$,`t��;����<U��8��h�5zJ�sh[z!�����J9���r�n(Lc<�y.��&�T����U����?ĉ��vM�]�`g`��d:Anh��d �TW"�d"7y]ټ8��9b��k|��.�Rس�	��#�C�eҺ�?��zS�j���g��zFc�!ݠ��Zw�vHٌ5��D�J����OT����@�� �ļ<����<�.,��[Վ�����z�Ƀy|�Nƥ�w����ո�D9�{�z{ �",/�)�Ż6>�>E�\��T�*j~����^,9_W�ֆ�լ�P���E�30�=M`'�đ�\�囇ȣ�|�g;ʑlxvY,��b7pY�$��\hG�nU��
t+Kk��(W�� �U�2�r�VG�Gn\]��|?�M�E�ȗ��6�^�j5ZvV�>�H�dӠ��=�H��J)4-۬�UÁ�EP��t���)a�D���[V���5��G�L&�l�(30 M�g<I�:wZ�5�_�>�h1���JR9��/H�@S+���g��Q���C�	�b)ұJ��i&p;I|���#�Jt�<_ʪRV�5��G�p���8��,R�D��טN�e���̳��wH�!u��������B�;|��K=����jgje�w��u��e�����g�$�l޹c�@�&��Cy4��"�kIAvf�����c�(���ş�>JZ��C��|��m�-���u;�����Y=9{���P�>�x�6��L`�
o�_k�ʧ��
����#G�����U *'�����V���Qi�y���3����H�A������X�_a�	@kǃ���]T��u}|(���I��8tː0���1�)�*w��6�uy��G��u����=9��,�J�]�žu
uŠ"K��W���il~��4k��$��Fp<tg4��M��g� ^����@:tԨ[�?��6���}~M^���ϕ'U�:���YK ���A3׀��E�u��M+i1_��Ur�����i�dB����֠��j����������q�\��q�h�q�!�H�N��P���x�2�n0��i�$��ץ
��?�S*͐�}	�G��Z��{��J\�:,����U��FL��{[�:���u|gIa��AcV4��;��g9a�u��#���$���f�,d�w��Ov��x�َ���#���ڮ6���,p���7����bҹ��5��.�v��7�T\�y�����k2�|�5�^�6���z=�_��L�*9��o�5���B�7�u8�����|P�A��x|]A����.���^';�v3��Y?����v���RCl�e�#�����byb0T䩹fyO#�����b@J�����4yrl.HD�qESx��Ts��"�L��P]�4�b@����XfV��^4�O���a+�;���s1l���w�Q��<\��k�B�r�Dٴ���T��lU���%M� IA�ߘi��t��qm���=�"�hPC^VHO���"y������#��w?M~����BL��>��&����Y6i�j��ۦf'�ۧ%?^��ƅ�s��MG�\{�`La^�_8�>:�K���!T4@&�П�<㡈'	C��o�5$&�4QՌ�סGN�>"e�ܹc��{]-
���s��ފd�۷,N��ڬN�����5tgA�C[���=��=�4l�ڞ$�͔�6>�ዖ��-j���Ϙ1gR U!�%��p:��=�ܑ}�ǻ���׻ zF�$h��1���~k�{�	�rKGM��Z�PDWnu�����0�^O�<6���!څ#��j�)$�HyuW$�B��%ߥ�X�pTh�����-�+�Mk���k&?:t�9/�nu܆9V�HV��R�BGY)N�{�^|:��k0���˜��2�̣5�f���X���W��ӑ��>���*3��|	��n6�#�$�%��q�����@��'_��-�?�I�Vk>k���YG{,1��߫#@T�'�ks-�����a��N4��U�����c�/�Ͷ�.��EeOB�����D�~�ͪ��yO��W��� s�],��e�e�,l�m�㙿u�	?�a�K|Τ����v���0�j�3-��G9�Z�p�F
��P-�-�_�D`��;9��2��+��쿾[FxR�g�-:o���{V�$Ý�Gҍ�� �Z>綌�1E���T2������qJ#���-c@�sV`������Y�7�!*��K���|�?��U��W�0�}��h������Bo�j��փ,r�e�(��wQ/g4�;\U�O�x>��,�|����;��Ҝ���7w�G�����HrNh0vP�>}n��Ƥ�KU*���&S���$}h���y�Nu���R��+�o_���|J�^�����/NG;��e�:0�� ?�z)��>���"�fjɷ?J��>/�<�����	��%Q�%j6U^���gKH}!5(ɮG��h%] <iaV^�fL*e	�#�K��h�A����*M5�n�׏�b���>#�����:���qy_���W�&�&7��n;���H�E�Q������q�����5�Injf���˱�^x?m�^�7��&C��S��_$kk[u���.�Rf��m7ܒ#�V���V��~H`}��3��U��Ղ�� ��\�����"�q� >�i7�cƂ�ł����鬭Z���=����4�܍�����D�|MˁXO*�P�, A<��,����"�l��@Y��ԯuTא�Am�㩴�[#����l�Ϭ_d5��(Te�O��Ib��i���7˂�m�9�FwA>�$O��E��[�"�vj��
0n��YZ���c����d� ��죰���\t���f��ʓC���$ˀ����ec�1N��Q-"�����{_%6w��{��{�q��J����2��U�4�ˎZ��xp���hR�CNs2�r�B��)l!;��C�Y$����5�[�+d]�t]��d�X��򤝣H�&#1����|TqK��B�_��%ͪ���0!i�R_�:8ηk�~
�Y ��i�4����ˁ-k��	�q��Hi���?����Y�f�I�y����b�6V[UǸRI-��ZO�#���+kG4���q�H�@�D�K]	���RB>�Qgu�m���iG t50�Ht	B��s�5LWټv���T��`1�����7�VPZ��q! �)��XK,}U��ć� ���*���YE[	��L�ۊ��S�0Ǩ4�W6[�u�E_���Os�i�s�؝�4����r��n�*�&��K�xN.5Heq i�ğc��ǘ*XAAvt�\��w;�`�vSG���� I�z�,���d�&9�|���
����?x��BY���  >vH�CY��9ˢI�w�4A!%�Ryo��i�EE�S.v��!�%ӷ���>}|��nXnG0~)p���*N���zS`���ҷ|Ĥl�O��k�*�E�^�M����Z@�`k�`���z�D}6������H@U���>S�Ⱥ�)���V�G#��{HK�=�Mr�ĸ��'P�HҼ��q�\p��D�gNe?�s&1�H,O�^��N%.l^_�3�#5�{���z+9F��'�`'p(�Cu8Tf:r���n�!��'�t��Cߺw/J�=9,[�H�?AAl�een�6�:&��N�� �����N �R��_F�L�c��î�oB����G@��� |��/����jnt����/�a4br�L2�A�a,E��e���Kt&�΋W���<\`��������$%�J��1�){�'���<A�������� f�	���X�="w|�-�\�v4<ڃ)�}���B�鏲D9�6>�_V����
W(�HZ��m��Z��>�ީ�"}zi�������{[�j���uof��!��F频����C�Ĵ��G����ms>�{�Bc�S��∝Ll�1zO��U�f���ްV>�髦H���]�L���EH�j��?�s�J0�.S�dC�n�1��ǉ.����l��xQh;���K�i%:�WȦ(k���jb�S?O�i���Ǚ۾X�g��P�{����������Y�'��~����R!����jjj_�M��ų[��+�����0�TU�D��*���PԸ]�/�h�j�)u��_�Ƚ���Ǘ=�B=,��"cƆ/5�7���-���f��uCe���Z�H&&~��C�D��gݤ���������HPK�����-�E(b�'���fkS�/J��-�� �\�0�_m"��#.�NF��vc��Z$,����s��B�- �a��o{��#���A*/0g)|X�`��sP�����d�w�r��G��k\����w� f��:����k�����M3s�v���&!�ҵt��g�;� �m�� u�[x��Nr8�tv��]Cem��~���	}n'4�PWS4QH;�CN��l�;�֋4ÿP"��(��	d1S�X�ii.��..B���SS	�b�\����x��3���	��VJQ�o��t3B�UWn�pk�-�-�]�Β�����m�"as���ilw��@)�Q��#}3���m��_`^$sw�=\���/;�Y7�8�8�����($@7OQ�����Fl�O�@�&J@<�tߣ���H@-��u��!;~hʎ�V�Pya>)� �S�-a������p���"e��]�	ӢD��L%�~r���S�'1�V��:��Nr;m���FSZ�7�o�x��޿�o��GS�$���><�G�ye6z�4���[N�X��?m�ˎ���z漎薏%�!�K}��jJPyݎ8�z��.LŗU��&p��_
?6�29��$�a7�Dy�R:�Pr�3N:%���.	T[�X-spba�za!�q8ٜe=��s!RM β�N�j�����Ee��k�T��跴J�F��1{v)#�R>ۃ���F���Q��~$'���/�ˎ�F�t�X�+ȌJ�a�2�,�=9�%�z\�u��\�^ܯ�TpK]5@9�cj��LU�%&�Խ��g��x���	�j��exo������s^Bt>_�P�h};�k=���|�k����l]�z[�����k/���:�j��$|�=Z �Q*r�7?1�A�4f��њY�1�"	n7�KZߐa�3����j@g�U�V�����nx��8*l�ߏ��fqh��'�a#�ն��J���.BV�Hv睘T8N7�}�bf4x�j,ܔ��g}�C���-3hM��	��YRb� �>[�塤w/���>)�}�����k�,�߂I�̙�L���� ^���-��ɲ� ������1��ʍ^���X���3zƬZԯ��f�����BL�ۈ���O�nz)��4�"~e0s��������ӡ��mֶIܽ�_�Q
����ٹ����~��ΐ殺d@��8c� �
)�	�zOp�TÍ��e'��毯��,�Y�!��{e&
��KNM!�Z\C�G��r��~�mN'=S��3l������W|����><�^MV�����D8���F���� ���N.�b����s�ִ�v�reX�2OjOICx��+�3����i�@/���GR������Aa��!����.Ѹ�I3�,�>ߝJ,�qs�7�E.��&�ⱓΨ:���#-�+��@���l�?��s7�I�%�F���<јy`)c����"�)�
�-�Vl\HS����"��T)v�!��e��{����^�Z��x�|�6��b,]��D���4�|.\
7x!Աm>�_vO���6�<yB�.j�g|n�nK��r��U�J�a2����Ѳ�T��%�p6��\�ʮ�/�ۇn�I�uQ�d�l�)�Es-Q>��۔ذ��F�yο��eK.N�9�Ґd"��z�%wP�$�I���ʕ:�mO���/��n/ϳ�D3^���=���x^������F'^Ek���M�՘5=�=���=��+-$�7�~N�g��'{^���z�C���B�m��f���ۼf�	%������ًWU��ǭ��O�ت���ٕ̒7*\_3r���;�xi4h�ŉ�t{�DB�(d�R���_�)dq�%Խm�`����yl�a*1��[�]�����z�1�?^[?����-DBD��efK}�z~�[ %����=00����?k�����6����GoH`�%��g�������1]��3%�^i�S�E���)9{�:uu4^ �IhEE\�͝����"X\u-� ���.�Ӏp?�)�����rF ��DH0�N.G����..j��M�9�;E��t1Q��Avˬ�����E�p�R-�p�˸~�	��6ޘ�\G�"a����k�Ș_ɍz�+�2�w#n���![(�j@��w�f!�y��7�����P�H�W�RU_%;͊��"戮2LY�B���!�{����K�ې:��皻����n:�9Ğo?O�wML%��� ��d¨��ͭ�yg�`�z³�[�S��Oo����'O;1�qwᑱj��(/Ur�Y�H�@ZH�3/w�ZH�֔q��X��lLJo�e_��>�-j�#��ҧ���E�#va��j�z�G-���4"G��K)\^�W��f���&����~�&���glD��S�����k�E<𩮎x`���_^&�R@��~e;>"�o/��>��V�Q�K��K�DS��z��(�NK�>�3h}�����ԛ��caf*/�<L��מ�L �r��� �ex�E�����F��v<�7|���}��˟$�դ;I}�&���hN�o�u�Dq�
�͓р[0�{S�fi�a�jZA/�Z��t3�pR2�U��י6à�\���z�,��H�F.���DR�ڧp;Ux��e���o�S�MJ���~/�*P�MRqѹDV:�<$���_^��0�1ۗ|��J��6?�vA�U�6��K�ʇk���+�X:m&�˽k�TS
�DLx�����v�S��������p�k��L�ǊOĩ���QB&�O�lQdݒ���?yd��n-�.�Mt`E�9���^�Rdα-��j�^^����5Q�`�T2"y� �$V&`b�׾����߄�`�������D{ǵ�������2ߪv�Ca&║����lPzO	�����g�hH��o�f	�ܘ��&��@�:�A�.��gb�'[�:ڶ�e{��Jb�
���������C��jP�]C�7ȝ�����?v�Qt=�78��Y,6��*�[5��M�<��T_�g��$�W�����1�E~g齦���V������|�;���f�]�m�T ��g�R����=�����2�ǊVd��r�y'x�"��^��S�)M;:&��.�@��a��|�b�|:�`������Aa�W2��(%��֪db��O�ǎD�HտS�A�svF�W�*�|O��U�Ǧ��.�j�'�x�ym\��t��:���Ȃ���3[�J�䎊D.��X���Z���ہ�\%� �
�(mA��:�9�F�{@�u��1^�zUp���h�cR���56�0��eb0x��௖�W��"n��� ��Z#�8e�B�9M78�rC	�O"��US�B7 ����1��x��w!t�k~oA��<�n�oǒ�$�w6�A�;b���^�뤖��>�:;өTϒLph����HD� ��mҫ6�3M�sv��8ݹ�%h�h� W����Ne�bq�W�x�6Q
����F��Q��h5^FO���/��֒2*	��
����?Y0�{3k�Eo,�O�H�N%�z��Tz*�_��MM�T��X��&��y%wo\�	�V�C��p��b�[��D�u�TZ��� HIR ���E�����	\����ݭ�A�a	�9�����Nß�w�.l�Y�j�{������#=�ݵW�n�G1�b����������!{�@���D�S���sA��?�R{�߂Z��si��d
#N=֜�ݹD��e��O�O�ly
1U�����;�y	��J���x����d��O�~}��S��tea�s��:�+;T�ˀ�aTf:0x��7|�%�?�3>�e�R-:��V��E���=Mk�c�����G���E$�$�p��"ђ����Cq��a�W�����k(Z�%ώ�u�rM[�&���P����9��lA�7������]�p][�rA��������B%
V��F4���D��GO"+ NK�ecA	�`"���ts�*��l���Y�WMg���:NP�hOF���be�}�[
��ϐ���/h��GVF�e��@V��\�& Ȗ�d5{�K[��X�|m|\�Ї�����,�D�� �V��h�*x�u��n5�g��s��se(�iZG�BՠS�!C��g��eU׹�z%%�&��/�����/��1���.DiL�����64�*ͪwݰg��;+�i5�X���a^y=(2,�L$���;��!���yJ�Y�>�Xt�7���oLQYf���p~��	G&W�����t���}�4	�s�,�c鞊�c����݄E��4���2�'2�P�z��o"�BO��9�tڇ��\�t#.X:%�NeIko��}��(���Z����P��qݝL��ɗ��m��\i�$�g��S�R�k��`mܧ�8��(GF�_����0�:�:+櫫�l�GN��<�܏���������Nl1��t-cKU�}L�e��<��3DliA�D��P��H����2k���5��J~���m��@��B0�C�(�s�?H?�O?��	s�2&Z�ݲ�4��0���*a\W7*FS0Ľ��A���4��&8}�Ċނ�K�[JU;�T�{%��O�q���{o� eܒ����A�ۉ�4䅇1��G�\�b�a�B��$ <~@B��?�$�y���!��'�%�#��z��Ѷ"&lH�?aL���)s>�3���E=���w��8������P�7���'ڊQW���!G͊b�l�Ԫ��`����[h�2��1����)��3���0v
Ajz2�PͿ%zRMZ���yF�4xRR۬�ߋ�o'w:?ZY��-lg������z���e�:n
�p���'ϨPTV�.	u�����RM�{��{�Ŋ�X!Iт�,�J�Q*�!�	=�k	��Mku(%d�g�̾��i Hv�F���H�TW���G��	c~x[P�@��V���Fo��ʶL3�B�����<�5s�bJF��p���^܊��\^�3��8��6��ȉY1�sy�K�n�aH��Pئ�]Z������-� �͍�|ۉy�Y��D(�~_|-�Ѐ��^��!d�>m���`���,�M}Y���}���xm����_�ڝ𺀲�	K :���L������O��h�͢v�mb�l�雂o�)�#��
k��ËH��� �&R� I�XK��|�8���O���	A�蒷��na�|t�!�6�C �Y���V���'G�g�Lu^yDM~����g��B�򧿧��v�Ow�ƴ��$
����`�.�������r(2����:�����m6do��Y}������\�i�b���ۚ���:\�cT��!�&2��Ra$+ŢuچvhЫ*�٨5t�F�ފ&�%f����h���-1n7�1^<x&���V�:[�Lo�.�)��9L�6�m���"�\���M��t�Mv$�Umg1gټ��  �<�?���~a�J�SK�!7��� SivWtʀ�^\]1��MD�$�U�F��g��ɀ��Y*~SR��c5ݧ���һ�fn��F�Bk����y�_��;�̰��7�U��X�\�\���W�CUVu��V�L���TY|��wnc�#�_��g���u�L)���M��\ta��#j�H��]�ȹ	��m�Y��{��b�i�����)�DR4,Pq��"��]��$4v�ڨ��Hж��A� ���iH�H���ٷ.��O��<y��w/�-��f���_�k�����E�����Q�׼!"�͐U���;���`گ*��}w�}��awX9V���83�m@�VH,���OM�Ϗ��)�J�j�vV��d%b���=��̦�g��G���sl� 6aJ����0S�(xQ��,	B��*Q0�����;��ˑF�D!�;��a� M�{�֥5?2Y�����/F��E���%u��Ns�nh���T9�
��.w�\;4�#�μ��X�b}�}L�Җ0�K��M�oZE�IӠ˘NHSkJ�Z:��a:<7= .&����ZwF��yoW^��B,��57d�E�y���B�.��U���ʗL���,4굯m�m'G;�/�B3�o�S���p�N&���=�/�
�9�I����𷭇냧��<u�ף�✷�F�6�ɔ"�ߠ�/�������~A;�%��X���Gw�I~�AbȘ=�J�ˠeT�LpZ'�M4b��e���K-� �RH�+���]R�?E(#��m�JL��[ѝr@6,ϚZ�3�0���մrQ��`�5P��WB�<�>�C+XW��Y�����ZQ��>?�q\�.���}�Nm�I9�ޡ������I��I���O�Ymt.�J����O�$ՖΨ���+i��).��	�߈#1��oMD^�lB�M��#�(�j��B�V��~�TО�"���L5<���o̓��|H�#R��D���K��1�QS�L�/L���(Q�oV�^CfB�l����]a;$�iM��W��C��>�e^)��%Ld�R9�xA���;� (X�b��.�'����ȢsKs�-:_J(�3;�PO�ɍ�7D$�n�@;���f�Pj"���w���#i4=�O�6�_��`����ܹ~D���P~�6V�	�M�L]'I |�}j\Z� ���[��=_�\���<��q�h�%���4O#����֢�">�|��5�i��C���p��X�*c�G3"�[�4�M{6u�V$�B�I�:֣�yQ%�7�y�:����DEe�ӊ��v��#��%:�� �� L���� B�����b;���Z|��N�;,�(�����bxD�/����0�\���l�(�Sv��^T9aL�ō
�>�J:֡¾V�A�o�-�п���O����oѫ�ڸ�'�:I��ed�#����qL�0+���7�~3�VĖ�蕫W!�b&�"~�n֚�a̙@���_'ǹ�ZÒ���2S��<7�νP�r5I��9	�����\��m}��r��Ί��f��M���'�����F�w���� s�I&��M�v{$'���V
zB��(YVUn�^JXO����9*�g��)���=��b��󸋮p
��a�0
��Z�U؉��fZ F���I9!v��x@U&�t�d/n�ӫ쫭��F�������¯|�Jg�4!Y�Yz+&$�K{E�����W����w��8lAܭu���5z��X��.�A��D²��ݭOVs��%Ɓ^��G�$�A�/�p2D��l���i��9s]xA�T ��x�rF�A�&������BN?.���g�i!s.��	���QGj���ߓ��n�����{���+���,xJ��r��!"�`yt��j�+�Q�#t@k��M�GH�}tI����d�Si�-]�����=*��X�ds�)����կ8\ɇv]KD���6��>�@�^|����#%�A*ː�ШD�����c�R>�vF2�AU6,�Y'p�w�J`���l7�_�Mn;���e���۪��Ԩ���2Ǐg��Ab�_i֝2���[��Vۿ��ɣ�u�B�}D�И&�!��Af�����=�]'�ո�?�$��n1Mϔc��o�.�b����2��ͼf�@��b+�ŧ� ��%�P
������Co�r=��d�p#����)�p�k��}�l�V[���&%�s{�8�Ky��H�����xN��'��u�V�O8�~e^j�܌��J��ov7G���{g�q9�CͿ~ƽ�8d��z�o�PA�$�^��͗Hܳ���Va�OM�t� v	�|W��~���+A�](�5�&D���%�x���P��2��Tv�S�OF�>W���[E1��ϝ��4J4���b�X�.&&Kڡf�#pD2�ۤ�_Р��	�~��J���ڥ����t@�$���4���4*��O�ZH'pu���}ͺ�B�%���\�(	����P��]I�#g�]'�gUI�O�#lq�z�G\�}�XL��1���G��6���x���s�32�H�ӗ�c�X�_�|��!ژ�v�%���]�����0�N�!P���b� ����G� ���p�������7W2trfL;WM����X��ђw���&��i��_�����4>/��gJu�/�UJ73p��v0�PY4��S!��P�����4~ǗQ��(h�IZ��͏�=�n("���ۢ0��1�;6sW	��L�V�s��z��i�2��#�	6�T0�^5%!3�p�L�Ry
�H��h���������[ۛ/$R�S�M:�}w�.�c�n�I�N%V9����&B:����;w�I���O��A��k�ڌ������ ��rWJ��}P�.(�U!a(�c/?�>:p D��?Ēe�A4�J�b�@F��)���%��<x��X[�1�o�}��L��&�9E�����,��'ENO�����#@'����%�Y���n��^�П�w�b	$ߤ��|�IM�\��
%+���W�{��\�s��ƒ:K�k6�`��=9�,qt��FM����6�n���)��p��\5��+nxjA���\� bki�d>,��ϐy�W����sIX��.jV�"���)��S�����i��'�zlƵWBr�ٮ�����>�x�e�>��a�ܟ2'����D�a��J^v<�7�iij��u�g��чЭU����ܖ2Y�ZX{?��S�[��y0ypĨ�m�9C7�ʹq�)��0�U��e& +�t�h�K���/ȱ,�����]���6����A��M�*�W����Y��t�,��$ 
��"yD�bPB�*�ޮ�(iC���HlE��R��O��/2V�XN˽7z:M��ɭ��$C��]0l�DVr�
F���uW�f'-�����#�
�k���W�jj9�v_+��*�B�pe�׆x�/�ǟ �̎��ηѧ���7�k��e�qF�	���-)�B�L`�j�ِ��>8�� .ce�Svc��ٯ��/����M��a��r�������2�8(�#�<�YG�ٴ���c�����TU�}�,�ϱ��C��$|�m@u�58wVks��8�5z�j˙��[���K�ہ����COkR��>�<t���i���7k�I��:vu�n������(c�.b|�j6�[Џ�2$T��"r*.Lچ��U#/��Y/���
���|ҙ��è��W��̈́�m��o*H��`r���M�I�`�*:����<���f��\�)����ۮZ��������Zj>�yl��]�0�
�5�Y�9�ie�D!�`a�t�J��2�㕵*����nh80��2m�U)(I2� u�	B�Fj@p�K+8���,D��/8��<Xft����<�obn��u{O4=pǁ������8>Gt�X���V�j �YƼY�&5ZՅd�^
K���WH1�/nk�S��W�I ��}�gKg