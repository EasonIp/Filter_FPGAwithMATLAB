��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�x�W��$�oC�Lw�S
�,h�eԀ)�CQ�_���o�E�'+��l�����qz%�[LըMū��ş��Yz�g�#Vz���E���_�����/��'�w|g>ѐ�=dC6����	NwJ!�
�PΙq����F�<hŚx��#��aT��R��`v����*>wEb�3�4��	ηto��b���RQX_�?+��M���C�ӛ��/�7X�FՃ�Bq���F����9��	X�\|(�-��:j��ۏ�,���$��,�Y
��c��9r�?�1���\G��L�T���|Q�CN�0���cJ�H.��3`�H�:sz�+�+�:	r9r+AY�[����9'�|�]�wy�WX6>���S��:O�0��fӭ��ҍ֞���gUbo�����`"�jyᛁ����Qy�J�k� a�q^���;��u|���܃Dq�� t��֨P�����<w?%X��̮T�\��i�n#�3̓g�`DcP��J�*M�*R̺	�+',C#�ڎ�>Pm����gE�Zқ84ud��Z��LmQ_+�f��sW��|�7��rX�\J�'q���v)-�0�t��Z|~3����~$���}����,�\IW'����X`��#�l�bJ�h�U�MͽӟVӎ6�Jg\��y���3��`t5w��?.�����~�Q�D�Oϭ�x�fZ;{��ǔ�J�	���;e�e����e���X���m�p�H�<�-�OBo)�<�P�X�m��ט��}�ƃ�V� ���k{������:΍�Ɗv`_�pQ���?K�z9�\��N�����p�_R��F��X�>DZ���B�{�7<ȁ�F��L�=��QI����e/mf�sW؊�H�s����4�#7��}V�w���,�x�#�ꅤ7�����0�7k+�~�O�8�Ry̶�C���M��kd��E��1�'�E/K|Μ�Ty������U�$�߉��LO#U�y�s�qdg�r�Ȫj�q|F2O��y�3kHo$\QЋe�t�D�F���%��.��>x;��8?ol:6��u��6������xL�×Z`ό�,�j�L��Nΐ���l����T5�
�%�'0:*��S>���f��vc��f�+J&W7�"v��o.�^�t�"��Y/��Jc�.�_�0sh��#��"?�He��ƹov����86�4�mW�:�z`�^���^���;&�>V�Ў��#� et�ͥ�!�����ml����=����N%``�9��})����&����3�B�
�c/h���.Ӎ��=~�:���	=V�]���hIb焕��TԺ�����SU�9��z�Bsއ�lS�w"nq���`��)��P�׊�Ļ��}s�h�@�����v���h�H���Tk
���㽇���Z�7�=E��r,ܠ;�q0-��Re���W�,r�pꄑb	��qD�6��z�F�X9����2zb(��V�+�����>��e���(ѡbM�6��(�V@�fߠu�Ə���WD�m�߱�$Y�u[#h�z~/G�?dgʙ�����_�UY����<R����|�`�$1[��"�F� C|ۭ4�N���L�sW���fW��X��y�b^�_+��gC曊�E�Wt��1>���;0���߂b+�²A����\&3,�YsJF��P���lq��ɇ��v������
}=���*�'�"� ����y�z?׻٢��7ʋ�mb���`���������ɡ�G�&Q�ʺ_�3�� n4n�&��n�il���&fy��O�K0���cK��Ǟ�OwVF}��^�6�ӣt����3EsR��̪M��g��d��m���FDZs��>-�-����T]�ʨ� *����.E�!�>�A
ݜM�p,	&�x���Z�&NʹX(vr��i��3 ��PJ����V|®��<��0��dh���p8�+��R��Ԉ��lO�i�0e��`�`�a�]�N��V�FK&�?�VD�.U�n���76!aA��T?�<E�)4���J��`�Vl`�wEk�H�e�7
^��ޣ���m=�/"���L#� G���p�P�c�mm� ݈ꝯ�@<�S��������������ī�:�|�8/�z{�a*�:�e��IE�.�v��L���P&�� G�|öHEH��sܞd�G�!�+�c�ܢ�wCe�*�#VxW��?�*��_B���o.3
_��<��_�F��+*�qx��Vy��a�1?e⋅]3�`z����w��a�biH��6���4d.��?�Wh� ��syY	���ܖ=������?��K8�oױ= q��X)f����	��䓑�#);1�X����@��b�Pn�U[��v����w�
ݛ�sD���)LNT�N���fp�S����0�4̍3i�֕�3�:��m5n(�N��4R������tpc��iL�yz���Б�)���ô�	�-�*u$$�|����aĭvYR@���)pH�L��X�{Ԍj�`��n?CV*����Tf�'�S�/�5`���b�}`�caFF�g�MFF5[�{���;%{^*�79�&��8.�`��AY+��4�މ�����«:W��_6*���bD�"��Ƈ�F��p�$���S$����F���E�_��[rsBQ���>x���IAe�fT�M��Z�qO�
�փ���a��qǉ��M�<�7LY�Q�Q�"E�tq� �h�Z��Z�F��uE�#��Z��G<�|��d�b�걹���!���'��Hyb���ÜF|�f�h�u��b�7D�hr"sd>�t�)��\3�;oŠO�½.5������X��p�^�+��6j[��l�o���:}�/�����}�ک�Z<d�	M���*����`Q%A"��R�+�(�^��i}D��tٽ�~�iQO���I����e��3D\����6Y�v~I֕t���z��W��od�^��l��M^I���k�;���wC1��O`�E/1G�3[g*��ed�l
 ��؊�O�S�(]�|q�l�v�Ʋ<�^�M���phb��4+��~R#�oY�f�|A]\��$I��2ȽL��O�[�e��*/�����M���Z��@�w&�,uT��%�� �i�K���xp;��&�t<�Mz�lΉ!�����oyfvK;���a׿��2i g�P��7s�ja��@;�gk`�A1�k��V�}��%���[z�K��ڰ#����n�H��
Iz�=��tD]��v�#+�F�>qc%s���bZ�?ռG2�Lb�y�p�*���Ն�D�`1��&�g =�|U\��\O�q� ���]Y�(�9�T�Z������,�8D��!$b������顕+�A�ْ�ŕ��"P�i�ȫ��e�Vډ����W^�v]&?����:�}���	8���V�F�o��Y{���1��;�G��d64#x�K�c����>�<�����O@�Z�գ����@pY ��u��=?�GC.�����X�S="�|[2��j��\{��G�?��5hZ�����$ܲum��ϧD^t1/~���*��d��Mp�7A���uy�{�l?����������ɻj��r:��*SF��\�J��U��K�z)i\��<��3�i�`/W�^ǛҖn�oRI��&���h����Ǯ�)�sye᪌o�ϵ�k�^��3�R�;�<�̣F�6�(�Kf5����i�4N����=$YD�
k�a��R��}:/�U��<��W;i�$h�٢�!z�$-5�ꔀk����.|H#����{v���#�)Kl��^ͺ0��	aty����7zʡ�^ZtdaS�a�Ǥ+�*�R+��3��"�1�l��p���"������x�r���^���������ͅS����~����ѣhڍ�0]��"��˫6��p�)-܂ �Yq�,,�\H]�i�&�h��� `�-g<�T\���ll�j.�n�ಲI��k��_�zv�������M	�^�%;�^�$�]�;D�GR�֯sRQSB�I!�.o/��3V�R��<��?�c��1���g_O��i���A{�`8HJy$�c-���:�n�����1Ǳ~��Y�6&{����7�wX_�.����f�e�x�]>]�����&z���Fr��j<�殢ҷ��"�!�-�o��MY 1����"�2��T�l�̬�.*�vf�3���4;l��
$C�2�M�G��	��
i)�$#{Ϲ�������G/�1�W=��4���H����3�s,������N���A��P�Q�49�
M
܍�ъ�������z�?��9R�*f���y^���͎N�:�L�.�y�F�������v��_�W<} \�����$��{�!�=�����z��'y�D�ɛ�K�̈�uL�3�m�N7�PD ���;���	,���r�b�����>�gm�>~|�ђ�@Y�\"��&�L�KfC����)f�h���L���y	�[�����e�Ц�����3�Þ�R���T��A��2�7����|2�0KQ��rnAm'��䋶t�J�L��I�|"mmIn�a��9����09мߚ�Ϩ�>��~��+�κ&�/<|�j�@���y��i\HS���a8�V�|�xỊ>S�<1e�����u�����2ڏ�a���^1�y��yGo�ve$*+OH�_�	�]��
/d�vi����U��L�c� �#�a�-��{=a����F�LD���_��S�9d���&_�!b���FMJ,����Y�<�L��oNuf�4��)�A�G^�"��v%�q-}�?q&]� -( �+Q/lI�@�w�+D1��})��GB�k+H7^�V[n3@�i��x���l���{c��V_�80�o6���8�mlJ��$��vF2����^�����j�LP����;��e���\8f�9Ÿ]�D�b�8/:�o3��b6}I�ý��s.�6�g�.�ה�,�����[�ӭ�2����A����.�9D�c�d
M��H�5W���"Jx��W�=�{F�uS\�f�n�C�Wь�� bIT�}��@t����+[˛z�̬��,ӌ3�����Q���T]�A�����HZ^G���^��Bs<%����qr�LR��-m���~���T��c�ɉV5!�^`����/}K�����,o�G]pT��т�'l����bNӪ:U�'9P����s��!���'���KI.�UڄZZ���׋�K�!p��MnUcFg��F� Px^��o���Mz�E &�k�s���$E0EO���ѓ�h��b-}��K�;��-�6"7��@?%�񂠥Br!��]�<����y���?��ɨ�	'��U�$��� �P"�P'N&lS|���������d�^����L*;Y���<�7���N��vO�m�k/d]ZI��=�(�D)��祸��6iɺy��Azr:H?C�	x�r�z�W2`��&��˚]AjA������E�A�-{"-�g�T ��PM���3��25�!;];����3�M'͛-|�5=����ܦ�鸱t)٤$j �a��\6%����4�{Ow���s�$O�e	
�$g��9��)�~L #d����5��1�{�� �`AP$:]��.��o�p������H)��㝢�1�����f�Z����'D
jr6�ls�B��7MfMo��4X=c�%��x��1�[�i�	��en���Ky�]�M�H˨��'�S���<�B����j�^>(֘ad��!1�Q)"����X���2;J�����^��]���Ś�$�餒0�r��.�\\^N�t�W=���,�_�u�s��![I�0`4�o?�6���y�l1��-Q��B�O�4�c?��l�#�B�9��5���q��}'�k7'� ��o��q�3��WX.K��
rx]/��nϯ*o,��oH��
<�"���� c<'���j�q�Nd��wAE*�.�(n�Ha��F�PF��$��\�zvdΚ�D�8�]g&�}G�v�6�I�sZb�\`�x_��ii90�p�'���� ��S�Tk�ږ�_����UZN��8p0F��c�@���v�}���%���Ό��xJ�Yn�P���P	sm����Y��ZLX��YD��v8*˧KE�H�C��&�-�\��pEGY��t��F^ՙoY�l]��Ϊ�T/+�(��/��mi_��Gyy����A��AX�M��\
��C����°L5I��H��u�>H�8SU�v�%����6`'}�>��y�?�y%��Lʢ�w�׬����| Nṥ�"� ����j�`��k<��n������S%G�^�4�q��xl��GAm[?�V�y�(T��iIJir�:�@<l��%��ЕeπB7ڢ
.p/}�rJ��|�,����J�$��yq��?T���&7l%�2Z,��I���A۽~M�����_I��H�Ay�ZǢ�>C�)�Պd���I�o]�K��>��G(zj�������&	 ���}�w��R؆8q�q��7{ֺ8+���S e�]]�]-Y iAsI�:-��c��\�K�D�i���n��F5��"\;q˽1?q�F�����2ƹ����6�;|/%�y^��V���T���/�ĚTA�P-�e8�/7+�8]Aa-X�Ĩ��7�;;�\�����j�bEG���[��c��a�����x�$�t�>똤���U>�ف��� �l�;$���dͩ�~�+�|�tg(B5S��^į*�>���m��q�?� �ή�A�I�J�Aԫ��,�)&�$�p�q��B�v��H5���C#]X�햷´->�2����霦����_�p��'d�4��ø�X�Qcl:d7vV�YhG���B�;4�R
-���Ni�<�s)�R�yᔺ�P`��<�!�z���^���ڡ�c�*�s�	�$�Z���?˛�`�L���キE^��I�\A��^��N��'�����? DЙ�>��Nje�,q|A���!�4�XZ�qgǭ����F��"h���}%���F����	t���7��X|�.\�{���vנX��߭�XU���LV��t	�o���A��R���˚��5hC��ٽ��(.P(V��WF���{�/c74C^a�3W�a߸jf��d=���нH�r�&0)�=Ɍ���OV4�M�K�V�C�)o��qT��X1�Rx��AB�3gO!��+DS��b�A�Ni�~`�t9�v�~j>�ٻU�Ap�XX�q���+�������rLr��~��
�^v���.�h����'\��|`�Nei�?�P�;k���Ś�ar.#�����
�y *�^
�R_����0IkI5�	�v��L��Q��6P���2D���E�P~~�>�#�V�]w��,�S&oO�n���Uaa�H�J�9�H�7~��ͅa�WG�$����sVpH׿�)^��b�KE<��.Z��U�6��|����erʌ�l^/Q�&TS.ڜ�4�p1�ȱg�5�2�q��ƀ��5���z���ب�b��2������v�T4��,"]����oL&Kv�n,r��A@Գ�����&V�Ș/)]��?�ZIhY$=UЃ�u�_0(߬�$��f~�Y�����t-�=W/=6D�=���S�س�[P���cZgk�9�⥐�lD��?⺦_읏�,:]�N.V�"��{��t؀"�2;���k�i%��6H�-Q4�\7���p��#2�ECe z-gAad�|>���K��h�� ��m��E�9+b��R)j
$�e�i�t�-v��Φ�p$uL{.߻��5�(괤������KKb.����~U�YBK%���S�"��;m��t&yU�6�Rqri�H�̇%��_ѝK���4lQ(%P!�)�iXwͭC��m.�f	�^)~]P�i���y��־��_+��Iu�eH4@�e�x��5;��{MRy�cW��G5-�j_��䅙�@�R4On�Dο��D6���������T�iIb;�=���D��b�\?E+`�%�]�?��E+�t�ۑ�XI�d#�1��WL>�U�Nv�}@�S-��4�[��Rl���4�5h�TH��i��++F[�t�A��Y�Rd�6UyК��m�?B��nS��c.!®�8ڲ�|���\��Fg���MUh���W��B33��
�Q��9%���,� �����k��b�#�ߔ]A�2hu��&z[��c������n�.M�e�T>l}Lj6�fwg��*w���By��iC���?KqU(�/��V�H%��o��N�c�����\��P!"oIߵ�FE��G-�) 9�M��k����'VbG���\�����S�P��Ŵ�s^y�O��<R�\C���Wv��K�B~�&V��Y	�Br�|�r�}>:�?̻�*J�=nW����3ψ��/A�� Oqh�W� ]Qn�K��F2wώ����̙L����͜�V<ƹ^7{���X�g�z�Q�d�`�o�0����՝(Ԩ�]?�,��
�8%��|+������2i��蛧��ۥ�E�(�3�K��#��}O8	]3Nx�Z艀��z���Oyd����bc�R :u�ܫ��?��)��<ۑ��-��B�Z�sUH ���w5v�ڟ"�?�O鑚v�9��"�K�KZ�C����q$