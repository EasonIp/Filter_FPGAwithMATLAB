��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�P�;�{��3�OT����n/\�@���V�F�	G�V��]� z�`t���y[q����a2��;��i�t��,-��1�� pz�jI;�"<i����#{���<�G�N�3�mŬ�#�:����(U-6��K��j�'��Y�}'	T�(L��ag�=���`m%5�|Nq�Y;�:�|���Q@Y遀 ץ1X�q��j�%|�H�����la�IKA�w��H�=0z �y���Ʀ#��au��#E*��p��c��>�$0i8Y=�P���(�]hϽ�8��1���y���*��V]�t����śvrs�C[o�3W�{�ZИMm���P�K ��L�:xv���U��M�X�[��:��p���C#[�̚�/���o0l����%8Qh+>U>A�G�r8!t��/��$�ѳ�yqO}�^.�q�k�_�:Ҏ�GBe��*�b�?�h�Z��3��T^���jL]|��s������ٗڳJ:�%`
��(#���gx�A��s�P(������v�[�q�� Vz
Ђ�x��M�3Ǣ��\I��ҷF#��_4`�E�J��<HK{0��?U(��B�Ȳ��b�w���n��xX<��|t��!�.u��#��հUEl��ݩ}O���*	"n��Bh�LXo���jT{�ׄF�_��C��1���%f��#��Y0	J^T
����/|<�69���u��I �A~�d�.�b�p��:\��m�E�/�̮�4�_s8��F	��ճ�)9��O�߱��{#�U-�4EQQ�2�s�jE������z��^��	EB����!6o`;�1ͽ���0����,�I�YBwN�����D@oM�OK�Y��8������"X=���y�8&�R�;<DD:b����D���djx��p�	��=#Pv�x~�[s�1�a�U�6���v�:��ZՁ-��%<�G�V�8E��/_8���� vҲ�N��FR�/g`���>l:�D��1V)Oa�)��ѿ,.���)t鬵���y8��b%�NA��QdC$p+�N����F�aC]($�w�1{�XW���2N࿀����(&�!�!�N3&����PӸ-n�lw�,�K���sD6'�:1����3p�iJ�S6�k�I)"S���L4گ����	��8d�Y����oqդHb}H���{MeX����~�������NS����%��ꬎ(V�R}��N�9۟#|v�yi�A#6~��:� �o,Ht`���Z�(Z(���yیV��P�8ͅȞmV��׎�;Nu��C�"s�����m�i�JYE��{*�o�-��z�>�ɀn����Z,�w�)���PC[�w���t�9x��@��T��D�7�C�
R��S��B�G �KxZ�`���@~ �Xo4œ�g��ozr�h�Sϯ�|���乨g}�Ba{�k��{SUN-^�7xR���=sU�r�k�ϧ�%+�0�0�,fCrw������_���Pm��|�ؠ2JR}N�m�:#����4e�
j����eգ+D5,�����Ec�H�L�D\��N�bN�/@�{_]9�P�#$�@��3��/'�=�ްs!A���>�Sp_�L|�5�*{!~�� ����֕���H�/��_/�R'I��sZ5������<�h*�@��!B�YrBW��cv�⣳_��M?p����W�ʆ���Ayf�J�w�2�$�S���&��A�*@��k-t��~�����Q)v��cʗ.*Nt��T@6�M�c
���:�͇.[��Ѕ���'J�wB�rz���Ij$�)�9T�Cy�B�~9D>|!+�~�s��C�̉�)wn>!@���ǌ2��`���ҋci�𻀗>Şo��w"�u��L��?��4�6�	�<R<���I���f�$���'�)S$�𯩫�0��kb�4E�8]&O+n�l�$��u�p�	��[��}�#��'dV�zƘ^B�X_=uJ,	�e��XÁy�V���e_]���rV��z�3!\\�o5aUf�j)��(��x{�P�_�z��͇ȣ*�-:����tCV'L�����M"K��Y���hUv!~
�,��cpe��t���1��L����0�aD[;�p,�M\�?GGF���E�W��m�\2� @�9�(u�:ܶ�N�����cw����eЅ[-���������p��OW������=VM5F�&W$�'�-Yف���u����	�Y`/�5���J
��B�ึQD��$ᰙr\6g�g	�ʍ%��dur�aG�tn&rq���}�=�RLK������>{��w��L�'��`9����id>G�K�E�y��"�a%Ұە�9.QW����@��������R���w���A��eo�	Ʈny��\{��QkdZJ�d�yp#I#�P���x-9Z����Z(ȟ%�Ǐ)���Y	S�_(uE��ݦ�	�1�W�0����X��q�V<pur��������0��X�:��;}��d%�\�%�g@�2A���
^��6�W]��x���ĸNBџ��J�m����nM�ȏ�۱97^<yXB&�4��	��(���}��>r|·���q��&4X�	��?N��L�)5��ԥ�4+L��f���A}���Ʀ�������u��h<�Bd14\�UD�ԝ�v���|���R��A��gr0��D��+� 
K8:��a8/݌��`�ѭm��[A:ѭi����X~�8sʘ������)M���>%& �w8u����;��<ŕߨq�{݃Y��`��3��]!@+�%�^��i�/�i�
��p���ú*N;E�������>�H$4ʡ��
�y�Y��E�߱Ի����{苧��]��Nidd֛���$ۼ#_m�1�v�f��}��O`��s��@b�t�����!o{�ž*]�kJ�]��Ì�L��`�a/����g�K�i�#h���[{�����mp�U��@��O�����r��s���A� )�E�`�����O�(Igo��Mr�!=��7��N���Cn1�;{:���s����
<\d#!Wod
�t���$ql�� F��é1'��!�9��?����a�7p�����/�w��N�i��=�I�E�֩4�r��� U�ѩ�/�l�ӧ��U0`gNL�܌q�@9oJ@IU�' ~{w�c5���K���M��Q���F�E�e����H����Y2F��%Mc���`�R6E�呸�Wd���)���PuJ�U�cҩ��Ȫ���C��!?j���k��M;w�ME���9깟��#:���"���;`�~�
��6�:��Rxۣ�ˊ��(�0�Y���r�x�����"�;����<!qV���E���sm����X���W+�����Q&�'�p=E:�.���^�(hF���+�Uu��Y�W��H�,gDS&��~��F���C�o�[�ϡh̢�i*�)J�����ϖ���i�����/��fk\�k ���x3ǒ=d����C�����sNu��$�9�3����"�"�|�UI����NY��K��z�jЪ�M���A��&�TSInkn`���lҎ4W��s�D����%�6qO��9���v�c���@�`�d�D�/��UG���� �3}�h]N�J��\BJ���٬4ѿ�tvt,|�S�ϴW�ΊGV���6���Uq���#0��E_��
�	�'�P��N�5�8�M�f�E9���ri�Z7�ײ�m���9�Ѽ�T'Gy�"���8�J+*w��l]��&�	+j���%��T��qחa:@�����pCzvk�Y��� �^�S�2�)�����Aj�c Hr�٢y~�kG�]1�A�7��4lu��'�z	}�,��y��7�[����0�������!9?���+���<���1~���a$������U�X]�h|����&����_ێ�5#��g�qg����=y��%�[���^���L����AH�?�>����d���j�֑�1��<6ݭ,`]�!����D`M~�l� }�$��n��Ѐ6
L_�	L��-��Ά}k~zavnPVv��&��Yqg������rE�d�SC[�~ʙj��e9�I�ɢ/Q�;�\}���=�D�t�5#c��l�Ϝ��T�\�Y^��t��ԣ��	ȏs�z�+�*
+�-y�- �
h9r��_��PwBjl�|�F�9��EUSZ.��@�Z���C+4"�;�a�AT<��aK�fέzE �Q-w��~&\[��D�1�c]�S��wf�pu���I�$���t�� ��M��Z��	���w�S��Tf�J�ÃC�:
4&1&��).8�kQ7���*��*�В{����}2���ȕ�Id�D�B��ܐ����i��p1Wc�	��^�pR��f�9��U���Pʦ}�w���7d>�>�~Cq���R��L�c������A��k�h?iNb~Ɛ��)�ֱs�������Wtk��t_ױ�^?��:t�ʕ�%Ժ��.�]���A��e�ǑD'���%N�Ϭ�^�K��S"R+�xU~aH�������J��R�m��2e֣�}�$�7��,�������x�6J���)�T��B�[\��=I��.y �T��M���Y�͊��e�K��q��Yr[�*/6�� -�m�a��Hs��:�[����\��hn�Sa�V���rGU�_�unK��- �>|oG���8�1����@)R�Ycg�#���^Z�:�[�D��B�|l�2���<�?���6^R,P<����K�t7���k�r��+΁�^,7��`v�%9Ұ��a7�|�?�5z�b%�6x�As��@�:�s��1
���Y+>9�(�TG�Uz�{Yr�˗�
��-����<���4}m��NoPN��s��pϳՊʁZt5��ۺyPT�#����xv2҄�^m�5H[b��t����W����Y �dA�յ���:���2�HO�$�qºEZ����~^6'���6�m>GL��W.�I_a��v���-��>�^&� Z��^�~����xL?�ٸ���BL��	�Bg��|#��Ҏ�C�K0Y��olF�>z�Bv%�����.2!L׭4��v �
h>ET;�"!2����Yh1&3\�kL��]j>ӞۈXPp�@O���ǰA1	P?"ǌRet���Cm4=�W�];�xN�E��B��s�Tb��f�e��'��p��Hīi0�������$Xk� Ks��U4Ӽo�M��p�_�����2�b@����$���k�_�@��0"�J���<ߓD�dZ�������<�2e�P���N ����D�4�:k`=9㮜XL��J��_ȀO,�vQy����1�<�c��@���п⒭3����'��-�=��V�"hH9sh��Nr'�@�u�õ\�"i��%��	��&b�}�I�()��}�ڴ;BBk����_�ސ�.�b�-�(~Uy}���tV�"D��j�ft�8�i?9�T�*� �X݄2�s��df�n�����]qo@9�fc3��z$��>L��=+h��In���.9kR5л2n������z���J�d���'���z!^����HF-P���o�,'��[�e�OA��f�u��#��Asj0�<`�y������K���@UՎt�g��mGf�{�F�[�9�j��R�s��uw��eS�?0�@�nc��}k�qb�(��G���΀���$7/P9�i�β�!� }1��<9Y�Ld��I� ����L<�аK��MQ\�w��:7ȃ*Zb��`"�$�Sp} �a�es�|���֮�)Z��M�N�@Ԅ�(�?Vxv�p�E�%qV�E��0X�gM�J;� 9n�:��|l������D�c�"Ԑ�u�<��nE1���٧i��i�����#�q2���"�|�Wq'
˂��`)2���s���N�b���h��|)U���k���StF%��krS_e��4nrs翰$���L�y��C5�M���EN㇓����^6_�K��jl���!��J|��'�0�"�R���� *5@��j=I��is�}��N�` .Cu����UƘ]�aY�W���-�nQs�N����u�Z�H��a&� �у��a����3���b��J�Q�c:�uq�tO]��\o�����N��iW�(t�s����7v�f�\��~z��
/���g0��9㽸�KTh� �`N}ȱ��Rb�������_�p���h�{F���T�G��g7��蔓�}2�k�p"�'��w��ɻ�Wb1���IZ���YպEX8���ф8��x�"��%�8���:��˟vC�Ҩ𡔏�z!��L�/�Q&H���<��ü��?��7w�g�?�ڬ��syd^9�U`=[*k�?����%楧o7�zo:.؋뇘˳ge�i}�)ۡΡh&ϥC�k��us%�R���/�K���� �ͷ�#uYߎ�彎�	�ڼ��X}�׎�<�,�X���f���eh_O;b��J�{���(�nf�R&`�����c(lGk�W�9X��_ep���Vc�b��Y�����Tu#�C�d�b���|D;i��^&����oa��EТ���;��`쳉�y�4��'Q{�+�����" Y�o`�T4����,��a�<�kU.��SR��u��7��}hc�H�EȐ��ݓs�#��Pҟ�{Q��:��k���D���v��܇8������:��	W
Ļ�@/�^5��mE�2P�K�F��y�u��Slu�A�^|��oSϰM�7��S����f.d��&'��^��$�VWB�_��_Ń}�:Ş��}nܴk Q'PY7��+?3"#=a/۹���8$���{��1�2��pc�~��˽�&���"~�97�M�89�2��֒tGaI�X�I�U�/���<�=� ����i	�HT��<�;��Z���1�)�I�(�xH���%��p���5r�B���;jy�	��Di;�&�T4�s����l̛�� ��� _�#ԍ����L>�㸝.�x�n'X�CO��[$��	hc��H�2�]�U�iT�ղ���� 20XN�)L��^PG�+��F�;�m��rc��+"��d��Z����dNC;|t=�!�Y�O3^�+@��v�
�*"ьů����l��H|t"*��ɞ������,+P\S��>�7��d�� B���y��@jpAظ�+�臂�bs�nt����D�%��a��=�2��tX��v�M��}���%��x�U�X�9eԹ��UP���O1������*�x@�d+��E� �P�;pD������g���N�Z�u�T��7!���TW@[t��5@�KmIr� ��\��$5��FuD�FB�}ݤ~i�3����b��U`A�!����&e���E;��o�������d�&���|�`�;�w�B<��y�Vo�*:�]���ᷱz{]�������8�b6�l��$e2e\7���#4^�ӧI� �����c�O��F�c�b�q	@"�Bx<��{ &��SP.Z��O�6����r[��y�䚸�C�;����j���H�����^d��������E��s���*������4s�qQ�Fy
 x�I�[K9�}5�`JE�1c �Ϯ�N/���yZnV2��+�yaR5��g�(o�Y�B���y�
�Tҟ{s8�r��}gY[L3�.y����DN���y��TQc��5&ap��\J P�l,%��~�Vٔ=| �o싦���bʎcA��eJ�4sg|c���-e2�tH�u5� �����M��u5�vM��G$,��nD�r�f�n� �}ή!�t�Rq�lxu r����;Eh��������B%��᭙��ؐ2������U���������TY��G�oׂC��gђWj_�'z"��'���+ct�A�]x���6�:�Õi�4�Q�n���)��R�``c&O�n_Di���F��,����ʀ>�����܋l4�;+��V`�[��tT���J�����o�_��H�I�9�bk�-����3���ȱc�ѡ����ox�VKͳ��>?�|Z1�KV��1�W������I6�k*_�Mb��7�*c������T���у&�E�A��\��#N�!{��x	)�T|���h�!�� S�JsCYF}X��^�m�Ō�۸q�����ϾyNͨT��^�L�h�S�ԓ�12��/e.D=�.V��P+�2�-��~���P6��%����b�9�.��7mZ�kJ�슷S��R���i'&锾��]�|��s�h��qZ��[z!Z־�� �::�K�$r���E[�3�S��F���N�K��RT�+��k���`TA��z ��hЕuV��l2��0�@c��#��D/��A#�:T!Ige��G�bO~�5�F�#4Beh�����d3Ww$+P�&�c]P.�v%�"��L��&��N�mh�j���2�d/�6$|D�)�E�L��Fӻ�b�_�b
�ȭ�G���SO���(1%^!=��R��c��j� "�4]S�d�ת�8з���v��3,��oAZ��,��S�u�?�t�0����1�~��;�M��Tl;�%�
�����K� ���T�������ݯ4�+zM$������E��9O6�RqMyt���.�ՐK�8'&����*���{�)�$X�:�6�
��^���jL����X�"�9�)�Z<*뉗ŀ��KxԶcp�+��k�Oҁ�,��0�!�Ҍ$ea�)NB��,�:h�b)��Њ��B�D~��r��Z��z{�3''�	����nx�0�;�_��D��{y�S�j��n|���`4�i����G%��Q��?E�Έ_���(fQw. ��L�M��aG���V�XaJ��+0��rc���6JŐ�D��
�,vY�K/&Y����Ł�Qs��Z�ݧC!��6-��c;�'�!Ω�8q�r�4.�IH������,�̨i�h��l�p��l�z�BI�)��wn���sT_˓����eȇ|P�����ݬI��K��0"y�1�ۨ�%��׺�q�?���k[S-O���(����!�b���ŸH0�L<O�C�Լ#�iLm�	ݫ��JCZ�<YUc��zٳ�.[�!@�K5�:#�W��d�ZA�)��^H��!����D�Ɵ�j#|/�x�n�N�^[���$�T;������MN0�O��O��"�x��t�Ҋ�|��|4*�)7,��������`G�Q����Z��[�����9��� A�KT�-łf#�oPIa:�cv5o(�1BZ��΍q��Dc�Yc�ē�5�:�a�3�`q��=	Gn�'V�A~m~�)��,�ө���������u�c��Ά^�C*�rәm�~q+�sE��Ԧ�dF&���f� =�B�)��������Э�Hw%�F\�R;���@��t�(��Z�\@^�h� g�?BEe5�����l�KG���)ڋ]g��n��po��v|]JލK���nKz�g�sh�� ��M�9I���[G΄�ҥ�qj�K������GF���L�	��]�������ĉ�Ǭ���iQ��M���� �-�<;���I�	�PD>W��MbL��| ۓJ(�4,�ueQ}*faz�����R���rHw�HbS����_�Rz��k�z��!*�*���W�wș�/˲)[DǑ�W��=�t�G���e�I�Т�LUD
����we�sɞ�;{��N $|�]��6N������!��v^�a�n��TXL	B�һl �}��l��$�Rw�1P��u��H�##pxe����@^~�����C� *�HאC�ȱOۑ���I˺c��� f�6#� �l�{fJѵ����]7-����(S<���%Y�X�ؾ�SSͩx�����n��u����X+]���3բ���rBS�`�Bbw��{l�}�זc?p�{�{��';xŢ��s�4>���Xx�!�����\�D_�J#6�1���t$F�u;���n����Y�g���=��^+���Wq�F!��ռ���$��B���\vqm�y�彋�!���&˿s�ml�9܋qX�P���e2���x������U�i��-��"I�-�?_��C]	�v&��&� ���#�Bפ�j=�!�'N�� ����ć6����3�������������A�%>rU��W|��TS�2\)N>�/A�5r���҃��c�ϑ�(��U��~KԄ� m���Np	U\�By����է �����u�n�&&0F~��������f�j�jL��p��y����V���`$�y��v�����-7�Z�q��/ax��O��K�ߏXѮ8��?N�^\�=ü��zD��:K�	�B�df�h�o��
�k�~���#����"	o��@��^6%_fe��X���c;��x'��jh�~��8������R2�8��j����E�4Pe��B��2�1:�*��Gq� ?T+�i�%Y�&=��dZ�Չ�Y:��bG����<̥�S�~2�V��~*�1��%���nvUs(|M)�/��F��֥��f�ꐴ� ��ơU]L*@�:�̃��;�S��z~�v��tC�����Ve�p._�J��U��1X�W�������g��oaĳ�4�I��(��kq�+\�9H���iǈ��k�5�p��0��8W�+���?;����Ԩ�A�� .��@���jC�C�K��J|��җ?��Oo�Yh�ߑ�N]���>4Ş����/7e���ur�{�1,�	v�
Z��Yܽ%�����Ih|��mX28�v�[�b�5�B	V����Ӂ:��������� f���/�ʵݕ6cC���K��,���	���Z1��oު,��P����p(CX>`X��[�(,{�3�n�.h��\�ˇ��K �韌/c*�%��T�����5I9�:���i¢S��
�[��DH<�nX՝6(���*��� I�z��U�B�rvV4�?�I<2�U����:�+i����MM�Oz��(��5T�yU�!���	�	NM[G��'"���.����3s|RH5C9�Ƚv��8�ھ]�Ȏ�t$#J���U�-��q�laJ���JZ���<�z��u�a+T���T�Ⳮ�o�i�x��{�%T ��y�{dÌ�I�?�{�6`[�T���}tlo��Ӎ�������X�4 �gp��%�3�lͷ@+���B�G��=@(R2��bg��ƞ�_�qNRHޣ����'��`������nb��j�L�쌶[H������?!�d��a�7[#b�� r�G|�GL-�`�C0ϓ���s�5�WUh�ӟɉ�[�~l���)3N6���k�1�;sp� �̶
�}&�d����χ�C�t��2&�X��2Κ6��t�G�����J�!�[�_�-���w�#��0q3���mK"f`�_K
��,oiq�5ٿ�ا!��R%45��5$u���A>i��;}M��%�F���%��_7l�]�N�B�Uߚ{ܭ2��b=������Q��n�v���޹�WB@�䅺�o�m��ٽ���������&��I�z_�v�	���#$|%�b�wʁ�QT��`=>u�z"]TsI�NNE�uvf��%M/KƲ�Qc���!�:.#�w���K��u.�J9R6�*�b5ˣ�z;��wf�K�s�u���n�V9�}y��������n"P��(�[��z�W�0ʡ\X�ڒ�1����DI�b�}��Y�=�6v����V�hC���f-k�);�c�:�7^G�����-����®mC�D��8����H��g�3��֩�AO`#[�;%�"\��x(���xh��p�ףo�hk�˷�ԄU��d�������Q�Y*s��P'�L"kjd�/���(�S.g)"���a�����`P�,o�I�1O�k���x��v&���eؔ��oJS�D�̋T��Rb$[;���R'�Ӌ���{7��S�Θx��z7�*�*,7��uDSJ-h�r����H�6�BLJ����T�˶���$m<�^ρ6�|��<fD�L�t�����Z��,6K:���^B��$7�ߵ=�k�K/�b��K�*XraY�"d#�'���C�w!�9 �IƯ�4�\%�Gw+p��{+i6�+���Yp����I�!��,��RR�,s�{�];:s,a��)���Dň?�r4WU��_��Ps+)��9� ~y�Gm����qX�z|�*�x_rJ���������Z	';����Í%W�Uڗ��:
;�gʭ�o6pW�'\�&�m�6U4��Em	݋q/����1�f�b�lA�YK��"�-��0p �p�@�r��^�]���qO����������zF�ƒ��[55Q��D����Ȩ�P}�A��.7)ѝ�,y��;!	���Hdk�#r	]'���0I��d�������̈'�cm,�q�g;�x�>�ྭ��d����A������f����N4*g��lE�8�Oq�7�U�c0�h�t{���a���Ug|���N��b�Lg���n�SS�2Ɂ�.dueD{%4�(-yp|Qu��~�*#X��j.j�4 ��h���cF�]9a�w4[�T�d��3Qx��I8�$��ji��h��H·0=_�'n��7�(�$` u�sl�77�N���B#'�r�5���IC6��LM���!I�+l��q��N�@�Uu"��iY.�mD������`l�4�D��	��@Sc�`!q�0�iQ�Ƭ~��e��zX���@��G�����R4�A�'U��}[�t�? M���E�g@�mk��2��l �57�N(�D�p���Φ~��ވG(������ώ�@%Q�Y��o"G�?�@>���3S�h�|C`2�t�s� �]���9�̍j}1Q*Q)k�s4ś�ʛx��P�����Q=q<\"�^d/} o՟���w����ZX%���{!zѦ�j_f�%�������Ի�]|Z}a�%Sߨy�����S�8��������lN�H�����JJd���9��Ox"��Z1)��a[;�T�"ؒٙ��f�0{�V��L�����x�`����@N���E�e�@q�D~ulP��}��dX�L
�Dz9���!��x��i��F��w��c*��f���@���ܣZ�-�\�7�}r��Ӣ�:�s��s�^��j���y]H�SU�ã	�x�<��,6x�H�ӪY��z�k�~η*�:�l�|�Aǝ��~�v�"�h�V
ݑF����h���m�������	��@A�il>q�'�=٧s������J+p���+}R�f��g�#�k��@ I�1�6U�_� �;eIm�a_�}s7���~7�\������#�Y�:�]:���*,�_��UT��:�^��#W�`�ː�l���(�3��5�{I��0SW�(`�q�9����<��cO�b���ی��љ@̝ m��p4��d6~ |�ԖM��d�AKhNG�z�#����x?3eM7��yL��,Yn^�	+�H���n�w/�#���Ⱙ��3?]�d�D��J-�8`ؗ;0j�3�XQ�֩����tc��iy�cb�m�4�wt��B��d0��F�Yg氶�w������J��y�pnUB��`�����;��}Ij"c<-s�����[X�d>�'%��_W'�ӻ�H�ڹ�/?�BM�*(C߬{�����H(�zs V��ҷ%����Ҧ��R��9�p�oz�<,HD���A$�YP`�!V�W��a'���AX�\���&�
2f��㫄5N\ԍ>Y�I
���$	�J�9&�-�Z���L,�'ܣ4/�F6=�@�K�*p��g;f�7��Y��TFl���E���&��	���=�`g$)G����B6�;���Z���2�#����̒�{;RZ�Lg�sٍ�(�aboP��~Hu�Y�T�����k���?6T}�43�<4��w����� �o;�Ga����TK�IꀭzryUZfy}3a� 0'�N�-P�h����~6���4�W�a��f-P|6ߘ A
M1I���_O�P����F�`�r� �ۍ��Ф����J��.��F�`��9�Qx���"�6cHK��p�G�x�aގ���\
����>�~��{��Y��y��q_��O�}���^����*�öC�.�s]��'P��K+�����%��@���d��R����)����94�D(�������<|�)g�k��D��UAAŵ����ڃ\�yX$�@�	Nʔ�tA�Cy6�S+�i�f�/P |p>�v%�M�Ɵ^���.���*��Ӗ��Yu$��CI\��4��,={�.�=1Z��u8�(���G�fbm"K^�W��n5�C���4��8���)�&-������<	�}�+�N�h�{ܒ���/��S\��؂m�l���冞��ڨ�_ԋM[wLu z�@�ܘ��-P�ʩTt0�Ǐ�vp��;+����à/�G%HcYb$bR]�����k����l�B�Kw��<����W!�;���(~��>��b���MԦ��u1���rI_U���PQB6K'2�Uy	7���wE�M�xXZ)��cB�v��I�
�Î�(���w�k������]B��U��0I��HpQ�ˮ��}Xp
\R�{
��am�G�'H��\w�u�_���`^U;�=V���v��@@7��@İ�5+�ｼ�@ye�Eɐ12U�|8+���vS��]M�d�~gNk���O|���a J��b�?Bm`�yXD��R�*C����^kY�0(A�i��M�:S!� ���:��Q�"&:ʰlv��|7� mW�]� ��^2g�`jٳ�.�8'�13�<1�z���%E��$���'4}�r�팞��<�ˆ-:���z��(}A��<c�6dӾ�C4j��Q��.��䅝R�?��@�t�dQU��_�"b����ә�\����:��TlGW���ŗܟk����q�1��+�c'wJ��4�����?)%%�(���/�������2BM��0!g���6�ۿq�U�R>�G�b�� �a�1Efp#�e���t�F�U{�	L�f��V�щ\t��A���i�Q�r� �:~aAk:6`�(��z.�ޏ�6Ɉ�9�r�R $ZeU�!J�B�֕͟g�4
Qº#� j�8id�١+�.�����y����M>Ù\2��g�ב~�-��\����GrE��aN��wE(��֏���=���U�e0��f��g	JDP0�~�w��{� ��)�z��wP
l���t����8rP�ݽ�B��LQiaj�����R�~�XCC�-��Ԇ��h����E��{�_�g��2���L�m2䭚�it���<�T�w�$�-?��y1�֢
�*�T�����'8���5���)�IL(\��1WϠ*2ܠ�*�����P�o��h�-�}��w9f{5�։��4o�0Nb��)&�H��`�;��s(ye�M��:���j��j��N�N*kg��¢�u?)��tN�!G(�F�:C��2������W� ��9�*':�*eI�״4�Z�yě�3g�{�=�4a>��'L9�'X����_�#y*�#���}�s���I�A7��bc��Qm��e��rbAg�Y��X1Y�e�����AJB�V�]0��k՝#�VT��׽?�#.�6r�z���e� �[��g0I�D5�����,P�J���4Ҩ�����ི~<����&��H@��,�̣�s_k98r*�G��-Zh��q�SP���c�������[�G��O>O���?w�3��WA�������'�y����j�f.J��x�+�Pˏ��I��AO�pJ��""t$Hx�� �Q�v����U��P؊ ��tа
VK�����ğ�Q%����wQ:�s�^�$�0<o,Ҵ�I���m����z���PT�~^�U�r�&�h�A�d��nu�W����}�˖����mh�]�	�2=��%���ϟ�g�.ޛ����t�!�4�5U�������Mǁ��э��9~�L3G��R���Ʈ7\n^d�*�eT~���ZR�\Q�?l5�ӎ��~�~c�7����i93㌶�ג#�\ʱvc3��}>a���d�]�2�HDt�?����	�x���	��eRs;���0���%V
��o �P�|*t_�C���ʆk�����:tRd�'��Ȏ�&2��J�m�`n��T(��T�3�����9��Vy�LD3	��k �̮l6���+�N�o��J;s�m���A�2�A��M!9p�b������F�O����|]/c}�XV5�\�=qD�����'�����;A��(Wc����D逰W���U��
2Q�[PK����ت�,�$$��<7�S��G���\B������]�$�������
�V�k$Zn�^���B��>������B�>���Z�S� ��	ƍ����ɀh!�nV+�oɩ/�d1�\u<D��&uBp-����3b�	��z����E��v*�	`r�����h�����0���;>x�m��e��, n���)a����VINmvBa�Ħ����6w���Χ��"��&e.���Qi��Ҫ������g� N��;R�p%��SZ�,M��hq���p,R���g��D#t���v1�s��q�{�ņ;s��
��	�QއF���N�F���=\Ⴀ&ѻt�煴��Y��n���{�d8!�(ܽ���+q�ۏ��{P�3cC�a�a���q���x���O7���?�	��K(�yD�2�~��۲%��!�r�9�J.������F��)#�Iqwn�j��6��I���[�XI|���Wm���;��eU�����v�&Qh׾���k|@��)xLI͌��vnK��ukK�7�tx�2�V�i%�-�Y�#l����z��?RSh�e�ϡ�d&x�x�񕿤��7(�,U���t�B�l�	`�6�g1;O�ß'�\�(j�#J!_EF�]�r���R�`e`����]��ޫ�S�L��⚴��+x8AB���DmYH���'��+W�}�G����A rd�טT� ߏ�4i��_$`�h��,��g��l]���O�o	]̰�a���;�8��E�\n`h�4N�"J��7�4�t��Z�>�D��}��x���|�����?G���t|J��:��a=*%�;s5�1�Qi�z����5zf1�&�_V��5����R���Ѻ�6�>�8�߲*��2{�Q�l�r���C��P��u�c1�߉�.��|5-�)�t�0v��g�J�3�@�
2j�e����,^(@#�s�Q<bk�"%4ɇ�p5�?�@��R�P����x �(d*ў��	�5D$���Y�x<��DO4�8pC[h�S�kB���0M" ��&�hc$q5y��mnVG]�E+�ƞ~�)S2��+��	���|+�]���F
��pL:�"6D�:�%�a���W���� ?C�M�2$=�3��"6K���V�}�j��Ϗ��5��s�Z��Vp.�5�-��o87��,/=жg�y�S��Hk*�b/����v�f^\�`��!���."_�}ۜ����8S`f{c�J"�EI��sC=w�`�/�A���oT��؈�H���	�ᗥ���_��G�)	�Ҡ�/2)v*���S����-350&V!��'��[[��]���/Z` ��c����@��c����&.U���k�{��D+n�}�db&m��yX�6Ba���W�9@Mc�Y�(]v�����Y����� h����Mʦ ��oq�n�%�'ƪeq@�("=�"�kX�$����2u�q���Z���td �����h7������?Ҷ�	Iㅌk_��qm/`Am�
2����]1�/��i��5�.*Ј��-&�0k��)��(�#����~ݍ�Aܗ��wv��N
4;Xl�9zd$1"�*�9�ϫ��t�)P0�!�����*��	J
!D�c/���:�����]�yn��&��3�ƣl�-�NuA�1]��j�H!��[�^j����u��
Z���2G208ۍ f���kb&�`42r����ˮ���PE���nnuT>eR�Y36����.�����pW���������e�rG�$�ih���V�8�F�Z�?�Z�uOGZ��0��;(b� *i�+B�f |���2��e�XK�8n���^*Z���7.qU�s�&�p���!��I_�{^^�Zn��nh��F�����-i�;U2!����G�L_�C��d��$:������7�gM��7SJ�W���ieا%����s3��c18���kv��I�q��Oa���^��F��\1/qf/�	����P$��D��>�k�i���Pl�
���wda�/�R��U��.@�8H�c��;"�Ɂ�|v�U���S��cB�8�8!-���zk�}����J��12K��D�[@ӌ��T���Y�P�ѠQ��J�ErH�Z��r��k�V 	QAo(v�ٱ�¨%�dSDW�nS=Y���j�>9@�@tz���2G =�\ �wcn�s~?8�í�W��d'^m �i�wב����abƌn���ʔ�?��*�G=��T!���_���3��*�gx��sr��Ъ���]dC�>&��7���[u%C[z�3-No2Ufif��~�����=��7�HqS��Y61�i��p�ߦ/A�e#K	�RV}=Ǐ�����1��3�5��n^Pl��{ 7��"&7����ݬ̧���gN����R��틢ꘟ��qz�j�K�іD���Y�1W/6�%�y-�������$w��9"� UV$[w�Fs)��X~�u0�\\�N
����u��pF��B4a�,r4��i�5M��E�yۮn�.v��6��/yP�����FZ?HY�N�ngJ��o��,�cY$�-I��l��46}�r�a�B!���p�1�AR��+��" ��v0@����Ɗ:��F m܀�I�Z�\�H��{��g���%w��ϐ+�8u5?�$�-����v&F/�vN3R��#c�-�p�`�8�6܃*����?aQY,f�՛a�P�'�OaÀ(��HHvAwL?�]2�[Px4��dD��՗�RP�vON� ���M=�:��
J��2	��Ә,��!���1�43cM^g������}�����1��һŜ��h�h�2�	0�R塀t\p�@ϝay 	?N;�j�5�J�������</]����V򝇳4�3�1�V���I���Nv�t�}P����V�HX����h
�ok����a�)��_� G�v��[���ިsk0�pG��'�K6���:���D�\Vi��Ɓ�\D����S}���q�� �}P>�|uds�0��]"QPu�A��X�˞`NPW�rW"�Ib8 �Di��d��w�nӒa�=;�d��Q��G���_�*���A�F���Ȭ��ڼ�=R�]�O"i�rsN<�{u<����T!G&�=G�J��W�1�@d7���e8��Rφ��c����?�I4����#����r���ikg��f���5��K�)C��wn�V��5����!��Ch�)�A�e���&~]�����'r�2��{X�m�����guJƮ�'e�~`)c�}�a̲v����䏐[�SfӒ��x,z7I���<���{�@��UCm�`�A�Q߲���
�Μ�����EURr���G�4WkD�M�!S��*��%Ϡ{�MCOb��pO��*�pP%�ݍ&�#������)�������}H���9f@cɪ=�&�l�-���6��G��+~~� ���Ky>�.�Z���ƚ���l�N�RrH˼���7h(���)���nsƾ�2,����&]���I��5�⁒�u��/s�ԙ�ZB�l����m��C~;O,ݶ3@C>��-el�<�2`3�3` \��`5UtG�_�e�!͞��䑰!����k���o&���"��y�?	*���! 5j��G�����Rk�ps�;�Ԏ{U�:.C�. ��a���� ��6���y�s���eC:䧤V@�T���b�Ё���M��T�g��TH�,��S�����������s��ì}I���?Yj�7�S�o�G� MMwr���_=���9�:��ݝS������Ht7D��F��!���`�R�WCD�����gʨ�f�|���jR��>��v56�.	ʍ�>��A�����x���~��`�yr�#��r��+}�e��Աz�vk�T�١��;5Hӱ�&%n� �h�f�I��A$�I����?��f7�Ԅ]C�:*��G>�DiJ��3:���k�eG�"��Fz���o��/:%��!d��MK��g~@wʲN�T�y�br%tY{��%��p
2�|��|�0�
�M�}����nr�M7Y�7}�<_7���9h�YD��u���>�05����L�qN���$^��W^p�;ⱄ�Q�F�0]n���bH�s6�`������Nך����1���;L����4;
����<&l��F�M
BgN����v�g+Eܣ�{bm���
j���ת�	@�&K��L�X�j!�ΐ�_��u1�e�v-=y�����$�K�lD��+b`���ydW��uf��=0� ��Vi��<���6��
�9A��DCkTp�yr �r%<<M4��{<nN�,�0let�$�����i��EY�U�7�w0s���� 3i�����/̰ub�wmԹ	
g��J�d�VXN�D���z&�l��y�]�O�R�u�7����\}���r;t�GZ�I�%{rS����#�r��PÕ��c�"~���f'<�;��$�$�TTA�0kO�O��3h\����3HYt!�,�V�ތ��ʈ}���ge�}��ѝ a�Q}��DJA���)=��u�G%^{��Q��*{��	�ذ�W�.���C�^�#�	!��g�w=��-F|QYuˌi�����d�g�� Ȗf���N?ŶD���Ҁ��y���O�Y�������喺�As󶳌E���M��Ӳ+�g�U�佹O%GۤUBjQ���ޅ�b�$$4_
#f�m,�ۛ����߉��1�G�{�Vd%!�]N~�6�c$��W��'O�]�XC�UhEHjQ��*��=�vIՊDg��B1�,3\C��(a�&1U34���� �9�<�'��i�{��yer։p�7�ﮉts�q#�v��#�������*�w�^l�¼�� gX�|Ay&���
�
�	�S�Js���:���S��wI�ي {Nsf� @8�m����@61����{�!-�m�|���Z|圲F�䍷H����|ﺥ	Q<��]��)Á��Ei�������e��ddp�����Fϗ�`SLPe�w��!�`۩��"� 3���g��a����a���?�0�݁��K���3z�i�PG����M��?���׽�{�=�%
\p�A��4=�U~r`�Wz��.�-X����Z���ӏ����։u�̲�K6�K{���.�I�ĉ�(~Ҝ���㐵A��^ČgrUX����h���/ݗ�2�J9�7 �5�m֞8騚�������a�B+�����LN�k��}�pC�h�S��C��[,�U�wXq0qk��'�	�_`n�&�;Г|Z`�0���Y1'U����S�g�Bȴ�\w�3Eѽs5��-����`��0�N}�!��^���frШ܃}_��[_��7ezq������3���4
_as2% ��|j���*h�$�$lY{����M�Į����ߐ��(����w������^��x�B�8�b%c����lV��0l;�ЎsH��66�N��Ҿn��R��<�S�e�r�#�f�4�W�h��5{��}hi��y�β����\�����_���Q8�@yM/D�C؃s��y}d�j�h���G���vd����Z�Q�VF>���AXs�yJ&OQ��<�Y[j�.��L�e^�=$�}�ޫ)���.s7Au�;����.U�(��'��39�H2��"��V��}�i.��˨��� g��{cƌ(A��Ԋ�'��Y�l!Nw�����/�����������p��lN�nS���Z,u$��T��v1�&dyb�M��5�bH(Qf�q��{}�*���瞙�"�N�q�e��qZY~ZE�v��&�9�?.�9Md��
�hR�r����d��0-~sJ��Qs{}�D·���&������IO-&�k �]�hu -5���YC�
�Z����(�`���0fR-��p�by�.��]��o~$b�}���`�V� �ݒeѺ3O~�+����5Te6�&�u�={Bg(	>O��W��U�2hDɸ��0E���9l��6:2�]���O�J��d��]�o
��>���Xd]��}�"�	u	֤���ЊV�-����i���g7v-?��	ǒ�*V�:�責��A'p��i�)(꬛��W�Pih�HJ�=�g��p�-WDb������-䔐	�5|t��k�L7
�I����ʣ�r�D��)*l�iqq�;.���~R*X���7"i{*&�K�VO`�@���G:!)�3d���
-��V�ҽQe��1���  �풢�T��q��*`�+O��j�E���Bu�?@
q����D)��k�~Y�\9�w*��xm������?{��qOғ�1��[�}�� �)��>D�W��E�L���;��뇛����Y>qޅrˮ�쌘��K��Ȧ�U�}�F#@[���t���+�l���9��'l&uIR��U�whuT��jn�0��v��鋗xRʄ!"w��T�D}�N�Xqװm�D,��� ���3bM̓��4�E�Y�����3��/3`�)�c۟���Z�M"r3L����h�c�"�5JB�����c�Va�2���J���͸��q��%�{\��r�=�@�坻���F6f$�DmAñ���&7�	U�ĞslX��a��!�z�������&��+�.l�����q�}��)���Z�m��C`� l&�����g�[z��a/�_�e�ZO�������D�X1ݮ=ֿ��G�m�F��� ��R@�)oc{j$�ɂ/�V�2k�2�����и1�����v�6x��=ϰ6�Ĝ�X�<��T�:�2g�bf�VNs�ǅ�~�\+|a$��;�>��
j�jB�#�q]���~=�D3��օ%������$�ms�q��V��(^ٛ�q�A$�A�Tq���ui1q��όA��W��0�x�, r�
�2tʗE� �������-���I����$�c�����(K��e��i�����7# �/���rO�cfg�0�G��=���8��� ���Y��pG]�s��f�@lGDk˅�Z�-�7*�Z����Y�ߏ�ѳ��� �!� {_#�v�6�7���Sw�'&�#�QQ�f��P��pcr_���R_�[g8J��9_���x������)��\�B����t�kp��g݀��1�ѦnI�2/f��Cm8��=v��udp��d`ʡ2�h�<��H�U��끶�b����E97]�~̄ĩ�e�����91�l9F%��s8�=t�N'�|�;N�>�g��S���%��}6EML�U��UiN���+��+�e[|cN3�֥ڻ�4���#JBO\x	Ef����������k�>^oH��j���6[x�LÊO�̶�$A��;M��Җ
��d_@�*�Cݮ�7�_�0ux[!q���0H"�N�����.5�E�S�[���W~��
V1�n.p�*\)3���y_޲��xx�5�/,��R#�}۠�����e2�G>w�-�
�!gr���o�R,8�J�Fz�-�}�^�Dk����ϡ�4�������_��9FH�
d��S,�,7L�֐��s��c�)���{=G����$s�K��{)&���4-'\JB�@�I:,+>ڡ������+�������Iڑm����� L �T_���D�ʕ��ZG���kL)�b^J>�%/���݆Ϭ��	��$X@E��b��aM�qhOGܒ�F�C�ݣ����a#4�!�Q�:���18��y� ����0�D%3&�K��C���O<evC.M��
�܃?���ݣ���D*R�gLӿ��?V��?�:J݅|���*6>�r����G�1���6{� ���6��H_(߉�b��Ws��ͧ���♌��SSٰv�8o=j�S���
��h��ĠG+b��I�cDw���-R0�}]���֬��9q�H�C��A�٫�V�T�!%��g�nBc��DQ�p�,���J�e��SNꮻ���0h@=)�s��8슆i:�iϲL�_!7�U�v�5ɦULS���
���M�}�i"�F��I1�����·:�'
���$P;9Ǔ9�0��/��'[���"�����xV|�G+�XG�:|��<iN'|�o�Q�wsI@*�B�{R�Hdͨ#��]���� rc�UlV sZ�c��`yQ���U�Ż��w�YH8Zn���n�
j� �! ���n&����O*����:9*4;R􀢲�W����Qi�6�v�)o2�|9� à���7x��o���1r��]!�,��b!)_`��ҁ(���A2�c���v���]�ry��C�H����p+�����p����P{�e���?�	Rm�A� ������L'�--��
?��K�|'4]���OB���1>��[�˞�~[]J;�@����@1^�0�Ɇ�����gB�Ǝ�x�#���CQX�Gq���R�!�!����mD�3�P]��A|�o� ���i�}/nm����>K�f7�?̇A��.Zl�K
}�'���i�6^B�da��`����5t� �YL:s�;�n��?�\��zrzwg�aJ��B��9����89Fv��ӱ�ө��2���K����~�g<[==#��M�}� W�@t���t������^�t�'gH	8'iv�YjQgn[D}�C�As�%%�������J��X@����'�v1q2v����=���.L��Ԡ:��N�`ќ�|���3(��v��Tn�$����v��0V~��x�m�� "I�
�|d��I�����g�1Y���Gq�S1g�D"\��RLc�ҭ"}��Uq&'��ԭ�F)��m(��&��X?Z�m�U:`�'������@�G�� Rf_�MR?o/*��^U�t��6��Dⲡ�W���Tr������[?,	9}n&����x��K��xKm�!E�5w@7e,B48Xg>��EB��(���1���}-*�h���WB��W�bD�������}��1�. ��g���om�2�VΒ���'+��9�+�n�RO#�N^�jq2S�YoqVA�[9�5U�V���r��~��葧o�`,Y��mr.�fa{�ft]s����p$�F�J$�VC5�`<�-H�&������%s*Q�d�$����s/���N�����9>�����a}�أ���=�2��#4O�Fa�T�qs32������z�T4�z�Kn-<�o����X��m��2����&��Ϊ��&����|8@�[ �ڇ�̴��K�HT�r�!q��؟�J?t�}�&�)�}�9��`��i�ݮ�w}��(��r�]0��s@C���4�����k���@�m��:�3��[�܂��_]^��j�Ujb�o��CO���۽c%�,�D'����Zr�6h�����&p��H<2M�����jRuT�`�ؒ`Q��l�,��ײR?��C�#�[w�}8v����������|}R~�[�?��r�+�tǾk�.�h��%�j���5��������j����S�F�es�f�����1�R˸,4����IM mN*�dՇ�"�;����
L����PC)�HL��}Ia��� �U#��.=�L�~�lĝf��V����e�e�c�}�A�F�c@���V"�6v�H�<�S9�c���.��:���'� q��K�M��p�6A����p\}��sK���}����|j��0�,��#p7m^�v�˽��~�]�U1&: 3g;Jֽ]�������D��L �*�y�G#�2��X+? ��N������=pܵ+�����FG��W�F`��<��;�WA�Ƃ~_]4d�v���P�	��p;���%�y8Z����N�h��k��]3ݟ)��E-W�b������Hm�{��-Xz������D�%d<�do�68��%V,�k%o���m]�R�nSEL�nO=2����E�3�0�*����s�m�1��}��jj^<�|�� �>�,_S�Gn��}�.#I�M�t��}2慪Ik������p�/������?fS1�y��tS��dC�ss���CS7):��p����|Tܣm�jLcj��[�6�� Nx+9�,��wL�j�!r.w�#��s��651As]:2��1�{��S��5VQ����\�xZ�f󙊳���';�����-���3����1O�H�f9f��[�/+�u�{�t
s��d�~�L��l��8���wTZT���-����Yp���6����Y�3cR@B�,���{��[�����uD*=�oH��+��������8��޽�%�Z�,�/V�����M�v��b_�!vF	}��f1]/����i�5;�?�,�[��"�������p�\���d��2�C+g���D��(��o�bp��,4%�A���h�"m�o�����y0�Le@\.h��6�N�W�$Rw��N��dhP=@����A����mVΩ!���hv�8��&[kKZ��y.�H�>���9̙y�c�h�p��ˏ�e}i�# �����чKmo,-���utYG7*�C�_��R@��	�}���f���L�[ ��8��!)L�7��Ҁ���t[�pc�+O���?��p�z�j[��F@�� S@4��N�1��M��󾳯�Xu��i-2$2bF\S�.c���4бd���ѯ��)����}1mO㠌�Iv��B!��7��v~k�Y{��CK$V5��=r�����hf+&�@�Rb�͆�	I�j�d��l��$���$�g�F�μ���I����I��ȿB��l��p9���ta�F*��=�����WtbF�Um����D{1*�S^��{+ЛIo|g"<$�X-<�M�y�4Mb�0�y���c��7�(��"���L�\�b�E|uޜ�;K�%܁���}� �Wnq�4)�r@7�P���F�$����\PU��@'�P��K�b�Q�h[v��l�)ۿ�PIpR���{eu��;%��܈����5?�,P;F-Q��t��'��F����+�]�O��ǚ�Q|؂�Y U�Ow�H�Ѽ��:-���p��`����
��%i�-�����X���eZ*<���˪kR_'�M�`�jJy���S�&���n�f�rC�ǉ�.&gf	T�Šg���C{������񮚻GL[��"��d�]U�Ә�.���Qnlx���`niw�A���?%������i�n���S'�4T���;��F	�o	5b�eCCH��sm��݆,.Ͱ)���� !�Pվ%y8�|88�iE_6'v���iJb��7��M�w���}[Hɾ;���0肓��l�a
�'�O��,��]s�7��}QX/ M�ŧ? �1�yv] ���ck�.�8|��4
�� �QVv����2�	�j�i�.�1ԣ��t�JWg6����6�Y��gEc,�ӕ�����e ��zFK�����pD=��Ν�och���q)m3ٙ.��*r�,2-��*����L�j��F-m���i��I<������(Ih�ؼZ���|��:n6�A��IY�lD�� �iH�%26��\�B�k&Q���C�|�A�2��
99�]$g�'T���Ysm�qQtڷ}��>h�r���b�d�����g1�J���\\���ꮽd�����-�Q�����ڰ bH��_�<�����5�$؊��D�h؍���_`�u`��E�K���k����(�Mx�ͽ��b�;�� E���O5�~�Z]9�)植!�$˲2��@L�'՞�t�$2��1�t�8�d �/sYx�q��^��'*����F�&��X�w�bYg{�m]��P����TxNXkd  	��K��}����sl������&�\O�bߩ �����u��pѵAr֛��*ː�f:a�h��4j�����J0J��6��:��Tb�k��`݄I#�e�ȟՁ��}��U�.�彪�U�V^6f�)��yO�D����F9Y�:�y�&���bF���/4�]����`�e�w t�u�����&��Y�3���@	���f��	Dh>&K��ڃ�������M9���_�*���zw�� 0�>ݐ!݀�I�C���b�y�QW?�;����hD�~�s�CPf9���I��#nҺ��@�}Ԇ�n�r�8��^ΰ����2$%�f[+�!ѣaT�:�V82 P�=�8��8h���W0l�3RV¯��[�.�g�>LO<�h~���@%#.�ڲ �c��<~�gk�ݵ�s�#���=�)g�si���-�����7�;��i�N|Ý�9�C	��ֳt!�w�z�MJF���c8F���}���V/�R�%�q��<�E�~d�n���V��Z�ݚ�
ަV��P��i�l��O���T1�a��b�g�)������;O�}�SK/��M8aT�H_�(�X�|G$+1���TT�=#��E�I��$8�p��RY��܀	�@��Cg�'�����9Mڪ�1s�r�۫l�pR��Hm���81��w�Ɔ�D�c���a��}�_�B�W}8q��0.%��X�c�-�>La/�.�@�i�����%�9:It���a��a¨Brb�)ȳ�C�&&��Ag򸚴Ǡ�o��y�F�C����Ү;����J��X{+�ެ["KXE6���jL�o者�Y���#�k8^�V�9��(��6{/�E]�1Qd�������"�,��5IzW#� j:F����a�4�Y-7�s�7	�4�Qb���"\Tj��s��Y�h��)ثh����D�A� bCPGS�Џ�\)�^H����h�	��NT�������'�U7O>!`1k[3RM��5�"��0|��o?�� ��+�� �]kY�6�n��K=�ox�!lv�������N���=q\��A���%%��g��4��|le}���f�G�u�UZ�1�e}5+یQ�gi��Ȼ�M���̼6��8dB%�;'4Xz�:�VB;('9|I����� Q�`QYh����}�#�0��Ҏ���;ʜ7r���#�R�}>��w��1;�TY7�N85�N{�JֹV�#�:�8$7O���'�0��^��I����rBU �<{�yȥ���|�ݼ��I�9?]W ��;��wpI�Z`�� ��תo�� .V�O��;�I�U����9T�%Eh�q�� ��/��� 7��5��
���]�����I����p͜~���w �K+�p��?�:դ�~I���8sO�����w�R]#��,[Güɫ���L1��e��b���>W�D5��n�S��+��������-U,p{�l��(���Ծz5G2����B�	��p�v�\���0��o�U����3Ҍ���&o�2�-t52�M��T���tw��!��6���i�E���Λ+�:j�X����3���X5AS�WR���Y�xͣ�H��ɸ[������f���+\�Tu��6��٤��}��MO������V"�΄QS�kbބCa�8x_7C��)g���A#��SPՕ��@�_�T��H�WMx1C���&|u�0�#�Y�~zY-vW}E�S哂o�6�e�-�Q��uœ����3��Y���������4^'�0��x��A00�z������SZ�~	
��z�P��L&0�C?v ��}8l����@��z���;�R�\�
���ɿ� =g����X�ڥ���	�O�:������oz�v	W�@�����;B��������N�!Kh"��{}��i$���.��C;萒���!���]�Ǔ��,>`�5�tD���E{��l��LMy���b�ANP�h�}��B5#�hyx�D��uJ(�Q7�����N&qc�d	��u��;}�e}�ײ������}"�E4��c�asH�|â���5��,��뭟"/���>I@�ڱ ���G�ԭy���l��'�R�u�p
E�9���X}�9k�����bK6�3�Ļ��Vݦ���6�]>�b����ql��E��!'ǽU���I���\�Ś{9<L��v��������.�њn��2���Kq�C��LJ�q{I�fn�Q3$8�����Pnn#E���B��Kaj�X쇗��H���e"�6bbWz��a>Q�.�'���e��>ON�����_��xZ+�ﾉ�6A,/BT����|B#�vq�V���$�<�AN^��6�����k����N?�i����ď�?�]��\H�2�:{>�8&\~TŁy�����R~�([|Щ�t7V�n�-�-r�?���Чf�<�?��[I��	����I�Sk� /�?��#�0�ő��vYQ���+��:�G��Bf�A+�>�N�t�����Ř��qk�?'gUՂ��0��
jI�9p	�p��q��AG4Ur���ܵI����&v�W��V �J>r�3�k��#������*��һT�~@=�8m�'w�.�h�I��n��K�� ��B��p<�lo�j�7��l#�����F<R��"aB�sI<d��X@��&��LH ��91
��Ђ���
�視f�(��vu)8vo�7����J(������&���'x���^Z��VS<�7���C��h	��~���p��?2�&T�֔U�2R�&�g?��Y���ڃ��s��)z1��[0���7���m��<�l���&h�!� �n�{�0}G��F�뗎_���zk>$���]�̅:�	�,M [j��O�65�Kqϼ ��X�~��D���Yg��+>k���Re��:����������X�%6���{��tuW���L�8���@��J�6}6
g�l BW�)�~�s4`X����W�'��ꋹ:�_�Rd��a��2�Q@_
�F�|����Q}A� ������Jn��?/��ҎC�V�/$������v�C���U@Eб�v߯w-��%~���\ec�D48���T��CL�AܶS�F<3O��2��W2~++�F/�J�Y];��ZY�6e��*퇖N+A�ʲ�d���r(�̚{.��E���6�2��1�`�9n��&ȁ����h��Q�ZR��]̑�Z�7*ҿZ5{��B�� ���a�aM}�{^!��Xwc_�u9*i�"��&o�&YްD�74M���R�~��A4�o��a��n��i�>�����1��ě��F����9gߵ�#�ƣ*�8��㱸%AVjO�(��!xMh�/�������"�נ�B���V�\{�e�E��	������v��b�[�ѥ'��g�����i���EY~�ܔ�����+^��&R�I?T�c�#4i:_�� e]f�r�g���HbD�
�N�����
;(e�q=����3#�Ypw~�p�mwn�@ܙR+5zd~�B�����][��ݏ�X"�:�e�uڎ��w��~� p%�z����+��>d��50--�0N>�=Z�ž����o�O���j�6R#g��މ�����W!χE��^\�8f	�����W���R���Ϯ�,�*)���0:�����}X� ��g��#�P�ط����5Y�+4�6,ϸu��mVA UMr�����j6��O�{�S�u��p���b�:	6$2��xtAT���o�;�QN�����:�<�t�$&�(|��B0Ӡ{O���N�H[ 8/ �N���`�g���˺
��e�첸���.��3��2��⢉��K@c��vM���������� �P+��Kw��}=�"���I7[�k�ǳ[���6.��m{oG�e*D���� �4�Z���I�2� oB2��JP�G������cU�ɘ��1v>o5 ��]"�wV���.B15���#���
Dw�t�t)W8�p�T�ӓO��9��}�۴��M�<��Q��1�2��p:mlWf{ޫ��2�I�LV�[��_����A��&�W�,4o<�J�@
m�C�_�n�B��[��ʡ�Ԕ(�ƣ0���.�qx?H:+2��M~����߸q�Y�h�6+Ai�W��_�nU���0i�|a����m ~�|'}�8���d��f��:�����l��v��JS�М:�g,C0� Ћ���W�No�׶K���#�3
K�fǝ��)�O�ח��4q@�*s\4.�"Π���)ڃ���Yp�Vu�W'	���z���Kh,� V��VWȄ��+	�X��ȥ�j����b�7����{��� �ì<��
��L@p@��1 ��~Fh�N<�����%qS+4�*^-\r���:λ������� D©�~��j�5J������7t)����Dy+� `u��l�)�/O�~��35��3�S�Mܼ�}��K�1�q�$�s�tȦ}D���WNi��!�6V�}�/W�1,	(���E&~a�K�Ʋĭ���C�ѝ�d�I���ө�:c��U�k�<�M}*��U��!��)6b���5jɥ=&Jt���#٣8�Lk��cfN��g��=���߰T����42k\����s�C�@Ha�1��|�~����GԄ	.���������@����r��9����houU��sȺ/�n�X&kI/ek� T���pV���/L��RP'鹂��z�! T�Ďl�L�zq~C�[ $�J�G_�Y ��*�2��B_D���^�w�9��D�.�9��ڬ��n�R4'5�S�f��uk`U��?��(�i	L�)�5��a�\\1�D�P��y�� �]��{�NM��j���I��i.�]_�y~̸S� d�!×������f�����%m�#	�M&B������G��r�t�R��#fY������h�z��`�B˕?�GX:�L2A�K�ıƐ�`l���޾��lsu�������B$�I(��>��C��f����]�(ps�c��S��|:i&�7�����t��wBG�:�,�^
K��J�M�/�,�9�Y���չ�Py�8>��`�%��~��^`�(A;S��=܉��(�v����I�3�o´V�GA;�~v�H,�Z�^4)�,f�:����B��ބ��I �aK��6��9�c��ɔ������Xވ]еC������4
���MXN&-����\Y����g�GgP��rF����⣼��ʠwY����`>�D9"k����VT��H%!��B.�_\gZ����C���0K\pc������sa����t��ߥc���*�����\1����x��-?	�I�O�YD/�8G��Q��y-9�N5���p#�Y%��](�g�-�$�<J�3IՌ�3P]r���������|���b�=_d�u���	;`?O���ӑ�ef��P#��y���)�g�L}�Tv���{�E�Z�Ic�$E
6��Bz��/���%9���[��*�����[�w���+��9[SI"�R�LU,�*0Ħr_&X�û�>�؈��vLt�!��P,�MG��S�:�9�06�R�R�Imu����b�|�H�9.�7�d���^��y��>8oC6�3co�
/�4���a�I�kߪ�����]�Y`�`�����G�0D
W(��K���.Y�O��1C2�ފ�Ŋ\�7u�x�Z$<���d��c�4�h�)R�
�W����(Y9kχz�-�3:s�MX�lk6���$g����Գ�F�}y؟�z���Iڂ-=G��D��vHq2���?r'��v-��ql1��XV9j[ӫ3�GE�R7��GKd1���Jk�����i)�Ǐϊ|+[q,�y� �F�_����N{���ؐ�Q�e�`��z���%O7����@\��>�����u<���j�,d
̑|婏%[��ֽB��D*��vxeh���%ce�APM����/74�s۸��|����]��5M;��zJ^y5a���:�=� �N��E���4��G�U^�u�a��|ACx���,e���g����S6�:綺R�)�7�H�-�MZ֖�ۧA��g����:8 �x�z���E���(.�}��&-,���G�w,T�/���Q�V��T 5���=���!��o� �i�
O�i�Yh]�?��hk��Oy�V��m?�a9E����&�E�
Lݿep}0f���7����2����ۤU͂���R��ʼ��zL�"�����I�������(ު'�%Z������U"�)Sz�% f��&T"YchN�s�G�������KAF���'ҥ��1q�|e[�-z��&���`�k�ѲZ`g�0��Ϲ5U�=�RF���lS@����F:�7��(��vj�V�j���cR\��<��w� G�`:���|:��wC����ۣ�[���"�%�,�a�u�i����C!Z.�6@�d�F�9���m��L:k��+�K�+x��>L�2T���#G�$�#A��p�5���`�����3�m�ߛ��.��S�%����)��w~ϭ	Bj�Be�<�|��v&���4b���=��~�!Y.3�1nq��;$޷��Q���	�y�������R��u@ߛot�Ӻ�Y|�-�$�*Sr'�y���U�F��0��<��E8ߡ��B#�3�I���F�Y�@��*F �|��4㏝������0���+�5�[�?d���gq�hQ�:�H���W@�ks��$5�H�$%���~�K*�-��ݩ���|�}z�x��|��}G�VSh���a��1�(��n6��x����G�G.pKi&�kle�|9,�aI6l����y��i���F���,��
��q�u+I��vI�����꺟����*�YJ��	���\D&}���v���J�v|0���2I�Q;x��/���D�����)k��#�c�~Q�qG�̋����
;�"��K��P�.H����_}�qऒx8BJ�!8Ռ5 ��'�Ep 5��'O(��y���	�+��H�-}sZ����6��CV���J����$<y7��� ,"J��iʃԡU�����;hGX!=£�|�+y/w�S��X}�>v��?�h�g�U��ՉW)V2��<�?�y�b3@�ܽ"� ��V �_qxr�0���XS��3�C��s��[�"�q}W�W�sql�J����~_�s��N�I�z��d���V�I�`���孔6e  �/۷V}z�Z�Lm��K�+�d��+����P>���g&�ܮ%�c;	�o"(��$�l��Γg�<$��(A�0�D�>l6��z1td��ϳPj�o8�I�:d��6ALhg��PQn؃��&+l��ا	��tz�*��.�C�l�Z*H��U����-�ބ��?��Q�������\?�Z���$��)��Z�!��h:����*�ĭ.:��P����ìC�����=��B��a���	�^r�/R��0�$:�Z��xPN��_��ثb��Xff:���H�H8^V.K�Zi�ݣBS���
����r��0Q�"R�X#�yP����E��*9Y�������������oj�����I�03(�#�6KNd�y1�(ې�w�p q��]Z�J53;�Sf,�dF�y��d"DV�J�b}c�( ��2Ѡ� M0��d�u���Vl���-����qφ�ѵf(���.!`�m1�nX�:4��'����& M��)�B�M�������/�������+�H�?V�zK�O;�DV��$���G��\
yr�]*��&�ڤ��͏^����'��. 2y�1-�������Ԍ��~�Qk6�㝤u�{f	`5���)��@���>�*����T-����$�q���ŝ L{΁j�n�r��?o��jbOq5�="Oaâ��2jN��X��ǳ��@M��1�ˆ��X!'DIK��aiS���7d�4CoXg�w���u����CQq�m�V���{��-�^���z	�j�\-m0�	����NG��mF��uv8�^�pS`Y���{��K�5��>�l)�';�=��ŕ�11�U��<)������B�עJfwN Ӈ�1r��=iO��q���C�H����Ԉ�id��r<v���r�h�prb��Wn�S{�V�m��y�����A��%����|s������`E�f�U߶�,w�1q������^�-�7=�x^U(�5$����>@����,*�G��n��iq��D�R�2u��Jr�9���w��.}@*-�|����^ء�Y��?_���4M�^��y80%�)�`&㨠x��ݯ�6�?˖Y�Lc����3aV� �N�42��ߤT2�WnV ��ʞ��O������ ���3[h}�*L@W��e8�LR_j
�@�f�|..��^���u�0��:���~H"�7,ϟ���3NWDf�\;�-uY֨���6�ȶ��R|p�U�?,��܂��3,�F�QBgٞ��m�u�2ΰ�+
�M��gs����(J�դ�B��gJ�]f��IQdT�b���d�k���Q��C O����B{k.Xp�R}ܛ��6��\U�Y�"(>�G����~N���Q ��H`K����j���,!���T�?��ґ$���s���kAS�3����zN�  z)qP�/c�8>#ҕ��:H��K|�~=�qU"���Ҡ�:�-�4t���!�W�uȟ�	�)���?uuC�S��0�i���B�	�m��,	 �5Ҝ_㝌�����XGsN,�ڨ��\��-s�����Nc�I��5;ח��jp�a��Aw`E�.��ӸS�^��GcǖfJ;�Ʋ�X��������J!�J�6$y`����;���~2�� �IԺI�x�d}݊/�f9�h�.�V����o��^�PPm�?sḂ���ES�-۶WEB*U��3��@Sp#�ÕS����g^@�&���EU_��@�T\�c"�%��,x���cs�c��U�B�5솚�gcO[�C`�,K��tY��:+h>N5ʵ}y>�����-�m��#������&[d�&W��!��:�_����W�*�������L��B��Õ�u�s��5-�e�*��s���(�)>�1�xkshwM�;�;"ys��0�A�S��{ CH�~��x�g��*�J�d�m2d��''�dH��|��4؞%�e��s�>�d��������� c��5�!��PG��Hm:*�9h��{���7�&�_qР�^"'��^#P�������D`�|�p�R�����x�i~Jv�;��i��C�v�Qa��1ݖ�K{+R�� eQ�N�&&�v��ben29�xY7���цS�����<FRM�O�A��Z�$�<aʏho�Y� ���p� .�c� �c}�g��J��&��Pȣ�R|��A_���=���p�,a�BT2\����H-T��[]����F�Y�$�gk��j��c)&lS�'׆7�AlO\���\�j�Ԍ8�萨�ؘvp�T��҈�*,H屌���EQl����E��w��U�ԷC�����R�i�p1�j	o߼�u	e�E�o\eы ����/a�|�ȵ~A�y�>lh�.�����݂>FB~��/��V�h���7\X� ⱔ�D�U�b0\_h�Tr��/t��-l�_������{��z�H]_��6r�m��J��`_$Hvz9@N`�,��6Θ2Vhi�YT�*#
gZ��P!.�b�ǟ�n��_7LԲOsI�Cن!R�AR����kv{��N�֊~���e] ߝ&�/�5��\��֖˄[��\"��?v���;6Jb(�����,5X�2s�)j��JNq�������f��W�mY��Gx&�[���ٺ/a�(���	�5���X8r�V*�G<�e�%~*XL� 	|߆�n��M�	~��=���m�(��;�
	��_��GI�,?zY0�s�WC��qM'��KĲ��� �����ۤׯ�@^�R�Wx)Yk�Ռ#|��E i��DX�c�g��?i<�qB�Z��xeM�ģ=�^t�	RU���C�T�*����|a�nZ+qo/�9+75n��-�C'��+��e��.�m�I��C]���N<2-[u`���2h���+�e�P G��v����w�+��),3F�@����a�]�!�yd��Q_	�#*;�ߙv_�z��ą�O'�\���X��3����4���EB�
�����R;�W�6��m�]`FH��Y�Vx[�(�`��Mkx�X��Л�Qi��s�b�Y��8u*�[�-�ආ�2��Mx�����
: ���*���	�eOzി����5e/��4���rd{�0
���UR(�+���v/���Y���v��<|)���`�lgm,�z���e����I}̟$�D�*�	�K�β���%O�U�z�������HN�#�j�<`ͤх������G�&��9�� ��ÖQ���S�@LS
d�����7�޺���e^j���*�{�[�y3W��i�q�i�I��}
�2V�^ضoե��7�,��xB�56��]n��i�շOE����ܬ(7mĽ�:��8����a��W�9h�v����"���c�6�pLAp�Ǹ��xpƦ�π�u"t�(ء�S�pMc���Zy��kU�s:�X闢F����;��gb���(����j��^s�c��L�4F�u����h��X�ˢ\/��Y���t��(�s�����7*�u�! h�K>�老�ގ�K�\RD��D¡z�dО&Ù��b���r3��	� 	z�Xl�Q�ܓ׫m`\oY%[�5�LM��v5bJQ`u��>.��4@��%���/
��^�pL\8q*�[���} ��̩��^���#�g��]�:gf����c�A�BmJ���m��ã�#�Ђ��rKg���p?Clg°�JV2��0�wL[b�G�2E���y �0'�J���9�C��IGv�+z&�"�1��S5$`oj�e�q �o���|B͌�S&�q8�&���y�I{��һ(R�ز/�:���_ȪS��FA��o��:��߽���n��5��|xFaO:�]������4c!��Z�b���3b�bk�t���6��.V�ǵ۰�B���)�U�ml#�8G+R��΀��)7݊�&���u�tڊ����}e �>�#~�xuZ�Q\��I\���_��_���; Fΐ��v|�c������Ǟ752����o�S���X���g璶y��Dфf����O�1!X"��L;D�J�Ԛ� �
�G_ň�G�������\\�kV�Ƨi��AM��k)3�i�N�s� VC}�٬`�"0~؎̜��8z��|��|�v������'8P'��w߁A�Ҷ�.��^���L����J1h�Dv�FM�hvt�*o6![���3b�:���LC�K�Y��T��*%SdҊWW�X_� 5�#3z*��I{N���l�� Fh��w�B=������F��nʽ���E"\.m,QHSs�U�!`���=����q�@���R5 ��@7�;X�*"�n՜m����w%���ɜ��W[VV-�A�Q�郖�p����u�:/-Yyϻ:���-P�Y�q������A.	�-���v��\*���.�l���ƺ˝ϰC��z�jA��8R�I>_K���H�+t_j4?&;�ͪ���L�K�j�{�DL/���Ž���y@�����q �����Y�=��:5�b�Y��ֺ�]���~��Z�h�|T��]V�U[x!�!�ҩN���֦��-�+�Y��Č�>�c4�eV1v�d��E���dٰ���G�c�f�����mpԒ:��'z�ܹ+��jT�/F���hR]��U#�����j���jf�#@8�*�ޥkV�(�[YǴT�-Ԕa��0�U�r�Hb�[$���u��Eu]l�����Jp>�_�f���sȂ_~�";�����r��X�S�>UHHӔ�o><���κ���oc�a�VL��b �(,-�e3v��@�.����-]����7��k%�0��5&��a�s�{�p�#)�=�Y�GznD���J����w���a���-�{��W�n�0�)��M��s0�F0業ㄋ��<�Q���$OD[[H�a^dH��Y���`w��B�s�5�ѹcb#��&��`ş�M�*P��x�����˫�E�:N��5�%d���=�ޝ��� �ɽrA��qe�t��EA����A��S�"�����#�k���Q~gTa��/G���r������jO4��������}� u�,����S'y7�b �À���~��5�i�&�em�Ps�Y[ɼQg����m��M%Γ6iz��1�h xB�M|68��4ė�GR�H�VGj�.	�, �VhQ���?�/&Z��iS\��<|�� Q1�Ob�䯇.�71������U�(��]^ H6o� "W1��_Ņ�$�e9�#�ÓHǅK�����'��F,�l�$�L��� �4��c����1�LZ�^����v%�6~K(8�ϏiN�R%�dSi�'�D��/��I����i\�x��̩�؂x�Δa/G��(𐃟�M׫��� �hE|�����6g��B``ފ�.��!���lr
� Mk*oS��?�@j��eרEkӫ�һ���z��J4��`�Ӂ����j0���O����u��Z�=����X}0�����N��a��};=>6���Cs	�N����P՘\��^D^�	�G����N���C�ز�D^u�)�Ӝp�񘮜����b�6�p�"6o�B.���N	�s^\o*;	�%=�Gv-\3��3��A
�-yR5S�p҆7/�')k<�F��n�#����d��$�o���X�G�Gj�Ȼ���Kr�-���wDB�S�2Zߴ�n��t�ܞ#��QY�7�� +� �n��<��e)}$���Ò8����2�w0��G�Ħ����o�z�3Key
@�}i�&�׌���X0=�u�������&\���B�&�rD-��lZ����������)�'>l�7�"D�i�s@��9I;E�^Go�}���������40_�*&�@� ��q>��7�/*�\�tQƒi�����Ų���0픥���
�X($���.���f6�㘀���F��Z����8!�5��f4e?u{�&R_��E����hڥϮ��7:��Юз`I�A0���2���cԥ	�1���<�e8GƣlE���uN�;ӓU5��~�a=�sI� ^�C��|� Xۼ=l��?������B/zc��v|�1nnĹKARj�"qٚ,ĺz�4�rw��^�����3�7��k��S���}���0#C9��l6O[2�Y��"A(B����\�t�������(�<�أN��SS�6#�#!qE�}���xibEc=���?���\�2D�?*�ⰶn�U�4��u�,L�/ȡ>����cE�	#l�y,������H���f�4��ƶr�_�l����M����¾j^J�h�]����KKd���W����uV=��KI��(C�HË[�u�b�6���\�a�R�* ����-N)A�{�ԜU�$�5ך��X��?��n��2��Ėa����!`�V��a�9�b����h�+Q*���(���$Sx.����<h	2Cՠ�bhzGMGp������@{���я#�` fb�q%��[	m���X�4�l͚��/�����F��gӋ���J��'�l.�y7�ŭm3[�2	בt�l5ZP^��[�,�O�ZJ)v�{0�+��@]&���� l���{�������]��QV#YW��L^����lvZ�S��.�ڿ�"�^�zG��V�<0l����]i����<�P��=��sE6nb�J��>U�m�Ko��إ�)oO����?�Td!������}��%u�xx`��3��C�T�jr�j�*�렏���u͈��7��i��$��ܘ2��~3�j@͚;�`����� �nŐ�n3��Eb�q(����/����i3%ؖ!�zoP��(lb}��hے�O:�_�5'7���G[0��n~�>�Gd��h�z�L����G/RxD�d���Ɗ+5�~Ծ�0w���@�齝���jE����W�*���"ܬ��n�f*~�Bb��/v���]Z��ܛ^�ˌ�4�3BG�ץ�V(7��`�k��n0��'M�"���@_A�n�q[-�tj����d�]!Z��3�ڙ�a��Bӱ�)��9Nˍ�~J��| �Y���m~%D�d��]>����:󜨀@խKxcX1�zLj���U����A+�r��s�[�s�^�~���[x��wd��|W��zA�3�q
=2=pd]�k�}��	>�[3U[!��p/N�?�+��o�fފVM����j�RH�����\q���g��ިr�4g(��u����X� ����J$���w�D.��/m�w=�"-!�N����gt����Q`�aK9������^���8e�L7<=@]�M��5t�D��,�Q=�~�d���W��˕�1�k�s��gDjП�H�uP-su�Q�Pj�87^q�"_YM��/��*�Âgabt�:��d2;��SA���!u� ��ܑ8��\B�;�݂�׺�gn�h/"C�-E���!UM:��qtL������V&T�=��e�&��Nh�iԣ��^��/�v)_����t�$D�*�:��R[k�&
rݐ�<��d�2�([M[[H�Ü���!�#��c�D3���V������BȲWG�4��o^׈�ԟ�K��":ns�;{��E�h}���QB9�s��Ѫ���t�ղ�&��
d_��<0��o�f�g�,L�6p�M=.#�.Ob�d��RP�Z:��6���Ofز��Q}Ԩc/��l%�u<���՛�OYd�r��DD�-��*^�����:Ċm�p`��((qG�o*T!Sۅ�����o��X�����i6ш����^�ʱ�؄_�`ՕX��~��qxD#C	]qJ�ޕZ����e06?�Oi�6�ط�)1����KK��A�����
.�ly*��~;�`�����P~��[u�JB�����d9a�C��1��0t��p��V���?�������QCg���Z��?ifZ#�U%�Tq��U�EWd	&yL��:Y���к��PD_�ɵ�K�|f��M�dU�q�D�*�5�؅�(�9��:�����`��7�z�=��ƹyZI����g�;
9^Taj@z61����u�"��L���C�ݤ�d`�Uv=���SQ����x���h �+]��`��]���,��Wk=G<F�Z�s��{���b?e��`ܻ���Bͯ��ސjJ&��B�v_���r���Y��ŮK�]@�52�.S`V�ĝ�WB�L�rͽ���!�����`����{�`�矚4)sP����r[���o�h��P����������BO������%�q5 ��� �ʨL9��c���<�r!��`���¡����?7c�6�j����4�G ���d����t��^(gc���2�+(��\��f&�$��1�1S��d>�~�1��P�L�_����D��>��;�R���s�T�����'m���q ����XFy���^�l�K锧#�t(��U��Ů�O�+v4��U�.ܿ�(i��=2S�������O}�idOW\��|��p�8Ӛj}��I&�X���?sx$�Z
Ni<�Ӥ�G�r��U7d����(����]�ۈ<�����/��A�~"�G�za���^�6z�A�A���ER[QB�U�d*�y�7� P/~탆e2ɩU9�����~~���a���H}H�D���j�dk��ݭy7F��&�����?��W�̹\��|s�/�d���P���8X��˂���h�v-�lCG���fH���x�[	�O�I��d�s�ɳ%ӉU��0��?���7�8�_W^H!R��8�0ͨ�+�