// Copyright (C) 1991-2012 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II 32-bit"
// VERSION "Version 12.1 Build 177 11/07/2012 SJ Full Version"

// DATE "08/08/2014 20:53:47"

// 
// Device: Altera EP4CE6F17C6 Package FBGA256
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module fft256 (
	clk,
	reset_n,
	inverse,
	sink_valid,
	sink_sop,
	sink_eop,
	sink_real,
	sink_imag,
	sink_error,
	source_ready,
	sink_ready,
	source_error,
	source_sop,
	source_eop,
	source_valid,
	source_exp,
	source_real,
	source_imag)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	inverse;
input 	sink_valid;
input 	sink_sop;
input 	sink_eop;
input 	[15:0] sink_real;
input 	[15:0] sink_imag;
input 	[1:0] sink_error;
input 	source_ready;
output 	sink_ready;
output 	[1:0] source_error;
output 	source_sop;
output 	source_eop;
output 	source_valid;
output 	[5:0] source_exp;
output 	[15:0] source_real;
output 	[15:0] source_imag;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_sink_1|at_sink_ready_s~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_error[0]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_error[1]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_sop_s~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_eop_s~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_valid_s~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[0]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[1]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[2]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[3]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[4]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[5]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[22]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[23]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[24]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[25]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[26]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[27]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[28]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[29]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[30]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[31]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[32]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[33]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[34]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[35]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[36]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[37]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[6]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[7]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[8]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[9]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[10]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[11]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[12]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[13]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[14]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[15]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[16]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[17]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[18]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[19]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[20]~q ;
wire \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[21]~q ;
wire \~GND~combout ;
wire \clk~input_o ;
wire \reset_n~input_o ;
wire \source_ready~input_o ;
wire \sink_valid~input_o ;
wire \sink_sop~input_o ;
wire \sink_eop~input_o ;
wire \sink_error[0]~input_o ;
wire \sink_error[1]~input_o ;
wire \inverse~input_o ;
wire \sink_real[0]~input_o ;
wire \sink_imag[0]~input_o ;
wire \sink_real[1]~input_o ;
wire \sink_imag[1]~input_o ;
wire \sink_real[2]~input_o ;
wire \sink_imag[2]~input_o ;
wire \sink_real[3]~input_o ;
wire \sink_imag[3]~input_o ;
wire \sink_real[4]~input_o ;
wire \sink_imag[4]~input_o ;
wire \sink_real[5]~input_o ;
wire \sink_imag[5]~input_o ;
wire \sink_real[6]~input_o ;
wire \sink_imag[6]~input_o ;
wire \sink_real[7]~input_o ;
wire \sink_imag[7]~input_o ;
wire \sink_real[8]~input_o ;
wire \sink_imag[8]~input_o ;
wire \sink_real[9]~input_o ;
wire \sink_imag[9]~input_o ;
wire \sink_real[10]~input_o ;
wire \sink_imag[10]~input_o ;
wire \sink_real[11]~input_o ;
wire \sink_imag[11]~input_o ;
wire \sink_real[12]~input_o ;
wire \sink_imag[12]~input_o ;
wire \sink_real[13]~input_o ;
wire \sink_imag[13]~input_o ;
wire \sink_real[14]~input_o ;
wire \sink_imag[14]~input_o ;
wire \sink_real[15]~input_o ;
wire \sink_imag[15]~input_o ;


fft256_asj_fft_si_sose_so_b_fft_121 asj_fft_si_sose_so_b_fft_121_inst(
	.at_sink_ready_s(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_sink_1|at_sink_ready_s~q ),
	.at_source_error_0(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_error[0]~q ),
	.at_source_error_1(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_error[1]~q ),
	.at_source_sop_s(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_sop_s~q ),
	.at_source_eop_s(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_eop_s~q ),
	.at_source_valid_s(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_valid_s~q ),
	.at_source_data_0(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[0]~q ),
	.at_source_data_1(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[1]~q ),
	.at_source_data_2(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[2]~q ),
	.at_source_data_3(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[3]~q ),
	.at_source_data_4(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[4]~q ),
	.at_source_data_5(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[5]~q ),
	.at_source_data_22(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[22]~q ),
	.at_source_data_23(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[23]~q ),
	.at_source_data_24(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[24]~q ),
	.at_source_data_25(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[25]~q ),
	.at_source_data_26(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[26]~q ),
	.at_source_data_27(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[27]~q ),
	.at_source_data_28(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[28]~q ),
	.at_source_data_29(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[29]~q ),
	.at_source_data_30(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[30]~q ),
	.at_source_data_31(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[31]~q ),
	.at_source_data_32(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[32]~q ),
	.at_source_data_33(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[33]~q ),
	.at_source_data_34(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[34]~q ),
	.at_source_data_35(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[35]~q ),
	.at_source_data_36(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[36]~q ),
	.at_source_data_37(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[37]~q ),
	.at_source_data_6(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[6]~q ),
	.at_source_data_7(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[7]~q ),
	.at_source_data_8(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[8]~q ),
	.at_source_data_9(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[9]~q ),
	.at_source_data_10(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[10]~q ),
	.at_source_data_11(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[11]~q ),
	.at_source_data_12(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[12]~q ),
	.at_source_data_13(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[13]~q ),
	.at_source_data_14(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[14]~q ),
	.at_source_data_15(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[15]~q ),
	.at_source_data_16(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[16]~q ),
	.at_source_data_17(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[17]~q ),
	.at_source_data_18(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[18]~q ),
	.at_source_data_19(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[19]~q ),
	.at_source_data_20(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[20]~q ),
	.at_source_data_21(\asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[21]~q ),
	.GND_port(\~GND~combout ),
	.clk(\clk~input_o ),
	.reset_n(\reset_n~input_o ),
	.source_ready(\source_ready~input_o ),
	.sink_valid(\sink_valid~input_o ),
	.sink_sop(\sink_sop~input_o ),
	.sink_eop(\sink_eop~input_o ),
	.sink_error_0(\sink_error[0]~input_o ),
	.sink_error_1(\sink_error[1]~input_o ),
	.inverse(\inverse~input_o ),
	.sink_real({\sink_real[15]~input_o ,\sink_real[14]~input_o ,\sink_real[13]~input_o ,\sink_real[12]~input_o ,\sink_real[11]~input_o ,\sink_real[10]~input_o ,\sink_real[9]~input_o ,\sink_real[8]~input_o ,\sink_real[7]~input_o ,\sink_real[6]~input_o ,\sink_real[5]~input_o ,
\sink_real[4]~input_o ,\sink_real[3]~input_o ,\sink_real[2]~input_o ,\sink_real[1]~input_o ,\sink_real[0]~input_o }),
	.sink_imag({\sink_imag[15]~input_o ,\sink_imag[14]~input_o ,\sink_imag[13]~input_o ,\sink_imag[12]~input_o ,\sink_imag[11]~input_o ,\sink_imag[10]~input_o ,\sink_imag[9]~input_o ,\sink_imag[8]~input_o ,\sink_imag[7]~input_o ,\sink_imag[6]~input_o ,\sink_imag[5]~input_o ,
\sink_imag[4]~input_o ,\sink_imag[3]~input_o ,\sink_imag[2]~input_o ,\sink_imag[1]~input_o ,\sink_imag[0]~input_o }));

cycloneive_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~GND~combout ),
	.cout());
defparam \~GND .lut_mask = 16'h0000;
defparam \~GND .sum_lutc_input = "datac";

assign \clk~input_o  = clk;

assign \reset_n~input_o  = reset_n;

assign \source_ready~input_o  = source_ready;

assign \sink_valid~input_o  = sink_valid;

assign \sink_sop~input_o  = sink_sop;

assign \sink_eop~input_o  = sink_eop;

assign \sink_error[0]~input_o  = sink_error[0];

assign \sink_error[1]~input_o  = sink_error[1];

assign \inverse~input_o  = inverse;

assign \sink_real[0]~input_o  = sink_real[0];

assign \sink_imag[0]~input_o  = sink_imag[0];

assign \sink_real[1]~input_o  = sink_real[1];

assign \sink_imag[1]~input_o  = sink_imag[1];

assign \sink_real[2]~input_o  = sink_real[2];

assign \sink_imag[2]~input_o  = sink_imag[2];

assign \sink_real[3]~input_o  = sink_real[3];

assign \sink_imag[3]~input_o  = sink_imag[3];

assign \sink_real[4]~input_o  = sink_real[4];

assign \sink_imag[4]~input_o  = sink_imag[4];

assign \sink_real[5]~input_o  = sink_real[5];

assign \sink_imag[5]~input_o  = sink_imag[5];

assign \sink_real[6]~input_o  = sink_real[6];

assign \sink_imag[6]~input_o  = sink_imag[6];

assign \sink_real[7]~input_o  = sink_real[7];

assign \sink_imag[7]~input_o  = sink_imag[7];

assign \sink_real[8]~input_o  = sink_real[8];

assign \sink_imag[8]~input_o  = sink_imag[8];

assign \sink_real[9]~input_o  = sink_real[9];

assign \sink_imag[9]~input_o  = sink_imag[9];

assign \sink_real[10]~input_o  = sink_real[10];

assign \sink_imag[10]~input_o  = sink_imag[10];

assign \sink_real[11]~input_o  = sink_real[11];

assign \sink_imag[11]~input_o  = sink_imag[11];

assign \sink_real[12]~input_o  = sink_real[12];

assign \sink_imag[12]~input_o  = sink_imag[12];

assign \sink_real[13]~input_o  = sink_real[13];

assign \sink_imag[13]~input_o  = sink_imag[13];

assign \sink_real[14]~input_o  = sink_real[14];

assign \sink_imag[14]~input_o  = sink_imag[14];

assign \sink_real[15]~input_o  = sink_real[15];

assign \sink_imag[15]~input_o  = sink_imag[15];

assign sink_ready = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_sink_1|at_sink_ready_s~q ;

assign source_error[0] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_error[0]~q ;

assign source_error[1] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_error[1]~q ;

assign source_sop = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_sop_s~q ;

assign source_eop = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_eop_s~q ;

assign source_valid = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_valid_s~q ;

assign source_exp[0] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[0]~q ;

assign source_exp[1] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[1]~q ;

assign source_exp[2] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[2]~q ;

assign source_exp[3] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[3]~q ;

assign source_exp[4] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[4]~q ;

assign source_exp[5] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[5]~q ;

assign source_real[0] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[22]~q ;

assign source_real[1] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[23]~q ;

assign source_real[2] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[24]~q ;

assign source_real[3] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[25]~q ;

assign source_real[4] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[26]~q ;

assign source_real[5] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[27]~q ;

assign source_real[6] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[28]~q ;

assign source_real[7] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[29]~q ;

assign source_real[8] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[30]~q ;

assign source_real[9] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[31]~q ;

assign source_real[10] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[32]~q ;

assign source_real[11] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[33]~q ;

assign source_real[12] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[34]~q ;

assign source_real[13] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[35]~q ;

assign source_real[14] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[36]~q ;

assign source_real[15] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[37]~q ;

assign source_imag[0] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[6]~q ;

assign source_imag[1] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[7]~q ;

assign source_imag[2] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[8]~q ;

assign source_imag[3] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[9]~q ;

assign source_imag[4] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[10]~q ;

assign source_imag[5] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[11]~q ;

assign source_imag[6] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[12]~q ;

assign source_imag[7] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[13]~q ;

assign source_imag[8] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[14]~q ;

assign source_imag[9] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[15]~q ;

assign source_imag[10] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[16]~q ;

assign source_imag[11] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[17]~q ;

assign source_imag[12] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[18]~q ;

assign source_imag[13] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[19]~q ;

assign source_imag[14] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[20]~q ;

assign source_imag[15] = \asj_fft_si_sose_so_b_fft_121_inst|auk_dsp_atlantic_source_1|at_source_data[21]~q ;

endmodule

module fft256_asj_fft_si_sose_so_b_fft_121 (
	at_sink_ready_s,
	at_source_error_0,
	at_source_error_1,
	at_source_sop_s,
	at_source_eop_s,
	at_source_valid_s,
	at_source_data_0,
	at_source_data_1,
	at_source_data_2,
	at_source_data_3,
	at_source_data_4,
	at_source_data_5,
	at_source_data_22,
	at_source_data_23,
	at_source_data_24,
	at_source_data_25,
	at_source_data_26,
	at_source_data_27,
	at_source_data_28,
	at_source_data_29,
	at_source_data_30,
	at_source_data_31,
	at_source_data_32,
	at_source_data_33,
	at_source_data_34,
	at_source_data_35,
	at_source_data_36,
	at_source_data_37,
	at_source_data_6,
	at_source_data_7,
	at_source_data_8,
	at_source_data_9,
	at_source_data_10,
	at_source_data_11,
	at_source_data_12,
	at_source_data_13,
	at_source_data_14,
	at_source_data_15,
	at_source_data_16,
	at_source_data_17,
	at_source_data_18,
	at_source_data_19,
	at_source_data_20,
	at_source_data_21,
	GND_port,
	clk,
	reset_n,
	source_ready,
	sink_valid,
	sink_sop,
	sink_eop,
	sink_error_0,
	sink_error_1,
	inverse,
	sink_real,
	sink_imag)/* synthesis synthesis_greybox=1 */;
output 	at_sink_ready_s;
output 	at_source_error_0;
output 	at_source_error_1;
output 	at_source_sop_s;
output 	at_source_eop_s;
output 	at_source_valid_s;
output 	at_source_data_0;
output 	at_source_data_1;
output 	at_source_data_2;
output 	at_source_data_3;
output 	at_source_data_4;
output 	at_source_data_5;
output 	at_source_data_22;
output 	at_source_data_23;
output 	at_source_data_24;
output 	at_source_data_25;
output 	at_source_data_26;
output 	at_source_data_27;
output 	at_source_data_28;
output 	at_source_data_29;
output 	at_source_data_30;
output 	at_source_data_31;
output 	at_source_data_32;
output 	at_source_data_33;
output 	at_source_data_34;
output 	at_source_data_35;
output 	at_source_data_36;
output 	at_source_data_37;
output 	at_source_data_6;
output 	at_source_data_7;
output 	at_source_data_8;
output 	at_source_data_9;
output 	at_source_data_10;
output 	at_source_data_11;
output 	at_source_data_12;
output 	at_source_data_13;
output 	at_source_data_14;
output 	at_source_data_15;
output 	at_source_data_16;
output 	at_source_data_17;
output 	at_source_data_18;
output 	at_source_data_19;
output 	at_source_data_20;
output 	at_source_data_21;
input 	GND_port;
input 	clk;
input 	reset_n;
input 	source_ready;
input 	sink_valid;
input 	sink_sop;
input 	sink_eop;
input 	sink_error_0;
input 	sink_error_1;
input 	inverse;
input 	[15:0] sink_real;
input 	[15:0] sink_imag;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \master_sink_ena~q ;
wire \data_count_sig[6]~q ;
wire \data_count_sig[4]~q ;
wire \data_count_sig[0]~q ;
wire \data_count_sig[5]~q ;
wire \data_count_sig[1]~q ;
wire \data_count_sig[7]~q ;
wire \data_count_sig[3]~q ;
wire \data_count_sig[2]~q ;
wire \fft_s1_cur.WAIT_FOR_INPUT~q ;
wire \fft_s1_cur.WRITE_INPUT~q ;
wire \data_count_sig[0]~9 ;
wire \data_count_sig[0]~8_combout ;
wire \data_count_sig[1]~11 ;
wire \data_count_sig[1]~10_combout ;
wire \data_count_sig[2]~13 ;
wire \data_count_sig[2]~12_combout ;
wire \data_count_sig[3]~15 ;
wire \data_count_sig[3]~14_combout ;
wire \data_count_sig[4]~17 ;
wire \data_count_sig[4]~16_combout ;
wire \data_count_sig[5]~19 ;
wire \data_count_sig[5]~18_combout ;
wire \data_count_sig[6]~21 ;
wire \data_count_sig[6]~20_combout ;
wire \data_count_sig[7]~25_combout ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[16] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[17] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[18] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[19] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[20] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[21] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[22] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[23] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[24] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[25] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[26] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[27] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[28] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[29] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[30] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ;
wire \gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[31] ;
wire \writer|disable_wr~q ;
wire \fft_s1_cur.FFT_PROCESS_A~q ;
wire \fft_s2_cur.LPP_OUTPUT_RDY~q ;
wire \fft_s2_cur.WAIT_FOR_LPP_INPUT~q ;
wire \fft_s2_cur.START_LPP~q ;
wire \fft_s1_cur.NO_WRITE~q ;
wire \output_count[1]~q ;
wire \output_count[2]~q ;
wire \output_count[3]~q ;
wire \output_count[0]~q ;
wire \output_count[4]~q ;
wire \output_count[5]~q ;
wire \output_count[6]~q ;
wire \output_count[7]~q ;
wire \writer|rdy_for_next_block~q ;
wire \fft_s1_cur.EARLY_DONE~q ;
wire \fft_s1_cur.DONE_WRITING~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~q ;
wire \output_count[0]~9 ;
wire \output_count[0]~8_combout ;
wire \output_count[1]~11 ;
wire \output_count[1]~10_combout ;
wire \output_count[2]~13 ;
wire \output_count[2]~12_combout ;
wire \output_count[3]~15 ;
wire \output_count[3]~14_combout ;
wire \output_count[4]~17 ;
wire \output_count[4]~16_combout ;
wire \output_count[5]~19 ;
wire \output_count[5]~18_combout ;
wire \output_count[6]~21 ;
wire \output_count[6]~20_combout ;
wire \output_count[7]~22_combout ;
wire \del_sop_cnt[0]~q ;
wire \del_sop_cnt[1]~q ;
wire \del_sop_cnt[2]~q ;
wire \del_sop_cnt[4]~q ;
wire \del_sop_cnt[3]~q ;
wire \core_imag_in[0]~q ;
wire \core_real_in[0]~q ;
wire \core_imag_in[1]~q ;
wire \core_real_in[1]~q ;
wire \core_imag_in[2]~q ;
wire \core_real_in[2]~q ;
wire \core_imag_in[3]~q ;
wire \core_real_in[3]~q ;
wire \core_imag_in[4]~q ;
wire \core_real_in[4]~q ;
wire \core_imag_in[5]~q ;
wire \core_real_in[5]~q ;
wire \core_imag_in[6]~q ;
wire \core_real_in[6]~q ;
wire \core_imag_in[7]~q ;
wire \core_real_in[7]~q ;
wire \core_imag_in[8]~q ;
wire \core_real_in[8]~q ;
wire \core_imag_in[9]~q ;
wire \core_real_in[9]~q ;
wire \core_imag_in[10]~q ;
wire \core_real_in[10]~q ;
wire \core_imag_in[11]~q ;
wire \core_real_in[11]~q ;
wire \core_imag_in[12]~q ;
wire \core_real_in[12]~q ;
wire \core_imag_in[13]~q ;
wire \core_real_in[13]~q ;
wire \core_imag_in[14]~q ;
wire \core_real_in[14]~q ;
wire \core_imag_in[15]~q ;
wire \core_real_in[15]~q ;
wire \del_sop_cnt[0]~6 ;
wire \del_sop_cnt[0]~5_combout ;
wire \del_sop_cnt[1]~8 ;
wire \del_sop_cnt[1]~7_combout ;
wire \del_sop_cnt[2]~10 ;
wire \del_sop_cnt[2]~9_combout ;
wire \del_sop_cnt[3]~12 ;
wire \del_sop_cnt[3]~11_combout ;
wire \del_sop_cnt[4]~13_combout ;
wire \k_count_wr[2]~q ;
wire \k_count_wr[0]~q ;
wire \k_count_wr[6]~q ;
wire \k_count_wr[3]~q ;
wire \k_count_wr[1]~q ;
wire \k_count_wr[7]~q ;
wire \k_count_wr[4]~q ;
wire \k_count_wr[5]~q ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \k_count_wr[0]~9 ;
wire \k_count_wr[0]~8_combout ;
wire \k_count_wr[1]~11 ;
wire \k_count_wr[1]~10_combout ;
wire \k_count_wr[2]~13 ;
wire \k_count_wr[2]~12_combout ;
wire \k_count_wr_en~q ;
wire \k_count_wr[3]~15 ;
wire \k_count_wr[3]~14_combout ;
wire \k_count_wr[4]~17 ;
wire \k_count_wr[4]~16_combout ;
wire \k_count_wr[5]~19 ;
wire \k_count_wr[5]~18_combout ;
wire \k_count_wr[6]~21 ;
wire \k_count_wr[6]~20_combout ;
wire \k_count_wr[7]~22_combout ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[22] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[23] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[24] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[25] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[26] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[27] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[28] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[29] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[30] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[31] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \writer|data_rdy_int~q ;
wire \twiddle_data_real[0]~q ;
wire \twiddle_data_real[15]~q ;
wire \twiddle_data_imag[1]~q ;
wire \twiddle_data_imag[2]~q ;
wire \twiddle_data_imag[3]~q ;
wire \twiddle_data_imag[4]~q ;
wire \twiddle_data_imag[5]~q ;
wire \twiddle_data_imag[6]~q ;
wire \twiddle_data_imag[7]~q ;
wire \twiddle_data_imag[8]~q ;
wire \twiddle_data_imag[9]~q ;
wire \twiddle_data_imag[10]~q ;
wire \twiddle_data_imag[11]~q ;
wire \twiddle_data_imag[12]~q ;
wire \twiddle_data_imag[13]~q ;
wire \twiddle_data_imag[14]~q ;
wire \twiddle_data_imag[15]~q ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[0] ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[0] ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[1] ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[1] ;
wire \Add2~1_cout ;
wire \Add2~3 ;
wire \Add2~2_combout ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[2] ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[2] ;
wire \Add2~5 ;
wire \Add2~4_combout ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[3] ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[3] ;
wire \Add2~7 ;
wire \Add2~6_combout ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[4] ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[4] ;
wire \Add2~9 ;
wire \Add2~8_combout ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[5] ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[5] ;
wire \Add2~11 ;
wire \Add2~10_combout ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[6] ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[6] ;
wire \Add2~13 ;
wire \Add2~12_combout ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[7] ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[7] ;
wire \Add2~15 ;
wire \Add2~14_combout ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[8] ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[8] ;
wire \Add2~17 ;
wire \Add2~16_combout ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[9] ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[9] ;
wire \Add2~19 ;
wire \Add2~18_combout ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[10] ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[10] ;
wire \Add2~21 ;
wire \Add2~20_combout ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[11] ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[11] ;
wire \Add2~23 ;
wire \Add2~22_combout ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[12] ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[12] ;
wire \Add2~25 ;
wire \Add2~24_combout ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[13] ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[13] ;
wire \Add2~27 ;
wire \Add2~26_combout ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[14] ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[14] ;
wire \Add2~29 ;
wire \Add2~28_combout ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[15] ;
wire \gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[15] ;
wire \Add2~30_combout ;
wire \twiddle_data_imag[1]~0_combout ;
wire \Add3~1_cout ;
wire \Add3~3 ;
wire \Add3~2_combout ;
wire \twiddle_data_imag[2]~1_combout ;
wire \Add3~5 ;
wire \Add3~4_combout ;
wire \twiddle_data_imag[3]~2_combout ;
wire \Add3~7 ;
wire \Add3~6_combout ;
wire \twiddle_data_imag[4]~3_combout ;
wire \Add3~9 ;
wire \Add3~8_combout ;
wire \twiddle_data_imag[5]~4_combout ;
wire \Add3~11 ;
wire \Add3~10_combout ;
wire \twiddle_data_imag[6]~5_combout ;
wire \Add3~13 ;
wire \Add3~12_combout ;
wire \twiddle_data_imag[7]~6_combout ;
wire \Add3~15 ;
wire \Add3~14_combout ;
wire \twiddle_data_imag[8]~7_combout ;
wire \Add3~17 ;
wire \Add3~16_combout ;
wire \twiddle_data_imag[9]~8_combout ;
wire \Add3~19 ;
wire \Add3~18_combout ;
wire \twiddle_data_imag[10]~9_combout ;
wire \Add3~21 ;
wire \Add3~20_combout ;
wire \twiddle_data_imag[11]~10_combout ;
wire \Add3~23 ;
wire \Add3~22_combout ;
wire \twiddle_data_imag[12]~11_combout ;
wire \Add3~25 ;
wire \Add3~24_combout ;
wire \twiddle_data_imag[13]~12_combout ;
wire \Add3~27 ;
wire \Add3~26_combout ;
wire \twiddle_data_imag[14]~13_combout ;
wire \Add3~29 ;
wire \Add3~28_combout ;
wire \Add3~30_combout ;
wire \gen_se:gen_new:twid_factors|twad_tempo[0]~q ;
wire \gen_se:gen_new:twid_factors|twad_tempe[1]~q ;
wire \gen_se:gen_new:twid_factors|twad_tempe[2]~q ;
wire \gen_se:gen_new:twid_factors|twad_tempe[3]~q ;
wire \gen_se:gen_new:twid_factors|twad_tempe[4]~q ;
wire \gen_se:gen_new:twid_factors|twad_tempe[5]~q ;
wire \gen_se:gen_new:twid_factors|twad_tempo[1]~q ;
wire \gen_se:gen_new:twid_factors|twad_tempo[2]~q ;
wire \gen_se:gen_new:twid_factors|twad_tempo[3]~q ;
wire \gen_se:gen_new:twid_factors|twad_tempo[4]~q ;
wire \gen_se:gen_new:twid_factors|twad_tempo[5]~q ;
wire \k_count_tw[0]~q ;
wire \k_count_tw[2]~q ;
wire \k_count_tw[1]~q ;
wire \k_count_tw[3]~q ;
wire \k_count_tw[5]~q ;
wire \k_count_tw[4]~q ;
wire \k_count_tw[7]~q ;
wire \k_count_tw[6]~q ;
wire \k_count_tw[0]~9 ;
wire \k_count_tw[0]~8_combout ;
wire \k_count_tw_en~q ;
wire \k_count_tw[1]~11 ;
wire \k_count_tw[1]~10_combout ;
wire \k_count_tw[2]~13 ;
wire \k_count_tw[2]~12_combout ;
wire \k_count_tw[3]~15 ;
wire \k_count_tw[3]~14_combout ;
wire \k_count_tw[4]~17 ;
wire \k_count_tw[4]~16_combout ;
wire \k_count_tw[5]~19 ;
wire \k_count_tw[5]~18_combout ;
wire \k_count_tw[6]~21 ;
wire \k_count_tw[6]~20_combout ;
wire \k_count_tw[7]~22_combout ;
wire \auk_dsp_interface_controller_1|source_packet_error[0]~q ;
wire \auk_dsp_interface_controller_1|source_packet_error[1]~q ;
wire \auk_dsp_interface_controller_1|source_stall_reg~q ;
wire \auk_dsp_interface_controller_1|sink_stall_reg~q ;
wire \auk_dsp_interface_controller_1|sink_ready_ctrl~0_combout ;
wire \auk_dsp_atlantic_sink_1|sink_start~q ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|empty_dff~q ;
wire \auk_dsp_atlantic_sink_1|sink_stall~combout ;
wire \auk_dsp_atlantic_sink_1|packet_error_s[0]~q ;
wire \auk_dsp_atlantic_sink_1|packet_error_s[1]~q ;
wire \master_source_ena~q ;
wire \sink_ready_ctrl_d~q ;
wire \auk_dsp_atlantic_sink_1|send_sop_s~q ;
wire \sop~q ;
wire \source_valid_ctrl_sop~0_combout ;
wire \source_valid_ctrl_sop~1_combout ;
wire \auk_dsp_interface_controller_1|stall_reg~q ;
wire \auk_dsp_atlantic_source_1|source_stall_int_d~q ;
wire \exponent_out[0]~q ;
wire \exponent_out[1]~q ;
wire \exponent_out[2]~q ;
wire \exponent_out[3]~q ;
wire \exponent_out[4]~q ;
wire \exponent_out[5]~q ;
wire \fft_real_out[0]~q ;
wire \fft_real_out[1]~q ;
wire \fft_real_out[2]~q ;
wire \fft_real_out[3]~q ;
wire \fft_real_out[4]~q ;
wire \fft_real_out[5]~q ;
wire \fft_real_out[6]~q ;
wire \fft_real_out[7]~q ;
wire \fft_real_out[8]~q ;
wire \fft_real_out[9]~q ;
wire \fft_real_out[10]~q ;
wire \fft_real_out[11]~q ;
wire \fft_real_out[12]~q ;
wire \fft_real_out[13]~q ;
wire \fft_real_out[14]~q ;
wire \fft_real_out[15]~q ;
wire \fft_imag_out[0]~q ;
wire \fft_imag_out[1]~q ;
wire \fft_imag_out[2]~q ;
wire \fft_imag_out[3]~q ;
wire \fft_imag_out[4]~q ;
wire \fft_imag_out[5]~q ;
wire \fft_imag_out[6]~q ;
wire \fft_imag_out[7]~q ;
wire \fft_imag_out[8]~q ;
wire \fft_imag_out[9]~q ;
wire \fft_imag_out[10]~q ;
wire \fft_imag_out[11]~q ;
wire \fft_imag_out[12]~q ;
wire \fft_imag_out[13]~q ;
wire \fft_imag_out[14]~q ;
wire \fft_imag_out[15]~q ;
wire \fft_s1_cur.IDLE~q ;
wire \WideOr3~0_combout ;
wire \global_clock_enable~0_combout ;
wire \auk_dsp_atlantic_source_1|Mux0~1_combout ;
wire \val_out~q ;
wire \master_source_ena~0_combout ;
wire \auk_dsp_atlantic_sink_1|send_eop_s~q ;
wire \sop~0_combout ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \master_source_sop~q ;
wire \data_count_sig[1]~22_combout ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \data_count_sig[1]~23_combout ;
wire \data_count_sig[6]~24_combout ;
wire \gen_se:bfpc|blk_exp[0]~q ;
wire \exponent_out~0_combout ;
wire \gen_se:bfpc|blk_exp[1]~q ;
wire \exponent_out~1_combout ;
wire \gen_se:bfpc|blk_exp[2]~q ;
wire \exponent_out~2_combout ;
wire \gen_se:bfpc|blk_exp[3]~q ;
wire \exponent_out~3_combout ;
wire \gen_se:bfpc|blk_exp[4]~q ;
wire \exponent_out~4_combout ;
wire \gen_se:bfpc|blk_exp[5]~q ;
wire \exponent_out~5_combout ;
wire \fft_dirn~q ;
wire \fft_real_out~0_combout ;
wire \fft_real_out~1_combout ;
wire \fft_real_out~2_combout ;
wire \fft_real_out~3_combout ;
wire \fft_real_out~4_combout ;
wire \fft_real_out~5_combout ;
wire \fft_real_out~6_combout ;
wire \fft_real_out~7_combout ;
wire \fft_real_out~8_combout ;
wire \fft_real_out~9_combout ;
wire \fft_real_out~10_combout ;
wire \fft_real_out~11_combout ;
wire \fft_real_out~12_combout ;
wire \fft_real_out~13_combout ;
wire \fft_real_out~14_combout ;
wire \fft_real_out~15_combout ;
wire \fft_imag_out~0_combout ;
wire \fft_imag_out~1_combout ;
wire \fft_imag_out~2_combout ;
wire \fft_imag_out~3_combout ;
wire \fft_imag_out~4_combout ;
wire \fft_imag_out~5_combout ;
wire \fft_imag_out~6_combout ;
wire \fft_imag_out~7_combout ;
wire \fft_imag_out~8_combout ;
wire \fft_imag_out~9_combout ;
wire \fft_imag_out~10_combout ;
wire \fft_imag_out~11_combout ;
wire \fft_imag_out~12_combout ;
wire \fft_imag_out~13_combout ;
wire \fft_imag_out~14_combout ;
wire \fft_imag_out~15_combout ;
wire \Selector5~0_combout ;
wire \Selector6~0_combout ;
wire \eop_out~q ;
wire \fft_s1_cur.IDLE~0_combout ;
wire \fft_s2_cur.IDLE~q ;
wire \fft_s2_cur.FIRST_LPP~q ;
wire \fft_s2_cur.LPP_DONE~q ;
wire \val_out~0_combout ;
wire \val_out~1_combout ;
wire \sop_out~q ;
wire \master_source_sop~0_combout ;
wire \sop_d~q ;
wire \wren_a~q ;
wire \ccc|a_ram_data_in_bus[0]~q ;
wire \ccc|wraddress_a_bus[0]~q ;
wire \ccc|wraddress_a_bus[1]~q ;
wire \ccc|wraddress_a_bus[2]~q ;
wire \ccc|wraddress_a_bus[3]~q ;
wire \ccc|wraddress_a_bus[4]~q ;
wire \ccc|wraddress_a_bus[5]~q ;
wire \ccc|wraddress_a_bus[6]~q ;
wire \ccc|wraddress_a_bus[7]~q ;
wire \ccc|rdaddress_a_bus[0]~q ;
wire \ccc|rdaddress_a_bus[1]~q ;
wire \ccc|rdaddress_a_bus[2]~q ;
wire \ccc|rdaddress_a_bus[3]~q ;
wire \ccc|rdaddress_a_bus[4]~q ;
wire \ccc|rdaddress_a_bus[5]~q ;
wire \ccc|rdaddress_a_bus[6]~q ;
wire \ccc|rdaddress_a_bus[7]~q ;
wire \ccc|a_ram_data_in_bus[16]~q ;
wire \fft_dirn~0_combout ;
wire \ccc|a_ram_data_in_bus[1]~q ;
wire \ccc|a_ram_data_in_bus[17]~q ;
wire \ccc|a_ram_data_in_bus[2]~q ;
wire \ccc|a_ram_data_in_bus[18]~q ;
wire \ccc|a_ram_data_in_bus[3]~q ;
wire \ccc|a_ram_data_in_bus[19]~q ;
wire \ccc|a_ram_data_in_bus[4]~q ;
wire \ccc|a_ram_data_in_bus[20]~q ;
wire \ccc|a_ram_data_in_bus[5]~q ;
wire \ccc|a_ram_data_in_bus[21]~q ;
wire \ccc|a_ram_data_in_bus[6]~q ;
wire \ccc|a_ram_data_in_bus[22]~q ;
wire \ccc|a_ram_data_in_bus[7]~q ;
wire \ccc|a_ram_data_in_bus[23]~q ;
wire \ccc|a_ram_data_in_bus[8]~q ;
wire \ccc|a_ram_data_in_bus[24]~q ;
wire \ccc|a_ram_data_in_bus[9]~q ;
wire \ccc|a_ram_data_in_bus[25]~q ;
wire \ccc|a_ram_data_in_bus[10]~q ;
wire \ccc|a_ram_data_in_bus[26]~q ;
wire \ccc|a_ram_data_in_bus[11]~q ;
wire \ccc|a_ram_data_in_bus[27]~q ;
wire \ccc|a_ram_data_in_bus[12]~q ;
wire \ccc|a_ram_data_in_bus[28]~q ;
wire \ccc|a_ram_data_in_bus[13]~q ;
wire \ccc|a_ram_data_in_bus[29]~q ;
wire \ccc|a_ram_data_in_bus[14]~q ;
wire \ccc|a_ram_data_in_bus[30]~q ;
wire \ccc|a_ram_data_in_bus[15]~q ;
wire \ccc|a_ram_data_in_bus[31]~q ;
wire \data_rdy_vec[24]~q ;
wire \Selector10~0_combout ;
wire \fft_s2_cur~8_combout ;
wire \Equal9~0_combout ;
wire \Equal9~1_combout ;
wire \Selector2~0_combout ;
wire \fft_s2_cur~9_combout ;
wire \ctrl|blk_done~q ;
wire \Selector0~0_combout ;
wire \Selector1~0_combout ;
wire \gen_se:bfpdft|bfp_detect|slb_i[0]~q ;
wire \gen_se:bfpdft|bfp_detect|Mux2~0_combout ;
wire \gen_se:bfpdft|bfp_detect|lut_out[0]~0_combout ;
wire \gen_se:bfpc|gen_so_crtl:gen_se_so:delay_next_pass_2|tdl_arr[0]~q ;
wire \sop_de~q ;
wire \gen_se:bfpdft|bfp_detect|Mux1~0_combout ;
wire \gen_se:bfpdft|bfp_detect|lut_out[1]~1_combout ;
wire \gen_se:bfpdft|bfp_detect|lut_out[2]~2_combout ;
wire \gen_se:bfpdft|bfp_detect|lut_out[2]~3_combout ;
wire \writer|gen_soe:delay_swd|tdl_arr[0]~q ;
wire \wren_a~2_combout ;
wire \data_rdy_vec[21]~q ;
wire \wren_a~3_combout ;
wire \wren_a~4_combout ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[0]~q ;
wire \writer|data_in_i[0]~q ;
wire \sel_ram_in~q ;
wire \wraddress_a_bus_ctrl_i[0]~q ;
wire \writer|wr_address_i_int[0]~q ;
wire \wraddress_a_bus_ctrl_i[1]~q ;
wire \writer|wr_address_i_int[1]~q ;
wire \wraddress_a_bus_ctrl_i[2]~q ;
wire \writer|wr_address_i_int[2]~q ;
wire \wraddress_a_bus_ctrl_i[3]~q ;
wire \writer|wr_address_i_int[3]~q ;
wire \wraddress_a_bus_ctrl_i[4]~q ;
wire \writer|wr_address_i_int[4]~q ;
wire \wraddress_a_bus_ctrl_i[5]~q ;
wire \writer|wr_address_i_int[5]~q ;
wire \wraddress_a_bus_ctrl_i[6]~q ;
wire \writer|wr_address_i_int[6]~q ;
wire \wraddress_a_bus_ctrl_i[7]~q ;
wire \writer|wr_address_i_int[7]~q ;
wire \rd_adgen|rd_addr_a[0]~q ;
wire \rd_adgen|rd_addr_a[1]~q ;
wire \rd_adgen|rd_addr_a[2]~q ;
wire \rd_adgen|rd_addr_a[3]~q ;
wire \rd_adgen|rd_addr_a[4]~q ;
wire \rd_adgen|rd_addr_a[5]~q ;
wire \rd_adgen|rd_addr_a[6]~q ;
wire \rd_adgen|rd_addr_a[7]~q ;
wire \writer|data_in_r[0]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[1]~q ;
wire \writer|data_in_i[1]~q ;
wire \writer|data_in_r[1]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[2]~q ;
wire \writer|data_in_i[2]~q ;
wire \writer|data_in_r[2]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[3]~q ;
wire \writer|data_in_i[3]~q ;
wire \writer|data_in_r[3]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[4]~q ;
wire \writer|data_in_i[4]~q ;
wire \writer|data_in_r[4]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[5]~q ;
wire \writer|data_in_i[5]~q ;
wire \writer|data_in_r[5]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[6]~q ;
wire \writer|data_in_i[6]~q ;
wire \writer|data_in_r[6]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[7]~q ;
wire \writer|data_in_i[7]~q ;
wire \writer|data_in_r[7]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[8]~q ;
wire \writer|data_in_i[8]~q ;
wire \writer|data_in_r[8]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[9]~q ;
wire \writer|data_in_i[9]~q ;
wire \writer|data_in_r[9]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[10]~q ;
wire \writer|data_in_i[10]~q ;
wire \writer|data_in_r[10]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[11]~q ;
wire \writer|data_in_i[11]~q ;
wire \writer|data_in_r[11]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[12]~q ;
wire \writer|data_in_i[12]~q ;
wire \writer|data_in_r[12]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[13]~q ;
wire \writer|data_in_i[13]~q ;
wire \writer|data_in_r[13]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[14]~q ;
wire \writer|data_in_i[14]~q ;
wire \writer|data_in_r[14]~q ;
wire \gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[15]~q ;
wire \writer|data_in_i[15]~q ;
wire \writer|data_in_r[15]~q ;
wire \writer|counter_i~0_combout ;
wire \data_rdy_vec[23]~q ;
wire \data_rdy_vec~0_combout ;
wire \no_del_input_blk:delay_next_block|tdl_arr[0]~q ;
wire \Selector9~0_combout ;
wire \output_sample_counter~0_combout ;
wire \ctrl|p[2]~q ;
wire \ctrl|p[0]~q ;
wire \ctrl|p[1]~q ;
wire \rd_adgen|rd_addr_a[0]~0_combout ;
wire \delay_swd|tdl_arr[9]~q ;
wire \sop_de~0_combout ;
wire \sop_de~1_combout ;
wire \Selector7~0_combout ;
wire \Selector8~0_combout ;
wire \data_rdy_vec[20]~q ;
wire \data_rdy_vec~1_combout ;
wire \sel_ram_in~0_combout ;
wire \gen_wraddr_se:wr_adgen|rd_addr_a[0]~q ;
wire \gen_wraddr_se:wr_adgen|rd_addr_a[1]~q ;
wire \gen_wraddr_se:wr_adgen|rd_addr_a[2]~q ;
wire \gen_wraddr_se:wr_adgen|rd_addr_a[3]~q ;
wire \gen_wraddr_se:wr_adgen|rd_addr_a[4]~q ;
wire \gen_wraddr_se:wr_adgen|rd_addr_a[5]~q ;
wire \gen_wraddr_se:wr_adgen|rd_addr_a[6]~q ;
wire \gen_wraddr_se:wr_adgen|rd_addr_a[7]~q ;
wire \ctrl|k_count[2]~q ;
wire \ctrl|k_count[0]~q ;
wire \ctrl|k_count[6]~q ;
wire \ctrl|k_count[3]~q ;
wire \ctrl|k_count[1]~q ;
wire \ctrl|k_count[7]~q ;
wire \ctrl|k_count[4]~q ;
wire \ctrl|k_count[5]~q ;
wire \data_rdy_vec[22]~q ;
wire \data_rdy_vec~2_combout ;
wire \data_rdy_vec[4]~q ;
wire \ctrl|next_pass_i~q ;
wire \data_rdy_vec[19]~q ;
wire \data_rdy_vec~3_combout ;
wire \data_real_in_reg[0]~q ;
wire \data_imag_in_reg[0]~q ;
wire \core_imag_in~0_combout ;
wire \p_tdl[18][0]~q ;
wire \p_tdl[18][1]~q ;
wire \p_tdl[18][2]~q ;
wire \core_real_in~0_combout ;
wire \data_real_in_reg[1]~q ;
wire \data_imag_in_reg[1]~q ;
wire \core_imag_in~1_combout ;
wire \core_real_in~1_combout ;
wire \data_real_in_reg[2]~q ;
wire \data_imag_in_reg[2]~q ;
wire \core_imag_in~2_combout ;
wire \core_real_in~2_combout ;
wire \data_real_in_reg[3]~q ;
wire \data_imag_in_reg[3]~q ;
wire \core_imag_in~3_combout ;
wire \core_real_in~3_combout ;
wire \data_real_in_reg[4]~q ;
wire \data_imag_in_reg[4]~q ;
wire \core_imag_in~4_combout ;
wire \core_real_in~4_combout ;
wire \data_real_in_reg[5]~q ;
wire \data_imag_in_reg[5]~q ;
wire \core_imag_in~5_combout ;
wire \core_real_in~5_combout ;
wire \data_real_in_reg[6]~q ;
wire \data_imag_in_reg[6]~q ;
wire \core_imag_in~6_combout ;
wire \core_real_in~6_combout ;
wire \data_real_in_reg[7]~q ;
wire \data_imag_in_reg[7]~q ;
wire \core_imag_in~7_combout ;
wire \core_real_in~7_combout ;
wire \data_real_in_reg[8]~q ;
wire \data_imag_in_reg[8]~q ;
wire \core_imag_in~8_combout ;
wire \core_real_in~8_combout ;
wire \data_real_in_reg[9]~q ;
wire \data_imag_in_reg[9]~q ;
wire \core_imag_in~9_combout ;
wire \core_real_in~9_combout ;
wire \data_real_in_reg[10]~q ;
wire \data_imag_in_reg[10]~q ;
wire \core_imag_in~10_combout ;
wire \core_real_in~10_combout ;
wire \data_real_in_reg[11]~q ;
wire \data_imag_in_reg[11]~q ;
wire \core_imag_in~11_combout ;
wire \core_real_in~11_combout ;
wire \data_real_in_reg[12]~q ;
wire \data_imag_in_reg[12]~q ;
wire \core_imag_in~12_combout ;
wire \core_real_in~12_combout ;
wire \data_real_in_reg[13]~q ;
wire \data_imag_in_reg[13]~q ;
wire \core_imag_in~13_combout ;
wire \core_real_in~13_combout ;
wire \data_real_in_reg[14]~q ;
wire \data_imag_in_reg[14]~q ;
wire \core_imag_in~14_combout ;
wire \core_real_in~14_combout ;
wire \data_real_in_reg[15]~q ;
wire \data_imag_in_reg[15]~q ;
wire \core_imag_in~15_combout ;
wire \core_real_in~15_combout ;
wire \data_rdy_vec~4_combout ;
wire \data_rdy_vec[3]~q ;
wire \data_rdy_vec~5_combout ;
wire \data_rdy_vec[18]~q ;
wire \data_rdy_vec~6_combout ;
wire \data_real_in_reg~0_combout ;
wire \data_imag_in_reg~0_combout ;
wire \p_tdl[17][0]~q ;
wire \p_tdl~0_combout ;
wire \p_tdl[17][1]~q ;
wire \p_tdl~1_combout ;
wire \p_tdl[17][2]~q ;
wire \p_tdl~2_combout ;
wire \data_real_in_reg~1_combout ;
wire \data_imag_in_reg~1_combout ;
wire \data_real_in_reg~2_combout ;
wire \data_imag_in_reg~2_combout ;
wire \data_real_in_reg~3_combout ;
wire \data_imag_in_reg~3_combout ;
wire \data_real_in_reg~4_combout ;
wire \data_imag_in_reg~4_combout ;
wire \data_real_in_reg~5_combout ;
wire \data_imag_in_reg~5_combout ;
wire \data_real_in_reg~6_combout ;
wire \data_imag_in_reg~6_combout ;
wire \data_real_in_reg~7_combout ;
wire \data_imag_in_reg~7_combout ;
wire \data_real_in_reg~8_combout ;
wire \data_imag_in_reg~8_combout ;
wire \data_real_in_reg~9_combout ;
wire \data_imag_in_reg~9_combout ;
wire \data_real_in_reg~10_combout ;
wire \data_imag_in_reg~10_combout ;
wire \data_real_in_reg~11_combout ;
wire \data_imag_in_reg~11_combout ;
wire \data_real_in_reg~12_combout ;
wire \data_imag_in_reg~12_combout ;
wire \data_real_in_reg~13_combout ;
wire \data_imag_in_reg~13_combout ;
wire \data_real_in_reg~14_combout ;
wire \data_imag_in_reg~14_combout ;
wire \data_real_in_reg~15_combout ;
wire \data_imag_in_reg~15_combout ;
wire \data_rdy_vec[2]~q ;
wire \data_rdy_vec~7_combout ;
wire \data_rdy_vec[17]~q ;
wire \data_rdy_vec~8_combout ;
wire \Equal5~0_combout ;
wire \Equal5~1_combout ;
wire \k_count_wr_en~0_combout ;
wire \Equal4~0_combout ;
wire \Equal4~1_combout ;
wire \k_count_wr_en~1_combout ;
wire \p_tdl[16][0]~q ;
wire \p_tdl~3_combout ;
wire \p_tdl[16][1]~q ;
wire \p_tdl~4_combout ;
wire \p_tdl[16][2]~q ;
wire \p_tdl~5_combout ;
wire \data_rdy_vec[1]~q ;
wire \data_rdy_vec~9_combout ;
wire \data_rdy_vec[16]~q ;
wire \data_rdy_vec~10_combout ;
wire \p_tdl[15][0]~q ;
wire \p_tdl~6_combout ;
wire \p_tdl[15][1]~q ;
wire \p_tdl~7_combout ;
wire \p_tdl[15][2]~q ;
wire \p_tdl~8_combout ;
wire \data_rdy_vec[0]~q ;
wire \data_rdy_vec~11_combout ;
wire \data_rdy_vec[15]~q ;
wire \data_rdy_vec~12_combout ;
wire \p_tdl[14][0]~q ;
wire \p_tdl~9_combout ;
wire \p_tdl[14][1]~q ;
wire \p_tdl~10_combout ;
wire \p_tdl[14][2]~q ;
wire \p_tdl~11_combout ;
wire \data_rdy_vec~13_combout ;
wire \data_rdy_vec[14]~q ;
wire \data_rdy_vec~14_combout ;
wire \twiddle_data_real[1]~q ;
wire \twiddle_data_real[2]~q ;
wire \twiddle_data_real[3]~q ;
wire \twiddle_data_real[4]~q ;
wire \twiddle_data_real[5]~q ;
wire \twiddle_data_real[6]~q ;
wire \twiddle_data_real[7]~q ;
wire \twiddle_data_real[8]~q ;
wire \twiddle_data_real[9]~q ;
wire \twiddle_data_real[10]~q ;
wire \twiddle_data_real[11]~q ;
wire \twiddle_data_real[12]~q ;
wire \twiddle_data_real[13]~q ;
wire \twiddle_data_real[14]~q ;
wire \twiddle_data_imag[0]~q ;
wire \p_tdl[13][0]~q ;
wire \p_tdl~12_combout ;
wire \p_tdl[13][1]~q ;
wire \p_tdl~13_combout ;
wire \p_tdl[13][2]~q ;
wire \p_tdl~14_combout ;
wire \data_rdy_vec[13]~q ;
wire \data_rdy_vec~15_combout ;
wire \quad_del_1[2]~q ;
wire \quad_del_1[0]~q ;
wire \quad_del_1[1]~q ;
wire \Mux15~0_combout ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \twiddle_data_imag~14_combout ;
wire \twiddle_data_imag[14]~15_combout ;
wire \twiddle_data_imag~16_combout ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \p_tdl[12][0]~q ;
wire \p_tdl~15_combout ;
wire \p_tdl[12][1]~q ;
wire \p_tdl~16_combout ;
wire \p_tdl[12][2]~q ;
wire \p_tdl~17_combout ;
wire \data_rdy_vec[12]~q ;
wire \data_rdy_vec~16_combout ;
wire \quad_del_0[2]~q ;
wire \quad_del_1~0_combout ;
wire \quad_del_0[0]~q ;
wire \quad_del_1~1_combout ;
wire \quad_del_0[1]~q ;
wire \quad_del_1~2_combout ;
wire \p_tdl[11][0]~q ;
wire \p_tdl~18_combout ;
wire \p_tdl[11][1]~q ;
wire \p_tdl~19_combout ;
wire \p_tdl[11][2]~q ;
wire \p_tdl~20_combout ;
wire \data_rdy_vec[11]~q ;
wire \data_rdy_vec~17_combout ;
wire \gen_se:gen_new:twid_factors|quad_reg[2]~q ;
wire \quad_del_0~0_combout ;
wire \gen_se:gen_new:twid_factors|quad_reg[0]~q ;
wire \quad_del_0~1_combout ;
wire \gen_se:gen_new:twid_factors|quad_reg[1]~q ;
wire \quad_del_0~2_combout ;
wire \p_tdl[10][0]~q ;
wire \p_tdl~21_combout ;
wire \p_tdl[10][1]~q ;
wire \p_tdl~22_combout ;
wire \p_tdl[10][2]~q ;
wire \p_tdl~23_combout ;
wire \data_rdy_vec[27]~q ;
wire \next_pass~combout ;
wire \data_rdy_vec[10]~q ;
wire \data_rdy_vec~18_combout ;
wire \p_tdl[9][0]~q ;
wire \p_tdl~24_combout ;
wire \p_tdl[9][1]~q ;
wire \p_tdl~25_combout ;
wire \p_tdl[9][2]~q ;
wire \p_tdl~26_combout ;
wire \data_rdy_vec[26]~q ;
wire \data_rdy_vec~19_combout ;
wire \data_rdy_vec[9]~q ;
wire \data_rdy_vec~20_combout ;
wire \gen_se:gen_new:twid_factors|data_addr_held_by1~0_combout ;
wire \gen_se:gen_new:twid_factors|data_addr_held_by2~0_combout ;
wire \p_tdl[8][0]~q ;
wire \p_tdl~27_combout ;
wire \p_tdl[8][1]~q ;
wire \p_tdl~28_combout ;
wire \p_tdl[8][2]~q ;
wire \p_tdl~29_combout ;
wire \data_rdy_vec[25]~q ;
wire \data_rdy_vec~21_combout ;
wire \data_rdy_vec[8]~q ;
wire \data_rdy_vec~22_combout ;
wire \ccc|ram_data_out[0]~q ;
wire \ccc|ram_data_out[2]~q ;
wire \gen_se:bfpc|slb_last[1]~q ;
wire \ccc|ram_data_out[1]~q ;
wire \gen_se:bfpc|slb_last[0]~q ;
wire \gen_se:bfpc|slb_last[2]~q ;
wire \ccc|ram_data_out[14]~q ;
wire \ccc|ram_data_out[12]~q ;
wire \ccc|ram_data_out[13]~q ;
wire \ccc|ram_data_out[15]~q ;
wire \ccc|ram_data_out[11]~q ;
wire \ccc|ram_data_out[10]~q ;
wire \ccc|ram_data_out[9]~q ;
wire \ccc|ram_data_out[8]~q ;
wire \ccc|ram_data_out[7]~q ;
wire \ccc|ram_data_out[6]~q ;
wire \ccc|ram_data_out[5]~q ;
wire \ccc|ram_data_out[4]~q ;
wire \ccc|ram_data_out[3]~q ;
wire \ccc|ram_data_out[16]~q ;
wire \ccc|ram_data_out[18]~q ;
wire \ccc|ram_data_out[17]~q ;
wire \ccc|ram_data_out[28]~q ;
wire \ccc|ram_data_out[29]~q ;
wire \ccc|ram_data_out[30]~q ;
wire \ccc|ram_data_out[31]~q ;
wire \ccc|ram_data_out[27]~q ;
wire \ccc|ram_data_out[26]~q ;
wire \ccc|ram_data_out[25]~q ;
wire \ccc|ram_data_out[24]~q ;
wire \ccc|ram_data_out[23]~q ;
wire \ccc|ram_data_out[22]~q ;
wire \ccc|ram_data_out[21]~q ;
wire \ccc|ram_data_out[20]~q ;
wire \ccc|ram_data_out[19]~q ;
wire \p_tdl[7][0]~q ;
wire \p_tdl~30_combout ;
wire \p_tdl[7][1]~q ;
wire \p_tdl~31_combout ;
wire \p_tdl[7][2]~q ;
wire \p_tdl~32_combout ;
wire \data_rdy_vec~23_combout ;
wire \data_rdy_vec[7]~q ;
wire \data_rdy_vec~24_combout ;
wire \Equal7~0_combout ;
wire \k_count_tw_en~0_combout ;
wire \Equal6~0_combout ;
wire \k_count_tw_en~1_combout ;
wire \p_tdl[6][0]~q ;
wire \p_tdl~33_combout ;
wire \p_tdl[6][1]~q ;
wire \p_tdl~34_combout ;
wire \p_tdl[6][2]~q ;
wire \p_tdl~35_combout ;
wire \data_rdy_vec[6]~q ;
wire \data_rdy_vec~25_combout ;
wire \p_tdl[5][0]~q ;
wire \p_tdl~36_combout ;
wire \p_tdl[5][1]~q ;
wire \p_tdl~37_combout ;
wire \p_tdl[5][2]~q ;
wire \p_tdl~38_combout ;
wire \data_rdy_vec[5]~q ;
wire \data_rdy_vec~26_combout ;
wire \p_tdl[4][0]~q ;
wire \p_tdl~39_combout ;
wire \p_tdl[4][1]~q ;
wire \p_tdl~40_combout ;
wire \p_tdl[4][2]~q ;
wire \p_tdl~41_combout ;
wire \data_rdy_vec~27_combout ;
wire \p_tdl[3][0]~q ;
wire \p_tdl~42_combout ;
wire \p_tdl[3][1]~q ;
wire \p_tdl~43_combout ;
wire \p_tdl[3][2]~q ;
wire \p_tdl~44_combout ;
wire \p_tdl[2][0]~q ;
wire \p_tdl~45_combout ;
wire \p_tdl[2][1]~q ;
wire \p_tdl~46_combout ;
wire \p_tdl[2][2]~q ;
wire \p_tdl~47_combout ;
wire \p_tdl[1][0]~q ;
wire \p_tdl~48_combout ;
wire \p_tdl[1][1]~q ;
wire \p_tdl~49_combout ;
wire \p_tdl[1][2]~q ;
wire \p_tdl~50_combout ;
wire \p_tdl[0][0]~q ;
wire \p_tdl~51_combout ;
wire \p_tdl[0][1]~q ;
wire \p_tdl~52_combout ;
wire \p_tdl[0][2]~q ;
wire \p_tdl~53_combout ;
wire \p_tdl~54_combout ;
wire \p_tdl~55_combout ;
wire \p_tdl~56_combout ;
wire \twiddle_data_real~5_combout ;
wire \twiddle_data_real~6_combout ;
wire \twiddle_data_real~100_combout ;
wire \twiddle_data_real~12_combout ;
wire \twiddle_data_real~13_combout ;
wire \twiddle_data_real~101_combout ;
wire \twiddle_data_real~19_combout ;
wire \twiddle_data_real~20_combout ;
wire \twiddle_data_real~102_combout ;
wire \twiddle_data_real~26_combout ;
wire \twiddle_data_real~27_combout ;
wire \twiddle_data_real~103_combout ;
wire \twiddle_data_real~33_combout ;
wire \twiddle_data_real~34_combout ;
wire \twiddle_data_real~104_combout ;
wire \twiddle_data_real~40_combout ;
wire \twiddle_data_real~41_combout ;
wire \twiddle_data_real~105_combout ;
wire \twiddle_data_real~47_combout ;
wire \twiddle_data_real~48_combout ;
wire \twiddle_data_real~106_combout ;
wire \twiddle_data_real~54_combout ;
wire \twiddle_data_real~55_combout ;
wire \twiddle_data_real~107_combout ;
wire \twiddle_data_real~61_combout ;
wire \twiddle_data_real~62_combout ;
wire \twiddle_data_real~108_combout ;
wire \twiddle_data_real~68_combout ;
wire \twiddle_data_real~69_combout ;
wire \twiddle_data_real~109_combout ;
wire \twiddle_data_real~75_combout ;
wire \twiddle_data_real~76_combout ;
wire \twiddle_data_real~110_combout ;
wire \twiddle_data_real~82_combout ;
wire \twiddle_data_real~83_combout ;
wire \twiddle_data_real~111_combout ;
wire \twiddle_data_real~89_combout ;
wire \twiddle_data_real~90_combout ;
wire \twiddle_data_real~112_combout ;
wire \twiddle_data_real~96_combout ;
wire \twiddle_data_real~97_combout ;
wire \twiddle_data_real~113_combout ;


fft256_auk_dspip_avalon_streaming_sink_fft_121 auk_dsp_atlantic_sink_1(
	.master_sink_ena(\master_sink_ena~q ),
	.q_b_16(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.q_b_0(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_17(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.q_b_1(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_18(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.q_b_2(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_19(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.q_b_3(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_20(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.q_b_4(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_21(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.q_b_5(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_22(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.q_b_6(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_23(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[23] ),
	.q_b_7(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_24(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[24] ),
	.q_b_8(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.q_b_25(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[25] ),
	.q_b_9(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.q_b_26(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[26] ),
	.q_b_10(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.q_b_27(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[27] ),
	.q_b_11(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_28(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[28] ),
	.q_b_12(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_29(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[29] ),
	.q_b_13(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.q_b_30(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[30] ),
	.q_b_14(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_31(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[31] ),
	.q_b_15(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.at_sink_ready_s1(at_sink_ready_s),
	.source_stall_reg(\auk_dsp_interface_controller_1|source_stall_reg~q ),
	.sink_stall_reg(\auk_dsp_interface_controller_1|sink_stall_reg~q ),
	.sink_ready_ctrl(\auk_dsp_interface_controller_1|sink_ready_ctrl~0_combout ),
	.sink_start1(\auk_dsp_atlantic_sink_1|sink_start~q ),
	.empty_dff(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|empty_dff~q ),
	.sink_stall1(\auk_dsp_atlantic_sink_1|sink_stall~combout ),
	.packet_error_s_0(\auk_dsp_atlantic_sink_1|packet_error_s[0]~q ),
	.packet_error_s_1(\auk_dsp_atlantic_sink_1|packet_error_s[1]~q ),
	.send_sop_s1(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.send_eop_s1(\auk_dsp_atlantic_sink_1|send_eop_s~q ),
	.clk(clk),
	.reset_n(reset_n),
	.sink_valid(sink_valid),
	.sink_sop(sink_sop),
	.sink_eop(sink_eop),
	.sink_error_0(sink_error_0),
	.sink_error_1(sink_error_1),
	.at_sink_data({sink_real[15],sink_real[14],sink_real[13],sink_real[12],sink_real[11],sink_real[10],sink_real[9],sink_real[8],sink_real[7],sink_real[6],sink_real[5],sink_real[4],sink_real[3],sink_real[2],sink_real[1],sink_real[0],sink_imag[15],sink_imag[14],sink_imag[13],sink_imag[12],sink_imag[11],sink_imag[10],sink_imag[9],sink_imag[8],sink_imag[7],sink_imag[6],sink_imag[5],sink_imag[4],
sink_imag[3],sink_imag[2],sink_imag[1],sink_imag[0]}));

fft256_asj_fft_tdl_bit_fft_121_3 \no_del_input_blk:delay_next_block (
	.data_in(\writer|rdy_for_next_block~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.tdl_arr_0(\no_del_input_blk:delay_next_block|tdl_arr[0]~q ),
	.clk(clk));

fft256_asj_fft_1tdp_rom_fft_121 \gen_se:gen_new:twrom (
	.q_a_0(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[0] ),
	.q_b_0(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[0] ),
	.q_a_1(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[1] ),
	.q_b_1(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[1] ),
	.q_a_2(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[2] ),
	.q_b_2(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[2] ),
	.q_a_3(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[3] ),
	.q_b_3(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[3] ),
	.q_a_4(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[4] ),
	.q_b_4(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[4] ),
	.q_a_5(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[5] ),
	.q_b_5(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[5] ),
	.q_a_6(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[6] ),
	.q_b_6(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[6] ),
	.q_a_7(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[7] ),
	.q_b_7(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[7] ),
	.q_a_8(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[8] ),
	.q_b_8(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[8] ),
	.q_a_9(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[9] ),
	.q_b_9(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[9] ),
	.q_a_10(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[10] ),
	.q_b_10(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[10] ),
	.q_a_11(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[11] ),
	.q_b_11(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[11] ),
	.q_a_12(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[12] ),
	.q_b_12(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[12] ),
	.q_a_13(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[13] ),
	.q_b_13(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[13] ),
	.q_a_14(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[14] ),
	.q_b_14(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[14] ),
	.q_a_15(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[15] ),
	.q_b_15(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[15] ),
	.twad_tempo_0(\gen_se:gen_new:twid_factors|twad_tempo[0]~q ),
	.twad_tempe_1(\gen_se:gen_new:twid_factors|twad_tempe[1]~q ),
	.twad_tempe_2(\gen_se:gen_new:twid_factors|twad_tempe[2]~q ),
	.twad_tempe_3(\gen_se:gen_new:twid_factors|twad_tempe[3]~q ),
	.twad_tempe_4(\gen_se:gen_new:twid_factors|twad_tempe[4]~q ),
	.twad_tempe_5(\gen_se:gen_new:twid_factors|twad_tempe[5]~q ),
	.twad_tempo_1(\gen_se:gen_new:twid_factors|twad_tempo[1]~q ),
	.twad_tempo_2(\gen_se:gen_new:twid_factors|twad_tempo[2]~q ),
	.twad_tempo_3(\gen_se:gen_new:twid_factors|twad_tempo[3]~q ),
	.twad_tempo_4(\gen_se:gen_new:twid_factors|twad_tempo[4]~q ),
	.twad_tempo_5(\gen_se:gen_new:twid_factors|twad_tempo[5]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.GND_port(GND_port),
	.clk(clk));

fft256_asj_fft_twadsogen_q_fft_121 \gen_se:gen_new:twid_factors (
	.twad_tempo_0(\gen_se:gen_new:twid_factors|twad_tempo[0]~q ),
	.twad_tempe_1(\gen_se:gen_new:twid_factors|twad_tempe[1]~q ),
	.twad_tempe_2(\gen_se:gen_new:twid_factors|twad_tempe[2]~q ),
	.twad_tempe_3(\gen_se:gen_new:twid_factors|twad_tempe[3]~q ),
	.twad_tempe_4(\gen_se:gen_new:twid_factors|twad_tempe[4]~q ),
	.twad_tempe_5(\gen_se:gen_new:twid_factors|twad_tempe[5]~q ),
	.twad_tempo_1(\gen_se:gen_new:twid_factors|twad_tempo[1]~q ),
	.twad_tempo_2(\gen_se:gen_new:twid_factors|twad_tempo[2]~q ),
	.twad_tempo_3(\gen_se:gen_new:twid_factors|twad_tempo[3]~q ),
	.twad_tempo_4(\gen_se:gen_new:twid_factors|twad_tempo[4]~q ),
	.twad_tempo_5(\gen_se:gen_new:twid_factors|twad_tempo[5]~q ),
	.k_count_tw_0(\k_count_tw[0]~q ),
	.k_count_tw_2(\k_count_tw[2]~q ),
	.k_count_tw_1(\k_count_tw[1]~q ),
	.k_count_tw_3(\k_count_tw[3]~q ),
	.k_count_tw_5(\k_count_tw[5]~q ),
	.k_count_tw_4(\k_count_tw[4]~q ),
	.k_count_tw_7(\k_count_tw[7]~q ),
	.k_count_tw_6(\k_count_tw[6]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.quad_reg_2(\gen_se:gen_new:twid_factors|quad_reg[2]~q ),
	.quad_reg_0(\gen_se:gen_new:twid_factors|quad_reg[0]~q ),
	.quad_reg_1(\gen_se:gen_new:twid_factors|quad_reg[1]~q ),
	.p_tdl_0_10(\p_tdl[10][0]~q ),
	.p_tdl_1_10(\p_tdl[10][1]~q ),
	.p_tdl_2_10(\p_tdl[10][2]~q ),
	.data_addr_held_by1(\gen_se:gen_new:twid_factors|data_addr_held_by1~0_combout ),
	.data_addr_held_by2(\gen_se:gen_new:twid_factors|data_addr_held_by2~0_combout ),
	.clk(clk));

fft256_asj_fft_bfp_ctrl_fft_121 \gen_se:bfpc (
	.rdy_for_next_block(\writer|rdy_for_next_block~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.blk_exp_0(\gen_se:bfpc|blk_exp[0]~q ),
	.blk_exp_1(\gen_se:bfpc|blk_exp[1]~q ),
	.blk_exp_2(\gen_se:bfpc|blk_exp[2]~q ),
	.blk_exp_3(\gen_se:bfpc|blk_exp[3]~q ),
	.blk_exp_4(\gen_se:bfpc|blk_exp[4]~q ),
	.blk_exp_5(\gen_se:bfpc|blk_exp[5]~q ),
	.sop_d(\sop_d~q ),
	.slb_i_0(\gen_se:bfpdft|bfp_detect|slb_i[0]~q ),
	.Mux2(\gen_se:bfpdft|bfp_detect|Mux2~0_combout ),
	.lut_out_0(\gen_se:bfpdft|bfp_detect|lut_out[0]~0_combout ),
	.tdl_arr_0(\gen_se:bfpc|gen_so_crtl:gen_se_so:delay_next_pass_2|tdl_arr[0]~q ),
	.Mux1(\gen_se:bfpdft|bfp_detect|Mux1~0_combout ),
	.lut_out_1(\gen_se:bfpdft|bfp_detect|lut_out[1]~1_combout ),
	.lut_out_2(\gen_se:bfpdft|bfp_detect|lut_out[2]~2_combout ),
	.lut_out_21(\gen_se:bfpdft|bfp_detect|lut_out[2]~3_combout ),
	.tdl_arr_9(\delay_swd|tdl_arr[9]~q ),
	.slb_last_1(\gen_se:bfpc|slb_last[1]~q ),
	.slb_last_0(\gen_se:bfpc|slb_last[0]~q ),
	.slb_last_2(\gen_se:bfpc|slb_last[2]~q ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

fft256_asj_fft_dft_bfp_sgl_fft_121 \gen_se:bfpdft (
	.pipeline_dffe_16(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_18(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_19(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_20(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_21(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_22(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_23(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~q ),
	.pipeline_dffe_24(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~q ),
	.pipeline_dffe_25(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~q ),
	.pipeline_dffe_26(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~q ),
	.pipeline_dffe_27(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_28(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_29(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_30(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_31(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~q ),
	.twiddle_data_real_0(\twiddle_data_real[0]~q ),
	.twiddle_data_real_15(\twiddle_data_real[15]~q ),
	.twiddle_data_imag_1(\twiddle_data_imag[1]~q ),
	.twiddle_data_imag_2(\twiddle_data_imag[2]~q ),
	.twiddle_data_imag_3(\twiddle_data_imag[3]~q ),
	.twiddle_data_imag_4(\twiddle_data_imag[4]~q ),
	.twiddle_data_imag_5(\twiddle_data_imag[5]~q ),
	.twiddle_data_imag_6(\twiddle_data_imag[6]~q ),
	.twiddle_data_imag_7(\twiddle_data_imag[7]~q ),
	.twiddle_data_imag_8(\twiddle_data_imag[8]~q ),
	.twiddle_data_imag_9(\twiddle_data_imag[9]~q ),
	.twiddle_data_imag_10(\twiddle_data_imag[10]~q ),
	.twiddle_data_imag_11(\twiddle_data_imag[11]~q ),
	.twiddle_data_imag_12(\twiddle_data_imag[12]~q ),
	.twiddle_data_imag_13(\twiddle_data_imag[13]~q ),
	.twiddle_data_imag_14(\twiddle_data_imag[14]~q ),
	.twiddle_data_imag_15(\twiddle_data_imag[15]~q ),
	.source_valid_ctrl_sop(\source_valid_ctrl_sop~1_combout ),
	.stall_reg(\auk_dsp_interface_controller_1|stall_reg~q ),
	.source_stall_int_d(\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.slb_i_0(\gen_se:bfpdft|bfp_detect|slb_i[0]~q ),
	.Mux2(\gen_se:bfpdft|bfp_detect|Mux2~0_combout ),
	.lut_out_0(\gen_se:bfpdft|bfp_detect|lut_out[0]~0_combout ),
	.tdl_arr_0(\gen_se:bfpc|gen_so_crtl:gen_se_so:delay_next_pass_2|tdl_arr[0]~q ),
	.Mux1(\gen_se:bfpdft|bfp_detect|Mux1~0_combout ),
	.lut_out_1(\gen_se:bfpdft|bfp_detect|lut_out[1]~1_combout ),
	.lut_out_2(\gen_se:bfpdft|bfp_detect|lut_out[2]~2_combout ),
	.lut_out_21(\gen_se:bfpdft|bfp_detect|lut_out[2]~3_combout ),
	.real_out_0(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[0]~q ),
	.real_out_1(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[1]~q ),
	.real_out_2(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[2]~q ),
	.real_out_3(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[3]~q ),
	.real_out_4(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[4]~q ),
	.real_out_5(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[5]~q ),
	.real_out_6(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[6]~q ),
	.real_out_7(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[7]~q ),
	.real_out_8(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[8]~q ),
	.real_out_9(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[9]~q ),
	.real_out_10(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[10]~q ),
	.real_out_11(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[11]~q ),
	.real_out_12(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[12]~q ),
	.real_out_13(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[13]~q ),
	.real_out_14(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[14]~q ),
	.real_out_15(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[15]~q ),
	.tdl_arr_01(\no_del_input_blk:delay_next_block|tdl_arr[0]~q ),
	.k_count_0(\ctrl|k_count[0]~q ),
	.k_count_1(\ctrl|k_count[1]~q ),
	.twiddle_data_real_1(\twiddle_data_real[1]~q ),
	.twiddle_data_real_2(\twiddle_data_real[2]~q ),
	.twiddle_data_real_3(\twiddle_data_real[3]~q ),
	.twiddle_data_real_4(\twiddle_data_real[4]~q ),
	.twiddle_data_real_5(\twiddle_data_real[5]~q ),
	.twiddle_data_real_6(\twiddle_data_real[6]~q ),
	.twiddle_data_real_7(\twiddle_data_real[7]~q ),
	.twiddle_data_real_8(\twiddle_data_real[8]~q ),
	.twiddle_data_real_9(\twiddle_data_real[9]~q ),
	.twiddle_data_real_10(\twiddle_data_real[10]~q ),
	.twiddle_data_real_11(\twiddle_data_real[11]~q ),
	.twiddle_data_real_12(\twiddle_data_real[12]~q ),
	.twiddle_data_real_13(\twiddle_data_real[13]~q ),
	.twiddle_data_real_14(\twiddle_data_real[14]~q ),
	.twiddle_data_imag_0(\twiddle_data_imag[0]~q ),
	.ram_data_out_0(\ccc|ram_data_out[0]~q ),
	.ram_data_out_2(\ccc|ram_data_out[2]~q ),
	.slb_last_1(\gen_se:bfpc|slb_last[1]~q ),
	.ram_data_out_1(\ccc|ram_data_out[1]~q ),
	.slb_last_0(\gen_se:bfpc|slb_last[0]~q ),
	.slb_last_2(\gen_se:bfpc|slb_last[2]~q ),
	.ram_data_out_14(\ccc|ram_data_out[14]~q ),
	.ram_data_out_12(\ccc|ram_data_out[12]~q ),
	.ram_data_out_13(\ccc|ram_data_out[13]~q ),
	.ram_data_out_15(\ccc|ram_data_out[15]~q ),
	.ram_data_out_11(\ccc|ram_data_out[11]~q ),
	.ram_data_out_10(\ccc|ram_data_out[10]~q ),
	.ram_data_out_9(\ccc|ram_data_out[9]~q ),
	.ram_data_out_8(\ccc|ram_data_out[8]~q ),
	.ram_data_out_7(\ccc|ram_data_out[7]~q ),
	.ram_data_out_6(\ccc|ram_data_out[6]~q ),
	.ram_data_out_5(\ccc|ram_data_out[5]~q ),
	.ram_data_out_4(\ccc|ram_data_out[4]~q ),
	.ram_data_out_3(\ccc|ram_data_out[3]~q ),
	.ram_data_out_16(\ccc|ram_data_out[16]~q ),
	.ram_data_out_18(\ccc|ram_data_out[18]~q ),
	.ram_data_out_17(\ccc|ram_data_out[17]~q ),
	.ram_data_out_28(\ccc|ram_data_out[28]~q ),
	.ram_data_out_29(\ccc|ram_data_out[29]~q ),
	.ram_data_out_30(\ccc|ram_data_out[30]~q ),
	.ram_data_out_31(\ccc|ram_data_out[31]~q ),
	.ram_data_out_27(\ccc|ram_data_out[27]~q ),
	.ram_data_out_26(\ccc|ram_data_out[26]~q ),
	.ram_data_out_25(\ccc|ram_data_out[25]~q ),
	.ram_data_out_24(\ccc|ram_data_out[24]~q ),
	.ram_data_out_23(\ccc|ram_data_out[23]~q ),
	.ram_data_out_22(\ccc|ram_data_out[22]~q ),
	.ram_data_out_21(\ccc|ram_data_out[21]~q ),
	.ram_data_out_20(\ccc|ram_data_out[20]~q ),
	.ram_data_out_19(\ccc|ram_data_out[19]~q ),
	.clk(clk),
	.reset(reset_n));

fft256_asj_fft_dataadgen_fft_121 \gen_wraddr_se:wr_adgen (
	.k_count_wr_2(\k_count_wr[2]~q ),
	.k_count_wr_0(\k_count_wr[0]~q ),
	.k_count_wr_6(\k_count_wr[6]~q ),
	.k_count_wr_3(\k_count_wr[3]~q ),
	.k_count_wr_1(\k_count_wr[1]~q ),
	.k_count_wr_7(\k_count_wr[7]~q ),
	.k_count_wr_4(\k_count_wr[4]~q ),
	.k_count_wr_5(\k_count_wr[5]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.rd_addr_a_0(\gen_wraddr_se:wr_adgen|rd_addr_a[0]~q ),
	.rd_addr_a_1(\gen_wraddr_se:wr_adgen|rd_addr_a[1]~q ),
	.rd_addr_a_2(\gen_wraddr_se:wr_adgen|rd_addr_a[2]~q ),
	.rd_addr_a_3(\gen_wraddr_se:wr_adgen|rd_addr_a[3]~q ),
	.rd_addr_a_4(\gen_wraddr_se:wr_adgen|rd_addr_a[4]~q ),
	.rd_addr_a_5(\gen_wraddr_se:wr_adgen|rd_addr_a[5]~q ),
	.rd_addr_a_6(\gen_wraddr_se:wr_adgen|rd_addr_a[6]~q ),
	.rd_addr_a_7(\gen_wraddr_se:wr_adgen|rd_addr_a[7]~q ),
	.p_tdl_0_18(\p_tdl[18][0]~q ),
	.p_tdl_1_18(\p_tdl[18][1]~q ),
	.p_tdl_2_18(\p_tdl[18][2]~q ),
	.clk(clk));

fft256_asj_fft_dataadgen_fft_121_1 rd_adgen(
	.global_clock_enable(\global_clock_enable~0_combout ),
	.rd_addr_a_0(\rd_adgen|rd_addr_a[0]~q ),
	.rd_addr_a_1(\rd_adgen|rd_addr_a[1]~q ),
	.rd_addr_a_2(\rd_adgen|rd_addr_a[2]~q ),
	.rd_addr_a_3(\rd_adgen|rd_addr_a[3]~q ),
	.rd_addr_a_4(\rd_adgen|rd_addr_a[4]~q ),
	.rd_addr_a_5(\rd_adgen|rd_addr_a[5]~q ),
	.rd_addr_a_6(\rd_adgen|rd_addr_a[6]~q ),
	.rd_addr_a_7(\rd_adgen|rd_addr_a[7]~q ),
	.p_2(\ctrl|p[2]~q ),
	.p_0(\ctrl|p[0]~q ),
	.p_1(\ctrl|p[1]~q ),
	.rd_addr_a_01(\rd_adgen|rd_addr_a[0]~0_combout ),
	.k_count_2(\ctrl|k_count[2]~q ),
	.k_count_0(\ctrl|k_count[0]~q ),
	.k_count_6(\ctrl|k_count[6]~q ),
	.k_count_3(\ctrl|k_count[3]~q ),
	.k_count_1(\ctrl|k_count[1]~q ),
	.k_count_7(\ctrl|k_count[7]~q ),
	.k_count_4(\ctrl|k_count[4]~q ),
	.k_count_5(\ctrl|k_count[5]~q ),
	.clk(clk));

fft256_asj_fft_1dp_ram_fft_121 \gen_1_ram:gen_M4K:dat_A (
	.q_b_0(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_16(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[16] ),
	.q_b_1(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_17(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[17] ),
	.q_b_2(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_18(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[18] ),
	.q_b_3(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_19(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[19] ),
	.q_b_4(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_20(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[20] ),
	.q_b_5(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_21(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[21] ),
	.q_b_6(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_22(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[22] ),
	.q_b_7(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_23(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[23] ),
	.q_b_8(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_24(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[24] ),
	.q_b_9(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_25(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[25] ),
	.q_b_10(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_26(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[26] ),
	.q_b_11(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_27(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[27] ),
	.q_b_12(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_28(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[28] ),
	.q_b_13(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_29(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[29] ),
	.q_b_14(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_30(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[30] ),
	.q_b_15(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_31(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[31] ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.wren_a(\wren_a~q ),
	.a_ram_data_in_bus_0(\ccc|a_ram_data_in_bus[0]~q ),
	.wraddress_a_bus_0(\ccc|wraddress_a_bus[0]~q ),
	.wraddress_a_bus_1(\ccc|wraddress_a_bus[1]~q ),
	.wraddress_a_bus_2(\ccc|wraddress_a_bus[2]~q ),
	.wraddress_a_bus_3(\ccc|wraddress_a_bus[3]~q ),
	.wraddress_a_bus_4(\ccc|wraddress_a_bus[4]~q ),
	.wraddress_a_bus_5(\ccc|wraddress_a_bus[5]~q ),
	.wraddress_a_bus_6(\ccc|wraddress_a_bus[6]~q ),
	.wraddress_a_bus_7(\ccc|wraddress_a_bus[7]~q ),
	.rdaddress_a_bus_0(\ccc|rdaddress_a_bus[0]~q ),
	.rdaddress_a_bus_1(\ccc|rdaddress_a_bus[1]~q ),
	.rdaddress_a_bus_2(\ccc|rdaddress_a_bus[2]~q ),
	.rdaddress_a_bus_3(\ccc|rdaddress_a_bus[3]~q ),
	.rdaddress_a_bus_4(\ccc|rdaddress_a_bus[4]~q ),
	.rdaddress_a_bus_5(\ccc|rdaddress_a_bus[5]~q ),
	.rdaddress_a_bus_6(\ccc|rdaddress_a_bus[6]~q ),
	.rdaddress_a_bus_7(\ccc|rdaddress_a_bus[7]~q ),
	.a_ram_data_in_bus_16(\ccc|a_ram_data_in_bus[16]~q ),
	.a_ram_data_in_bus_1(\ccc|a_ram_data_in_bus[1]~q ),
	.a_ram_data_in_bus_17(\ccc|a_ram_data_in_bus[17]~q ),
	.a_ram_data_in_bus_2(\ccc|a_ram_data_in_bus[2]~q ),
	.a_ram_data_in_bus_18(\ccc|a_ram_data_in_bus[18]~q ),
	.a_ram_data_in_bus_3(\ccc|a_ram_data_in_bus[3]~q ),
	.a_ram_data_in_bus_19(\ccc|a_ram_data_in_bus[19]~q ),
	.a_ram_data_in_bus_4(\ccc|a_ram_data_in_bus[4]~q ),
	.a_ram_data_in_bus_20(\ccc|a_ram_data_in_bus[20]~q ),
	.a_ram_data_in_bus_5(\ccc|a_ram_data_in_bus[5]~q ),
	.a_ram_data_in_bus_21(\ccc|a_ram_data_in_bus[21]~q ),
	.a_ram_data_in_bus_6(\ccc|a_ram_data_in_bus[6]~q ),
	.a_ram_data_in_bus_22(\ccc|a_ram_data_in_bus[22]~q ),
	.a_ram_data_in_bus_7(\ccc|a_ram_data_in_bus[7]~q ),
	.a_ram_data_in_bus_23(\ccc|a_ram_data_in_bus[23]~q ),
	.a_ram_data_in_bus_8(\ccc|a_ram_data_in_bus[8]~q ),
	.a_ram_data_in_bus_24(\ccc|a_ram_data_in_bus[24]~q ),
	.a_ram_data_in_bus_9(\ccc|a_ram_data_in_bus[9]~q ),
	.a_ram_data_in_bus_25(\ccc|a_ram_data_in_bus[25]~q ),
	.a_ram_data_in_bus_10(\ccc|a_ram_data_in_bus[10]~q ),
	.a_ram_data_in_bus_26(\ccc|a_ram_data_in_bus[26]~q ),
	.a_ram_data_in_bus_11(\ccc|a_ram_data_in_bus[11]~q ),
	.a_ram_data_in_bus_27(\ccc|a_ram_data_in_bus[27]~q ),
	.a_ram_data_in_bus_12(\ccc|a_ram_data_in_bus[12]~q ),
	.a_ram_data_in_bus_28(\ccc|a_ram_data_in_bus[28]~q ),
	.a_ram_data_in_bus_13(\ccc|a_ram_data_in_bus[13]~q ),
	.a_ram_data_in_bus_29(\ccc|a_ram_data_in_bus[29]~q ),
	.a_ram_data_in_bus_14(\ccc|a_ram_data_in_bus[14]~q ),
	.a_ram_data_in_bus_30(\ccc|a_ram_data_in_bus[30]~q ),
	.a_ram_data_in_bus_15(\ccc|a_ram_data_in_bus[15]~q ),
	.a_ram_data_in_bus_31(\ccc|a_ram_data_in_bus[31]~q ),
	.clk(clk));

fft256_asj_fft_unbburst_sose_ctrl_fft_121 ccc(
	.q_b_0(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.q_b_16(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[16] ),
	.q_b_1(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.q_b_17(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[17] ),
	.q_b_2(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.q_b_18(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[18] ),
	.q_b_3(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.q_b_19(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[19] ),
	.q_b_4(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.q_b_20(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[20] ),
	.q_b_5(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.q_b_21(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[21] ),
	.q_b_6(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.q_b_22(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[22] ),
	.q_b_7(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.q_b_23(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[23] ),
	.q_b_8(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.q_b_24(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[24] ),
	.q_b_9(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.q_b_25(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[25] ),
	.q_b_10(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.q_b_26(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[26] ),
	.q_b_11(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.q_b_27(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[27] ),
	.q_b_12(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.q_b_28(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[28] ),
	.q_b_13(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.q_b_29(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[29] ),
	.q_b_14(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.q_b_30(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[30] ),
	.q_b_15(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.q_b_31(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[31] ),
	.pipeline_dffe_16(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_18(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_19(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_20(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_21(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_22(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_23(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~q ),
	.pipeline_dffe_24(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~q ),
	.pipeline_dffe_25(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~q ),
	.pipeline_dffe_26(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~q ),
	.pipeline_dffe_27(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_28(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_29(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_30(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_31(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.a_ram_data_in_bus_0(\ccc|a_ram_data_in_bus[0]~q ),
	.wraddress_a_bus_0(\ccc|wraddress_a_bus[0]~q ),
	.wraddress_a_bus_1(\ccc|wraddress_a_bus[1]~q ),
	.wraddress_a_bus_2(\ccc|wraddress_a_bus[2]~q ),
	.wraddress_a_bus_3(\ccc|wraddress_a_bus[3]~q ),
	.wraddress_a_bus_4(\ccc|wraddress_a_bus[4]~q ),
	.wraddress_a_bus_5(\ccc|wraddress_a_bus[5]~q ),
	.wraddress_a_bus_6(\ccc|wraddress_a_bus[6]~q ),
	.wraddress_a_bus_7(\ccc|wraddress_a_bus[7]~q ),
	.rdaddress_a_bus_0(\ccc|rdaddress_a_bus[0]~q ),
	.rdaddress_a_bus_1(\ccc|rdaddress_a_bus[1]~q ),
	.rdaddress_a_bus_2(\ccc|rdaddress_a_bus[2]~q ),
	.rdaddress_a_bus_3(\ccc|rdaddress_a_bus[3]~q ),
	.rdaddress_a_bus_4(\ccc|rdaddress_a_bus[4]~q ),
	.rdaddress_a_bus_5(\ccc|rdaddress_a_bus[5]~q ),
	.rdaddress_a_bus_6(\ccc|rdaddress_a_bus[6]~q ),
	.rdaddress_a_bus_7(\ccc|rdaddress_a_bus[7]~q ),
	.a_ram_data_in_bus_16(\ccc|a_ram_data_in_bus[16]~q ),
	.a_ram_data_in_bus_1(\ccc|a_ram_data_in_bus[1]~q ),
	.a_ram_data_in_bus_17(\ccc|a_ram_data_in_bus[17]~q ),
	.a_ram_data_in_bus_2(\ccc|a_ram_data_in_bus[2]~q ),
	.a_ram_data_in_bus_18(\ccc|a_ram_data_in_bus[18]~q ),
	.a_ram_data_in_bus_3(\ccc|a_ram_data_in_bus[3]~q ),
	.a_ram_data_in_bus_19(\ccc|a_ram_data_in_bus[19]~q ),
	.a_ram_data_in_bus_4(\ccc|a_ram_data_in_bus[4]~q ),
	.a_ram_data_in_bus_20(\ccc|a_ram_data_in_bus[20]~q ),
	.a_ram_data_in_bus_5(\ccc|a_ram_data_in_bus[5]~q ),
	.a_ram_data_in_bus_21(\ccc|a_ram_data_in_bus[21]~q ),
	.a_ram_data_in_bus_6(\ccc|a_ram_data_in_bus[6]~q ),
	.a_ram_data_in_bus_22(\ccc|a_ram_data_in_bus[22]~q ),
	.a_ram_data_in_bus_7(\ccc|a_ram_data_in_bus[7]~q ),
	.a_ram_data_in_bus_23(\ccc|a_ram_data_in_bus[23]~q ),
	.a_ram_data_in_bus_8(\ccc|a_ram_data_in_bus[8]~q ),
	.a_ram_data_in_bus_24(\ccc|a_ram_data_in_bus[24]~q ),
	.a_ram_data_in_bus_9(\ccc|a_ram_data_in_bus[9]~q ),
	.a_ram_data_in_bus_25(\ccc|a_ram_data_in_bus[25]~q ),
	.a_ram_data_in_bus_10(\ccc|a_ram_data_in_bus[10]~q ),
	.a_ram_data_in_bus_26(\ccc|a_ram_data_in_bus[26]~q ),
	.a_ram_data_in_bus_11(\ccc|a_ram_data_in_bus[11]~q ),
	.a_ram_data_in_bus_27(\ccc|a_ram_data_in_bus[27]~q ),
	.a_ram_data_in_bus_12(\ccc|a_ram_data_in_bus[12]~q ),
	.a_ram_data_in_bus_28(\ccc|a_ram_data_in_bus[28]~q ),
	.a_ram_data_in_bus_13(\ccc|a_ram_data_in_bus[13]~q ),
	.a_ram_data_in_bus_29(\ccc|a_ram_data_in_bus[29]~q ),
	.a_ram_data_in_bus_14(\ccc|a_ram_data_in_bus[14]~q ),
	.a_ram_data_in_bus_30(\ccc|a_ram_data_in_bus[30]~q ),
	.a_ram_data_in_bus_15(\ccc|a_ram_data_in_bus[15]~q ),
	.a_ram_data_in_bus_31(\ccc|a_ram_data_in_bus[31]~q ),
	.data_rdy_vec_21(\data_rdy_vec[21]~q ),
	.real_out_0(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[0]~q ),
	.data_in_i_0(\writer|data_in_i[0]~q ),
	.sel_ram_in(\sel_ram_in~q ),
	.wraddress_a_bus_ctrl_i_0(\wraddress_a_bus_ctrl_i[0]~q ),
	.wr_address_i_int_0(\writer|wr_address_i_int[0]~q ),
	.wraddress_a_bus_ctrl_i_1(\wraddress_a_bus_ctrl_i[1]~q ),
	.wr_address_i_int_1(\writer|wr_address_i_int[1]~q ),
	.wraddress_a_bus_ctrl_i_2(\wraddress_a_bus_ctrl_i[2]~q ),
	.wr_address_i_int_2(\writer|wr_address_i_int[2]~q ),
	.wraddress_a_bus_ctrl_i_3(\wraddress_a_bus_ctrl_i[3]~q ),
	.wr_address_i_int_3(\writer|wr_address_i_int[3]~q ),
	.wraddress_a_bus_ctrl_i_4(\wraddress_a_bus_ctrl_i[4]~q ),
	.wr_address_i_int_4(\writer|wr_address_i_int[4]~q ),
	.wraddress_a_bus_ctrl_i_5(\wraddress_a_bus_ctrl_i[5]~q ),
	.wr_address_i_int_5(\writer|wr_address_i_int[5]~q ),
	.wraddress_a_bus_ctrl_i_6(\wraddress_a_bus_ctrl_i[6]~q ),
	.wr_address_i_int_6(\writer|wr_address_i_int[6]~q ),
	.wraddress_a_bus_ctrl_i_7(\wraddress_a_bus_ctrl_i[7]~q ),
	.wr_address_i_int_7(\writer|wr_address_i_int[7]~q ),
	.rd_addr_a_0(\rd_adgen|rd_addr_a[0]~q ),
	.rd_addr_a_1(\rd_adgen|rd_addr_a[1]~q ),
	.rd_addr_a_2(\rd_adgen|rd_addr_a[2]~q ),
	.rd_addr_a_3(\rd_adgen|rd_addr_a[3]~q ),
	.rd_addr_a_4(\rd_adgen|rd_addr_a[4]~q ),
	.rd_addr_a_5(\rd_adgen|rd_addr_a[5]~q ),
	.rd_addr_a_6(\rd_adgen|rd_addr_a[6]~q ),
	.rd_addr_a_7(\rd_adgen|rd_addr_a[7]~q ),
	.data_in_r_0(\writer|data_in_r[0]~q ),
	.real_out_1(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[1]~q ),
	.data_in_i_1(\writer|data_in_i[1]~q ),
	.data_in_r_1(\writer|data_in_r[1]~q ),
	.real_out_2(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[2]~q ),
	.data_in_i_2(\writer|data_in_i[2]~q ),
	.data_in_r_2(\writer|data_in_r[2]~q ),
	.real_out_3(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[3]~q ),
	.data_in_i_3(\writer|data_in_i[3]~q ),
	.data_in_r_3(\writer|data_in_r[3]~q ),
	.real_out_4(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[4]~q ),
	.data_in_i_4(\writer|data_in_i[4]~q ),
	.data_in_r_4(\writer|data_in_r[4]~q ),
	.real_out_5(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[5]~q ),
	.data_in_i_5(\writer|data_in_i[5]~q ),
	.data_in_r_5(\writer|data_in_r[5]~q ),
	.real_out_6(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[6]~q ),
	.data_in_i_6(\writer|data_in_i[6]~q ),
	.data_in_r_6(\writer|data_in_r[6]~q ),
	.real_out_7(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[7]~q ),
	.data_in_i_7(\writer|data_in_i[7]~q ),
	.data_in_r_7(\writer|data_in_r[7]~q ),
	.real_out_8(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[8]~q ),
	.data_in_i_8(\writer|data_in_i[8]~q ),
	.data_in_r_8(\writer|data_in_r[8]~q ),
	.real_out_9(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[9]~q ),
	.data_in_i_9(\writer|data_in_i[9]~q ),
	.data_in_r_9(\writer|data_in_r[9]~q ),
	.real_out_10(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[10]~q ),
	.data_in_i_10(\writer|data_in_i[10]~q ),
	.data_in_r_10(\writer|data_in_r[10]~q ),
	.real_out_11(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[11]~q ),
	.data_in_i_11(\writer|data_in_i[11]~q ),
	.data_in_r_11(\writer|data_in_r[11]~q ),
	.real_out_12(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[12]~q ),
	.data_in_i_12(\writer|data_in_i[12]~q ),
	.data_in_r_12(\writer|data_in_r[12]~q ),
	.real_out_13(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[13]~q ),
	.data_in_i_13(\writer|data_in_i[13]~q ),
	.data_in_r_13(\writer|data_in_r[13]~q ),
	.real_out_14(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[14]~q ),
	.data_in_i_14(\writer|data_in_i[14]~q ),
	.data_in_r_14(\writer|data_in_r[14]~q ),
	.real_out_15(\gen_se:bfpdft|gen_da0:gen_canonic:cm1|real_out[15]~q ),
	.data_in_i_15(\writer|data_in_i[15]~q ),
	.data_in_r_15(\writer|data_in_r[15]~q ),
	.ram_data_out_0(\ccc|ram_data_out[0]~q ),
	.ram_data_out_2(\ccc|ram_data_out[2]~q ),
	.ram_data_out_1(\ccc|ram_data_out[1]~q ),
	.ram_data_out_14(\ccc|ram_data_out[14]~q ),
	.ram_data_out_12(\ccc|ram_data_out[12]~q ),
	.ram_data_out_13(\ccc|ram_data_out[13]~q ),
	.ram_data_out_15(\ccc|ram_data_out[15]~q ),
	.ram_data_out_11(\ccc|ram_data_out[11]~q ),
	.ram_data_out_10(\ccc|ram_data_out[10]~q ),
	.ram_data_out_9(\ccc|ram_data_out[9]~q ),
	.ram_data_out_8(\ccc|ram_data_out[8]~q ),
	.ram_data_out_7(\ccc|ram_data_out[7]~q ),
	.ram_data_out_6(\ccc|ram_data_out[6]~q ),
	.ram_data_out_5(\ccc|ram_data_out[5]~q ),
	.ram_data_out_4(\ccc|ram_data_out[4]~q ),
	.ram_data_out_3(\ccc|ram_data_out[3]~q ),
	.ram_data_out_16(\ccc|ram_data_out[16]~q ),
	.ram_data_out_18(\ccc|ram_data_out[18]~q ),
	.ram_data_out_17(\ccc|ram_data_out[17]~q ),
	.ram_data_out_28(\ccc|ram_data_out[28]~q ),
	.ram_data_out_29(\ccc|ram_data_out[29]~q ),
	.ram_data_out_30(\ccc|ram_data_out[30]~q ),
	.ram_data_out_31(\ccc|ram_data_out[31]~q ),
	.ram_data_out_27(\ccc|ram_data_out[27]~q ),
	.ram_data_out_26(\ccc|ram_data_out[26]~q ),
	.ram_data_out_25(\ccc|ram_data_out[25]~q ),
	.ram_data_out_24(\ccc|ram_data_out[24]~q ),
	.ram_data_out_23(\ccc|ram_data_out[23]~q ),
	.ram_data_out_22(\ccc|ram_data_out[22]~q ),
	.ram_data_out_21(\ccc|ram_data_out[21]~q ),
	.ram_data_out_20(\ccc|ram_data_out[20]~q ),
	.ram_data_out_19(\ccc|ram_data_out[19]~q ),
	.clk(clk));

fft256_asj_fft_in_write_sgl_fft_121 writer(
	.disable_wr1(\writer|disable_wr~q ),
	.rdy_for_next_block1(\writer|rdy_for_next_block~q ),
	.core_imag_in_0(\core_imag_in[0]~q ),
	.core_real_in_0(\core_real_in[0]~q ),
	.core_imag_in_1(\core_imag_in[1]~q ),
	.core_real_in_1(\core_real_in[1]~q ),
	.core_imag_in_2(\core_imag_in[2]~q ),
	.core_real_in_2(\core_real_in[2]~q ),
	.core_imag_in_3(\core_imag_in[3]~q ),
	.core_real_in_3(\core_real_in[3]~q ),
	.core_imag_in_4(\core_imag_in[4]~q ),
	.core_real_in_4(\core_real_in[4]~q ),
	.core_imag_in_5(\core_imag_in[5]~q ),
	.core_real_in_5(\core_real_in[5]~q ),
	.core_imag_in_6(\core_imag_in[6]~q ),
	.core_real_in_6(\core_real_in[6]~q ),
	.core_imag_in_7(\core_imag_in[7]~q ),
	.core_real_in_7(\core_real_in[7]~q ),
	.core_imag_in_8(\core_imag_in[8]~q ),
	.core_real_in_8(\core_real_in[8]~q ),
	.core_imag_in_9(\core_imag_in[9]~q ),
	.core_real_in_9(\core_real_in[9]~q ),
	.core_imag_in_10(\core_imag_in[10]~q ),
	.core_real_in_10(\core_real_in[10]~q ),
	.core_imag_in_11(\core_imag_in[11]~q ),
	.core_real_in_11(\core_real_in[11]~q ),
	.core_imag_in_12(\core_imag_in[12]~q ),
	.core_real_in_12(\core_real_in[12]~q ),
	.core_imag_in_13(\core_imag_in[13]~q ),
	.core_real_in_13(\core_real_in[13]~q ),
	.core_imag_in_14(\core_imag_in[14]~q ),
	.core_real_in_14(\core_real_in[14]~q ),
	.core_imag_in_15(\core_imag_in[15]~q ),
	.core_real_in_15(\core_real_in[15]~q ),
	.data_rdy_int1(\writer|data_rdy_int~q ),
	.send_sop_s(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.blk_done(\ctrl|blk_done~q ),
	.tdl_arr_0(\writer|gen_soe:delay_swd|tdl_arr[0]~q ),
	.data_in_i_0(\writer|data_in_i[0]~q ),
	.wr_address_i_int_0(\writer|wr_address_i_int[0]~q ),
	.wr_address_i_int_1(\writer|wr_address_i_int[1]~q ),
	.wr_address_i_int_2(\writer|wr_address_i_int[2]~q ),
	.wr_address_i_int_3(\writer|wr_address_i_int[3]~q ),
	.wr_address_i_int_4(\writer|wr_address_i_int[4]~q ),
	.wr_address_i_int_5(\writer|wr_address_i_int[5]~q ),
	.wr_address_i_int_6(\writer|wr_address_i_int[6]~q ),
	.wr_address_i_int_7(\writer|wr_address_i_int[7]~q ),
	.data_in_r_0(\writer|data_in_r[0]~q ),
	.data_in_i_1(\writer|data_in_i[1]~q ),
	.data_in_r_1(\writer|data_in_r[1]~q ),
	.data_in_i_2(\writer|data_in_i[2]~q ),
	.data_in_r_2(\writer|data_in_r[2]~q ),
	.data_in_i_3(\writer|data_in_i[3]~q ),
	.data_in_r_3(\writer|data_in_r[3]~q ),
	.data_in_i_4(\writer|data_in_i[4]~q ),
	.data_in_r_4(\writer|data_in_r[4]~q ),
	.data_in_i_5(\writer|data_in_i[5]~q ),
	.data_in_r_5(\writer|data_in_r[5]~q ),
	.data_in_i_6(\writer|data_in_i[6]~q ),
	.data_in_r_6(\writer|data_in_r[6]~q ),
	.data_in_i_7(\writer|data_in_i[7]~q ),
	.data_in_r_7(\writer|data_in_r[7]~q ),
	.data_in_i_8(\writer|data_in_i[8]~q ),
	.data_in_r_8(\writer|data_in_r[8]~q ),
	.data_in_i_9(\writer|data_in_i[9]~q ),
	.data_in_r_9(\writer|data_in_r[9]~q ),
	.data_in_i_10(\writer|data_in_i[10]~q ),
	.data_in_r_10(\writer|data_in_r[10]~q ),
	.data_in_i_11(\writer|data_in_i[11]~q ),
	.data_in_r_11(\writer|data_in_r[11]~q ),
	.data_in_i_12(\writer|data_in_i[12]~q ),
	.data_in_r_12(\writer|data_in_r[12]~q ),
	.data_in_i_13(\writer|data_in_i[13]~q ),
	.data_in_r_13(\writer|data_in_r[13]~q ),
	.data_in_i_14(\writer|data_in_i[14]~q ),
	.data_in_r_14(\writer|data_in_r[14]~q ),
	.data_in_i_15(\writer|data_in_i[15]~q ),
	.data_in_r_15(\writer|data_in_r[15]~q ),
	.counter_i(\writer|counter_i~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

fft256_asj_fft_tdl_bit_rst_fft_121_2 delay_swd(
	.global_clock_enable(\global_clock_enable~0_combout ),
	.tdl_arr_9(\delay_swd|tdl_arr[9]~q ),
	.next_pass(\next_pass~combout ),
	.clk(clk),
	.reset_n(reset_n));

fft256_asj_fft_m_k_counter_fft_121 ctrl(
	.rdy_for_next_block(\writer|rdy_for_next_block~q ),
	.send_sop_s(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.blk_done1(\ctrl|blk_done~q ),
	.counter_i(\writer|counter_i~0_combout ),
	.p_2(\ctrl|p[2]~q ),
	.p_0(\ctrl|p[0]~q ),
	.p_1(\ctrl|p[1]~q ),
	.rd_addr_a_0(\rd_adgen|rd_addr_a[0]~0_combout ),
	.k_count_2(\ctrl|k_count[2]~q ),
	.k_count_0(\ctrl|k_count[0]~q ),
	.k_count_6(\ctrl|k_count[6]~q ),
	.k_count_3(\ctrl|k_count[3]~q ),
	.k_count_1(\ctrl|k_count[1]~q ),
	.k_count_7(\ctrl|k_count[7]~q ),
	.k_count_4(\ctrl|k_count[4]~q ),
	.k_count_5(\ctrl|k_count[5]~q ),
	.data_rdy_vec_4(\data_rdy_vec[4]~q ),
	.next_pass_i1(\ctrl|next_pass_i~q ),
	.clk(clk),
	.reset_n(reset_n));

fft256_auk_dspip_avalon_streaming_controller_fft_121 auk_dsp_interface_controller_1(
	.master_sink_ena(\master_sink_ena~q ),
	.source_packet_error_0(\auk_dsp_interface_controller_1|source_packet_error[0]~q ),
	.source_packet_error_1(\auk_dsp_interface_controller_1|source_packet_error[1]~q ),
	.source_stall_reg1(\auk_dsp_interface_controller_1|source_stall_reg~q ),
	.sink_stall_reg1(\auk_dsp_interface_controller_1|sink_stall_reg~q ),
	.sink_ready_ctrl(\auk_dsp_interface_controller_1|sink_ready_ctrl~0_combout ),
	.sink_start(\auk_dsp_atlantic_sink_1|sink_start~q ),
	.empty_dff(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|empty_dff~q ),
	.sink_stall(\auk_dsp_atlantic_sink_1|sink_stall~combout ),
	.packet_error_s_0(\auk_dsp_atlantic_sink_1|packet_error_s[0]~q ),
	.packet_error_s_1(\auk_dsp_atlantic_sink_1|packet_error_s[1]~q ),
	.stall_reg1(\auk_dsp_interface_controller_1|stall_reg~q ),
	.Mux0(\auk_dsp_atlantic_source_1|Mux0~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

fft256_auk_dspip_avalon_streaming_source_fft_121 auk_dsp_atlantic_source_1(
	.data_count({\data_count_sig[7]~q ,\data_count_sig[6]~q ,\data_count_sig[5]~q ,\data_count_sig[4]~q ,\data_count_sig[3]~q ,\data_count_sig[2]~q ,\data_count_sig[1]~q ,\data_count_sig[0]~q }),
	.at_source_error_0(at_source_error_0),
	.at_source_error_1(at_source_error_1),
	.at_source_sop_s1(at_source_sop_s),
	.at_source_eop_s1(at_source_eop_s),
	.at_source_valid_s1(at_source_valid_s),
	.at_source_data_0(at_source_data_0),
	.at_source_data_1(at_source_data_1),
	.at_source_data_2(at_source_data_2),
	.at_source_data_3(at_source_data_3),
	.at_source_data_4(at_source_data_4),
	.at_source_data_5(at_source_data_5),
	.at_source_data_22(at_source_data_22),
	.at_source_data_23(at_source_data_23),
	.at_source_data_24(at_source_data_24),
	.at_source_data_25(at_source_data_25),
	.at_source_data_26(at_source_data_26),
	.at_source_data_27(at_source_data_27),
	.at_source_data_28(at_source_data_28),
	.at_source_data_29(at_source_data_29),
	.at_source_data_30(at_source_data_30),
	.at_source_data_31(at_source_data_31),
	.at_source_data_32(at_source_data_32),
	.at_source_data_33(at_source_data_33),
	.at_source_data_34(at_source_data_34),
	.at_source_data_35(at_source_data_35),
	.at_source_data_36(at_source_data_36),
	.at_source_data_37(at_source_data_37),
	.at_source_data_6(at_source_data_6),
	.at_source_data_7(at_source_data_7),
	.at_source_data_8(at_source_data_8),
	.at_source_data_9(at_source_data_9),
	.at_source_data_10(at_source_data_10),
	.at_source_data_11(at_source_data_11),
	.at_source_data_12(at_source_data_12),
	.at_source_data_13(at_source_data_13),
	.at_source_data_14(at_source_data_14),
	.at_source_data_15(at_source_data_15),
	.at_source_data_16(at_source_data_16),
	.at_source_data_17(at_source_data_17),
	.at_source_data_18(at_source_data_18),
	.at_source_data_19(at_source_data_19),
	.at_source_data_20(at_source_data_20),
	.at_source_data_21(at_source_data_21),
	.source_packet_error_0(\auk_dsp_interface_controller_1|source_packet_error[0]~q ),
	.source_packet_error_1(\auk_dsp_interface_controller_1|source_packet_error[1]~q ),
	.source_stall_reg(\auk_dsp_interface_controller_1|source_stall_reg~q ),
	.master_source_ena(\master_source_ena~q ),
	.source_valid_ctrl_sop(\source_valid_ctrl_sop~0_combout ),
	.source_valid_ctrl_sop1(\source_valid_ctrl_sop~1_combout ),
	.stall_reg(\auk_dsp_interface_controller_1|stall_reg~q ),
	.source_stall_int_d1(\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.data({\fft_real_out[15]~q ,\fft_real_out[14]~q ,\fft_real_out[13]~q ,\fft_real_out[12]~q ,\fft_real_out[11]~q ,\fft_real_out[10]~q ,\fft_real_out[9]~q ,\fft_real_out[8]~q ,\fft_real_out[7]~q ,\fft_real_out[6]~q ,\fft_real_out[5]~q ,\fft_real_out[4]~q ,\fft_real_out[3]~q ,
\fft_real_out[2]~q ,\fft_real_out[1]~q ,\fft_real_out[0]~q ,\fft_imag_out[15]~q ,\fft_imag_out[14]~q ,\fft_imag_out[13]~q ,\fft_imag_out[12]~q ,\fft_imag_out[11]~q ,\fft_imag_out[10]~q ,\fft_imag_out[9]~q ,\fft_imag_out[8]~q ,\fft_imag_out[7]~q ,\fft_imag_out[6]~q ,
\fft_imag_out[5]~q ,\fft_imag_out[4]~q ,\fft_imag_out[3]~q ,\fft_imag_out[2]~q ,\fft_imag_out[1]~q ,\fft_imag_out[0]~q ,\exponent_out[5]~q ,\exponent_out[4]~q ,\exponent_out[3]~q ,\exponent_out[2]~q ,\exponent_out[1]~q ,\exponent_out[0]~q }),
	.Mux0(\auk_dsp_atlantic_source_1|Mux0~1_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.source_ready(source_ready));

dffeas master_sink_ena(
	.clk(clk),
	.d(\WideOr3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\master_sink_ena~q ),
	.prn(vcc));
defparam master_sink_ena.is_wysiwyg = "true";
defparam master_sink_ena.power_up = "low";

dffeas \data_count_sig[6] (
	.clk(clk),
	.d(\data_count_sig[6]~20_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[1]~23_combout ),
	.ena(\data_count_sig[6]~24_combout ),
	.q(\data_count_sig[6]~q ),
	.prn(vcc));
defparam \data_count_sig[6] .is_wysiwyg = "true";
defparam \data_count_sig[6] .power_up = "low";

dffeas \data_count_sig[4] (
	.clk(clk),
	.d(\data_count_sig[4]~16_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[1]~23_combout ),
	.ena(\data_count_sig[6]~24_combout ),
	.q(\data_count_sig[4]~q ),
	.prn(vcc));
defparam \data_count_sig[4] .is_wysiwyg = "true";
defparam \data_count_sig[4] .power_up = "low";

dffeas \data_count_sig[0] (
	.clk(clk),
	.d(\data_count_sig[0]~8_combout ),
	.asdata(\master_source_sop~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[1]~23_combout ),
	.ena(\data_count_sig[6]~24_combout ),
	.q(\data_count_sig[0]~q ),
	.prn(vcc));
defparam \data_count_sig[0] .is_wysiwyg = "true";
defparam \data_count_sig[0] .power_up = "low";

dffeas \data_count_sig[5] (
	.clk(clk),
	.d(\data_count_sig[5]~18_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[1]~23_combout ),
	.ena(\data_count_sig[6]~24_combout ),
	.q(\data_count_sig[5]~q ),
	.prn(vcc));
defparam \data_count_sig[5] .is_wysiwyg = "true";
defparam \data_count_sig[5] .power_up = "low";

dffeas \data_count_sig[1] (
	.clk(clk),
	.d(\data_count_sig[1]~10_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[1]~23_combout ),
	.ena(\data_count_sig[6]~24_combout ),
	.q(\data_count_sig[1]~q ),
	.prn(vcc));
defparam \data_count_sig[1] .is_wysiwyg = "true";
defparam \data_count_sig[1] .power_up = "low";

dffeas \data_count_sig[7] (
	.clk(clk),
	.d(\data_count_sig[7]~25_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[1]~23_combout ),
	.ena(\data_count_sig[6]~24_combout ),
	.q(\data_count_sig[7]~q ),
	.prn(vcc));
defparam \data_count_sig[7] .is_wysiwyg = "true";
defparam \data_count_sig[7] .power_up = "low";

dffeas \data_count_sig[3] (
	.clk(clk),
	.d(\data_count_sig[3]~14_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[1]~23_combout ),
	.ena(\data_count_sig[6]~24_combout ),
	.q(\data_count_sig[3]~q ),
	.prn(vcc));
defparam \data_count_sig[3] .is_wysiwyg = "true";
defparam \data_count_sig[3] .power_up = "low";

dffeas \data_count_sig[2] (
	.clk(clk),
	.d(\data_count_sig[2]~12_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[1]~23_combout ),
	.ena(\data_count_sig[6]~24_combout ),
	.q(\data_count_sig[2]~q ),
	.prn(vcc));
defparam \data_count_sig[2] .is_wysiwyg = "true";
defparam \data_count_sig[2] .power_up = "low";

dffeas \fft_s1_cur.WAIT_FOR_INPUT (
	.clk(clk),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_s1_cur.WAIT_FOR_INPUT~q ),
	.prn(vcc));
defparam \fft_s1_cur.WAIT_FOR_INPUT .is_wysiwyg = "true";
defparam \fft_s1_cur.WAIT_FOR_INPUT .power_up = "low";

dffeas \fft_s1_cur.WRITE_INPUT (
	.clk(clk),
	.d(\Selector6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_s1_cur.WRITE_INPUT~q ),
	.prn(vcc));
defparam \fft_s1_cur.WRITE_INPUT .is_wysiwyg = "true";
defparam \fft_s1_cur.WRITE_INPUT .power_up = "low";

cycloneive_lcell_comb \data_count_sig[0]~8 (
	.dataa(\data_count_sig[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\data_count_sig[0]~8_combout ),
	.cout(\data_count_sig[0]~9 ));
defparam \data_count_sig[0]~8 .lut_mask = 16'h55AA;
defparam \data_count_sig[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_count_sig[1]~10 (
	.dataa(\data_count_sig[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[0]~9 ),
	.combout(\data_count_sig[1]~10_combout ),
	.cout(\data_count_sig[1]~11 ));
defparam \data_count_sig[1]~10 .lut_mask = 16'h5A5F;
defparam \data_count_sig[1]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_count_sig[2]~12 (
	.dataa(\data_count_sig[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[1]~11 ),
	.combout(\data_count_sig[2]~12_combout ),
	.cout(\data_count_sig[2]~13 ));
defparam \data_count_sig[2]~12 .lut_mask = 16'h5AAF;
defparam \data_count_sig[2]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_count_sig[3]~14 (
	.dataa(\data_count_sig[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[2]~13 ),
	.combout(\data_count_sig[3]~14_combout ),
	.cout(\data_count_sig[3]~15 ));
defparam \data_count_sig[3]~14 .lut_mask = 16'h5A5F;
defparam \data_count_sig[3]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_count_sig[4]~16 (
	.dataa(\data_count_sig[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[3]~15 ),
	.combout(\data_count_sig[4]~16_combout ),
	.cout(\data_count_sig[4]~17 ));
defparam \data_count_sig[4]~16 .lut_mask = 16'h5AAF;
defparam \data_count_sig[4]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_count_sig[5]~18 (
	.dataa(\data_count_sig[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[4]~17 ),
	.combout(\data_count_sig[5]~18_combout ),
	.cout(\data_count_sig[5]~19 ));
defparam \data_count_sig[5]~18 .lut_mask = 16'h5A5F;
defparam \data_count_sig[5]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_count_sig[6]~20 (
	.dataa(\data_count_sig[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[5]~19 ),
	.combout(\data_count_sig[6]~20_combout ),
	.cout(\data_count_sig[6]~21 ));
defparam \data_count_sig[6]~20 .lut_mask = 16'h5AAF;
defparam \data_count_sig[6]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_count_sig[7]~25 (
	.dataa(\data_count_sig[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\data_count_sig[6]~21 ),
	.combout(\data_count_sig[7]~25_combout ),
	.cout());
defparam \data_count_sig[7]~25 .lut_mask = 16'h5A5A;
defparam \data_count_sig[7]~25 .sum_lutc_input = "cin";

dffeas \fft_s1_cur.FFT_PROCESS_A (
	.clk(clk),
	.d(\Selector10~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_s1_cur.FFT_PROCESS_A~q ),
	.prn(vcc));
defparam \fft_s1_cur.FFT_PROCESS_A .is_wysiwyg = "true";
defparam \fft_s1_cur.FFT_PROCESS_A .power_up = "low";

dffeas \fft_s2_cur.LPP_OUTPUT_RDY (
	.clk(clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_s2_cur.LPP_OUTPUT_RDY~q ),
	.prn(vcc));
defparam \fft_s2_cur.LPP_OUTPUT_RDY .is_wysiwyg = "true";
defparam \fft_s2_cur.LPP_OUTPUT_RDY .power_up = "low";

dffeas \fft_s2_cur.WAIT_FOR_LPP_INPUT (
	.clk(clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.prn(vcc));
defparam \fft_s2_cur.WAIT_FOR_LPP_INPUT .is_wysiwyg = "true";
defparam \fft_s2_cur.WAIT_FOR_LPP_INPUT .power_up = "low";

dffeas \fft_s2_cur.START_LPP (
	.clk(clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_s2_cur.START_LPP~q ),
	.prn(vcc));
defparam \fft_s2_cur.START_LPP .is_wysiwyg = "true";
defparam \fft_s2_cur.START_LPP .power_up = "low";

dffeas \fft_s1_cur.NO_WRITE (
	.clk(clk),
	.d(\Selector9~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_s1_cur.NO_WRITE~q ),
	.prn(vcc));
defparam \fft_s1_cur.NO_WRITE .is_wysiwyg = "true";
defparam \fft_s1_cur.NO_WRITE .power_up = "low";

dffeas \output_count[1] (
	.clk(clk),
	.d(\output_count[1]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\output_sample_counter~0_combout ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\output_count[1]~q ),
	.prn(vcc));
defparam \output_count[1] .is_wysiwyg = "true";
defparam \output_count[1] .power_up = "low";

dffeas \output_count[2] (
	.clk(clk),
	.d(\output_count[2]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\output_sample_counter~0_combout ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\output_count[2]~q ),
	.prn(vcc));
defparam \output_count[2] .is_wysiwyg = "true";
defparam \output_count[2] .power_up = "low";

dffeas \output_count[3] (
	.clk(clk),
	.d(\output_count[3]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\output_sample_counter~0_combout ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\output_count[3]~q ),
	.prn(vcc));
defparam \output_count[3] .is_wysiwyg = "true";
defparam \output_count[3] .power_up = "low";

dffeas \output_count[0] (
	.clk(clk),
	.d(\output_count[0]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\output_sample_counter~0_combout ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\output_count[0]~q ),
	.prn(vcc));
defparam \output_count[0] .is_wysiwyg = "true";
defparam \output_count[0] .power_up = "low";

dffeas \output_count[4] (
	.clk(clk),
	.d(\output_count[4]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\output_sample_counter~0_combout ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\output_count[4]~q ),
	.prn(vcc));
defparam \output_count[4] .is_wysiwyg = "true";
defparam \output_count[4] .power_up = "low";

dffeas \output_count[5] (
	.clk(clk),
	.d(\output_count[5]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\output_sample_counter~0_combout ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\output_count[5]~q ),
	.prn(vcc));
defparam \output_count[5] .is_wysiwyg = "true";
defparam \output_count[5] .power_up = "low";

dffeas \output_count[6] (
	.clk(clk),
	.d(\output_count[6]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\output_sample_counter~0_combout ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\output_count[6]~q ),
	.prn(vcc));
defparam \output_count[6] .is_wysiwyg = "true";
defparam \output_count[6] .power_up = "low";

dffeas \output_count[7] (
	.clk(clk),
	.d(\output_count[7]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\output_sample_counter~0_combout ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\output_count[7]~q ),
	.prn(vcc));
defparam \output_count[7] .is_wysiwyg = "true";
defparam \output_count[7] .power_up = "low";

dffeas \fft_s1_cur.EARLY_DONE (
	.clk(clk),
	.d(\Selector7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_s1_cur.EARLY_DONE~q ),
	.prn(vcc));
defparam \fft_s1_cur.EARLY_DONE .is_wysiwyg = "true";
defparam \fft_s1_cur.EARLY_DONE .power_up = "low";

dffeas \fft_s1_cur.DONE_WRITING (
	.clk(clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_s1_cur.DONE_WRITING~q ),
	.prn(vcc));
defparam \fft_s1_cur.DONE_WRITING .is_wysiwyg = "true";
defparam \fft_s1_cur.DONE_WRITING .power_up = "low";

cycloneive_lcell_comb \output_count[0]~8 (
	.dataa(\output_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\output_count[0]~8_combout ),
	.cout(\output_count[0]~9 ));
defparam \output_count[0]~8 .lut_mask = 16'h55AA;
defparam \output_count[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \output_count[1]~10 (
	.dataa(\output_count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_count[0]~9 ),
	.combout(\output_count[1]~10_combout ),
	.cout(\output_count[1]~11 ));
defparam \output_count[1]~10 .lut_mask = 16'h5A5F;
defparam \output_count[1]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_count[2]~12 (
	.dataa(\output_count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_count[1]~11 ),
	.combout(\output_count[2]~12_combout ),
	.cout(\output_count[2]~13 ));
defparam \output_count[2]~12 .lut_mask = 16'h5AAF;
defparam \output_count[2]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_count[3]~14 (
	.dataa(\output_count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_count[2]~13 ),
	.combout(\output_count[3]~14_combout ),
	.cout(\output_count[3]~15 ));
defparam \output_count[3]~14 .lut_mask = 16'h5A5F;
defparam \output_count[3]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_count[4]~16 (
	.dataa(\output_count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_count[3]~15 ),
	.combout(\output_count[4]~16_combout ),
	.cout(\output_count[4]~17 ));
defparam \output_count[4]~16 .lut_mask = 16'h5AAF;
defparam \output_count[4]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_count[5]~18 (
	.dataa(\output_count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_count[4]~17 ),
	.combout(\output_count[5]~18_combout ),
	.cout(\output_count[5]~19 ));
defparam \output_count[5]~18 .lut_mask = 16'h5A5F;
defparam \output_count[5]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_count[6]~20 (
	.dataa(\output_count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_count[5]~19 ),
	.combout(\output_count[6]~20_combout ),
	.cout(\output_count[6]~21 ));
defparam \output_count[6]~20 .lut_mask = 16'h5AAF;
defparam \output_count[6]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_count[7]~22 (
	.dataa(\output_count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\output_count[6]~21 ),
	.combout(\output_count[7]~22_combout ),
	.cout());
defparam \output_count[7]~22 .lut_mask = 16'h5A5A;
defparam \output_count[7]~22 .sum_lutc_input = "cin";

dffeas \del_sop_cnt[0] (
	.clk(clk),
	.d(\del_sop_cnt[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\fft_s2_cur.START_LPP~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\del_sop_cnt[0]~q ),
	.prn(vcc));
defparam \del_sop_cnt[0] .is_wysiwyg = "true";
defparam \del_sop_cnt[0] .power_up = "low";

dffeas \del_sop_cnt[1] (
	.clk(clk),
	.d(\del_sop_cnt[1]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\fft_s2_cur.START_LPP~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\del_sop_cnt[1]~q ),
	.prn(vcc));
defparam \del_sop_cnt[1] .is_wysiwyg = "true";
defparam \del_sop_cnt[1] .power_up = "low";

dffeas \del_sop_cnt[2] (
	.clk(clk),
	.d(\del_sop_cnt[2]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\fft_s2_cur.START_LPP~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\del_sop_cnt[2]~q ),
	.prn(vcc));
defparam \del_sop_cnt[2] .is_wysiwyg = "true";
defparam \del_sop_cnt[2] .power_up = "low";

dffeas \del_sop_cnt[4] (
	.clk(clk),
	.d(\del_sop_cnt[4]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\fft_s2_cur.START_LPP~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\del_sop_cnt[4]~q ),
	.prn(vcc));
defparam \del_sop_cnt[4] .is_wysiwyg = "true";
defparam \del_sop_cnt[4] .power_up = "low";

dffeas \del_sop_cnt[3] (
	.clk(clk),
	.d(\del_sop_cnt[3]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\fft_s2_cur.START_LPP~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\del_sop_cnt[3]~q ),
	.prn(vcc));
defparam \del_sop_cnt[3] .is_wysiwyg = "true";
defparam \del_sop_cnt[3] .power_up = "low";

dffeas \core_imag_in[0] (
	.clk(clk),
	.d(\core_imag_in~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[0]~q ),
	.prn(vcc));
defparam \core_imag_in[0] .is_wysiwyg = "true";
defparam \core_imag_in[0] .power_up = "low";

dffeas \core_real_in[0] (
	.clk(clk),
	.d(\core_real_in~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[0]~q ),
	.prn(vcc));
defparam \core_real_in[0] .is_wysiwyg = "true";
defparam \core_real_in[0] .power_up = "low";

dffeas \core_imag_in[1] (
	.clk(clk),
	.d(\core_imag_in~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[1]~q ),
	.prn(vcc));
defparam \core_imag_in[1] .is_wysiwyg = "true";
defparam \core_imag_in[1] .power_up = "low";

dffeas \core_real_in[1] (
	.clk(clk),
	.d(\core_real_in~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[1]~q ),
	.prn(vcc));
defparam \core_real_in[1] .is_wysiwyg = "true";
defparam \core_real_in[1] .power_up = "low";

dffeas \core_imag_in[2] (
	.clk(clk),
	.d(\core_imag_in~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[2]~q ),
	.prn(vcc));
defparam \core_imag_in[2] .is_wysiwyg = "true";
defparam \core_imag_in[2] .power_up = "low";

dffeas \core_real_in[2] (
	.clk(clk),
	.d(\core_real_in~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[2]~q ),
	.prn(vcc));
defparam \core_real_in[2] .is_wysiwyg = "true";
defparam \core_real_in[2] .power_up = "low";

dffeas \core_imag_in[3] (
	.clk(clk),
	.d(\core_imag_in~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[3]~q ),
	.prn(vcc));
defparam \core_imag_in[3] .is_wysiwyg = "true";
defparam \core_imag_in[3] .power_up = "low";

dffeas \core_real_in[3] (
	.clk(clk),
	.d(\core_real_in~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[3]~q ),
	.prn(vcc));
defparam \core_real_in[3] .is_wysiwyg = "true";
defparam \core_real_in[3] .power_up = "low";

dffeas \core_imag_in[4] (
	.clk(clk),
	.d(\core_imag_in~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[4]~q ),
	.prn(vcc));
defparam \core_imag_in[4] .is_wysiwyg = "true";
defparam \core_imag_in[4] .power_up = "low";

dffeas \core_real_in[4] (
	.clk(clk),
	.d(\core_real_in~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[4]~q ),
	.prn(vcc));
defparam \core_real_in[4] .is_wysiwyg = "true";
defparam \core_real_in[4] .power_up = "low";

dffeas \core_imag_in[5] (
	.clk(clk),
	.d(\core_imag_in~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[5]~q ),
	.prn(vcc));
defparam \core_imag_in[5] .is_wysiwyg = "true";
defparam \core_imag_in[5] .power_up = "low";

dffeas \core_real_in[5] (
	.clk(clk),
	.d(\core_real_in~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[5]~q ),
	.prn(vcc));
defparam \core_real_in[5] .is_wysiwyg = "true";
defparam \core_real_in[5] .power_up = "low";

dffeas \core_imag_in[6] (
	.clk(clk),
	.d(\core_imag_in~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[6]~q ),
	.prn(vcc));
defparam \core_imag_in[6] .is_wysiwyg = "true";
defparam \core_imag_in[6] .power_up = "low";

dffeas \core_real_in[6] (
	.clk(clk),
	.d(\core_real_in~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[6]~q ),
	.prn(vcc));
defparam \core_real_in[6] .is_wysiwyg = "true";
defparam \core_real_in[6] .power_up = "low";

dffeas \core_imag_in[7] (
	.clk(clk),
	.d(\core_imag_in~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[7]~q ),
	.prn(vcc));
defparam \core_imag_in[7] .is_wysiwyg = "true";
defparam \core_imag_in[7] .power_up = "low";

dffeas \core_real_in[7] (
	.clk(clk),
	.d(\core_real_in~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[7]~q ),
	.prn(vcc));
defparam \core_real_in[7] .is_wysiwyg = "true";
defparam \core_real_in[7] .power_up = "low";

dffeas \core_imag_in[8] (
	.clk(clk),
	.d(\core_imag_in~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[8]~q ),
	.prn(vcc));
defparam \core_imag_in[8] .is_wysiwyg = "true";
defparam \core_imag_in[8] .power_up = "low";

dffeas \core_real_in[8] (
	.clk(clk),
	.d(\core_real_in~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[8]~q ),
	.prn(vcc));
defparam \core_real_in[8] .is_wysiwyg = "true";
defparam \core_real_in[8] .power_up = "low";

dffeas \core_imag_in[9] (
	.clk(clk),
	.d(\core_imag_in~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[9]~q ),
	.prn(vcc));
defparam \core_imag_in[9] .is_wysiwyg = "true";
defparam \core_imag_in[9] .power_up = "low";

dffeas \core_real_in[9] (
	.clk(clk),
	.d(\core_real_in~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[9]~q ),
	.prn(vcc));
defparam \core_real_in[9] .is_wysiwyg = "true";
defparam \core_real_in[9] .power_up = "low";

dffeas \core_imag_in[10] (
	.clk(clk),
	.d(\core_imag_in~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[10]~q ),
	.prn(vcc));
defparam \core_imag_in[10] .is_wysiwyg = "true";
defparam \core_imag_in[10] .power_up = "low";

dffeas \core_real_in[10] (
	.clk(clk),
	.d(\core_real_in~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[10]~q ),
	.prn(vcc));
defparam \core_real_in[10] .is_wysiwyg = "true";
defparam \core_real_in[10] .power_up = "low";

dffeas \core_imag_in[11] (
	.clk(clk),
	.d(\core_imag_in~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[11]~q ),
	.prn(vcc));
defparam \core_imag_in[11] .is_wysiwyg = "true";
defparam \core_imag_in[11] .power_up = "low";

dffeas \core_real_in[11] (
	.clk(clk),
	.d(\core_real_in~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[11]~q ),
	.prn(vcc));
defparam \core_real_in[11] .is_wysiwyg = "true";
defparam \core_real_in[11] .power_up = "low";

dffeas \core_imag_in[12] (
	.clk(clk),
	.d(\core_imag_in~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[12]~q ),
	.prn(vcc));
defparam \core_imag_in[12] .is_wysiwyg = "true";
defparam \core_imag_in[12] .power_up = "low";

dffeas \core_real_in[12] (
	.clk(clk),
	.d(\core_real_in~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[12]~q ),
	.prn(vcc));
defparam \core_real_in[12] .is_wysiwyg = "true";
defparam \core_real_in[12] .power_up = "low";

dffeas \core_imag_in[13] (
	.clk(clk),
	.d(\core_imag_in~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[13]~q ),
	.prn(vcc));
defparam \core_imag_in[13] .is_wysiwyg = "true";
defparam \core_imag_in[13] .power_up = "low";

dffeas \core_real_in[13] (
	.clk(clk),
	.d(\core_real_in~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[13]~q ),
	.prn(vcc));
defparam \core_real_in[13] .is_wysiwyg = "true";
defparam \core_real_in[13] .power_up = "low";

dffeas \core_imag_in[14] (
	.clk(clk),
	.d(\core_imag_in~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[14]~q ),
	.prn(vcc));
defparam \core_imag_in[14] .is_wysiwyg = "true";
defparam \core_imag_in[14] .power_up = "low";

dffeas \core_real_in[14] (
	.clk(clk),
	.d(\core_real_in~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[14]~q ),
	.prn(vcc));
defparam \core_real_in[14] .is_wysiwyg = "true";
defparam \core_real_in[14] .power_up = "low";

dffeas \core_imag_in[15] (
	.clk(clk),
	.d(\core_imag_in~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_imag_in[15]~q ),
	.prn(vcc));
defparam \core_imag_in[15] .is_wysiwyg = "true";
defparam \core_imag_in[15] .power_up = "low";

dffeas \core_real_in[15] (
	.clk(clk),
	.d(\core_real_in~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\core_real_in[15]~q ),
	.prn(vcc));
defparam \core_real_in[15] .is_wysiwyg = "true";
defparam \core_real_in[15] .power_up = "low";

cycloneive_lcell_comb \del_sop_cnt[0]~5 (
	.dataa(\del_sop_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\del_sop_cnt[0]~5_combout ),
	.cout(\del_sop_cnt[0]~6 ));
defparam \del_sop_cnt[0]~5 .lut_mask = 16'h55AA;
defparam \del_sop_cnt[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \del_sop_cnt[1]~7 (
	.dataa(\del_sop_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_sop_cnt[0]~6 ),
	.combout(\del_sop_cnt[1]~7_combout ),
	.cout(\del_sop_cnt[1]~8 ));
defparam \del_sop_cnt[1]~7 .lut_mask = 16'h5A5F;
defparam \del_sop_cnt[1]~7 .sum_lutc_input = "cin";

cycloneive_lcell_comb \del_sop_cnt[2]~9 (
	.dataa(\del_sop_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_sop_cnt[1]~8 ),
	.combout(\del_sop_cnt[2]~9_combout ),
	.cout(\del_sop_cnt[2]~10 ));
defparam \del_sop_cnt[2]~9 .lut_mask = 16'h5AAF;
defparam \del_sop_cnt[2]~9 .sum_lutc_input = "cin";

cycloneive_lcell_comb \del_sop_cnt[3]~11 (
	.dataa(\del_sop_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_sop_cnt[2]~10 ),
	.combout(\del_sop_cnt[3]~11_combout ),
	.cout(\del_sop_cnt[3]~12 ));
defparam \del_sop_cnt[3]~11 .lut_mask = 16'h5A5F;
defparam \del_sop_cnt[3]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \del_sop_cnt[4]~13 (
	.dataa(\del_sop_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\del_sop_cnt[3]~12 ),
	.combout(\del_sop_cnt[4]~13_combout ),
	.cout());
defparam \del_sop_cnt[4]~13 .lut_mask = 16'h5A5A;
defparam \del_sop_cnt[4]~13 .sum_lutc_input = "cin";

dffeas \k_count_wr[2] (
	.clk(clk),
	.d(\k_count_wr[2]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_count_wr_en~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_wr[2]~q ),
	.prn(vcc));
defparam \k_count_wr[2] .is_wysiwyg = "true";
defparam \k_count_wr[2] .power_up = "low";

dffeas \k_count_wr[0] (
	.clk(clk),
	.d(\k_count_wr[0]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_count_wr_en~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_wr[0]~q ),
	.prn(vcc));
defparam \k_count_wr[0] .is_wysiwyg = "true";
defparam \k_count_wr[0] .power_up = "low";

dffeas \k_count_wr[6] (
	.clk(clk),
	.d(\k_count_wr[6]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_count_wr_en~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_wr[6]~q ),
	.prn(vcc));
defparam \k_count_wr[6] .is_wysiwyg = "true";
defparam \k_count_wr[6] .power_up = "low";

dffeas \k_count_wr[3] (
	.clk(clk),
	.d(\k_count_wr[3]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_count_wr_en~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_wr[3]~q ),
	.prn(vcc));
defparam \k_count_wr[3] .is_wysiwyg = "true";
defparam \k_count_wr[3] .power_up = "low";

dffeas \k_count_wr[1] (
	.clk(clk),
	.d(\k_count_wr[1]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_count_wr_en~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_wr[1]~q ),
	.prn(vcc));
defparam \k_count_wr[1] .is_wysiwyg = "true";
defparam \k_count_wr[1] .power_up = "low";

dffeas \k_count_wr[7] (
	.clk(clk),
	.d(\k_count_wr[7]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_count_wr_en~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_wr[7]~q ),
	.prn(vcc));
defparam \k_count_wr[7] .is_wysiwyg = "true";
defparam \k_count_wr[7] .power_up = "low";

dffeas \k_count_wr[4] (
	.clk(clk),
	.d(\k_count_wr[4]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_count_wr_en~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_wr[4]~q ),
	.prn(vcc));
defparam \k_count_wr[4] .is_wysiwyg = "true";
defparam \k_count_wr[4] .power_up = "low";

dffeas \k_count_wr[5] (
	.clk(clk),
	.d(\k_count_wr[5]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_count_wr_en~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_wr[5]~q ),
	.prn(vcc));
defparam \k_count_wr[5] .is_wysiwyg = "true";
defparam \k_count_wr[5] .power_up = "low";

cycloneive_lcell_comb \k_count_wr[0]~8 (
	.dataa(\k_count_wr[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\k_count_wr[0]~8_combout ),
	.cout(\k_count_wr[0]~9 ));
defparam \k_count_wr[0]~8 .lut_mask = 16'h55AA;
defparam \k_count_wr[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \k_count_wr[1]~10 (
	.dataa(\k_count_wr[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k_count_wr[0]~9 ),
	.combout(\k_count_wr[1]~10_combout ),
	.cout(\k_count_wr[1]~11 ));
defparam \k_count_wr[1]~10 .lut_mask = 16'h5A5F;
defparam \k_count_wr[1]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \k_count_wr[2]~12 (
	.dataa(\k_count_wr[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k_count_wr[1]~11 ),
	.combout(\k_count_wr[2]~12_combout ),
	.cout(\k_count_wr[2]~13 ));
defparam \k_count_wr[2]~12 .lut_mask = 16'h5AAF;
defparam \k_count_wr[2]~12 .sum_lutc_input = "cin";

dffeas k_count_wr_en(
	.clk(clk),
	.d(\k_count_wr_en~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_wr_en~q ),
	.prn(vcc));
defparam k_count_wr_en.is_wysiwyg = "true";
defparam k_count_wr_en.power_up = "low";

cycloneive_lcell_comb \k_count_wr[3]~14 (
	.dataa(\k_count_wr[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k_count_wr[2]~13 ),
	.combout(\k_count_wr[3]~14_combout ),
	.cout(\k_count_wr[3]~15 ));
defparam \k_count_wr[3]~14 .lut_mask = 16'h5A5F;
defparam \k_count_wr[3]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \k_count_wr[4]~16 (
	.dataa(\k_count_wr[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k_count_wr[3]~15 ),
	.combout(\k_count_wr[4]~16_combout ),
	.cout(\k_count_wr[4]~17 ));
defparam \k_count_wr[4]~16 .lut_mask = 16'h5AAF;
defparam \k_count_wr[4]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \k_count_wr[5]~18 (
	.dataa(\k_count_wr[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k_count_wr[4]~17 ),
	.combout(\k_count_wr[5]~18_combout ),
	.cout(\k_count_wr[5]~19 ));
defparam \k_count_wr[5]~18 .lut_mask = 16'h5A5F;
defparam \k_count_wr[5]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \k_count_wr[6]~20 (
	.dataa(\k_count_wr[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k_count_wr[5]~19 ),
	.combout(\k_count_wr[6]~20_combout ),
	.cout(\k_count_wr[6]~21 ));
defparam \k_count_wr[6]~20 .lut_mask = 16'h5AAF;
defparam \k_count_wr[6]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \k_count_wr[7]~22 (
	.dataa(\k_count_wr[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\k_count_wr[6]~21 ),
	.combout(\k_count_wr[7]~22_combout ),
	.cout());
defparam \k_count_wr[7]~22 .lut_mask = 16'h5A5A;
defparam \k_count_wr[7]~22 .sum_lutc_input = "cin";

dffeas \twiddle_data_real[0] (
	.clk(clk),
	.d(\Mux15~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_real[0]~q ),
	.prn(vcc));
defparam \twiddle_data_real[0] .is_wysiwyg = "true";
defparam \twiddle_data_real[0] .power_up = "low";

dffeas \twiddle_data_real[15] (
	.clk(clk),
	.d(\Mux0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_real[15]~q ),
	.prn(vcc));
defparam \twiddle_data_real[15] .is_wysiwyg = "true";
defparam \twiddle_data_real[15] .power_up = "low";

dffeas \twiddle_data_imag[1] (
	.clk(clk),
	.d(\twiddle_data_imag[1]~0_combout ),
	.asdata(\Add3~2_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\twiddle_data_imag[14]~15_combout ),
	.sload(\quad_del_1[2]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_imag[1]~q ),
	.prn(vcc));
defparam \twiddle_data_imag[1] .is_wysiwyg = "true";
defparam \twiddle_data_imag[1] .power_up = "low";

dffeas \twiddle_data_imag[2] (
	.clk(clk),
	.d(\twiddle_data_imag[2]~1_combout ),
	.asdata(\Add3~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\twiddle_data_imag[14]~15_combout ),
	.sload(\quad_del_1[2]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_imag[2]~q ),
	.prn(vcc));
defparam \twiddle_data_imag[2] .is_wysiwyg = "true";
defparam \twiddle_data_imag[2] .power_up = "low";

dffeas \twiddle_data_imag[3] (
	.clk(clk),
	.d(\twiddle_data_imag[3]~2_combout ),
	.asdata(\Add3~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\twiddle_data_imag[14]~15_combout ),
	.sload(\quad_del_1[2]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_imag[3]~q ),
	.prn(vcc));
defparam \twiddle_data_imag[3] .is_wysiwyg = "true";
defparam \twiddle_data_imag[3] .power_up = "low";

dffeas \twiddle_data_imag[4] (
	.clk(clk),
	.d(\twiddle_data_imag[4]~3_combout ),
	.asdata(\Add3~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\twiddle_data_imag[14]~15_combout ),
	.sload(\quad_del_1[2]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_imag[4]~q ),
	.prn(vcc));
defparam \twiddle_data_imag[4] .is_wysiwyg = "true";
defparam \twiddle_data_imag[4] .power_up = "low";

dffeas \twiddle_data_imag[5] (
	.clk(clk),
	.d(\twiddle_data_imag[5]~4_combout ),
	.asdata(\Add3~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\twiddle_data_imag[14]~15_combout ),
	.sload(\quad_del_1[2]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_imag[5]~q ),
	.prn(vcc));
defparam \twiddle_data_imag[5] .is_wysiwyg = "true";
defparam \twiddle_data_imag[5] .power_up = "low";

dffeas \twiddle_data_imag[6] (
	.clk(clk),
	.d(\twiddle_data_imag[6]~5_combout ),
	.asdata(\Add3~12_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\twiddle_data_imag[14]~15_combout ),
	.sload(\quad_del_1[2]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_imag[6]~q ),
	.prn(vcc));
defparam \twiddle_data_imag[6] .is_wysiwyg = "true";
defparam \twiddle_data_imag[6] .power_up = "low";

dffeas \twiddle_data_imag[7] (
	.clk(clk),
	.d(\twiddle_data_imag[7]~6_combout ),
	.asdata(\Add3~14_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\twiddle_data_imag[14]~15_combout ),
	.sload(\quad_del_1[2]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_imag[7]~q ),
	.prn(vcc));
defparam \twiddle_data_imag[7] .is_wysiwyg = "true";
defparam \twiddle_data_imag[7] .power_up = "low";

dffeas \twiddle_data_imag[8] (
	.clk(clk),
	.d(\twiddle_data_imag[8]~7_combout ),
	.asdata(\Add3~16_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\twiddle_data_imag[14]~15_combout ),
	.sload(\quad_del_1[2]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_imag[8]~q ),
	.prn(vcc));
defparam \twiddle_data_imag[8] .is_wysiwyg = "true";
defparam \twiddle_data_imag[8] .power_up = "low";

dffeas \twiddle_data_imag[9] (
	.clk(clk),
	.d(\twiddle_data_imag[9]~8_combout ),
	.asdata(\Add3~18_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\twiddle_data_imag[14]~15_combout ),
	.sload(\quad_del_1[2]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_imag[9]~q ),
	.prn(vcc));
defparam \twiddle_data_imag[9] .is_wysiwyg = "true";
defparam \twiddle_data_imag[9] .power_up = "low";

dffeas \twiddle_data_imag[10] (
	.clk(clk),
	.d(\twiddle_data_imag[10]~9_combout ),
	.asdata(\Add3~20_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\twiddle_data_imag[14]~15_combout ),
	.sload(\quad_del_1[2]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_imag[10]~q ),
	.prn(vcc));
defparam \twiddle_data_imag[10] .is_wysiwyg = "true";
defparam \twiddle_data_imag[10] .power_up = "low";

dffeas \twiddle_data_imag[11] (
	.clk(clk),
	.d(\twiddle_data_imag[11]~10_combout ),
	.asdata(\Add3~22_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\twiddle_data_imag[14]~15_combout ),
	.sload(\quad_del_1[2]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_imag[11]~q ),
	.prn(vcc));
defparam \twiddle_data_imag[11] .is_wysiwyg = "true";
defparam \twiddle_data_imag[11] .power_up = "low";

dffeas \twiddle_data_imag[12] (
	.clk(clk),
	.d(\twiddle_data_imag[12]~11_combout ),
	.asdata(\Add3~24_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\twiddle_data_imag[14]~15_combout ),
	.sload(\quad_del_1[2]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_imag[12]~q ),
	.prn(vcc));
defparam \twiddle_data_imag[12] .is_wysiwyg = "true";
defparam \twiddle_data_imag[12] .power_up = "low";

dffeas \twiddle_data_imag[13] (
	.clk(clk),
	.d(\twiddle_data_imag[13]~12_combout ),
	.asdata(\Add3~26_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\twiddle_data_imag[14]~15_combout ),
	.sload(\quad_del_1[2]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_imag[13]~q ),
	.prn(vcc));
defparam \twiddle_data_imag[13] .is_wysiwyg = "true";
defparam \twiddle_data_imag[13] .power_up = "low";

dffeas \twiddle_data_imag[14] (
	.clk(clk),
	.d(\twiddle_data_imag[14]~13_combout ),
	.asdata(\Add3~28_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\twiddle_data_imag[14]~15_combout ),
	.sload(\quad_del_1[2]~q ),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_imag[14]~q ),
	.prn(vcc));
defparam \twiddle_data_imag[14] .is_wysiwyg = "true";
defparam \twiddle_data_imag[14] .power_up = "low";

dffeas \twiddle_data_imag[15] (
	.clk(clk),
	.d(\Mux16~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_imag[15]~q ),
	.prn(vcc));
defparam \twiddle_data_imag[15] .is_wysiwyg = "true";
defparam \twiddle_data_imag[15] .power_up = "low";

cycloneive_lcell_comb \Add2~1 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[0] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\Add2~1_cout ));
defparam \Add2~1 .lut_mask = 16'h0055;
defparam \Add2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add2~2 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[1] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~1_cout ),
	.combout(\Add2~2_combout ),
	.cout(\Add2~3 ));
defparam \Add2~2 .lut_mask = 16'h5AAF;
defparam \Add2~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~4 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[2] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~3 ),
	.combout(\Add2~4_combout ),
	.cout(\Add2~5 ));
defparam \Add2~4 .lut_mask = 16'h5A5F;
defparam \Add2~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~6 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[3] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~5 ),
	.combout(\Add2~6_combout ),
	.cout(\Add2~7 ));
defparam \Add2~6 .lut_mask = 16'h5AAF;
defparam \Add2~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~8 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[4] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~7 ),
	.combout(\Add2~8_combout ),
	.cout(\Add2~9 ));
defparam \Add2~8 .lut_mask = 16'h5A5F;
defparam \Add2~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~10 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[5] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~9 ),
	.combout(\Add2~10_combout ),
	.cout(\Add2~11 ));
defparam \Add2~10 .lut_mask = 16'h5AAF;
defparam \Add2~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~12 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[6] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~11 ),
	.combout(\Add2~12_combout ),
	.cout(\Add2~13 ));
defparam \Add2~12 .lut_mask = 16'h5A5F;
defparam \Add2~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~14 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[7] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~13 ),
	.combout(\Add2~14_combout ),
	.cout(\Add2~15 ));
defparam \Add2~14 .lut_mask = 16'h5AAF;
defparam \Add2~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~16 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[8] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~15 ),
	.combout(\Add2~16_combout ),
	.cout(\Add2~17 ));
defparam \Add2~16 .lut_mask = 16'h5A5F;
defparam \Add2~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~18 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[9] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~17 ),
	.combout(\Add2~18_combout ),
	.cout(\Add2~19 ));
defparam \Add2~18 .lut_mask = 16'h5AAF;
defparam \Add2~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~20 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[10] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~19 ),
	.combout(\Add2~20_combout ),
	.cout(\Add2~21 ));
defparam \Add2~20 .lut_mask = 16'h5A5F;
defparam \Add2~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~22 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[11] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~21 ),
	.combout(\Add2~22_combout ),
	.cout(\Add2~23 ));
defparam \Add2~22 .lut_mask = 16'h5AAF;
defparam \Add2~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~24 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[12] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~23 ),
	.combout(\Add2~24_combout ),
	.cout(\Add2~25 ));
defparam \Add2~24 .lut_mask = 16'h5A5F;
defparam \Add2~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~26 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[13] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~25 ),
	.combout(\Add2~26_combout ),
	.cout(\Add2~27 ));
defparam \Add2~26 .lut_mask = 16'h5AAF;
defparam \Add2~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~28 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[14] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~27 ),
	.combout(\Add2~28_combout ),
	.cout(\Add2~29 ));
defparam \Add2~28 .lut_mask = 16'h5A5F;
defparam \Add2~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~30 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[15] ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add2~29 ),
	.combout(\Add2~30_combout ),
	.cout());
defparam \Add2~30 .lut_mask = 16'h5A5A;
defparam \Add2~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twiddle_data_imag[1]~0 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[1] ),
	.datab(\quad_del_1[1]~q ),
	.datac(gnd),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_imag[1]~0_combout ),
	.cout());
defparam \twiddle_data_imag[1]~0 .lut_mask = 16'hAACC;
defparam \twiddle_data_imag[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~1 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[0] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\Add3~1_cout ));
defparam \Add3~1 .lut_mask = 16'h0055;
defparam \Add3~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~2 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[1] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~1_cout ),
	.combout(\Add3~2_combout ),
	.cout(\Add3~3 ));
defparam \Add3~2 .lut_mask = 16'h5AAF;
defparam \Add3~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twiddle_data_imag[2]~1 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[2] ),
	.datab(\quad_del_1[1]~q ),
	.datac(gnd),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_imag[2]~1_combout ),
	.cout());
defparam \twiddle_data_imag[2]~1 .lut_mask = 16'hAACC;
defparam \twiddle_data_imag[2]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~4 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[2] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~3 ),
	.combout(\Add3~4_combout ),
	.cout(\Add3~5 ));
defparam \Add3~4 .lut_mask = 16'h5A5F;
defparam \Add3~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twiddle_data_imag[3]~2 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[3] ),
	.datab(\quad_del_1[1]~q ),
	.datac(gnd),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_imag[3]~2_combout ),
	.cout());
defparam \twiddle_data_imag[3]~2 .lut_mask = 16'hAACC;
defparam \twiddle_data_imag[3]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~6 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[3] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~5 ),
	.combout(\Add3~6_combout ),
	.cout(\Add3~7 ));
defparam \Add3~6 .lut_mask = 16'h5AAF;
defparam \Add3~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twiddle_data_imag[4]~3 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[4] ),
	.datab(\quad_del_1[1]~q ),
	.datac(gnd),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_imag[4]~3_combout ),
	.cout());
defparam \twiddle_data_imag[4]~3 .lut_mask = 16'hAACC;
defparam \twiddle_data_imag[4]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~8 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[4] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~7 ),
	.combout(\Add3~8_combout ),
	.cout(\Add3~9 ));
defparam \Add3~8 .lut_mask = 16'h5A5F;
defparam \Add3~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twiddle_data_imag[5]~4 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[5] ),
	.datab(\quad_del_1[1]~q ),
	.datac(gnd),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_imag[5]~4_combout ),
	.cout());
defparam \twiddle_data_imag[5]~4 .lut_mask = 16'hAACC;
defparam \twiddle_data_imag[5]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~10 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[5] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~9 ),
	.combout(\Add3~10_combout ),
	.cout(\Add3~11 ));
defparam \Add3~10 .lut_mask = 16'h5AAF;
defparam \Add3~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twiddle_data_imag[6]~5 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[6] ),
	.datab(\quad_del_1[1]~q ),
	.datac(gnd),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_imag[6]~5_combout ),
	.cout());
defparam \twiddle_data_imag[6]~5 .lut_mask = 16'hAACC;
defparam \twiddle_data_imag[6]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~12 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[6] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~11 ),
	.combout(\Add3~12_combout ),
	.cout(\Add3~13 ));
defparam \Add3~12 .lut_mask = 16'h5A5F;
defparam \Add3~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twiddle_data_imag[7]~6 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[7] ),
	.datab(\quad_del_1[1]~q ),
	.datac(gnd),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_imag[7]~6_combout ),
	.cout());
defparam \twiddle_data_imag[7]~6 .lut_mask = 16'hAACC;
defparam \twiddle_data_imag[7]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~14 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[7] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~13 ),
	.combout(\Add3~14_combout ),
	.cout(\Add3~15 ));
defparam \Add3~14 .lut_mask = 16'h5AAF;
defparam \Add3~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twiddle_data_imag[8]~7 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[8] ),
	.datab(\quad_del_1[1]~q ),
	.datac(gnd),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_imag[8]~7_combout ),
	.cout());
defparam \twiddle_data_imag[8]~7 .lut_mask = 16'hAACC;
defparam \twiddle_data_imag[8]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~16 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[8] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~15 ),
	.combout(\Add3~16_combout ),
	.cout(\Add3~17 ));
defparam \Add3~16 .lut_mask = 16'h5A5F;
defparam \Add3~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twiddle_data_imag[9]~8 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[9] ),
	.datab(\quad_del_1[1]~q ),
	.datac(gnd),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_imag[9]~8_combout ),
	.cout());
defparam \twiddle_data_imag[9]~8 .lut_mask = 16'hAACC;
defparam \twiddle_data_imag[9]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~18 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[9] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~17 ),
	.combout(\Add3~18_combout ),
	.cout(\Add3~19 ));
defparam \Add3~18 .lut_mask = 16'h5AAF;
defparam \Add3~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twiddle_data_imag[10]~9 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[10] ),
	.datab(\quad_del_1[1]~q ),
	.datac(gnd),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_imag[10]~9_combout ),
	.cout());
defparam \twiddle_data_imag[10]~9 .lut_mask = 16'hAACC;
defparam \twiddle_data_imag[10]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~20 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[10] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~19 ),
	.combout(\Add3~20_combout ),
	.cout(\Add3~21 ));
defparam \Add3~20 .lut_mask = 16'h5A5F;
defparam \Add3~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twiddle_data_imag[11]~10 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[11] ),
	.datab(\quad_del_1[1]~q ),
	.datac(gnd),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_imag[11]~10_combout ),
	.cout());
defparam \twiddle_data_imag[11]~10 .lut_mask = 16'hAACC;
defparam \twiddle_data_imag[11]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~22 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[11] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~21 ),
	.combout(\Add3~22_combout ),
	.cout(\Add3~23 ));
defparam \Add3~22 .lut_mask = 16'h5AAF;
defparam \Add3~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twiddle_data_imag[12]~11 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[12] ),
	.datab(\quad_del_1[1]~q ),
	.datac(gnd),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_imag[12]~11_combout ),
	.cout());
defparam \twiddle_data_imag[12]~11 .lut_mask = 16'hAACC;
defparam \twiddle_data_imag[12]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~24 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[12] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~23 ),
	.combout(\Add3~24_combout ),
	.cout(\Add3~25 ));
defparam \Add3~24 .lut_mask = 16'h5A5F;
defparam \Add3~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twiddle_data_imag[13]~12 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[13] ),
	.datab(\quad_del_1[1]~q ),
	.datac(gnd),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_imag[13]~12_combout ),
	.cout());
defparam \twiddle_data_imag[13]~12 .lut_mask = 16'hAACC;
defparam \twiddle_data_imag[13]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~26 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[13] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~25 ),
	.combout(\Add3~26_combout ),
	.cout(\Add3~27 ));
defparam \Add3~26 .lut_mask = 16'h5AAF;
defparam \Add3~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twiddle_data_imag[14]~13 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[14] ),
	.datab(\quad_del_1[1]~q ),
	.datac(gnd),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_imag[14]~13_combout ),
	.cout());
defparam \twiddle_data_imag[14]~13 .lut_mask = 16'hAACC;
defparam \twiddle_data_imag[14]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~28 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[14] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~27 ),
	.combout(\Add3~28_combout ),
	.cout(\Add3~29 ));
defparam \Add3~28 .lut_mask = 16'h5A5F;
defparam \Add3~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add3~30 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[15] ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add3~29 ),
	.combout(\Add3~30_combout ),
	.cout());
defparam \Add3~30 .lut_mask = 16'h5A5A;
defparam \Add3~30 .sum_lutc_input = "cin";

dffeas \k_count_tw[0] (
	.clk(clk),
	.d(\k_count_tw[0]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_count_tw_en~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_tw[0]~q ),
	.prn(vcc));
defparam \k_count_tw[0] .is_wysiwyg = "true";
defparam \k_count_tw[0] .power_up = "low";

dffeas \k_count_tw[2] (
	.clk(clk),
	.d(\k_count_tw[2]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_count_tw_en~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_tw[2]~q ),
	.prn(vcc));
defparam \k_count_tw[2] .is_wysiwyg = "true";
defparam \k_count_tw[2] .power_up = "low";

dffeas \k_count_tw[1] (
	.clk(clk),
	.d(\k_count_tw[1]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_count_tw_en~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_tw[1]~q ),
	.prn(vcc));
defparam \k_count_tw[1] .is_wysiwyg = "true";
defparam \k_count_tw[1] .power_up = "low";

dffeas \k_count_tw[3] (
	.clk(clk),
	.d(\k_count_tw[3]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_count_tw_en~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_tw[3]~q ),
	.prn(vcc));
defparam \k_count_tw[3] .is_wysiwyg = "true";
defparam \k_count_tw[3] .power_up = "low";

dffeas \k_count_tw[5] (
	.clk(clk),
	.d(\k_count_tw[5]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_count_tw_en~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_tw[5]~q ),
	.prn(vcc));
defparam \k_count_tw[5] .is_wysiwyg = "true";
defparam \k_count_tw[5] .power_up = "low";

dffeas \k_count_tw[4] (
	.clk(clk),
	.d(\k_count_tw[4]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_count_tw_en~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_tw[4]~q ),
	.prn(vcc));
defparam \k_count_tw[4] .is_wysiwyg = "true";
defparam \k_count_tw[4] .power_up = "low";

dffeas \k_count_tw[7] (
	.clk(clk),
	.d(\k_count_tw[7]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_count_tw_en~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_tw[7]~q ),
	.prn(vcc));
defparam \k_count_tw[7] .is_wysiwyg = "true";
defparam \k_count_tw[7] .power_up = "low";

dffeas \k_count_tw[6] (
	.clk(clk),
	.d(\k_count_tw[6]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_count_tw_en~q ),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_tw[6]~q ),
	.prn(vcc));
defparam \k_count_tw[6] .is_wysiwyg = "true";
defparam \k_count_tw[6] .power_up = "low";

cycloneive_lcell_comb \k_count_tw[0]~8 (
	.dataa(\k_count_tw[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\k_count_tw[0]~8_combout ),
	.cout(\k_count_tw[0]~9 ));
defparam \k_count_tw[0]~8 .lut_mask = 16'h55AA;
defparam \k_count_tw[0]~8 .sum_lutc_input = "datac";

dffeas k_count_tw_en(
	.clk(clk),
	.d(\k_count_tw_en~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\k_count_tw_en~q ),
	.prn(vcc));
defparam k_count_tw_en.is_wysiwyg = "true";
defparam k_count_tw_en.power_up = "low";

cycloneive_lcell_comb \k_count_tw[1]~10 (
	.dataa(\k_count_tw[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k_count_tw[0]~9 ),
	.combout(\k_count_tw[1]~10_combout ),
	.cout(\k_count_tw[1]~11 ));
defparam \k_count_tw[1]~10 .lut_mask = 16'h5A5F;
defparam \k_count_tw[1]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \k_count_tw[2]~12 (
	.dataa(\k_count_tw[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k_count_tw[1]~11 ),
	.combout(\k_count_tw[2]~12_combout ),
	.cout(\k_count_tw[2]~13 ));
defparam \k_count_tw[2]~12 .lut_mask = 16'h5AAF;
defparam \k_count_tw[2]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \k_count_tw[3]~14 (
	.dataa(\k_count_tw[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k_count_tw[2]~13 ),
	.combout(\k_count_tw[3]~14_combout ),
	.cout(\k_count_tw[3]~15 ));
defparam \k_count_tw[3]~14 .lut_mask = 16'h5A5F;
defparam \k_count_tw[3]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \k_count_tw[4]~16 (
	.dataa(\k_count_tw[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k_count_tw[3]~15 ),
	.combout(\k_count_tw[4]~16_combout ),
	.cout(\k_count_tw[4]~17 ));
defparam \k_count_tw[4]~16 .lut_mask = 16'h5AAF;
defparam \k_count_tw[4]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \k_count_tw[5]~18 (
	.dataa(\k_count_tw[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k_count_tw[4]~17 ),
	.combout(\k_count_tw[5]~18_combout ),
	.cout(\k_count_tw[5]~19 ));
defparam \k_count_tw[5]~18 .lut_mask = 16'h5A5F;
defparam \k_count_tw[5]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \k_count_tw[6]~20 (
	.dataa(\k_count_tw[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k_count_tw[5]~19 ),
	.combout(\k_count_tw[6]~20_combout ),
	.cout(\k_count_tw[6]~21 ));
defparam \k_count_tw[6]~20 .lut_mask = 16'h5AAF;
defparam \k_count_tw[6]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \k_count_tw[7]~22 (
	.dataa(\k_count_tw[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\k_count_tw[6]~21 ),
	.combout(\k_count_tw[7]~22_combout ),
	.cout());
defparam \k_count_tw[7]~22 .lut_mask = 16'h5A5A;
defparam \k_count_tw[7]~22 .sum_lutc_input = "cin";

dffeas master_source_ena(
	.clk(clk),
	.d(\master_source_ena~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\master_source_ena~q ),
	.prn(vcc));
defparam master_source_ena.is_wysiwyg = "true";
defparam master_source_ena.power_up = "low";

dffeas sink_ready_ctrl_d(
	.clk(clk),
	.d(\auk_dsp_interface_controller_1|sink_ready_ctrl~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_ready_ctrl_d~q ),
	.prn(vcc));
defparam sink_ready_ctrl_d.is_wysiwyg = "true";
defparam sink_ready_ctrl_d.power_up = "low";

dffeas sop(
	.clk(clk),
	.d(\sop~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sop~q ),
	.prn(vcc));
defparam sop.is_wysiwyg = "true";
defparam sop.power_up = "low";

cycloneive_lcell_comb \source_valid_ctrl_sop~0 (
	.dataa(\auk_dsp_interface_controller_1|sink_stall_reg~q ),
	.datab(\sink_ready_ctrl_d~q ),
	.datac(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datad(\sop~q ),
	.cin(gnd),
	.combout(\source_valid_ctrl_sop~0_combout ),
	.cout());
defparam \source_valid_ctrl_sop~0 .lut_mask = 16'hBFFF;
defparam \source_valid_ctrl_sop~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \source_valid_ctrl_sop~1 (
	.dataa(gnd),
	.datab(\sink_ready_ctrl_d~q ),
	.datac(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datad(\sop~q ),
	.cin(gnd),
	.combout(\source_valid_ctrl_sop~1_combout ),
	.cout());
defparam \source_valid_ctrl_sop~1 .lut_mask = 16'h3FFF;
defparam \source_valid_ctrl_sop~1 .sum_lutc_input = "datac";

dffeas \exponent_out[0] (
	.clk(clk),
	.d(\exponent_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\exponent_out[0]~q ),
	.prn(vcc));
defparam \exponent_out[0] .is_wysiwyg = "true";
defparam \exponent_out[0] .power_up = "low";

dffeas \exponent_out[1] (
	.clk(clk),
	.d(\exponent_out~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\exponent_out[1]~q ),
	.prn(vcc));
defparam \exponent_out[1] .is_wysiwyg = "true";
defparam \exponent_out[1] .power_up = "low";

dffeas \exponent_out[2] (
	.clk(clk),
	.d(\exponent_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\exponent_out[2]~q ),
	.prn(vcc));
defparam \exponent_out[2] .is_wysiwyg = "true";
defparam \exponent_out[2] .power_up = "low";

dffeas \exponent_out[3] (
	.clk(clk),
	.d(\exponent_out~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\exponent_out[3]~q ),
	.prn(vcc));
defparam \exponent_out[3] .is_wysiwyg = "true";
defparam \exponent_out[3] .power_up = "low";

dffeas \exponent_out[4] (
	.clk(clk),
	.d(\exponent_out~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\exponent_out[4]~q ),
	.prn(vcc));
defparam \exponent_out[4] .is_wysiwyg = "true";
defparam \exponent_out[4] .power_up = "low";

dffeas \exponent_out[5] (
	.clk(clk),
	.d(\exponent_out~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\exponent_out[5]~q ),
	.prn(vcc));
defparam \exponent_out[5] .is_wysiwyg = "true";
defparam \exponent_out[5] .power_up = "low";

dffeas \fft_real_out[0] (
	.clk(clk),
	.d(\fft_real_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[0]~q ),
	.prn(vcc));
defparam \fft_real_out[0] .is_wysiwyg = "true";
defparam \fft_real_out[0] .power_up = "low";

dffeas \fft_real_out[1] (
	.clk(clk),
	.d(\fft_real_out~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[1]~q ),
	.prn(vcc));
defparam \fft_real_out[1] .is_wysiwyg = "true";
defparam \fft_real_out[1] .power_up = "low";

dffeas \fft_real_out[2] (
	.clk(clk),
	.d(\fft_real_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[2]~q ),
	.prn(vcc));
defparam \fft_real_out[2] .is_wysiwyg = "true";
defparam \fft_real_out[2] .power_up = "low";

dffeas \fft_real_out[3] (
	.clk(clk),
	.d(\fft_real_out~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[3]~q ),
	.prn(vcc));
defparam \fft_real_out[3] .is_wysiwyg = "true";
defparam \fft_real_out[3] .power_up = "low";

dffeas \fft_real_out[4] (
	.clk(clk),
	.d(\fft_real_out~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[4]~q ),
	.prn(vcc));
defparam \fft_real_out[4] .is_wysiwyg = "true";
defparam \fft_real_out[4] .power_up = "low";

dffeas \fft_real_out[5] (
	.clk(clk),
	.d(\fft_real_out~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[5]~q ),
	.prn(vcc));
defparam \fft_real_out[5] .is_wysiwyg = "true";
defparam \fft_real_out[5] .power_up = "low";

dffeas \fft_real_out[6] (
	.clk(clk),
	.d(\fft_real_out~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[6]~q ),
	.prn(vcc));
defparam \fft_real_out[6] .is_wysiwyg = "true";
defparam \fft_real_out[6] .power_up = "low";

dffeas \fft_real_out[7] (
	.clk(clk),
	.d(\fft_real_out~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[7]~q ),
	.prn(vcc));
defparam \fft_real_out[7] .is_wysiwyg = "true";
defparam \fft_real_out[7] .power_up = "low";

dffeas \fft_real_out[8] (
	.clk(clk),
	.d(\fft_real_out~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[8]~q ),
	.prn(vcc));
defparam \fft_real_out[8] .is_wysiwyg = "true";
defparam \fft_real_out[8] .power_up = "low";

dffeas \fft_real_out[9] (
	.clk(clk),
	.d(\fft_real_out~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[9]~q ),
	.prn(vcc));
defparam \fft_real_out[9] .is_wysiwyg = "true";
defparam \fft_real_out[9] .power_up = "low";

dffeas \fft_real_out[10] (
	.clk(clk),
	.d(\fft_real_out~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[10]~q ),
	.prn(vcc));
defparam \fft_real_out[10] .is_wysiwyg = "true";
defparam \fft_real_out[10] .power_up = "low";

dffeas \fft_real_out[11] (
	.clk(clk),
	.d(\fft_real_out~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[11]~q ),
	.prn(vcc));
defparam \fft_real_out[11] .is_wysiwyg = "true";
defparam \fft_real_out[11] .power_up = "low";

dffeas \fft_real_out[12] (
	.clk(clk),
	.d(\fft_real_out~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[12]~q ),
	.prn(vcc));
defparam \fft_real_out[12] .is_wysiwyg = "true";
defparam \fft_real_out[12] .power_up = "low";

dffeas \fft_real_out[13] (
	.clk(clk),
	.d(\fft_real_out~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[13]~q ),
	.prn(vcc));
defparam \fft_real_out[13] .is_wysiwyg = "true";
defparam \fft_real_out[13] .power_up = "low";

dffeas \fft_real_out[14] (
	.clk(clk),
	.d(\fft_real_out~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[14]~q ),
	.prn(vcc));
defparam \fft_real_out[14] .is_wysiwyg = "true";
defparam \fft_real_out[14] .power_up = "low";

dffeas \fft_real_out[15] (
	.clk(clk),
	.d(\fft_real_out~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_real_out[15]~q ),
	.prn(vcc));
defparam \fft_real_out[15] .is_wysiwyg = "true";
defparam \fft_real_out[15] .power_up = "low";

dffeas \fft_imag_out[0] (
	.clk(clk),
	.d(\fft_imag_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[0]~q ),
	.prn(vcc));
defparam \fft_imag_out[0] .is_wysiwyg = "true";
defparam \fft_imag_out[0] .power_up = "low";

dffeas \fft_imag_out[1] (
	.clk(clk),
	.d(\fft_imag_out~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[1]~q ),
	.prn(vcc));
defparam \fft_imag_out[1] .is_wysiwyg = "true";
defparam \fft_imag_out[1] .power_up = "low";

dffeas \fft_imag_out[2] (
	.clk(clk),
	.d(\fft_imag_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[2]~q ),
	.prn(vcc));
defparam \fft_imag_out[2] .is_wysiwyg = "true";
defparam \fft_imag_out[2] .power_up = "low";

dffeas \fft_imag_out[3] (
	.clk(clk),
	.d(\fft_imag_out~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[3]~q ),
	.prn(vcc));
defparam \fft_imag_out[3] .is_wysiwyg = "true";
defparam \fft_imag_out[3] .power_up = "low";

dffeas \fft_imag_out[4] (
	.clk(clk),
	.d(\fft_imag_out~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[4]~q ),
	.prn(vcc));
defparam \fft_imag_out[4] .is_wysiwyg = "true";
defparam \fft_imag_out[4] .power_up = "low";

dffeas \fft_imag_out[5] (
	.clk(clk),
	.d(\fft_imag_out~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[5]~q ),
	.prn(vcc));
defparam \fft_imag_out[5] .is_wysiwyg = "true";
defparam \fft_imag_out[5] .power_up = "low";

dffeas \fft_imag_out[6] (
	.clk(clk),
	.d(\fft_imag_out~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[6]~q ),
	.prn(vcc));
defparam \fft_imag_out[6] .is_wysiwyg = "true";
defparam \fft_imag_out[6] .power_up = "low";

dffeas \fft_imag_out[7] (
	.clk(clk),
	.d(\fft_imag_out~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[7]~q ),
	.prn(vcc));
defparam \fft_imag_out[7] .is_wysiwyg = "true";
defparam \fft_imag_out[7] .power_up = "low";

dffeas \fft_imag_out[8] (
	.clk(clk),
	.d(\fft_imag_out~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[8]~q ),
	.prn(vcc));
defparam \fft_imag_out[8] .is_wysiwyg = "true";
defparam \fft_imag_out[8] .power_up = "low";

dffeas \fft_imag_out[9] (
	.clk(clk),
	.d(\fft_imag_out~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[9]~q ),
	.prn(vcc));
defparam \fft_imag_out[9] .is_wysiwyg = "true";
defparam \fft_imag_out[9] .power_up = "low";

dffeas \fft_imag_out[10] (
	.clk(clk),
	.d(\fft_imag_out~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[10]~q ),
	.prn(vcc));
defparam \fft_imag_out[10] .is_wysiwyg = "true";
defparam \fft_imag_out[10] .power_up = "low";

dffeas \fft_imag_out[11] (
	.clk(clk),
	.d(\fft_imag_out~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[11]~q ),
	.prn(vcc));
defparam \fft_imag_out[11] .is_wysiwyg = "true";
defparam \fft_imag_out[11] .power_up = "low";

dffeas \fft_imag_out[12] (
	.clk(clk),
	.d(\fft_imag_out~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[12]~q ),
	.prn(vcc));
defparam \fft_imag_out[12] .is_wysiwyg = "true";
defparam \fft_imag_out[12] .power_up = "low";

dffeas \fft_imag_out[13] (
	.clk(clk),
	.d(\fft_imag_out~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[13]~q ),
	.prn(vcc));
defparam \fft_imag_out[13] .is_wysiwyg = "true";
defparam \fft_imag_out[13] .power_up = "low";

dffeas \fft_imag_out[14] (
	.clk(clk),
	.d(\fft_imag_out~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[14]~q ),
	.prn(vcc));
defparam \fft_imag_out[14] .is_wysiwyg = "true";
defparam \fft_imag_out[14] .power_up = "low";

dffeas \fft_imag_out[15] (
	.clk(clk),
	.d(\fft_imag_out~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_imag_out[15]~q ),
	.prn(vcc));
defparam \fft_imag_out[15] .is_wysiwyg = "true";
defparam \fft_imag_out[15] .power_up = "low";

dffeas \fft_s1_cur.IDLE (
	.clk(clk),
	.d(\fft_s1_cur.IDLE~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_s1_cur.IDLE~q ),
	.prn(vcc));
defparam \fft_s1_cur.IDLE .is_wysiwyg = "true";
defparam \fft_s1_cur.IDLE .power_up = "low";

cycloneive_lcell_comb \WideOr3~0 (
	.dataa(\fft_s1_cur.WAIT_FOR_INPUT~q ),
	.datab(\fft_s1_cur.WRITE_INPUT~q ),
	.datac(gnd),
	.datad(\fft_s1_cur.IDLE~q ),
	.cin(gnd),
	.combout(\WideOr3~0_combout ),
	.cout());
defparam \WideOr3~0 .lut_mask = 16'hEEFF;
defparam \WideOr3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \global_clock_enable~0 (
	.dataa(\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.datab(\source_valid_ctrl_sop~1_combout ),
	.datac(gnd),
	.datad(\auk_dsp_interface_controller_1|stall_reg~q ),
	.cin(gnd),
	.combout(\global_clock_enable~0_combout ),
	.cout());
defparam \global_clock_enable~0 .lut_mask = 16'hDD11;
defparam \global_clock_enable~0 .sum_lutc_input = "datac";

dffeas val_out(
	.clk(clk),
	.d(\val_out~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\val_out~q ),
	.prn(vcc));
defparam val_out.is_wysiwyg = "true";
defparam val_out.power_up = "low";

cycloneive_lcell_comb \master_source_ena~0 (
	.dataa(reset_n),
	.datab(\val_out~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\master_source_ena~0_combout ),
	.cout());
defparam \master_source_ena~0 .lut_mask = 16'hEEEE;
defparam \master_source_ena~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sop~0 (
	.dataa(\auk_dsp_atlantic_sink_1|send_eop_s~q ),
	.datab(\sink_ready_ctrl_d~q ),
	.datac(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datad(\sop~q ),
	.cin(gnd),
	.combout(\sop~0_combout ),
	.cout());
defparam \sop~0 .lut_mask = 16'hF7D5;
defparam \sop~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \LessThan0~0 (
	.dataa(\data_count_sig[6]~q ),
	.datab(\data_count_sig[0]~q ),
	.datac(\data_count_sig[5]~q ),
	.datad(\data_count_sig[4]~q ),
	.cin(gnd),
	.combout(\LessThan0~0_combout ),
	.cout());
defparam \LessThan0~0 .lut_mask = 16'h7FFF;
defparam \LessThan0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \LessThan0~1 (
	.dataa(\data_count_sig[3]~q ),
	.datab(\data_count_sig[1]~q ),
	.datac(\data_count_sig[7]~q ),
	.datad(\data_count_sig[2]~q ),
	.cin(gnd),
	.combout(\LessThan0~1_combout ),
	.cout());
defparam \LessThan0~1 .lut_mask = 16'h7FFF;
defparam \LessThan0~1 .sum_lutc_input = "datac";

dffeas master_source_sop(
	.clk(clk),
	.d(\master_source_sop~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\master_source_sop~q ),
	.prn(vcc));
defparam master_source_sop.is_wysiwyg = "true";
defparam master_source_sop.power_up = "low";

cycloneive_lcell_comb \data_count_sig[1]~22 (
	.dataa(\LessThan0~0_combout ),
	.datab(\LessThan0~1_combout ),
	.datac(gnd),
	.datad(\master_source_sop~q ),
	.cin(gnd),
	.combout(\data_count_sig[1]~22_combout ),
	.cout());
defparam \data_count_sig[1]~22 .lut_mask = 16'hEEFF;
defparam \data_count_sig[1]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\data_count_sig[6]~q ),
	.datab(\data_count_sig[0]~q ),
	.datac(\data_count_sig[5]~q ),
	.datad(\data_count_sig[4]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h7FFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\data_count_sig[3]~q ),
	.datab(\data_count_sig[1]~q ),
	.datac(\data_count_sig[7]~q ),
	.datad(\data_count_sig[2]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h7FFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_count_sig[1]~23 (
	.dataa(\data_count_sig[1]~22_combout ),
	.datab(gnd),
	.datac(\Equal0~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\data_count_sig[1]~23_combout ),
	.cout());
defparam \data_count_sig[1]~23 .lut_mask = 16'hFFF5;
defparam \data_count_sig[1]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_count_sig[6]~24 (
	.dataa(\global_clock_enable~0_combout ),
	.datab(\data_count_sig[1]~22_combout ),
	.datac(\Equal0~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\data_count_sig[6]~24_combout ),
	.cout());
defparam \data_count_sig[6]~24 .lut_mask = 16'hBFFF;
defparam \data_count_sig[6]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \exponent_out~0 (
	.dataa(reset_n),
	.datab(\val_out~q ),
	.datac(\gen_se:bfpc|blk_exp[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~0_combout ),
	.cout());
defparam \exponent_out~0 .lut_mask = 16'hFEFE;
defparam \exponent_out~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \exponent_out~1 (
	.dataa(reset_n),
	.datab(\val_out~q ),
	.datac(\gen_se:bfpc|blk_exp[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~1_combout ),
	.cout());
defparam \exponent_out~1 .lut_mask = 16'hFEFE;
defparam \exponent_out~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \exponent_out~2 (
	.dataa(reset_n),
	.datab(\val_out~q ),
	.datac(\gen_se:bfpc|blk_exp[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~2_combout ),
	.cout());
defparam \exponent_out~2 .lut_mask = 16'hFEFE;
defparam \exponent_out~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \exponent_out~3 (
	.dataa(reset_n),
	.datab(\val_out~q ),
	.datac(\gen_se:bfpc|blk_exp[3]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~3_combout ),
	.cout());
defparam \exponent_out~3 .lut_mask = 16'hFEFE;
defparam \exponent_out~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \exponent_out~4 (
	.dataa(reset_n),
	.datab(\val_out~q ),
	.datac(\gen_se:bfpc|blk_exp[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~4_combout ),
	.cout());
defparam \exponent_out~4 .lut_mask = 16'hFEFE;
defparam \exponent_out~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \exponent_out~5 (
	.dataa(reset_n),
	.datab(\val_out~q ),
	.datac(\gen_se:bfpc|blk_exp[5]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~5_combout ),
	.cout());
defparam \exponent_out~5 .lut_mask = 16'hFEFE;
defparam \exponent_out~5 .sum_lutc_input = "datac";

dffeas fft_dirn(
	.clk(clk),
	.d(\fft_dirn~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fft_dirn~q ),
	.prn(vcc));
defparam fft_dirn.is_wysiwyg = "true";
defparam fft_dirn.power_up = "low";

cycloneive_lcell_comb \fft_real_out~0 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[16] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~0_combout ),
	.cout());
defparam \fft_real_out~0 .lut_mask = 16'hFAFC;
defparam \fft_real_out~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~1 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[17] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~1_combout ),
	.cout());
defparam \fft_real_out~1 .lut_mask = 16'hFAFC;
defparam \fft_real_out~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~2 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[18] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~2_combout ),
	.cout());
defparam \fft_real_out~2 .lut_mask = 16'hFAFC;
defparam \fft_real_out~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~3 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[19] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~3_combout ),
	.cout());
defparam \fft_real_out~3 .lut_mask = 16'hFAFC;
defparam \fft_real_out~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~4 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[20] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~4_combout ),
	.cout());
defparam \fft_real_out~4 .lut_mask = 16'hFAFC;
defparam \fft_real_out~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~5 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[21] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~5_combout ),
	.cout());
defparam \fft_real_out~5 .lut_mask = 16'hFAFC;
defparam \fft_real_out~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~6 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[22] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~6_combout ),
	.cout());
defparam \fft_real_out~6 .lut_mask = 16'hFAFC;
defparam \fft_real_out~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~7 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[23] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~7_combout ),
	.cout());
defparam \fft_real_out~7 .lut_mask = 16'hFAFC;
defparam \fft_real_out~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~8 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[24] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~8_combout ),
	.cout());
defparam \fft_real_out~8 .lut_mask = 16'hFAFC;
defparam \fft_real_out~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~9 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[25] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~9_combout ),
	.cout());
defparam \fft_real_out~9 .lut_mask = 16'hFAFC;
defparam \fft_real_out~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~10 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[26] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~10_combout ),
	.cout());
defparam \fft_real_out~10 .lut_mask = 16'hFAFC;
defparam \fft_real_out~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~11 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[27] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~11_combout ),
	.cout());
defparam \fft_real_out~11 .lut_mask = 16'hFAFC;
defparam \fft_real_out~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~12 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[28] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~12_combout ),
	.cout());
defparam \fft_real_out~12 .lut_mask = 16'hFAFC;
defparam \fft_real_out~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~13 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[29] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~13_combout ),
	.cout());
defparam \fft_real_out~13 .lut_mask = 16'hFAFC;
defparam \fft_real_out~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~14 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[30] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~14_combout ),
	.cout());
defparam \fft_real_out~14 .lut_mask = 16'hFAFC;
defparam \fft_real_out~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~15 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[31] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~15_combout ),
	.cout());
defparam \fft_real_out~15 .lut_mask = 16'hFAFC;
defparam \fft_real_out~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~0 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[16] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[0] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~0_combout ),
	.cout());
defparam \fft_imag_out~0 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~1 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[17] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[1] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~1_combout ),
	.cout());
defparam \fft_imag_out~1 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~2 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[18] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[2] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~2_combout ),
	.cout());
defparam \fft_imag_out~2 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~3 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[19] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[3] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~3_combout ),
	.cout());
defparam \fft_imag_out~3 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~4 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[20] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[4] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~4_combout ),
	.cout());
defparam \fft_imag_out~4 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~5 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[21] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[5] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~5_combout ),
	.cout());
defparam \fft_imag_out~5 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~6 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[22] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[6] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~6_combout ),
	.cout());
defparam \fft_imag_out~6 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~7 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[23] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[7] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~7_combout ),
	.cout());
defparam \fft_imag_out~7 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~8 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[24] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[8] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~8_combout ),
	.cout());
defparam \fft_imag_out~8 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~9 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[25] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[9] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~9_combout ),
	.cout());
defparam \fft_imag_out~9 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~10 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[26] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[10] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~10_combout ),
	.cout());
defparam \fft_imag_out~10 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~11 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[27] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[11] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~11_combout ),
	.cout());
defparam \fft_imag_out~11 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~12 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[28] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[12] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~12_combout ),
	.cout());
defparam \fft_imag_out~12 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~13 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[29] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[13] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~13_combout ),
	.cout());
defparam \fft_imag_out~13 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~14 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[30] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[14] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~14_combout ),
	.cout());
defparam \fft_imag_out~14 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~15 (
	.dataa(\master_source_ena~0_combout ),
	.datab(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[31] ),
	.datac(\gen_1_ram:gen_M4K:dat_A|dat_A|gen_M4K:altsyncram_component|auto_generated|q_b[15] ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~15_combout ),
	.cout());
defparam \fft_imag_out~15 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector5~0 (
	.dataa(\fft_s1_cur.WAIT_FOR_INPUT~q ),
	.datab(gnd),
	.datac(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datad(\fft_s1_cur.IDLE~q ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hAFFF;
defparam \Selector5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector6~0 (
	.dataa(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datab(\fft_s1_cur.WAIT_FOR_INPUT~q ),
	.datac(\fft_s1_cur.WRITE_INPUT~q ),
	.datad(\writer|disable_wr~q ),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
defparam \Selector6~0 .lut_mask = 16'hFEFF;
defparam \Selector6~0 .sum_lutc_input = "datac";

dffeas eop_out(
	.clk(clk),
	.d(\fft_s2_cur.LPP_DONE~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\eop_out~q ),
	.prn(vcc));
defparam eop_out.is_wysiwyg = "true";
defparam eop_out.power_up = "low";

cycloneive_lcell_comb \fft_s1_cur.IDLE~0 (
	.dataa(\eop_out~q ),
	.datab(\fft_s1_cur.FFT_PROCESS_A~q ),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\fft_s1_cur.IDLE~0_combout ),
	.cout());
defparam \fft_s1_cur.IDLE~0 .lut_mask = 16'hFF77;
defparam \fft_s1_cur.IDLE~0 .sum_lutc_input = "datac";

dffeas \fft_s2_cur.IDLE (
	.clk(clk),
	.d(reset_n),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_s2_cur.IDLE~q ),
	.prn(vcc));
defparam \fft_s2_cur.IDLE .is_wysiwyg = "true";
defparam \fft_s2_cur.IDLE .power_up = "low";

dffeas \fft_s2_cur.FIRST_LPP (
	.clk(clk),
	.d(\fft_s2_cur~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_s2_cur.FIRST_LPP~q ),
	.prn(vcc));
defparam \fft_s2_cur.FIRST_LPP .is_wysiwyg = "true";
defparam \fft_s2_cur.FIRST_LPP .power_up = "low";

dffeas \fft_s2_cur.LPP_DONE (
	.clk(clk),
	.d(\fft_s2_cur~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\fft_s2_cur.LPP_DONE~q ),
	.prn(vcc));
defparam \fft_s2_cur.LPP_DONE .is_wysiwyg = "true";
defparam \fft_s2_cur.LPP_DONE .power_up = "low";

cycloneive_lcell_comb \val_out~0 (
	.dataa(\fft_s2_cur.IDLE~q ),
	.datab(\fft_s2_cur.FIRST_LPP~q ),
	.datac(\fft_s2_cur.LPP_OUTPUT_RDY~q ),
	.datad(\fft_s2_cur.LPP_DONE~q ),
	.cin(gnd),
	.combout(\val_out~0_combout ),
	.cout());
defparam \val_out~0 .lut_mask = 16'hFFFE;
defparam \val_out~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \val_out~1 (
	.dataa(\val_out~0_combout ),
	.datab(gnd),
	.datac(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datad(\fft_s2_cur.START_LPP~q ),
	.cin(gnd),
	.combout(\val_out~1_combout ),
	.cout());
defparam \val_out~1 .lut_mask = 16'hAFFF;
defparam \val_out~1 .sum_lutc_input = "datac";

dffeas sop_out(
	.clk(clk),
	.d(\fft_s2_cur.FIRST_LPP~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\sop_out~q ),
	.prn(vcc));
defparam sop_out.is_wysiwyg = "true";
defparam sop_out.power_up = "low";

cycloneive_lcell_comb \master_source_sop~0 (
	.dataa(reset_n),
	.datab(\val_out~q ),
	.datac(\sop_out~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\master_source_sop~0_combout ),
	.cout());
defparam \master_source_sop~0 .lut_mask = 16'hFEFE;
defparam \master_source_sop~0 .sum_lutc_input = "datac";

dffeas sop_d(
	.clk(clk),
	.d(\sop_de~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\sop_d~q ),
	.prn(vcc));
defparam sop_d.is_wysiwyg = "true";
defparam sop_d.power_up = "low";

dffeas wren_a(
	.clk(clk),
	.d(\wren_a~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wren_a~q ),
	.prn(vcc));
defparam wren_a.is_wysiwyg = "true";
defparam wren_a.power_up = "low";

cycloneive_lcell_comb \fft_dirn~0 (
	.dataa(\fft_dirn~q ),
	.datab(inverse),
	.datac(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datad(\global_clock_enable~0_combout ),
	.cin(gnd),
	.combout(\fft_dirn~0_combout ),
	.cout());
defparam \fft_dirn~0 .lut_mask = 16'hEFFE;
defparam \fft_dirn~0 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[24] (
	.clk(clk),
	.d(\data_rdy_vec~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[24]~q ),
	.prn(vcc));
defparam \data_rdy_vec[24] .is_wysiwyg = "true";
defparam \data_rdy_vec[24] .power_up = "low";

cycloneive_lcell_comb \Selector10~0 (
	.dataa(\data_rdy_vec[24]~q ),
	.datab(\fft_s1_cur.NO_WRITE~q ),
	.datac(\fft_s1_cur.FFT_PROCESS_A~q ),
	.datad(\eop_out~q ),
	.cin(gnd),
	.combout(\Selector10~0_combout ),
	.cout());
defparam \Selector10~0 .lut_mask = 16'hFEFF;
defparam \Selector10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s2_cur~8 (
	.dataa(reset_n),
	.datab(\fft_s2_cur.START_LPP~q ),
	.datac(\sop_d~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\fft_s2_cur~8_combout ),
	.cout());
defparam \fft_s2_cur~8 .lut_mask = 16'hFEFE;
defparam \fft_s2_cur~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal9~0 (
	.dataa(\output_count[1]~q ),
	.datab(\output_count[2]~q ),
	.datac(\output_count[3]~q ),
	.datad(\output_count[0]~q ),
	.cin(gnd),
	.combout(\Equal9~0_combout ),
	.cout());
defparam \Equal9~0 .lut_mask = 16'hFEFF;
defparam \Equal9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal9~1 (
	.dataa(\output_count[4]~q ),
	.datab(\output_count[5]~q ),
	.datac(\output_count[6]~q ),
	.datad(\output_count[7]~q ),
	.cin(gnd),
	.combout(\Equal9~1_combout ),
	.cout());
defparam \Equal9~1 .lut_mask = 16'hFFFE;
defparam \Equal9~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~0 (
	.dataa(\fft_s2_cur.FIRST_LPP~q ),
	.datab(\fft_s2_cur.LPP_OUTPUT_RDY~q ),
	.datac(\Equal9~0_combout ),
	.datad(\Equal9~1_combout ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hEFFF;
defparam \Selector2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s2_cur~9 (
	.dataa(reset_n),
	.datab(\fft_s2_cur.LPP_OUTPUT_RDY~q ),
	.datac(\Equal9~0_combout ),
	.datad(\Equal9~1_combout ),
	.cin(gnd),
	.combout(\fft_s2_cur~9_combout ),
	.cout());
defparam \fft_s2_cur~9 .lut_mask = 16'hFFFE;
defparam \fft_s2_cur~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector0~0 (
	.dataa(\fft_s2_cur.LPP_DONE~q ),
	.datab(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datac(\ctrl|blk_done~q ),
	.datad(\fft_s2_cur.IDLE~q ),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hEFFF;
defparam \Selector0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~0 (
	.dataa(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datab(\ctrl|blk_done~q ),
	.datac(\fft_s2_cur.START_LPP~q ),
	.datad(\sop_d~q ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hFEFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

dffeas sop_de(
	.clk(clk),
	.d(\sop_de~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\sop_de~q ),
	.prn(vcc));
defparam sop_de.is_wysiwyg = "true";
defparam sop_de.power_up = "low";

cycloneive_lcell_comb \wren_a~2 (
	.dataa(\writer|gen_soe:delay_swd|tdl_arr[0]~q ),
	.datab(\fft_s1_cur.WRITE_INPUT~q ),
	.datac(\fft_s1_cur.EARLY_DONE~q ),
	.datad(\fft_s1_cur.DONE_WRITING~q ),
	.cin(gnd),
	.combout(\wren_a~2_combout ),
	.cout());
defparam \wren_a~2 .lut_mask = 16'hFFFE;
defparam \wren_a~2 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[21] (
	.clk(clk),
	.d(\data_rdy_vec~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[21]~q ),
	.prn(vcc));
defparam \data_rdy_vec[21] .is_wysiwyg = "true";
defparam \data_rdy_vec[21] .power_up = "low";

cycloneive_lcell_comb \wren_a~3 (
	.dataa(\data_rdy_vec[21]~q ),
	.datab(\fft_s1_cur.WRITE_INPUT~q ),
	.datac(\fft_s1_cur.EARLY_DONE~q ),
	.datad(\fft_s1_cur.DONE_WRITING~q ),
	.cin(gnd),
	.combout(\wren_a~3_combout ),
	.cout());
defparam \wren_a~3 .lut_mask = 16'hBFFF;
defparam \wren_a~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wren_a~4 (
	.dataa(\fft_s1_cur.IDLE~q ),
	.datab(\wren_a~2_combout ),
	.datac(\wren_a~3_combout ),
	.datad(\fft_s1_cur.NO_WRITE~q ),
	.cin(gnd),
	.combout(\wren_a~4_combout ),
	.cout());
defparam \wren_a~4 .lut_mask = 16'hFEFF;
defparam \wren_a~4 .sum_lutc_input = "datac";

dffeas sel_ram_in(
	.clk(clk),
	.d(\sel_ram_in~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\sel_ram_in~q ),
	.prn(vcc));
defparam sel_ram_in.is_wysiwyg = "true";
defparam sel_ram_in.power_up = "low";

dffeas \wraddress_a_bus_ctrl_i[0] (
	.clk(clk),
	.d(\gen_wraddr_se:wr_adgen|rd_addr_a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wraddress_a_bus_ctrl_i[0]~q ),
	.prn(vcc));
defparam \wraddress_a_bus_ctrl_i[0] .is_wysiwyg = "true";
defparam \wraddress_a_bus_ctrl_i[0] .power_up = "low";

dffeas \wraddress_a_bus_ctrl_i[1] (
	.clk(clk),
	.d(\gen_wraddr_se:wr_adgen|rd_addr_a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wraddress_a_bus_ctrl_i[1]~q ),
	.prn(vcc));
defparam \wraddress_a_bus_ctrl_i[1] .is_wysiwyg = "true";
defparam \wraddress_a_bus_ctrl_i[1] .power_up = "low";

dffeas \wraddress_a_bus_ctrl_i[2] (
	.clk(clk),
	.d(\gen_wraddr_se:wr_adgen|rd_addr_a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wraddress_a_bus_ctrl_i[2]~q ),
	.prn(vcc));
defparam \wraddress_a_bus_ctrl_i[2] .is_wysiwyg = "true";
defparam \wraddress_a_bus_ctrl_i[2] .power_up = "low";

dffeas \wraddress_a_bus_ctrl_i[3] (
	.clk(clk),
	.d(\gen_wraddr_se:wr_adgen|rd_addr_a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wraddress_a_bus_ctrl_i[3]~q ),
	.prn(vcc));
defparam \wraddress_a_bus_ctrl_i[3] .is_wysiwyg = "true";
defparam \wraddress_a_bus_ctrl_i[3] .power_up = "low";

dffeas \wraddress_a_bus_ctrl_i[4] (
	.clk(clk),
	.d(\gen_wraddr_se:wr_adgen|rd_addr_a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wraddress_a_bus_ctrl_i[4]~q ),
	.prn(vcc));
defparam \wraddress_a_bus_ctrl_i[4] .is_wysiwyg = "true";
defparam \wraddress_a_bus_ctrl_i[4] .power_up = "low";

dffeas \wraddress_a_bus_ctrl_i[5] (
	.clk(clk),
	.d(\gen_wraddr_se:wr_adgen|rd_addr_a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wraddress_a_bus_ctrl_i[5]~q ),
	.prn(vcc));
defparam \wraddress_a_bus_ctrl_i[5] .is_wysiwyg = "true";
defparam \wraddress_a_bus_ctrl_i[5] .power_up = "low";

dffeas \wraddress_a_bus_ctrl_i[6] (
	.clk(clk),
	.d(\gen_wraddr_se:wr_adgen|rd_addr_a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wraddress_a_bus_ctrl_i[6]~q ),
	.prn(vcc));
defparam \wraddress_a_bus_ctrl_i[6] .is_wysiwyg = "true";
defparam \wraddress_a_bus_ctrl_i[6] .power_up = "low";

dffeas \wraddress_a_bus_ctrl_i[7] (
	.clk(clk),
	.d(\gen_wraddr_se:wr_adgen|rd_addr_a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\wraddress_a_bus_ctrl_i[7]~q ),
	.prn(vcc));
defparam \wraddress_a_bus_ctrl_i[7] .is_wysiwyg = "true";
defparam \wraddress_a_bus_ctrl_i[7] .power_up = "low";

dffeas \data_rdy_vec[23] (
	.clk(clk),
	.d(\data_rdy_vec~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[23]~q ),
	.prn(vcc));
defparam \data_rdy_vec[23] .is_wysiwyg = "true";
defparam \data_rdy_vec[23] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~0 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[23]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~0_combout ),
	.cout());
defparam \data_rdy_vec~0 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector9~0 (
	.dataa(\fft_s1_cur.DONE_WRITING~q ),
	.datab(\no_del_input_blk:delay_next_block|tdl_arr[0]~q ),
	.datac(\fft_s1_cur.NO_WRITE~q ),
	.datad(\data_rdy_vec[24]~q ),
	.cin(gnd),
	.combout(\Selector9~0_combout ),
	.cout());
defparam \Selector9~0 .lut_mask = 16'hFEFF;
defparam \Selector9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \output_sample_counter~0 (
	.dataa(\fft_s2_cur.FIRST_LPP~q ),
	.datab(\fft_s2_cur.LPP_OUTPUT_RDY~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\output_sample_counter~0_combout ),
	.cout());
defparam \output_sample_counter~0 .lut_mask = 16'h7777;
defparam \output_sample_counter~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sop_de~0 (
	.dataa(\fft_s2_cur.START_LPP~q ),
	.datab(\del_sop_cnt[0]~q ),
	.datac(\del_sop_cnt[1]~q ),
	.datad(\del_sop_cnt[2]~q ),
	.cin(gnd),
	.combout(\sop_de~0_combout ),
	.cout());
defparam \sop_de~0 .lut_mask = 16'hFEFF;
defparam \sop_de~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sop_de~1 (
	.dataa(\sop_de~0_combout ),
	.datab(\del_sop_cnt[4]~q ),
	.datac(gnd),
	.datad(\del_sop_cnt[3]~q ),
	.cin(gnd),
	.combout(\sop_de~1_combout ),
	.cout());
defparam \sop_de~1 .lut_mask = 16'hEEFF;
defparam \sop_de~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector7~0 (
	.dataa(\fft_s1_cur.WRITE_INPUT~q ),
	.datab(\writer|disable_wr~q ),
	.datac(\fft_s1_cur.EARLY_DONE~q ),
	.datad(\writer|rdy_for_next_block~q ),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
defparam \Selector7~0 .lut_mask = 16'hFEFF;
defparam \Selector7~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector8~0 (
	.dataa(\writer|rdy_for_next_block~q ),
	.datab(\fft_s1_cur.EARLY_DONE~q ),
	.datac(\fft_s1_cur.DONE_WRITING~q ),
	.datad(\no_del_input_blk:delay_next_block|tdl_arr[0]~q ),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
defparam \Selector8~0 .lut_mask = 16'hFEFF;
defparam \Selector8~0 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[20] (
	.clk(clk),
	.d(\data_rdy_vec~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[20]~q ),
	.prn(vcc));
defparam \data_rdy_vec[20] .is_wysiwyg = "true";
defparam \data_rdy_vec[20] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~1 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~1_combout ),
	.cout());
defparam \data_rdy_vec~1 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sel_ram_in~0 (
	.dataa(\fft_s1_cur.WRITE_INPUT~q ),
	.datab(\fft_s1_cur.EARLY_DONE~q ),
	.datac(\fft_s1_cur.DONE_WRITING~q ),
	.datad(\fft_s1_cur.IDLE~q ),
	.cin(gnd),
	.combout(\sel_ram_in~0_combout ),
	.cout());
defparam \sel_ram_in~0 .lut_mask = 16'hFF7F;
defparam \sel_ram_in~0 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[22] (
	.clk(clk),
	.d(\data_rdy_vec~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[22]~q ),
	.prn(vcc));
defparam \data_rdy_vec[22] .is_wysiwyg = "true";
defparam \data_rdy_vec[22] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~2 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[22]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~2_combout ),
	.cout());
defparam \data_rdy_vec~2 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~2 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[4] (
	.clk(clk),
	.d(\data_rdy_vec~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[4]~q ),
	.prn(vcc));
defparam \data_rdy_vec[4] .is_wysiwyg = "true";
defparam \data_rdy_vec[4] .power_up = "low";

dffeas \data_rdy_vec[19] (
	.clk(clk),
	.d(\data_rdy_vec~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[19]~q ),
	.prn(vcc));
defparam \data_rdy_vec[19] .is_wysiwyg = "true";
defparam \data_rdy_vec[19] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~3 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[19]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~3_combout ),
	.cout());
defparam \data_rdy_vec~3 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~3 .sum_lutc_input = "datac";

dffeas \data_real_in_reg[0] (
	.clk(clk),
	.d(\data_real_in_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[0]~q ),
	.prn(vcc));
defparam \data_real_in_reg[0] .is_wysiwyg = "true";
defparam \data_real_in_reg[0] .power_up = "low";

dffeas \data_imag_in_reg[0] (
	.clk(clk),
	.d(\data_imag_in_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[0]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[0] .is_wysiwyg = "true";
defparam \data_imag_in_reg[0] .power_up = "low";

cycloneive_lcell_comb \core_imag_in~0 (
	.dataa(\data_real_in_reg[0]~q ),
	.datab(\data_imag_in_reg[0]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~0_combout ),
	.cout());
defparam \core_imag_in~0 .lut_mask = 16'hAACC;
defparam \core_imag_in~0 .sum_lutc_input = "datac";

dffeas \p_tdl[18][0] (
	.clk(clk),
	.d(\p_tdl~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[18][0]~q ),
	.prn(vcc));
defparam \p_tdl[18][0] .is_wysiwyg = "true";
defparam \p_tdl[18][0] .power_up = "low";

dffeas \p_tdl[18][1] (
	.clk(clk),
	.d(\p_tdl~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[18][1]~q ),
	.prn(vcc));
defparam \p_tdl[18][1] .is_wysiwyg = "true";
defparam \p_tdl[18][1] .power_up = "low";

dffeas \p_tdl[18][2] (
	.clk(clk),
	.d(\p_tdl~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[18][2]~q ),
	.prn(vcc));
defparam \p_tdl[18][2] .is_wysiwyg = "true";
defparam \p_tdl[18][2] .power_up = "low";

cycloneive_lcell_comb \core_real_in~0 (
	.dataa(\data_imag_in_reg[0]~q ),
	.datab(\data_real_in_reg[0]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~0_combout ),
	.cout());
defparam \core_real_in~0 .lut_mask = 16'hAACC;
defparam \core_real_in~0 .sum_lutc_input = "datac";

dffeas \data_real_in_reg[1] (
	.clk(clk),
	.d(\data_real_in_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[1]~q ),
	.prn(vcc));
defparam \data_real_in_reg[1] .is_wysiwyg = "true";
defparam \data_real_in_reg[1] .power_up = "low";

dffeas \data_imag_in_reg[1] (
	.clk(clk),
	.d(\data_imag_in_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[1]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[1] .is_wysiwyg = "true";
defparam \data_imag_in_reg[1] .power_up = "low";

cycloneive_lcell_comb \core_imag_in~1 (
	.dataa(\data_real_in_reg[1]~q ),
	.datab(\data_imag_in_reg[1]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~1_combout ),
	.cout());
defparam \core_imag_in~1 .lut_mask = 16'hAACC;
defparam \core_imag_in~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_real_in~1 (
	.dataa(\data_imag_in_reg[1]~q ),
	.datab(\data_real_in_reg[1]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~1_combout ),
	.cout());
defparam \core_real_in~1 .lut_mask = 16'hAACC;
defparam \core_real_in~1 .sum_lutc_input = "datac";

dffeas \data_real_in_reg[2] (
	.clk(clk),
	.d(\data_real_in_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[2]~q ),
	.prn(vcc));
defparam \data_real_in_reg[2] .is_wysiwyg = "true";
defparam \data_real_in_reg[2] .power_up = "low";

dffeas \data_imag_in_reg[2] (
	.clk(clk),
	.d(\data_imag_in_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[2]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[2] .is_wysiwyg = "true";
defparam \data_imag_in_reg[2] .power_up = "low";

cycloneive_lcell_comb \core_imag_in~2 (
	.dataa(\data_real_in_reg[2]~q ),
	.datab(\data_imag_in_reg[2]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~2_combout ),
	.cout());
defparam \core_imag_in~2 .lut_mask = 16'hAACC;
defparam \core_imag_in~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_real_in~2 (
	.dataa(\data_imag_in_reg[2]~q ),
	.datab(\data_real_in_reg[2]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~2_combout ),
	.cout());
defparam \core_real_in~2 .lut_mask = 16'hAACC;
defparam \core_real_in~2 .sum_lutc_input = "datac";

dffeas \data_real_in_reg[3] (
	.clk(clk),
	.d(\data_real_in_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[3]~q ),
	.prn(vcc));
defparam \data_real_in_reg[3] .is_wysiwyg = "true";
defparam \data_real_in_reg[3] .power_up = "low";

dffeas \data_imag_in_reg[3] (
	.clk(clk),
	.d(\data_imag_in_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[3]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[3] .is_wysiwyg = "true";
defparam \data_imag_in_reg[3] .power_up = "low";

cycloneive_lcell_comb \core_imag_in~3 (
	.dataa(\data_real_in_reg[3]~q ),
	.datab(\data_imag_in_reg[3]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~3_combout ),
	.cout());
defparam \core_imag_in~3 .lut_mask = 16'hAACC;
defparam \core_imag_in~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_real_in~3 (
	.dataa(\data_imag_in_reg[3]~q ),
	.datab(\data_real_in_reg[3]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~3_combout ),
	.cout());
defparam \core_real_in~3 .lut_mask = 16'hAACC;
defparam \core_real_in~3 .sum_lutc_input = "datac";

dffeas \data_real_in_reg[4] (
	.clk(clk),
	.d(\data_real_in_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[4]~q ),
	.prn(vcc));
defparam \data_real_in_reg[4] .is_wysiwyg = "true";
defparam \data_real_in_reg[4] .power_up = "low";

dffeas \data_imag_in_reg[4] (
	.clk(clk),
	.d(\data_imag_in_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[4]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[4] .is_wysiwyg = "true";
defparam \data_imag_in_reg[4] .power_up = "low";

cycloneive_lcell_comb \core_imag_in~4 (
	.dataa(\data_real_in_reg[4]~q ),
	.datab(\data_imag_in_reg[4]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~4_combout ),
	.cout());
defparam \core_imag_in~4 .lut_mask = 16'hAACC;
defparam \core_imag_in~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_real_in~4 (
	.dataa(\data_imag_in_reg[4]~q ),
	.datab(\data_real_in_reg[4]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~4_combout ),
	.cout());
defparam \core_real_in~4 .lut_mask = 16'hAACC;
defparam \core_real_in~4 .sum_lutc_input = "datac";

dffeas \data_real_in_reg[5] (
	.clk(clk),
	.d(\data_real_in_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[5]~q ),
	.prn(vcc));
defparam \data_real_in_reg[5] .is_wysiwyg = "true";
defparam \data_real_in_reg[5] .power_up = "low";

dffeas \data_imag_in_reg[5] (
	.clk(clk),
	.d(\data_imag_in_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[5]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[5] .is_wysiwyg = "true";
defparam \data_imag_in_reg[5] .power_up = "low";

cycloneive_lcell_comb \core_imag_in~5 (
	.dataa(\data_real_in_reg[5]~q ),
	.datab(\data_imag_in_reg[5]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~5_combout ),
	.cout());
defparam \core_imag_in~5 .lut_mask = 16'hAACC;
defparam \core_imag_in~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_real_in~5 (
	.dataa(\data_imag_in_reg[5]~q ),
	.datab(\data_real_in_reg[5]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~5_combout ),
	.cout());
defparam \core_real_in~5 .lut_mask = 16'hAACC;
defparam \core_real_in~5 .sum_lutc_input = "datac";

dffeas \data_real_in_reg[6] (
	.clk(clk),
	.d(\data_real_in_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[6]~q ),
	.prn(vcc));
defparam \data_real_in_reg[6] .is_wysiwyg = "true";
defparam \data_real_in_reg[6] .power_up = "low";

dffeas \data_imag_in_reg[6] (
	.clk(clk),
	.d(\data_imag_in_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[6]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[6] .is_wysiwyg = "true";
defparam \data_imag_in_reg[6] .power_up = "low";

cycloneive_lcell_comb \core_imag_in~6 (
	.dataa(\data_real_in_reg[6]~q ),
	.datab(\data_imag_in_reg[6]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~6_combout ),
	.cout());
defparam \core_imag_in~6 .lut_mask = 16'hAACC;
defparam \core_imag_in~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_real_in~6 (
	.dataa(\data_imag_in_reg[6]~q ),
	.datab(\data_real_in_reg[6]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~6_combout ),
	.cout());
defparam \core_real_in~6 .lut_mask = 16'hAACC;
defparam \core_real_in~6 .sum_lutc_input = "datac";

dffeas \data_real_in_reg[7] (
	.clk(clk),
	.d(\data_real_in_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[7]~q ),
	.prn(vcc));
defparam \data_real_in_reg[7] .is_wysiwyg = "true";
defparam \data_real_in_reg[7] .power_up = "low";

dffeas \data_imag_in_reg[7] (
	.clk(clk),
	.d(\data_imag_in_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[7]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[7] .is_wysiwyg = "true";
defparam \data_imag_in_reg[7] .power_up = "low";

cycloneive_lcell_comb \core_imag_in~7 (
	.dataa(\data_real_in_reg[7]~q ),
	.datab(\data_imag_in_reg[7]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~7_combout ),
	.cout());
defparam \core_imag_in~7 .lut_mask = 16'hAACC;
defparam \core_imag_in~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_real_in~7 (
	.dataa(\data_imag_in_reg[7]~q ),
	.datab(\data_real_in_reg[7]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~7_combout ),
	.cout());
defparam \core_real_in~7 .lut_mask = 16'hAACC;
defparam \core_real_in~7 .sum_lutc_input = "datac";

dffeas \data_real_in_reg[8] (
	.clk(clk),
	.d(\data_real_in_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[8]~q ),
	.prn(vcc));
defparam \data_real_in_reg[8] .is_wysiwyg = "true";
defparam \data_real_in_reg[8] .power_up = "low";

dffeas \data_imag_in_reg[8] (
	.clk(clk),
	.d(\data_imag_in_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[8]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[8] .is_wysiwyg = "true";
defparam \data_imag_in_reg[8] .power_up = "low";

cycloneive_lcell_comb \core_imag_in~8 (
	.dataa(\data_real_in_reg[8]~q ),
	.datab(\data_imag_in_reg[8]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~8_combout ),
	.cout());
defparam \core_imag_in~8 .lut_mask = 16'hAACC;
defparam \core_imag_in~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_real_in~8 (
	.dataa(\data_imag_in_reg[8]~q ),
	.datab(\data_real_in_reg[8]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~8_combout ),
	.cout());
defparam \core_real_in~8 .lut_mask = 16'hAACC;
defparam \core_real_in~8 .sum_lutc_input = "datac";

dffeas \data_real_in_reg[9] (
	.clk(clk),
	.d(\data_real_in_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[9]~q ),
	.prn(vcc));
defparam \data_real_in_reg[9] .is_wysiwyg = "true";
defparam \data_real_in_reg[9] .power_up = "low";

dffeas \data_imag_in_reg[9] (
	.clk(clk),
	.d(\data_imag_in_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[9]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[9] .is_wysiwyg = "true";
defparam \data_imag_in_reg[9] .power_up = "low";

cycloneive_lcell_comb \core_imag_in~9 (
	.dataa(\data_real_in_reg[9]~q ),
	.datab(\data_imag_in_reg[9]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~9_combout ),
	.cout());
defparam \core_imag_in~9 .lut_mask = 16'hAACC;
defparam \core_imag_in~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_real_in~9 (
	.dataa(\data_imag_in_reg[9]~q ),
	.datab(\data_real_in_reg[9]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~9_combout ),
	.cout());
defparam \core_real_in~9 .lut_mask = 16'hAACC;
defparam \core_real_in~9 .sum_lutc_input = "datac";

dffeas \data_real_in_reg[10] (
	.clk(clk),
	.d(\data_real_in_reg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[10]~q ),
	.prn(vcc));
defparam \data_real_in_reg[10] .is_wysiwyg = "true";
defparam \data_real_in_reg[10] .power_up = "low";

dffeas \data_imag_in_reg[10] (
	.clk(clk),
	.d(\data_imag_in_reg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[10]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[10] .is_wysiwyg = "true";
defparam \data_imag_in_reg[10] .power_up = "low";

cycloneive_lcell_comb \core_imag_in~10 (
	.dataa(\data_real_in_reg[10]~q ),
	.datab(\data_imag_in_reg[10]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~10_combout ),
	.cout());
defparam \core_imag_in~10 .lut_mask = 16'hAACC;
defparam \core_imag_in~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_real_in~10 (
	.dataa(\data_imag_in_reg[10]~q ),
	.datab(\data_real_in_reg[10]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~10_combout ),
	.cout());
defparam \core_real_in~10 .lut_mask = 16'hAACC;
defparam \core_real_in~10 .sum_lutc_input = "datac";

dffeas \data_real_in_reg[11] (
	.clk(clk),
	.d(\data_real_in_reg~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[11]~q ),
	.prn(vcc));
defparam \data_real_in_reg[11] .is_wysiwyg = "true";
defparam \data_real_in_reg[11] .power_up = "low";

dffeas \data_imag_in_reg[11] (
	.clk(clk),
	.d(\data_imag_in_reg~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[11]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[11] .is_wysiwyg = "true";
defparam \data_imag_in_reg[11] .power_up = "low";

cycloneive_lcell_comb \core_imag_in~11 (
	.dataa(\data_real_in_reg[11]~q ),
	.datab(\data_imag_in_reg[11]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~11_combout ),
	.cout());
defparam \core_imag_in~11 .lut_mask = 16'hAACC;
defparam \core_imag_in~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_real_in~11 (
	.dataa(\data_imag_in_reg[11]~q ),
	.datab(\data_real_in_reg[11]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~11_combout ),
	.cout());
defparam \core_real_in~11 .lut_mask = 16'hAACC;
defparam \core_real_in~11 .sum_lutc_input = "datac";

dffeas \data_real_in_reg[12] (
	.clk(clk),
	.d(\data_real_in_reg~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[12]~q ),
	.prn(vcc));
defparam \data_real_in_reg[12] .is_wysiwyg = "true";
defparam \data_real_in_reg[12] .power_up = "low";

dffeas \data_imag_in_reg[12] (
	.clk(clk),
	.d(\data_imag_in_reg~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[12]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[12] .is_wysiwyg = "true";
defparam \data_imag_in_reg[12] .power_up = "low";

cycloneive_lcell_comb \core_imag_in~12 (
	.dataa(\data_real_in_reg[12]~q ),
	.datab(\data_imag_in_reg[12]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~12_combout ),
	.cout());
defparam \core_imag_in~12 .lut_mask = 16'hAACC;
defparam \core_imag_in~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_real_in~12 (
	.dataa(\data_imag_in_reg[12]~q ),
	.datab(\data_real_in_reg[12]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~12_combout ),
	.cout());
defparam \core_real_in~12 .lut_mask = 16'hAACC;
defparam \core_real_in~12 .sum_lutc_input = "datac";

dffeas \data_real_in_reg[13] (
	.clk(clk),
	.d(\data_real_in_reg~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[13]~q ),
	.prn(vcc));
defparam \data_real_in_reg[13] .is_wysiwyg = "true";
defparam \data_real_in_reg[13] .power_up = "low";

dffeas \data_imag_in_reg[13] (
	.clk(clk),
	.d(\data_imag_in_reg~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[13]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[13] .is_wysiwyg = "true";
defparam \data_imag_in_reg[13] .power_up = "low";

cycloneive_lcell_comb \core_imag_in~13 (
	.dataa(\data_real_in_reg[13]~q ),
	.datab(\data_imag_in_reg[13]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~13_combout ),
	.cout());
defparam \core_imag_in~13 .lut_mask = 16'hAACC;
defparam \core_imag_in~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_real_in~13 (
	.dataa(\data_imag_in_reg[13]~q ),
	.datab(\data_real_in_reg[13]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~13_combout ),
	.cout());
defparam \core_real_in~13 .lut_mask = 16'hAACC;
defparam \core_real_in~13 .sum_lutc_input = "datac";

dffeas \data_real_in_reg[14] (
	.clk(clk),
	.d(\data_real_in_reg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[14]~q ),
	.prn(vcc));
defparam \data_real_in_reg[14] .is_wysiwyg = "true";
defparam \data_real_in_reg[14] .power_up = "low";

dffeas \data_imag_in_reg[14] (
	.clk(clk),
	.d(\data_imag_in_reg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[14]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[14] .is_wysiwyg = "true";
defparam \data_imag_in_reg[14] .power_up = "low";

cycloneive_lcell_comb \core_imag_in~14 (
	.dataa(\data_real_in_reg[14]~q ),
	.datab(\data_imag_in_reg[14]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~14_combout ),
	.cout());
defparam \core_imag_in~14 .lut_mask = 16'hAACC;
defparam \core_imag_in~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_real_in~14 (
	.dataa(\data_imag_in_reg[14]~q ),
	.datab(\data_real_in_reg[14]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~14_combout ),
	.cout());
defparam \core_real_in~14 .lut_mask = 16'hAACC;
defparam \core_real_in~14 .sum_lutc_input = "datac";

dffeas \data_real_in_reg[15] (
	.clk(clk),
	.d(\data_real_in_reg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[15]~q ),
	.prn(vcc));
defparam \data_real_in_reg[15] .is_wysiwyg = "true";
defparam \data_real_in_reg[15] .power_up = "low";

dffeas \data_imag_in_reg[15] (
	.clk(clk),
	.d(\data_imag_in_reg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[15]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[15] .is_wysiwyg = "true";
defparam \data_imag_in_reg[15] .power_up = "low";

cycloneive_lcell_comb \core_imag_in~15 (
	.dataa(\data_real_in_reg[15]~q ),
	.datab(\data_imag_in_reg[15]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~15_combout ),
	.cout());
defparam \core_imag_in~15 .lut_mask = 16'hAACC;
defparam \core_imag_in~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_real_in~15 (
	.dataa(\data_imag_in_reg[15]~q ),
	.datab(\data_real_in_reg[15]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~15_combout ),
	.cout());
defparam \core_real_in~15 .lut_mask = 16'hAACC;
defparam \core_real_in~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_rdy_vec~4 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[21]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~4_combout ),
	.cout());
defparam \data_rdy_vec~4 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~4 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[3] (
	.clk(clk),
	.d(\data_rdy_vec~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[3]~q ),
	.prn(vcc));
defparam \data_rdy_vec[3] .is_wysiwyg = "true";
defparam \data_rdy_vec[3] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~5 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~5_combout ),
	.cout());
defparam \data_rdy_vec~5 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~5 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[18] (
	.clk(clk),
	.d(\data_rdy_vec~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[18]~q ),
	.prn(vcc));
defparam \data_rdy_vec[18] .is_wysiwyg = "true";
defparam \data_rdy_vec[18] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~6 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[18]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~6_combout ),
	.cout());
defparam \data_rdy_vec~6 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~0 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~0_combout ),
	.cout());
defparam \data_real_in_reg~0 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~0 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~0_combout ),
	.cout());
defparam \data_imag_in_reg~0 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~0 .sum_lutc_input = "datac";

dffeas \p_tdl[17][0] (
	.clk(clk),
	.d(\p_tdl~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[17][0]~q ),
	.prn(vcc));
defparam \p_tdl[17][0] .is_wysiwyg = "true";
defparam \p_tdl[17][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~0 (
	.dataa(reset_n),
	.datab(\p_tdl[17][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~0_combout ),
	.cout());
defparam \p_tdl~0 .lut_mask = 16'hEEEE;
defparam \p_tdl~0 .sum_lutc_input = "datac";

dffeas \p_tdl[17][1] (
	.clk(clk),
	.d(\p_tdl~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[17][1]~q ),
	.prn(vcc));
defparam \p_tdl[17][1] .is_wysiwyg = "true";
defparam \p_tdl[17][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~1 (
	.dataa(reset_n),
	.datab(\p_tdl[17][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~1_combout ),
	.cout());
defparam \p_tdl~1 .lut_mask = 16'hEEEE;
defparam \p_tdl~1 .sum_lutc_input = "datac";

dffeas \p_tdl[17][2] (
	.clk(clk),
	.d(\p_tdl~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[17][2]~q ),
	.prn(vcc));
defparam \p_tdl[17][2] .is_wysiwyg = "true";
defparam \p_tdl[17][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~2 (
	.dataa(reset_n),
	.datab(\p_tdl[17][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~2_combout ),
	.cout());
defparam \p_tdl~2 .lut_mask = 16'hEEEE;
defparam \p_tdl~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~1 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~1_combout ),
	.cout());
defparam \data_real_in_reg~1 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~1 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~1_combout ),
	.cout());
defparam \data_imag_in_reg~1 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~2 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~2_combout ),
	.cout());
defparam \data_real_in_reg~2 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~2 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~2_combout ),
	.cout());
defparam \data_imag_in_reg~2 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~3 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~3_combout ),
	.cout());
defparam \data_real_in_reg~3 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~3 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~3_combout ),
	.cout());
defparam \data_imag_in_reg~3 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~4 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~4_combout ),
	.cout());
defparam \data_real_in_reg~4 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~4 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~4_combout ),
	.cout());
defparam \data_imag_in_reg~4 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~5 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~5_combout ),
	.cout());
defparam \data_real_in_reg~5 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~5 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~5_combout ),
	.cout());
defparam \data_imag_in_reg~5 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~6 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~6_combout ),
	.cout());
defparam \data_real_in_reg~6 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~6 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~6_combout ),
	.cout());
defparam \data_imag_in_reg~6 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~7 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[23] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~7_combout ),
	.cout());
defparam \data_real_in_reg~7 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~7 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~7_combout ),
	.cout());
defparam \data_imag_in_reg~7 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~8 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[24] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~8_combout ),
	.cout());
defparam \data_real_in_reg~8 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~8 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~8_combout ),
	.cout());
defparam \data_imag_in_reg~8 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~9 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[25] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~9_combout ),
	.cout());
defparam \data_real_in_reg~9 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~9 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~9_combout ),
	.cout());
defparam \data_imag_in_reg~9 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~10 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[26] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~10_combout ),
	.cout());
defparam \data_real_in_reg~10 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~10 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~10_combout ),
	.cout());
defparam \data_imag_in_reg~10 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~11 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[27] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~11_combout ),
	.cout());
defparam \data_real_in_reg~11 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~11 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~11_combout ),
	.cout());
defparam \data_imag_in_reg~11 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~12 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[28] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~12_combout ),
	.cout());
defparam \data_real_in_reg~12 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~12 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~12_combout ),
	.cout());
defparam \data_imag_in_reg~12 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~13 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[29] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~13_combout ),
	.cout());
defparam \data_real_in_reg~13 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~13 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~13_combout ),
	.cout());
defparam \data_imag_in_reg~13 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~14 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[30] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~14_combout ),
	.cout());
defparam \data_real_in_reg~14 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~14 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~14_combout ),
	.cout());
defparam \data_imag_in_reg~14 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~15 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[31] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~15_combout ),
	.cout());
defparam \data_real_in_reg~15 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~15 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~15_combout ),
	.cout());
defparam \data_imag_in_reg~15 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~15 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[2] (
	.clk(clk),
	.d(\data_rdy_vec~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[2]~q ),
	.prn(vcc));
defparam \data_rdy_vec[2] .is_wysiwyg = "true";
defparam \data_rdy_vec[2] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~7 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~7_combout ),
	.cout());
defparam \data_rdy_vec~7 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~7 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[17] (
	.clk(clk),
	.d(\data_rdy_vec~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[17]~q ),
	.prn(vcc));
defparam \data_rdy_vec[17] .is_wysiwyg = "true";
defparam \data_rdy_vec[17] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~8 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~8_combout ),
	.cout());
defparam \data_rdy_vec~8 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal5~0 (
	.dataa(\k_count_wr[6]~q ),
	.datab(\k_count_wr[2]~q ),
	.datac(\k_count_wr[0]~q ),
	.datad(\k_count_wr[7]~q ),
	.cin(gnd),
	.combout(\Equal5~0_combout ),
	.cout());
defparam \Equal5~0 .lut_mask = 16'hFFFE;
defparam \Equal5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal5~1 (
	.dataa(\k_count_wr[3]~q ),
	.datab(\k_count_wr[1]~q ),
	.datac(\k_count_wr[4]~q ),
	.datad(\k_count_wr[5]~q ),
	.cin(gnd),
	.combout(\Equal5~1_combout ),
	.cout());
defparam \Equal5~1 .lut_mask = 16'hFFFE;
defparam \Equal5~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \k_count_wr_en~0 (
	.dataa(\k_count_wr_en~q ),
	.datab(gnd),
	.datac(\Equal5~0_combout ),
	.datad(\Equal5~1_combout ),
	.cin(gnd),
	.combout(\k_count_wr_en~0_combout ),
	.cout());
defparam \k_count_wr_en~0 .lut_mask = 16'hAFFF;
defparam \k_count_wr_en~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal4~0 (
	.dataa(\ctrl|k_count[1]~q ),
	.datab(\ctrl|k_count[6]~q ),
	.datac(\ctrl|k_count[3]~q ),
	.datad(\ctrl|k_count[5]~q ),
	.cin(gnd),
	.combout(\Equal4~0_combout ),
	.cout());
defparam \Equal4~0 .lut_mask = 16'hBFFF;
defparam \Equal4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal4~1 (
	.dataa(\ctrl|k_count[4]~q ),
	.datab(gnd),
	.datac(\ctrl|k_count[2]~q ),
	.datad(\ctrl|k_count[0]~q ),
	.cin(gnd),
	.combout(\Equal4~1_combout ),
	.cout());
defparam \Equal4~1 .lut_mask = 16'hAFFF;
defparam \Equal4~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \k_count_wr_en~1 (
	.dataa(\k_count_wr_en~0_combout ),
	.datab(\Equal4~0_combout ),
	.datac(\Equal4~1_combout ),
	.datad(\ctrl|k_count[7]~q ),
	.cin(gnd),
	.combout(\k_count_wr_en~1_combout ),
	.cout());
defparam \k_count_wr_en~1 .lut_mask = 16'hFEFF;
defparam \k_count_wr_en~1 .sum_lutc_input = "datac";

dffeas \p_tdl[16][0] (
	.clk(clk),
	.d(\p_tdl~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[16][0]~q ),
	.prn(vcc));
defparam \p_tdl[16][0] .is_wysiwyg = "true";
defparam \p_tdl[16][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~3 (
	.dataa(reset_n),
	.datab(\p_tdl[16][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~3_combout ),
	.cout());
defparam \p_tdl~3 .lut_mask = 16'hEEEE;
defparam \p_tdl~3 .sum_lutc_input = "datac";

dffeas \p_tdl[16][1] (
	.clk(clk),
	.d(\p_tdl~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[16][1]~q ),
	.prn(vcc));
defparam \p_tdl[16][1] .is_wysiwyg = "true";
defparam \p_tdl[16][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~4 (
	.dataa(reset_n),
	.datab(\p_tdl[16][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~4_combout ),
	.cout());
defparam \p_tdl~4 .lut_mask = 16'hEEEE;
defparam \p_tdl~4 .sum_lutc_input = "datac";

dffeas \p_tdl[16][2] (
	.clk(clk),
	.d(\p_tdl~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[16][2]~q ),
	.prn(vcc));
defparam \p_tdl[16][2] .is_wysiwyg = "true";
defparam \p_tdl[16][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~5 (
	.dataa(reset_n),
	.datab(\p_tdl[16][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~5_combout ),
	.cout());
defparam \p_tdl~5 .lut_mask = 16'hEEEE;
defparam \p_tdl~5 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[1] (
	.clk(clk),
	.d(\data_rdy_vec~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[1]~q ),
	.prn(vcc));
defparam \data_rdy_vec[1] .is_wysiwyg = "true";
defparam \data_rdy_vec[1] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~9 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~9_combout ),
	.cout());
defparam \data_rdy_vec~9 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~9 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[16] (
	.clk(clk),
	.d(\data_rdy_vec~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[16]~q ),
	.prn(vcc));
defparam \data_rdy_vec[16] .is_wysiwyg = "true";
defparam \data_rdy_vec[16] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~10 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~10_combout ),
	.cout());
defparam \data_rdy_vec~10 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~10 .sum_lutc_input = "datac";

dffeas \p_tdl[15][0] (
	.clk(clk),
	.d(\p_tdl~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[15][0]~q ),
	.prn(vcc));
defparam \p_tdl[15][0] .is_wysiwyg = "true";
defparam \p_tdl[15][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~6 (
	.dataa(reset_n),
	.datab(\p_tdl[15][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~6_combout ),
	.cout());
defparam \p_tdl~6 .lut_mask = 16'hEEEE;
defparam \p_tdl~6 .sum_lutc_input = "datac";

dffeas \p_tdl[15][1] (
	.clk(clk),
	.d(\p_tdl~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[15][1]~q ),
	.prn(vcc));
defparam \p_tdl[15][1] .is_wysiwyg = "true";
defparam \p_tdl[15][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~7 (
	.dataa(reset_n),
	.datab(\p_tdl[15][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~7_combout ),
	.cout());
defparam \p_tdl~7 .lut_mask = 16'hEEEE;
defparam \p_tdl~7 .sum_lutc_input = "datac";

dffeas \p_tdl[15][2] (
	.clk(clk),
	.d(\p_tdl~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[15][2]~q ),
	.prn(vcc));
defparam \p_tdl[15][2] .is_wysiwyg = "true";
defparam \p_tdl[15][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~8 (
	.dataa(reset_n),
	.datab(\p_tdl[15][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~8_combout ),
	.cout());
defparam \p_tdl~8 .lut_mask = 16'hEEEE;
defparam \p_tdl~8 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[0] (
	.clk(clk),
	.d(\data_rdy_vec~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[0]~q ),
	.prn(vcc));
defparam \data_rdy_vec[0] .is_wysiwyg = "true";
defparam \data_rdy_vec[0] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~11 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~11_combout ),
	.cout());
defparam \data_rdy_vec~11 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~11 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[15] (
	.clk(clk),
	.d(\data_rdy_vec~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[15]~q ),
	.prn(vcc));
defparam \data_rdy_vec[15] .is_wysiwyg = "true";
defparam \data_rdy_vec[15] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~12 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~12_combout ),
	.cout());
defparam \data_rdy_vec~12 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~12 .sum_lutc_input = "datac";

dffeas \p_tdl[14][0] (
	.clk(clk),
	.d(\p_tdl~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[14][0]~q ),
	.prn(vcc));
defparam \p_tdl[14][0] .is_wysiwyg = "true";
defparam \p_tdl[14][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~9 (
	.dataa(reset_n),
	.datab(\p_tdl[14][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~9_combout ),
	.cout());
defparam \p_tdl~9 .lut_mask = 16'hEEEE;
defparam \p_tdl~9 .sum_lutc_input = "datac";

dffeas \p_tdl[14][1] (
	.clk(clk),
	.d(\p_tdl~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[14][1]~q ),
	.prn(vcc));
defparam \p_tdl[14][1] .is_wysiwyg = "true";
defparam \p_tdl[14][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~10 (
	.dataa(reset_n),
	.datab(\p_tdl[14][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~10_combout ),
	.cout());
defparam \p_tdl~10 .lut_mask = 16'hEEEE;
defparam \p_tdl~10 .sum_lutc_input = "datac";

dffeas \p_tdl[14][2] (
	.clk(clk),
	.d(\p_tdl~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[14][2]~q ),
	.prn(vcc));
defparam \p_tdl[14][2] .is_wysiwyg = "true";
defparam \p_tdl[14][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~11 (
	.dataa(reset_n),
	.datab(\p_tdl[14][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~11_combout ),
	.cout());
defparam \p_tdl~11 .lut_mask = 16'hEEEE;
defparam \p_tdl~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_rdy_vec~13 (
	.dataa(reset_n),
	.datab(\writer|data_rdy_int~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~13_combout ),
	.cout());
defparam \data_rdy_vec~13 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~13 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[14] (
	.clk(clk),
	.d(\data_rdy_vec~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[14]~q ),
	.prn(vcc));
defparam \data_rdy_vec[14] .is_wysiwyg = "true";
defparam \data_rdy_vec[14] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~14 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~14_combout ),
	.cout());
defparam \data_rdy_vec~14 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~14 .sum_lutc_input = "datac";

dffeas \twiddle_data_real[1] (
	.clk(clk),
	.d(\twiddle_data_real~109_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_real[1]~q ),
	.prn(vcc));
defparam \twiddle_data_real[1] .is_wysiwyg = "true";
defparam \twiddle_data_real[1] .power_up = "low";

dffeas \twiddle_data_real[2] (
	.clk(clk),
	.d(\twiddle_data_real~110_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_real[2]~q ),
	.prn(vcc));
defparam \twiddle_data_real[2] .is_wysiwyg = "true";
defparam \twiddle_data_real[2] .power_up = "low";

dffeas \twiddle_data_real[3] (
	.clk(clk),
	.d(\twiddle_data_real~111_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_real[3]~q ),
	.prn(vcc));
defparam \twiddle_data_real[3] .is_wysiwyg = "true";
defparam \twiddle_data_real[3] .power_up = "low";

dffeas \twiddle_data_real[4] (
	.clk(clk),
	.d(\twiddle_data_real~112_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_real[4]~q ),
	.prn(vcc));
defparam \twiddle_data_real[4] .is_wysiwyg = "true";
defparam \twiddle_data_real[4] .power_up = "low";

dffeas \twiddle_data_real[5] (
	.clk(clk),
	.d(\twiddle_data_real~100_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_real[5]~q ),
	.prn(vcc));
defparam \twiddle_data_real[5] .is_wysiwyg = "true";
defparam \twiddle_data_real[5] .power_up = "low";

dffeas \twiddle_data_real[6] (
	.clk(clk),
	.d(\twiddle_data_real~101_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_real[6]~q ),
	.prn(vcc));
defparam \twiddle_data_real[6] .is_wysiwyg = "true";
defparam \twiddle_data_real[6] .power_up = "low";

dffeas \twiddle_data_real[7] (
	.clk(clk),
	.d(\twiddle_data_real~102_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_real[7]~q ),
	.prn(vcc));
defparam \twiddle_data_real[7] .is_wysiwyg = "true";
defparam \twiddle_data_real[7] .power_up = "low";

dffeas \twiddle_data_real[8] (
	.clk(clk),
	.d(\twiddle_data_real~103_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_real[8]~q ),
	.prn(vcc));
defparam \twiddle_data_real[8] .is_wysiwyg = "true";
defparam \twiddle_data_real[8] .power_up = "low";

dffeas \twiddle_data_real[9] (
	.clk(clk),
	.d(\twiddle_data_real~104_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_real[9]~q ),
	.prn(vcc));
defparam \twiddle_data_real[9] .is_wysiwyg = "true";
defparam \twiddle_data_real[9] .power_up = "low";

dffeas \twiddle_data_real[10] (
	.clk(clk),
	.d(\twiddle_data_real~105_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_real[10]~q ),
	.prn(vcc));
defparam \twiddle_data_real[10] .is_wysiwyg = "true";
defparam \twiddle_data_real[10] .power_up = "low";

dffeas \twiddle_data_real[11] (
	.clk(clk),
	.d(\twiddle_data_real~106_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_real[11]~q ),
	.prn(vcc));
defparam \twiddle_data_real[11] .is_wysiwyg = "true";
defparam \twiddle_data_real[11] .power_up = "low";

dffeas \twiddle_data_real[12] (
	.clk(clk),
	.d(\twiddle_data_real~107_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_real[12]~q ),
	.prn(vcc));
defparam \twiddle_data_real[12] .is_wysiwyg = "true";
defparam \twiddle_data_real[12] .power_up = "low";

dffeas \twiddle_data_real[13] (
	.clk(clk),
	.d(\twiddle_data_real~108_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_real[13]~q ),
	.prn(vcc));
defparam \twiddle_data_real[13] .is_wysiwyg = "true";
defparam \twiddle_data_real[13] .power_up = "low";

dffeas \twiddle_data_real[14] (
	.clk(clk),
	.d(\twiddle_data_real~113_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_real[14]~q ),
	.prn(vcc));
defparam \twiddle_data_real[14] .is_wysiwyg = "true";
defparam \twiddle_data_real[14] .power_up = "low";

dffeas \twiddle_data_imag[0] (
	.clk(clk),
	.d(\twiddle_data_imag~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\twiddle_data_imag[0]~q ),
	.prn(vcc));
defparam \twiddle_data_imag[0] .is_wysiwyg = "true";
defparam \twiddle_data_imag[0] .power_up = "low";

dffeas \p_tdl[13][0] (
	.clk(clk),
	.d(\p_tdl~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[13][0]~q ),
	.prn(vcc));
defparam \p_tdl[13][0] .is_wysiwyg = "true";
defparam \p_tdl[13][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~12 (
	.dataa(reset_n),
	.datab(\p_tdl[13][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~12_combout ),
	.cout());
defparam \p_tdl~12 .lut_mask = 16'hEEEE;
defparam \p_tdl~12 .sum_lutc_input = "datac";

dffeas \p_tdl[13][1] (
	.clk(clk),
	.d(\p_tdl~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[13][1]~q ),
	.prn(vcc));
defparam \p_tdl[13][1] .is_wysiwyg = "true";
defparam \p_tdl[13][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~13 (
	.dataa(reset_n),
	.datab(\p_tdl[13][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~13_combout ),
	.cout());
defparam \p_tdl~13 .lut_mask = 16'hEEEE;
defparam \p_tdl~13 .sum_lutc_input = "datac";

dffeas \p_tdl[13][2] (
	.clk(clk),
	.d(\p_tdl~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[13][2]~q ),
	.prn(vcc));
defparam \p_tdl[13][2] .is_wysiwyg = "true";
defparam \p_tdl[13][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~14 (
	.dataa(reset_n),
	.datab(\p_tdl[13][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~14_combout ),
	.cout());
defparam \p_tdl~14 .lut_mask = 16'hEEEE;
defparam \p_tdl~14 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[13] (
	.clk(clk),
	.d(\data_rdy_vec~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[13]~q ),
	.prn(vcc));
defparam \data_rdy_vec[13] .is_wysiwyg = "true";
defparam \data_rdy_vec[13] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~15 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~15_combout ),
	.cout());
defparam \data_rdy_vec~15 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~15 .sum_lutc_input = "datac";

dffeas \quad_del_1[2] (
	.clk(clk),
	.d(\quad_del_1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\quad_del_1[2]~q ),
	.prn(vcc));
defparam \quad_del_1[2] .is_wysiwyg = "true";
defparam \quad_del_1[2] .power_up = "low";

dffeas \quad_del_1[0] (
	.clk(clk),
	.d(\quad_del_1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\quad_del_1[0]~q ),
	.prn(vcc));
defparam \quad_del_1[0] .is_wysiwyg = "true";
defparam \quad_del_1[0] .power_up = "low";

dffeas \quad_del_1[1] (
	.clk(clk),
	.d(\quad_del_1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\quad_del_1[1]~q ),
	.prn(vcc));
defparam \quad_del_1[1] .is_wysiwyg = "true";
defparam \quad_del_1[1] .power_up = "low";

cycloneive_lcell_comb \Mux15~0 (
	.dataa(\quad_del_1[2]~q ),
	.datab(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[0] ),
	.datac(\quad_del_1[0]~q ),
	.datad(\quad_del_1[1]~q ),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
defparam \Mux15~0 .lut_mask = 16'hEFFE;
defparam \Mux15~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\quad_del_1[0]~q ),
	.datad(\quad_del_1[2]~q ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'h0FFF;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~1 (
	.dataa(\quad_del_1[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\quad_del_1[1]~q ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hAAFF;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~2 (
	.dataa(\Mux0~0_combout ),
	.datab(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[15] ),
	.datac(\quad_del_1[1]~q ),
	.datad(\Add2~30_combout ),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
defparam \Mux0~2 .lut_mask = 16'hFFAC;
defparam \Mux0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~3 (
	.dataa(\Mux0~1_combout ),
	.datab(\quad_del_1[0]~q ),
	.datac(\Add2~30_combout ),
	.datad(\Mux0~2_combout ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
defparam \Mux0~3 .lut_mask = 16'hFFFE;
defparam \Mux0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_imag~14 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[0] ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[0]~q ),
	.datad(\quad_del_1[2]~q ),
	.cin(gnd),
	.combout(\twiddle_data_imag~14_combout ),
	.cout());
defparam \twiddle_data_imag~14 .lut_mask = 16'hEFFE;
defparam \twiddle_data_imag~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_imag[14]~15 (
	.dataa(\quad_del_1[2]~q ),
	.datab(\quad_del_1[0]~q ),
	.datac(\quad_del_1[1]~q ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data_imag[14]~15_combout ),
	.cout());
defparam \twiddle_data_imag[14]~15 .lut_mask = 16'hFEFF;
defparam \twiddle_data_imag[14]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_imag~16 (
	.dataa(\twiddle_data_imag~14_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\twiddle_data_imag[14]~15_combout ),
	.cin(gnd),
	.combout(\twiddle_data_imag~16_combout ),
	.cout());
defparam \twiddle_data_imag~16 .lut_mask = 16'hAAFF;
defparam \twiddle_data_imag~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~0 (
	.dataa(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_a[15] ),
	.datab(gnd),
	.datac(gnd),
	.datad(\quad_del_1[2]~q ),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
defparam \Mux16~0 .lut_mask = 16'hAAFF;
defparam \Mux16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~1 (
	.dataa(\Mux16~0_combout ),
	.datab(\Mux0~1_combout ),
	.datac(\Add3~30_combout ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
defparam \Mux16~1 .lut_mask = 16'hFEFF;
defparam \Mux16~1 .sum_lutc_input = "datac";

dffeas \p_tdl[12][0] (
	.clk(clk),
	.d(\p_tdl~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[12][0]~q ),
	.prn(vcc));
defparam \p_tdl[12][0] .is_wysiwyg = "true";
defparam \p_tdl[12][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~15 (
	.dataa(reset_n),
	.datab(\p_tdl[12][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~15_combout ),
	.cout());
defparam \p_tdl~15 .lut_mask = 16'hEEEE;
defparam \p_tdl~15 .sum_lutc_input = "datac";

dffeas \p_tdl[12][1] (
	.clk(clk),
	.d(\p_tdl~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[12][1]~q ),
	.prn(vcc));
defparam \p_tdl[12][1] .is_wysiwyg = "true";
defparam \p_tdl[12][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~16 (
	.dataa(reset_n),
	.datab(\p_tdl[12][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~16_combout ),
	.cout());
defparam \p_tdl~16 .lut_mask = 16'hEEEE;
defparam \p_tdl~16 .sum_lutc_input = "datac";

dffeas \p_tdl[12][2] (
	.clk(clk),
	.d(\p_tdl~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[12][2]~q ),
	.prn(vcc));
defparam \p_tdl[12][2] .is_wysiwyg = "true";
defparam \p_tdl[12][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~17 (
	.dataa(reset_n),
	.datab(\p_tdl[12][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~17_combout ),
	.cout());
defparam \p_tdl~17 .lut_mask = 16'hEEEE;
defparam \p_tdl~17 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[12] (
	.clk(clk),
	.d(\data_rdy_vec~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[12]~q ),
	.prn(vcc));
defparam \data_rdy_vec[12] .is_wysiwyg = "true";
defparam \data_rdy_vec[12] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~16 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~16_combout ),
	.cout());
defparam \data_rdy_vec~16 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~16 .sum_lutc_input = "datac";

dffeas \quad_del_0[2] (
	.clk(clk),
	.d(\quad_del_0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\quad_del_0[2]~q ),
	.prn(vcc));
defparam \quad_del_0[2] .is_wysiwyg = "true";
defparam \quad_del_0[2] .power_up = "low";

cycloneive_lcell_comb \quad_del_1~0 (
	.dataa(reset_n),
	.datab(\quad_del_0[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\quad_del_1~0_combout ),
	.cout());
defparam \quad_del_1~0 .lut_mask = 16'hEEEE;
defparam \quad_del_1~0 .sum_lutc_input = "datac";

dffeas \quad_del_0[0] (
	.clk(clk),
	.d(\quad_del_0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\quad_del_0[0]~q ),
	.prn(vcc));
defparam \quad_del_0[0] .is_wysiwyg = "true";
defparam \quad_del_0[0] .power_up = "low";

cycloneive_lcell_comb \quad_del_1~1 (
	.dataa(reset_n),
	.datab(\quad_del_0[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\quad_del_1~1_combout ),
	.cout());
defparam \quad_del_1~1 .lut_mask = 16'hEEEE;
defparam \quad_del_1~1 .sum_lutc_input = "datac";

dffeas \quad_del_0[1] (
	.clk(clk),
	.d(\quad_del_0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\quad_del_0[1]~q ),
	.prn(vcc));
defparam \quad_del_0[1] .is_wysiwyg = "true";
defparam \quad_del_0[1] .power_up = "low";

cycloneive_lcell_comb \quad_del_1~2 (
	.dataa(reset_n),
	.datab(\quad_del_0[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\quad_del_1~2_combout ),
	.cout());
defparam \quad_del_1~2 .lut_mask = 16'hEEEE;
defparam \quad_del_1~2 .sum_lutc_input = "datac";

dffeas \p_tdl[11][0] (
	.clk(clk),
	.d(\p_tdl~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[11][0]~q ),
	.prn(vcc));
defparam \p_tdl[11][0] .is_wysiwyg = "true";
defparam \p_tdl[11][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~18 (
	.dataa(reset_n),
	.datab(\p_tdl[11][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~18_combout ),
	.cout());
defparam \p_tdl~18 .lut_mask = 16'hEEEE;
defparam \p_tdl~18 .sum_lutc_input = "datac";

dffeas \p_tdl[11][1] (
	.clk(clk),
	.d(\p_tdl~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[11][1]~q ),
	.prn(vcc));
defparam \p_tdl[11][1] .is_wysiwyg = "true";
defparam \p_tdl[11][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~19 (
	.dataa(reset_n),
	.datab(\p_tdl[11][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~19_combout ),
	.cout());
defparam \p_tdl~19 .lut_mask = 16'hEEEE;
defparam \p_tdl~19 .sum_lutc_input = "datac";

dffeas \p_tdl[11][2] (
	.clk(clk),
	.d(\p_tdl~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[11][2]~q ),
	.prn(vcc));
defparam \p_tdl[11][2] .is_wysiwyg = "true";
defparam \p_tdl[11][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~20 (
	.dataa(reset_n),
	.datab(\p_tdl[11][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~20_combout ),
	.cout());
defparam \p_tdl~20 .lut_mask = 16'hEEEE;
defparam \p_tdl~20 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[11] (
	.clk(clk),
	.d(\data_rdy_vec~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[11]~q ),
	.prn(vcc));
defparam \data_rdy_vec[11] .is_wysiwyg = "true";
defparam \data_rdy_vec[11] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~17 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~17_combout ),
	.cout());
defparam \data_rdy_vec~17 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \quad_del_0~0 (
	.dataa(reset_n),
	.datab(\gen_se:gen_new:twid_factors|quad_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\quad_del_0~0_combout ),
	.cout());
defparam \quad_del_0~0 .lut_mask = 16'hEEEE;
defparam \quad_del_0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \quad_del_0~1 (
	.dataa(reset_n),
	.datab(\gen_se:gen_new:twid_factors|quad_reg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\quad_del_0~1_combout ),
	.cout());
defparam \quad_del_0~1 .lut_mask = 16'hEEEE;
defparam \quad_del_0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \quad_del_0~2 (
	.dataa(reset_n),
	.datab(\gen_se:gen_new:twid_factors|quad_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\quad_del_0~2_combout ),
	.cout());
defparam \quad_del_0~2 .lut_mask = 16'hEEEE;
defparam \quad_del_0~2 .sum_lutc_input = "datac";

dffeas \p_tdl[10][0] (
	.clk(clk),
	.d(\p_tdl~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[10][0]~q ),
	.prn(vcc));
defparam \p_tdl[10][0] .is_wysiwyg = "true";
defparam \p_tdl[10][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~21 (
	.dataa(reset_n),
	.datab(\p_tdl[10][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~21_combout ),
	.cout());
defparam \p_tdl~21 .lut_mask = 16'hEEEE;
defparam \p_tdl~21 .sum_lutc_input = "datac";

dffeas \p_tdl[10][1] (
	.clk(clk),
	.d(\p_tdl~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[10][1]~q ),
	.prn(vcc));
defparam \p_tdl[10][1] .is_wysiwyg = "true";
defparam \p_tdl[10][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~22 (
	.dataa(reset_n),
	.datab(\p_tdl[10][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~22_combout ),
	.cout());
defparam \p_tdl~22 .lut_mask = 16'hEEEE;
defparam \p_tdl~22 .sum_lutc_input = "datac";

dffeas \p_tdl[10][2] (
	.clk(clk),
	.d(\p_tdl~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[10][2]~q ),
	.prn(vcc));
defparam \p_tdl[10][2] .is_wysiwyg = "true";
defparam \p_tdl[10][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~23 (
	.dataa(reset_n),
	.datab(\p_tdl[10][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~23_combout ),
	.cout());
defparam \p_tdl~23 .lut_mask = 16'hEEEE;
defparam \p_tdl~23 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[27] (
	.clk(clk),
	.d(\data_rdy_vec~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[27]~q ),
	.prn(vcc));
defparam \data_rdy_vec[27] .is_wysiwyg = "true";
defparam \data_rdy_vec[27] .power_up = "low";

cycloneive_lcell_comb next_pass(
	.dataa(\ctrl|next_pass_i~q ),
	.datab(\data_rdy_vec[27]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pass~combout ),
	.cout());
defparam next_pass.lut_mask = 16'hEEEE;
defparam next_pass.sum_lutc_input = "datac";

dffeas \data_rdy_vec[10] (
	.clk(clk),
	.d(\data_rdy_vec~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[10]~q ),
	.prn(vcc));
defparam \data_rdy_vec[10] .is_wysiwyg = "true";
defparam \data_rdy_vec[10] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~18 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~18_combout ),
	.cout());
defparam \data_rdy_vec~18 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~18 .sum_lutc_input = "datac";

dffeas \p_tdl[9][0] (
	.clk(clk),
	.d(\p_tdl~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[9][0]~q ),
	.prn(vcc));
defparam \p_tdl[9][0] .is_wysiwyg = "true";
defparam \p_tdl[9][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~24 (
	.dataa(reset_n),
	.datab(\p_tdl[9][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~24_combout ),
	.cout());
defparam \p_tdl~24 .lut_mask = 16'hEEEE;
defparam \p_tdl~24 .sum_lutc_input = "datac";

dffeas \p_tdl[9][1] (
	.clk(clk),
	.d(\p_tdl~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[9][1]~q ),
	.prn(vcc));
defparam \p_tdl[9][1] .is_wysiwyg = "true";
defparam \p_tdl[9][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~25 (
	.dataa(reset_n),
	.datab(\p_tdl[9][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~25_combout ),
	.cout());
defparam \p_tdl~25 .lut_mask = 16'hEEEE;
defparam \p_tdl~25 .sum_lutc_input = "datac";

dffeas \p_tdl[9][2] (
	.clk(clk),
	.d(\p_tdl~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[9][2]~q ),
	.prn(vcc));
defparam \p_tdl[9][2] .is_wysiwyg = "true";
defparam \p_tdl[9][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~26 (
	.dataa(reset_n),
	.datab(\p_tdl[9][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~26_combout ),
	.cout());
defparam \p_tdl~26 .lut_mask = 16'hEEEE;
defparam \p_tdl~26 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[26] (
	.clk(clk),
	.d(\data_rdy_vec~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[26]~q ),
	.prn(vcc));
defparam \data_rdy_vec[26] .is_wysiwyg = "true";
defparam \data_rdy_vec[26] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~19 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[26]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~19_combout ),
	.cout());
defparam \data_rdy_vec~19 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~19 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[9] (
	.clk(clk),
	.d(\data_rdy_vec~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[9]~q ),
	.prn(vcc));
defparam \data_rdy_vec[9] .is_wysiwyg = "true";
defparam \data_rdy_vec[9] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~20 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~20_combout ),
	.cout());
defparam \data_rdy_vec~20 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~20 .sum_lutc_input = "datac";

dffeas \p_tdl[8][0] (
	.clk(clk),
	.d(\p_tdl~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[8][0]~q ),
	.prn(vcc));
defparam \p_tdl[8][0] .is_wysiwyg = "true";
defparam \p_tdl[8][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~27 (
	.dataa(reset_n),
	.datab(\p_tdl[8][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~27_combout ),
	.cout());
defparam \p_tdl~27 .lut_mask = 16'hEEEE;
defparam \p_tdl~27 .sum_lutc_input = "datac";

dffeas \p_tdl[8][1] (
	.clk(clk),
	.d(\p_tdl~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[8][1]~q ),
	.prn(vcc));
defparam \p_tdl[8][1] .is_wysiwyg = "true";
defparam \p_tdl[8][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~28 (
	.dataa(reset_n),
	.datab(\p_tdl[8][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~28_combout ),
	.cout());
defparam \p_tdl~28 .lut_mask = 16'hEEEE;
defparam \p_tdl~28 .sum_lutc_input = "datac";

dffeas \p_tdl[8][2] (
	.clk(clk),
	.d(\p_tdl~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[8][2]~q ),
	.prn(vcc));
defparam \p_tdl[8][2] .is_wysiwyg = "true";
defparam \p_tdl[8][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~29 (
	.dataa(reset_n),
	.datab(\p_tdl[8][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~29_combout ),
	.cout());
defparam \p_tdl~29 .lut_mask = 16'hEEEE;
defparam \p_tdl~29 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[25] (
	.clk(clk),
	.d(\data_rdy_vec~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[25]~q ),
	.prn(vcc));
defparam \data_rdy_vec[25] .is_wysiwyg = "true";
defparam \data_rdy_vec[25] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~21 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[25]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~21_combout ),
	.cout());
defparam \data_rdy_vec~21 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~21 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[8] (
	.clk(clk),
	.d(\data_rdy_vec~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[8]~q ),
	.prn(vcc));
defparam \data_rdy_vec[8] .is_wysiwyg = "true";
defparam \data_rdy_vec[8] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~22 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~22_combout ),
	.cout());
defparam \data_rdy_vec~22 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~22 .sum_lutc_input = "datac";

dffeas \p_tdl[7][0] (
	.clk(clk),
	.d(\p_tdl~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[7][0]~q ),
	.prn(vcc));
defparam \p_tdl[7][0] .is_wysiwyg = "true";
defparam \p_tdl[7][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~30 (
	.dataa(reset_n),
	.datab(\p_tdl[7][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~30_combout ),
	.cout());
defparam \p_tdl~30 .lut_mask = 16'hEEEE;
defparam \p_tdl~30 .sum_lutc_input = "datac";

dffeas \p_tdl[7][1] (
	.clk(clk),
	.d(\p_tdl~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[7][1]~q ),
	.prn(vcc));
defparam \p_tdl[7][1] .is_wysiwyg = "true";
defparam \p_tdl[7][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~31 (
	.dataa(reset_n),
	.datab(\p_tdl[7][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~31_combout ),
	.cout());
defparam \p_tdl~31 .lut_mask = 16'hEEEE;
defparam \p_tdl~31 .sum_lutc_input = "datac";

dffeas \p_tdl[7][2] (
	.clk(clk),
	.d(\p_tdl~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[7][2]~q ),
	.prn(vcc));
defparam \p_tdl[7][2] .is_wysiwyg = "true";
defparam \p_tdl[7][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~32 (
	.dataa(reset_n),
	.datab(\p_tdl[7][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~32_combout ),
	.cout());
defparam \p_tdl~32 .lut_mask = 16'hEEEE;
defparam \p_tdl~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_rdy_vec~23 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[24]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~23_combout ),
	.cout());
defparam \data_rdy_vec~23 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~23 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[7] (
	.clk(clk),
	.d(\data_rdy_vec~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[7]~q ),
	.prn(vcc));
defparam \data_rdy_vec[7] .is_wysiwyg = "true";
defparam \data_rdy_vec[7] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~24 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~24_combout ),
	.cout());
defparam \data_rdy_vec~24 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal7~0 (
	.dataa(\k_count_tw[7]~q ),
	.datab(\k_count_tw[6]~q ),
	.datac(\k_count_tw[5]~q ),
	.datad(\k_count_tw[4]~q ),
	.cin(gnd),
	.combout(\Equal7~0_combout ),
	.cout());
defparam \Equal7~0 .lut_mask = 16'hFFFE;
defparam \Equal7~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \k_count_tw_en~0 (
	.dataa(\k_count_tw_en~q ),
	.datab(\gen_se:gen_new:twid_factors|data_addr_held_by1~0_combout ),
	.datac(\gen_se:gen_new:twid_factors|data_addr_held_by2~0_combout ),
	.datad(\Equal7~0_combout ),
	.cin(gnd),
	.combout(\k_count_tw_en~0_combout ),
	.cout());
defparam \k_count_tw_en~0 .lut_mask = 16'hBFFF;
defparam \k_count_tw_en~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~0 (
	.dataa(\ctrl|k_count[2]~q ),
	.datab(\ctrl|k_count[0]~q ),
	.datac(gnd),
	.datad(\ctrl|k_count[4]~q ),
	.cin(gnd),
	.combout(\Equal6~0_combout ),
	.cout());
defparam \Equal6~0 .lut_mask = 16'hEEFF;
defparam \Equal6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \k_count_tw_en~1 (
	.dataa(\k_count_tw_en~0_combout ),
	.datab(\Equal4~0_combout ),
	.datac(\Equal6~0_combout ),
	.datad(\ctrl|k_count[7]~q ),
	.cin(gnd),
	.combout(\k_count_tw_en~1_combout ),
	.cout());
defparam \k_count_tw_en~1 .lut_mask = 16'hFEFF;
defparam \k_count_tw_en~1 .sum_lutc_input = "datac";

dffeas \p_tdl[6][0] (
	.clk(clk),
	.d(\p_tdl~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[6][0]~q ),
	.prn(vcc));
defparam \p_tdl[6][0] .is_wysiwyg = "true";
defparam \p_tdl[6][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~33 (
	.dataa(reset_n),
	.datab(\p_tdl[6][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~33_combout ),
	.cout());
defparam \p_tdl~33 .lut_mask = 16'hEEEE;
defparam \p_tdl~33 .sum_lutc_input = "datac";

dffeas \p_tdl[6][1] (
	.clk(clk),
	.d(\p_tdl~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[6][1]~q ),
	.prn(vcc));
defparam \p_tdl[6][1] .is_wysiwyg = "true";
defparam \p_tdl[6][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~34 (
	.dataa(reset_n),
	.datab(\p_tdl[6][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~34_combout ),
	.cout());
defparam \p_tdl~34 .lut_mask = 16'hEEEE;
defparam \p_tdl~34 .sum_lutc_input = "datac";

dffeas \p_tdl[6][2] (
	.clk(clk),
	.d(\p_tdl~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[6][2]~q ),
	.prn(vcc));
defparam \p_tdl[6][2] .is_wysiwyg = "true";
defparam \p_tdl[6][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~35 (
	.dataa(reset_n),
	.datab(\p_tdl[6][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~35_combout ),
	.cout());
defparam \p_tdl~35 .lut_mask = 16'hEEEE;
defparam \p_tdl~35 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[6] (
	.clk(clk),
	.d(\data_rdy_vec~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[6]~q ),
	.prn(vcc));
defparam \data_rdy_vec[6] .is_wysiwyg = "true";
defparam \data_rdy_vec[6] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~25 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~25_combout ),
	.cout());
defparam \data_rdy_vec~25 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~25 .sum_lutc_input = "datac";

dffeas \p_tdl[5][0] (
	.clk(clk),
	.d(\p_tdl~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[5][0]~q ),
	.prn(vcc));
defparam \p_tdl[5][0] .is_wysiwyg = "true";
defparam \p_tdl[5][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~36 (
	.dataa(reset_n),
	.datab(\p_tdl[5][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~36_combout ),
	.cout());
defparam \p_tdl~36 .lut_mask = 16'hEEEE;
defparam \p_tdl~36 .sum_lutc_input = "datac";

dffeas \p_tdl[5][1] (
	.clk(clk),
	.d(\p_tdl~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[5][1]~q ),
	.prn(vcc));
defparam \p_tdl[5][1] .is_wysiwyg = "true";
defparam \p_tdl[5][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~37 (
	.dataa(reset_n),
	.datab(\p_tdl[5][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~37_combout ),
	.cout());
defparam \p_tdl~37 .lut_mask = 16'hEEEE;
defparam \p_tdl~37 .sum_lutc_input = "datac";

dffeas \p_tdl[5][2] (
	.clk(clk),
	.d(\p_tdl~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[5][2]~q ),
	.prn(vcc));
defparam \p_tdl[5][2] .is_wysiwyg = "true";
defparam \p_tdl[5][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~38 (
	.dataa(reset_n),
	.datab(\p_tdl[5][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~38_combout ),
	.cout());
defparam \p_tdl~38 .lut_mask = 16'hEEEE;
defparam \p_tdl~38 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[5] (
	.clk(clk),
	.d(\data_rdy_vec~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[5]~q ),
	.prn(vcc));
defparam \data_rdy_vec[5] .is_wysiwyg = "true";
defparam \data_rdy_vec[5] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~26 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~26_combout ),
	.cout());
defparam \data_rdy_vec~26 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~26 .sum_lutc_input = "datac";

dffeas \p_tdl[4][0] (
	.clk(clk),
	.d(\p_tdl~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[4][0]~q ),
	.prn(vcc));
defparam \p_tdl[4][0] .is_wysiwyg = "true";
defparam \p_tdl[4][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~39 (
	.dataa(reset_n),
	.datab(\p_tdl[4][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~39_combout ),
	.cout());
defparam \p_tdl~39 .lut_mask = 16'hEEEE;
defparam \p_tdl~39 .sum_lutc_input = "datac";

dffeas \p_tdl[4][1] (
	.clk(clk),
	.d(\p_tdl~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[4][1]~q ),
	.prn(vcc));
defparam \p_tdl[4][1] .is_wysiwyg = "true";
defparam \p_tdl[4][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~40 (
	.dataa(reset_n),
	.datab(\p_tdl[4][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~40_combout ),
	.cout());
defparam \p_tdl~40 .lut_mask = 16'hEEEE;
defparam \p_tdl~40 .sum_lutc_input = "datac";

dffeas \p_tdl[4][2] (
	.clk(clk),
	.d(\p_tdl~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[4][2]~q ),
	.prn(vcc));
defparam \p_tdl[4][2] .is_wysiwyg = "true";
defparam \p_tdl[4][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~41 (
	.dataa(reset_n),
	.datab(\p_tdl[4][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~41_combout ),
	.cout());
defparam \p_tdl~41 .lut_mask = 16'hEEEE;
defparam \p_tdl~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_rdy_vec~27 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~27_combout ),
	.cout());
defparam \data_rdy_vec~27 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~27 .sum_lutc_input = "datac";

dffeas \p_tdl[3][0] (
	.clk(clk),
	.d(\p_tdl~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[3][0]~q ),
	.prn(vcc));
defparam \p_tdl[3][0] .is_wysiwyg = "true";
defparam \p_tdl[3][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~42 (
	.dataa(reset_n),
	.datab(\p_tdl[3][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~42_combout ),
	.cout());
defparam \p_tdl~42 .lut_mask = 16'hEEEE;
defparam \p_tdl~42 .sum_lutc_input = "datac";

dffeas \p_tdl[3][1] (
	.clk(clk),
	.d(\p_tdl~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[3][1]~q ),
	.prn(vcc));
defparam \p_tdl[3][1] .is_wysiwyg = "true";
defparam \p_tdl[3][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~43 (
	.dataa(reset_n),
	.datab(\p_tdl[3][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~43_combout ),
	.cout());
defparam \p_tdl~43 .lut_mask = 16'hEEEE;
defparam \p_tdl~43 .sum_lutc_input = "datac";

dffeas \p_tdl[3][2] (
	.clk(clk),
	.d(\p_tdl~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[3][2]~q ),
	.prn(vcc));
defparam \p_tdl[3][2] .is_wysiwyg = "true";
defparam \p_tdl[3][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~44 (
	.dataa(reset_n),
	.datab(\p_tdl[3][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~44_combout ),
	.cout());
defparam \p_tdl~44 .lut_mask = 16'hEEEE;
defparam \p_tdl~44 .sum_lutc_input = "datac";

dffeas \p_tdl[2][0] (
	.clk(clk),
	.d(\p_tdl~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[2][0]~q ),
	.prn(vcc));
defparam \p_tdl[2][0] .is_wysiwyg = "true";
defparam \p_tdl[2][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~45 (
	.dataa(reset_n),
	.datab(\p_tdl[2][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~45_combout ),
	.cout());
defparam \p_tdl~45 .lut_mask = 16'hEEEE;
defparam \p_tdl~45 .sum_lutc_input = "datac";

dffeas \p_tdl[2][1] (
	.clk(clk),
	.d(\p_tdl~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[2][1]~q ),
	.prn(vcc));
defparam \p_tdl[2][1] .is_wysiwyg = "true";
defparam \p_tdl[2][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~46 (
	.dataa(reset_n),
	.datab(\p_tdl[2][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~46_combout ),
	.cout());
defparam \p_tdl~46 .lut_mask = 16'hEEEE;
defparam \p_tdl~46 .sum_lutc_input = "datac";

dffeas \p_tdl[2][2] (
	.clk(clk),
	.d(\p_tdl~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[2][2]~q ),
	.prn(vcc));
defparam \p_tdl[2][2] .is_wysiwyg = "true";
defparam \p_tdl[2][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~47 (
	.dataa(reset_n),
	.datab(\p_tdl[2][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~47_combout ),
	.cout());
defparam \p_tdl~47 .lut_mask = 16'hEEEE;
defparam \p_tdl~47 .sum_lutc_input = "datac";

dffeas \p_tdl[1][0] (
	.clk(clk),
	.d(\p_tdl~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[1][0]~q ),
	.prn(vcc));
defparam \p_tdl[1][0] .is_wysiwyg = "true";
defparam \p_tdl[1][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~48 (
	.dataa(reset_n),
	.datab(\p_tdl[1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~48_combout ),
	.cout());
defparam \p_tdl~48 .lut_mask = 16'hEEEE;
defparam \p_tdl~48 .sum_lutc_input = "datac";

dffeas \p_tdl[1][1] (
	.clk(clk),
	.d(\p_tdl~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[1][1]~q ),
	.prn(vcc));
defparam \p_tdl[1][1] .is_wysiwyg = "true";
defparam \p_tdl[1][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~49 (
	.dataa(reset_n),
	.datab(\p_tdl[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~49_combout ),
	.cout());
defparam \p_tdl~49 .lut_mask = 16'hEEEE;
defparam \p_tdl~49 .sum_lutc_input = "datac";

dffeas \p_tdl[1][2] (
	.clk(clk),
	.d(\p_tdl~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[1][2]~q ),
	.prn(vcc));
defparam \p_tdl[1][2] .is_wysiwyg = "true";
defparam \p_tdl[1][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~50 (
	.dataa(reset_n),
	.datab(\p_tdl[1][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~50_combout ),
	.cout());
defparam \p_tdl~50 .lut_mask = 16'hEEEE;
defparam \p_tdl~50 .sum_lutc_input = "datac";

dffeas \p_tdl[0][0] (
	.clk(clk),
	.d(\p_tdl~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[0][0]~q ),
	.prn(vcc));
defparam \p_tdl[0][0] .is_wysiwyg = "true";
defparam \p_tdl[0][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~51 (
	.dataa(reset_n),
	.datab(\p_tdl[0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~51_combout ),
	.cout());
defparam \p_tdl~51 .lut_mask = 16'hEEEE;
defparam \p_tdl~51 .sum_lutc_input = "datac";

dffeas \p_tdl[0][1] (
	.clk(clk),
	.d(\p_tdl~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[0][1]~q ),
	.prn(vcc));
defparam \p_tdl[0][1] .is_wysiwyg = "true";
defparam \p_tdl[0][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~52 (
	.dataa(reset_n),
	.datab(\p_tdl[0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~52_combout ),
	.cout());
defparam \p_tdl~52 .lut_mask = 16'hEEEE;
defparam \p_tdl~52 .sum_lutc_input = "datac";

dffeas \p_tdl[0][2] (
	.clk(clk),
	.d(\p_tdl~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~0_combout ),
	.q(\p_tdl[0][2]~q ),
	.prn(vcc));
defparam \p_tdl[0][2] .is_wysiwyg = "true";
defparam \p_tdl[0][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~53 (
	.dataa(reset_n),
	.datab(\p_tdl[0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~53_combout ),
	.cout());
defparam \p_tdl~53 .lut_mask = 16'hEEEE;
defparam \p_tdl~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p_tdl~54 (
	.dataa(reset_n),
	.datab(\ctrl|p[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~54_combout ),
	.cout());
defparam \p_tdl~54 .lut_mask = 16'hEEEE;
defparam \p_tdl~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p_tdl~55 (
	.dataa(reset_n),
	.datab(\ctrl|p[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~55_combout ),
	.cout());
defparam \p_tdl~55 .lut_mask = 16'hEEEE;
defparam \p_tdl~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p_tdl~56 (
	.dataa(reset_n),
	.datab(\ctrl|p[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~56_combout ),
	.cout());
defparam \p_tdl~56 .lut_mask = 16'hEEEE;
defparam \p_tdl~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~5 (
	.dataa(\Add2~10_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~5_combout ),
	.cout());
defparam \twiddle_data_real~5 .lut_mask = 16'hEBBE;
defparam \twiddle_data_real~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~6 (
	.dataa(\Add2~10_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~6_combout ),
	.cout());
defparam \twiddle_data_real~6 .lut_mask = 16'hBEFF;
defparam \twiddle_data_real~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~100 (
	.dataa(\twiddle_data_real~5_combout ),
	.datab(\twiddle_data_real~6_combout ),
	.datac(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[5] ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data_real~100_combout ),
	.cout());
defparam \twiddle_data_real~100 .lut_mask = 16'hACFF;
defparam \twiddle_data_real~100 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~12 (
	.dataa(\Add2~12_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~12_combout ),
	.cout());
defparam \twiddle_data_real~12 .lut_mask = 16'hEBBE;
defparam \twiddle_data_real~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~13 (
	.dataa(\Add2~12_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~13_combout ),
	.cout());
defparam \twiddle_data_real~13 .lut_mask = 16'hBEFF;
defparam \twiddle_data_real~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~101 (
	.dataa(\twiddle_data_real~12_combout ),
	.datab(\twiddle_data_real~13_combout ),
	.datac(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[6] ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data_real~101_combout ),
	.cout());
defparam \twiddle_data_real~101 .lut_mask = 16'hACFF;
defparam \twiddle_data_real~101 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~19 (
	.dataa(\Add2~14_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~19_combout ),
	.cout());
defparam \twiddle_data_real~19 .lut_mask = 16'hEBBE;
defparam \twiddle_data_real~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~20 (
	.dataa(\Add2~14_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~20_combout ),
	.cout());
defparam \twiddle_data_real~20 .lut_mask = 16'hBEFF;
defparam \twiddle_data_real~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~102 (
	.dataa(\twiddle_data_real~19_combout ),
	.datab(\twiddle_data_real~20_combout ),
	.datac(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[7] ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data_real~102_combout ),
	.cout());
defparam \twiddle_data_real~102 .lut_mask = 16'hACFF;
defparam \twiddle_data_real~102 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~26 (
	.dataa(\Add2~16_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~26_combout ),
	.cout());
defparam \twiddle_data_real~26 .lut_mask = 16'hEBBE;
defparam \twiddle_data_real~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~27 (
	.dataa(\Add2~16_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~27_combout ),
	.cout());
defparam \twiddle_data_real~27 .lut_mask = 16'hBEFF;
defparam \twiddle_data_real~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~103 (
	.dataa(\twiddle_data_real~26_combout ),
	.datab(\twiddle_data_real~27_combout ),
	.datac(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[8] ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data_real~103_combout ),
	.cout());
defparam \twiddle_data_real~103 .lut_mask = 16'hACFF;
defparam \twiddle_data_real~103 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~33 (
	.dataa(\Add2~18_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~33_combout ),
	.cout());
defparam \twiddle_data_real~33 .lut_mask = 16'hEBBE;
defparam \twiddle_data_real~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~34 (
	.dataa(\Add2~18_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~34_combout ),
	.cout());
defparam \twiddle_data_real~34 .lut_mask = 16'hBEFF;
defparam \twiddle_data_real~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~104 (
	.dataa(\twiddle_data_real~33_combout ),
	.datab(\twiddle_data_real~34_combout ),
	.datac(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[9] ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data_real~104_combout ),
	.cout());
defparam \twiddle_data_real~104 .lut_mask = 16'hACFF;
defparam \twiddle_data_real~104 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~40 (
	.dataa(\Add2~20_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~40_combout ),
	.cout());
defparam \twiddle_data_real~40 .lut_mask = 16'hEBBE;
defparam \twiddle_data_real~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~41 (
	.dataa(\Add2~20_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~41_combout ),
	.cout());
defparam \twiddle_data_real~41 .lut_mask = 16'hBEFF;
defparam \twiddle_data_real~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~105 (
	.dataa(\twiddle_data_real~40_combout ),
	.datab(\twiddle_data_real~41_combout ),
	.datac(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[10] ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data_real~105_combout ),
	.cout());
defparam \twiddle_data_real~105 .lut_mask = 16'hACFF;
defparam \twiddle_data_real~105 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~47 (
	.dataa(\Add2~22_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~47_combout ),
	.cout());
defparam \twiddle_data_real~47 .lut_mask = 16'hEBBE;
defparam \twiddle_data_real~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~48 (
	.dataa(\Add2~22_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~48_combout ),
	.cout());
defparam \twiddle_data_real~48 .lut_mask = 16'hBEFF;
defparam \twiddle_data_real~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~106 (
	.dataa(\twiddle_data_real~47_combout ),
	.datab(\twiddle_data_real~48_combout ),
	.datac(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[11] ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data_real~106_combout ),
	.cout());
defparam \twiddle_data_real~106 .lut_mask = 16'hACFF;
defparam \twiddle_data_real~106 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~54 (
	.dataa(\Add2~24_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~54_combout ),
	.cout());
defparam \twiddle_data_real~54 .lut_mask = 16'hEBBE;
defparam \twiddle_data_real~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~55 (
	.dataa(\Add2~24_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~55_combout ),
	.cout());
defparam \twiddle_data_real~55 .lut_mask = 16'hBEFF;
defparam \twiddle_data_real~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~107 (
	.dataa(\twiddle_data_real~54_combout ),
	.datab(\twiddle_data_real~55_combout ),
	.datac(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[12] ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data_real~107_combout ),
	.cout());
defparam \twiddle_data_real~107 .lut_mask = 16'hACFF;
defparam \twiddle_data_real~107 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~61 (
	.dataa(\Add2~26_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~61_combout ),
	.cout());
defparam \twiddle_data_real~61 .lut_mask = 16'hEBBE;
defparam \twiddle_data_real~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~62 (
	.dataa(\Add2~26_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~62_combout ),
	.cout());
defparam \twiddle_data_real~62 .lut_mask = 16'hBEFF;
defparam \twiddle_data_real~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~108 (
	.dataa(\twiddle_data_real~61_combout ),
	.datab(\twiddle_data_real~62_combout ),
	.datac(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[13] ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data_real~108_combout ),
	.cout());
defparam \twiddle_data_real~108 .lut_mask = 16'hACFF;
defparam \twiddle_data_real~108 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~68 (
	.dataa(\quad_del_1[1]~q ),
	.datab(\quad_del_1[2]~q ),
	.datac(\quad_del_1[0]~q ),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\twiddle_data_real~68_combout ),
	.cout());
defparam \twiddle_data_real~68 .lut_mask = 16'hFF96;
defparam \twiddle_data_real~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~69 (
	.dataa(\quad_del_1[1]~q ),
	.datab(\quad_del_1[2]~q ),
	.datac(\quad_del_1[0]~q ),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\twiddle_data_real~69_combout ),
	.cout());
defparam \twiddle_data_real~69 .lut_mask = 16'hFF6F;
defparam \twiddle_data_real~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~109 (
	.dataa(\twiddle_data_real~68_combout ),
	.datab(\twiddle_data_real~69_combout ),
	.datac(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[1] ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data_real~109_combout ),
	.cout());
defparam \twiddle_data_real~109 .lut_mask = 16'hACFF;
defparam \twiddle_data_real~109 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~75 (
	.dataa(\quad_del_1[1]~q ),
	.datab(\quad_del_1[2]~q ),
	.datac(\quad_del_1[0]~q ),
	.datad(\Add2~4_combout ),
	.cin(gnd),
	.combout(\twiddle_data_real~75_combout ),
	.cout());
defparam \twiddle_data_real~75 .lut_mask = 16'hFF96;
defparam \twiddle_data_real~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~76 (
	.dataa(\quad_del_1[1]~q ),
	.datab(\quad_del_1[2]~q ),
	.datac(\quad_del_1[0]~q ),
	.datad(\Add2~4_combout ),
	.cin(gnd),
	.combout(\twiddle_data_real~76_combout ),
	.cout());
defparam \twiddle_data_real~76 .lut_mask = 16'hFF6F;
defparam \twiddle_data_real~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~110 (
	.dataa(\twiddle_data_real~75_combout ),
	.datab(\twiddle_data_real~76_combout ),
	.datac(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[2] ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data_real~110_combout ),
	.cout());
defparam \twiddle_data_real~110 .lut_mask = 16'hACFF;
defparam \twiddle_data_real~110 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~82 (
	.dataa(\quad_del_1[1]~q ),
	.datab(\quad_del_1[2]~q ),
	.datac(\quad_del_1[0]~q ),
	.datad(\Add2~6_combout ),
	.cin(gnd),
	.combout(\twiddle_data_real~82_combout ),
	.cout());
defparam \twiddle_data_real~82 .lut_mask = 16'hFF96;
defparam \twiddle_data_real~82 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~83 (
	.dataa(\quad_del_1[1]~q ),
	.datab(\quad_del_1[2]~q ),
	.datac(\quad_del_1[0]~q ),
	.datad(\Add2~6_combout ),
	.cin(gnd),
	.combout(\twiddle_data_real~83_combout ),
	.cout());
defparam \twiddle_data_real~83 .lut_mask = 16'hFF6F;
defparam \twiddle_data_real~83 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~111 (
	.dataa(\twiddle_data_real~82_combout ),
	.datab(\twiddle_data_real~83_combout ),
	.datac(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[3] ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data_real~111_combout ),
	.cout());
defparam \twiddle_data_real~111 .lut_mask = 16'hACFF;
defparam \twiddle_data_real~111 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~89 (
	.dataa(\quad_del_1[1]~q ),
	.datab(\quad_del_1[2]~q ),
	.datac(\quad_del_1[0]~q ),
	.datad(\Add2~8_combout ),
	.cin(gnd),
	.combout(\twiddle_data_real~89_combout ),
	.cout());
defparam \twiddle_data_real~89 .lut_mask = 16'hFF96;
defparam \twiddle_data_real~89 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~90 (
	.dataa(\quad_del_1[1]~q ),
	.datab(\quad_del_1[2]~q ),
	.datac(\quad_del_1[0]~q ),
	.datad(\Add2~8_combout ),
	.cin(gnd),
	.combout(\twiddle_data_real~90_combout ),
	.cout());
defparam \twiddle_data_real~90 .lut_mask = 16'hFF6F;
defparam \twiddle_data_real~90 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~112 (
	.dataa(\twiddle_data_real~89_combout ),
	.datab(\twiddle_data_real~90_combout ),
	.datac(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[4] ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data_real~112_combout ),
	.cout());
defparam \twiddle_data_real~112 .lut_mask = 16'hACFF;
defparam \twiddle_data_real~112 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~96 (
	.dataa(\Add2~28_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~96_combout ),
	.cout());
defparam \twiddle_data_real~96 .lut_mask = 16'hEBBE;
defparam \twiddle_data_real~96 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~97 (
	.dataa(\Add2~28_combout ),
	.datab(\quad_del_1[1]~q ),
	.datac(\quad_del_1[2]~q ),
	.datad(\quad_del_1[0]~q ),
	.cin(gnd),
	.combout(\twiddle_data_real~97_combout ),
	.cout());
defparam \twiddle_data_real~97 .lut_mask = 16'hBEFF;
defparam \twiddle_data_real~97 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data_real~113 (
	.dataa(\twiddle_data_real~96_combout ),
	.datab(\twiddle_data_real~97_combout ),
	.datac(\gen_se:gen_new:twrom|gen_auto:sin_1n|altsyncram_component|auto_generated|q_b[14] ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data_real~113_combout ),
	.cout());
defparam \twiddle_data_real~113 .lut_mask = 16'hACFF;
defparam \twiddle_data_real~113 .sum_lutc_input = "datac";

endmodule

module fft256_asj_fft_1dp_ram_fft_121 (
	q_b_0,
	q_b_16,
	q_b_1,
	q_b_17,
	q_b_2,
	q_b_18,
	q_b_3,
	q_b_19,
	q_b_4,
	q_b_20,
	q_b_5,
	q_b_21,
	q_b_6,
	q_b_22,
	q_b_7,
	q_b_23,
	q_b_8,
	q_b_24,
	q_b_9,
	q_b_25,
	q_b_10,
	q_b_26,
	q_b_11,
	q_b_27,
	q_b_12,
	q_b_28,
	q_b_13,
	q_b_29,
	q_b_14,
	q_b_30,
	q_b_15,
	q_b_31,
	global_clock_enable,
	wren_a,
	a_ram_data_in_bus_0,
	wraddress_a_bus_0,
	wraddress_a_bus_1,
	wraddress_a_bus_2,
	wraddress_a_bus_3,
	wraddress_a_bus_4,
	wraddress_a_bus_5,
	wraddress_a_bus_6,
	wraddress_a_bus_7,
	rdaddress_a_bus_0,
	rdaddress_a_bus_1,
	rdaddress_a_bus_2,
	rdaddress_a_bus_3,
	rdaddress_a_bus_4,
	rdaddress_a_bus_5,
	rdaddress_a_bus_6,
	rdaddress_a_bus_7,
	a_ram_data_in_bus_16,
	a_ram_data_in_bus_1,
	a_ram_data_in_bus_17,
	a_ram_data_in_bus_2,
	a_ram_data_in_bus_18,
	a_ram_data_in_bus_3,
	a_ram_data_in_bus_19,
	a_ram_data_in_bus_4,
	a_ram_data_in_bus_20,
	a_ram_data_in_bus_5,
	a_ram_data_in_bus_21,
	a_ram_data_in_bus_6,
	a_ram_data_in_bus_22,
	a_ram_data_in_bus_7,
	a_ram_data_in_bus_23,
	a_ram_data_in_bus_8,
	a_ram_data_in_bus_24,
	a_ram_data_in_bus_9,
	a_ram_data_in_bus_25,
	a_ram_data_in_bus_10,
	a_ram_data_in_bus_26,
	a_ram_data_in_bus_11,
	a_ram_data_in_bus_27,
	a_ram_data_in_bus_12,
	a_ram_data_in_bus_28,
	a_ram_data_in_bus_13,
	a_ram_data_in_bus_29,
	a_ram_data_in_bus_14,
	a_ram_data_in_bus_30,
	a_ram_data_in_bus_15,
	a_ram_data_in_bus_31,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_16;
output 	q_b_1;
output 	q_b_17;
output 	q_b_2;
output 	q_b_18;
output 	q_b_3;
output 	q_b_19;
output 	q_b_4;
output 	q_b_20;
output 	q_b_5;
output 	q_b_21;
output 	q_b_6;
output 	q_b_22;
output 	q_b_7;
output 	q_b_23;
output 	q_b_8;
output 	q_b_24;
output 	q_b_9;
output 	q_b_25;
output 	q_b_10;
output 	q_b_26;
output 	q_b_11;
output 	q_b_27;
output 	q_b_12;
output 	q_b_28;
output 	q_b_13;
output 	q_b_29;
output 	q_b_14;
output 	q_b_30;
output 	q_b_15;
output 	q_b_31;
input 	global_clock_enable;
input 	wren_a;
input 	a_ram_data_in_bus_0;
input 	wraddress_a_bus_0;
input 	wraddress_a_bus_1;
input 	wraddress_a_bus_2;
input 	wraddress_a_bus_3;
input 	wraddress_a_bus_4;
input 	wraddress_a_bus_5;
input 	wraddress_a_bus_6;
input 	wraddress_a_bus_7;
input 	rdaddress_a_bus_0;
input 	rdaddress_a_bus_1;
input 	rdaddress_a_bus_2;
input 	rdaddress_a_bus_3;
input 	rdaddress_a_bus_4;
input 	rdaddress_a_bus_5;
input 	rdaddress_a_bus_6;
input 	rdaddress_a_bus_7;
input 	a_ram_data_in_bus_16;
input 	a_ram_data_in_bus_1;
input 	a_ram_data_in_bus_17;
input 	a_ram_data_in_bus_2;
input 	a_ram_data_in_bus_18;
input 	a_ram_data_in_bus_3;
input 	a_ram_data_in_bus_19;
input 	a_ram_data_in_bus_4;
input 	a_ram_data_in_bus_20;
input 	a_ram_data_in_bus_5;
input 	a_ram_data_in_bus_21;
input 	a_ram_data_in_bus_6;
input 	a_ram_data_in_bus_22;
input 	a_ram_data_in_bus_7;
input 	a_ram_data_in_bus_23;
input 	a_ram_data_in_bus_8;
input 	a_ram_data_in_bus_24;
input 	a_ram_data_in_bus_9;
input 	a_ram_data_in_bus_25;
input 	a_ram_data_in_bus_10;
input 	a_ram_data_in_bus_26;
input 	a_ram_data_in_bus_11;
input 	a_ram_data_in_bus_27;
input 	a_ram_data_in_bus_12;
input 	a_ram_data_in_bus_28;
input 	a_ram_data_in_bus_13;
input 	a_ram_data_in_bus_29;
input 	a_ram_data_in_bus_14;
input 	a_ram_data_in_bus_30;
input 	a_ram_data_in_bus_15;
input 	a_ram_data_in_bus_31;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_asj_fft_data_ram_fft_121 dat_A(
	.q_b_0(q_b_0),
	.q_b_16(q_b_16),
	.q_b_1(q_b_1),
	.q_b_17(q_b_17),
	.q_b_2(q_b_2),
	.q_b_18(q_b_18),
	.q_b_3(q_b_3),
	.q_b_19(q_b_19),
	.q_b_4(q_b_4),
	.q_b_20(q_b_20),
	.q_b_5(q_b_5),
	.q_b_21(q_b_21),
	.q_b_6(q_b_6),
	.q_b_22(q_b_22),
	.q_b_7(q_b_7),
	.q_b_23(q_b_23),
	.q_b_8(q_b_8),
	.q_b_24(q_b_24),
	.q_b_9(q_b_9),
	.q_b_25(q_b_25),
	.q_b_10(q_b_10),
	.q_b_26(q_b_26),
	.q_b_11(q_b_11),
	.q_b_27(q_b_27),
	.q_b_12(q_b_12),
	.q_b_28(q_b_28),
	.q_b_13(q_b_13),
	.q_b_29(q_b_29),
	.q_b_14(q_b_14),
	.q_b_30(q_b_30),
	.q_b_15(q_b_15),
	.q_b_31(q_b_31),
	.global_clock_enable(global_clock_enable),
	.wren_a(wren_a),
	.a_ram_data_in_bus_0(a_ram_data_in_bus_0),
	.wraddress_a_bus_0(wraddress_a_bus_0),
	.wraddress_a_bus_1(wraddress_a_bus_1),
	.wraddress_a_bus_2(wraddress_a_bus_2),
	.wraddress_a_bus_3(wraddress_a_bus_3),
	.wraddress_a_bus_4(wraddress_a_bus_4),
	.wraddress_a_bus_5(wraddress_a_bus_5),
	.wraddress_a_bus_6(wraddress_a_bus_6),
	.wraddress_a_bus_7(wraddress_a_bus_7),
	.rdaddress_a_bus_0(rdaddress_a_bus_0),
	.rdaddress_a_bus_1(rdaddress_a_bus_1),
	.rdaddress_a_bus_2(rdaddress_a_bus_2),
	.rdaddress_a_bus_3(rdaddress_a_bus_3),
	.rdaddress_a_bus_4(rdaddress_a_bus_4),
	.rdaddress_a_bus_5(rdaddress_a_bus_5),
	.rdaddress_a_bus_6(rdaddress_a_bus_6),
	.rdaddress_a_bus_7(rdaddress_a_bus_7),
	.a_ram_data_in_bus_16(a_ram_data_in_bus_16),
	.a_ram_data_in_bus_1(a_ram_data_in_bus_1),
	.a_ram_data_in_bus_17(a_ram_data_in_bus_17),
	.a_ram_data_in_bus_2(a_ram_data_in_bus_2),
	.a_ram_data_in_bus_18(a_ram_data_in_bus_18),
	.a_ram_data_in_bus_3(a_ram_data_in_bus_3),
	.a_ram_data_in_bus_19(a_ram_data_in_bus_19),
	.a_ram_data_in_bus_4(a_ram_data_in_bus_4),
	.a_ram_data_in_bus_20(a_ram_data_in_bus_20),
	.a_ram_data_in_bus_5(a_ram_data_in_bus_5),
	.a_ram_data_in_bus_21(a_ram_data_in_bus_21),
	.a_ram_data_in_bus_6(a_ram_data_in_bus_6),
	.a_ram_data_in_bus_22(a_ram_data_in_bus_22),
	.a_ram_data_in_bus_7(a_ram_data_in_bus_7),
	.a_ram_data_in_bus_23(a_ram_data_in_bus_23),
	.a_ram_data_in_bus_8(a_ram_data_in_bus_8),
	.a_ram_data_in_bus_24(a_ram_data_in_bus_24),
	.a_ram_data_in_bus_9(a_ram_data_in_bus_9),
	.a_ram_data_in_bus_25(a_ram_data_in_bus_25),
	.a_ram_data_in_bus_10(a_ram_data_in_bus_10),
	.a_ram_data_in_bus_26(a_ram_data_in_bus_26),
	.a_ram_data_in_bus_11(a_ram_data_in_bus_11),
	.a_ram_data_in_bus_27(a_ram_data_in_bus_27),
	.a_ram_data_in_bus_12(a_ram_data_in_bus_12),
	.a_ram_data_in_bus_28(a_ram_data_in_bus_28),
	.a_ram_data_in_bus_13(a_ram_data_in_bus_13),
	.a_ram_data_in_bus_29(a_ram_data_in_bus_29),
	.a_ram_data_in_bus_14(a_ram_data_in_bus_14),
	.a_ram_data_in_bus_30(a_ram_data_in_bus_30),
	.a_ram_data_in_bus_15(a_ram_data_in_bus_15),
	.a_ram_data_in_bus_31(a_ram_data_in_bus_31),
	.clk(clk));

endmodule

module fft256_asj_fft_data_ram_fft_121 (
	q_b_0,
	q_b_16,
	q_b_1,
	q_b_17,
	q_b_2,
	q_b_18,
	q_b_3,
	q_b_19,
	q_b_4,
	q_b_20,
	q_b_5,
	q_b_21,
	q_b_6,
	q_b_22,
	q_b_7,
	q_b_23,
	q_b_8,
	q_b_24,
	q_b_9,
	q_b_25,
	q_b_10,
	q_b_26,
	q_b_11,
	q_b_27,
	q_b_12,
	q_b_28,
	q_b_13,
	q_b_29,
	q_b_14,
	q_b_30,
	q_b_15,
	q_b_31,
	global_clock_enable,
	wren_a,
	a_ram_data_in_bus_0,
	wraddress_a_bus_0,
	wraddress_a_bus_1,
	wraddress_a_bus_2,
	wraddress_a_bus_3,
	wraddress_a_bus_4,
	wraddress_a_bus_5,
	wraddress_a_bus_6,
	wraddress_a_bus_7,
	rdaddress_a_bus_0,
	rdaddress_a_bus_1,
	rdaddress_a_bus_2,
	rdaddress_a_bus_3,
	rdaddress_a_bus_4,
	rdaddress_a_bus_5,
	rdaddress_a_bus_6,
	rdaddress_a_bus_7,
	a_ram_data_in_bus_16,
	a_ram_data_in_bus_1,
	a_ram_data_in_bus_17,
	a_ram_data_in_bus_2,
	a_ram_data_in_bus_18,
	a_ram_data_in_bus_3,
	a_ram_data_in_bus_19,
	a_ram_data_in_bus_4,
	a_ram_data_in_bus_20,
	a_ram_data_in_bus_5,
	a_ram_data_in_bus_21,
	a_ram_data_in_bus_6,
	a_ram_data_in_bus_22,
	a_ram_data_in_bus_7,
	a_ram_data_in_bus_23,
	a_ram_data_in_bus_8,
	a_ram_data_in_bus_24,
	a_ram_data_in_bus_9,
	a_ram_data_in_bus_25,
	a_ram_data_in_bus_10,
	a_ram_data_in_bus_26,
	a_ram_data_in_bus_11,
	a_ram_data_in_bus_27,
	a_ram_data_in_bus_12,
	a_ram_data_in_bus_28,
	a_ram_data_in_bus_13,
	a_ram_data_in_bus_29,
	a_ram_data_in_bus_14,
	a_ram_data_in_bus_30,
	a_ram_data_in_bus_15,
	a_ram_data_in_bus_31,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_16;
output 	q_b_1;
output 	q_b_17;
output 	q_b_2;
output 	q_b_18;
output 	q_b_3;
output 	q_b_19;
output 	q_b_4;
output 	q_b_20;
output 	q_b_5;
output 	q_b_21;
output 	q_b_6;
output 	q_b_22;
output 	q_b_7;
output 	q_b_23;
output 	q_b_8;
output 	q_b_24;
output 	q_b_9;
output 	q_b_25;
output 	q_b_10;
output 	q_b_26;
output 	q_b_11;
output 	q_b_27;
output 	q_b_12;
output 	q_b_28;
output 	q_b_13;
output 	q_b_29;
output 	q_b_14;
output 	q_b_30;
output 	q_b_15;
output 	q_b_31;
input 	global_clock_enable;
input 	wren_a;
input 	a_ram_data_in_bus_0;
input 	wraddress_a_bus_0;
input 	wraddress_a_bus_1;
input 	wraddress_a_bus_2;
input 	wraddress_a_bus_3;
input 	wraddress_a_bus_4;
input 	wraddress_a_bus_5;
input 	wraddress_a_bus_6;
input 	wraddress_a_bus_7;
input 	rdaddress_a_bus_0;
input 	rdaddress_a_bus_1;
input 	rdaddress_a_bus_2;
input 	rdaddress_a_bus_3;
input 	rdaddress_a_bus_4;
input 	rdaddress_a_bus_5;
input 	rdaddress_a_bus_6;
input 	rdaddress_a_bus_7;
input 	a_ram_data_in_bus_16;
input 	a_ram_data_in_bus_1;
input 	a_ram_data_in_bus_17;
input 	a_ram_data_in_bus_2;
input 	a_ram_data_in_bus_18;
input 	a_ram_data_in_bus_3;
input 	a_ram_data_in_bus_19;
input 	a_ram_data_in_bus_4;
input 	a_ram_data_in_bus_20;
input 	a_ram_data_in_bus_5;
input 	a_ram_data_in_bus_21;
input 	a_ram_data_in_bus_6;
input 	a_ram_data_in_bus_22;
input 	a_ram_data_in_bus_7;
input 	a_ram_data_in_bus_23;
input 	a_ram_data_in_bus_8;
input 	a_ram_data_in_bus_24;
input 	a_ram_data_in_bus_9;
input 	a_ram_data_in_bus_25;
input 	a_ram_data_in_bus_10;
input 	a_ram_data_in_bus_26;
input 	a_ram_data_in_bus_11;
input 	a_ram_data_in_bus_27;
input 	a_ram_data_in_bus_12;
input 	a_ram_data_in_bus_28;
input 	a_ram_data_in_bus_13;
input 	a_ram_data_in_bus_29;
input 	a_ram_data_in_bus_14;
input 	a_ram_data_in_bus_30;
input 	a_ram_data_in_bus_15;
input 	a_ram_data_in_bus_31;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_altsyncram_1 \gen_M4K:altsyncram_component (
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.clocken0(global_clock_enable),
	.wren_a(wren_a),
	.data_a({a_ram_data_in_bus_31,a_ram_data_in_bus_30,a_ram_data_in_bus_29,a_ram_data_in_bus_28,a_ram_data_in_bus_27,a_ram_data_in_bus_26,a_ram_data_in_bus_25,a_ram_data_in_bus_24,a_ram_data_in_bus_23,a_ram_data_in_bus_22,a_ram_data_in_bus_21,a_ram_data_in_bus_20,
a_ram_data_in_bus_19,a_ram_data_in_bus_18,a_ram_data_in_bus_17,a_ram_data_in_bus_16,a_ram_data_in_bus_15,a_ram_data_in_bus_14,a_ram_data_in_bus_13,a_ram_data_in_bus_12,a_ram_data_in_bus_11,a_ram_data_in_bus_10,a_ram_data_in_bus_9,a_ram_data_in_bus_8,
a_ram_data_in_bus_7,a_ram_data_in_bus_6,a_ram_data_in_bus_5,a_ram_data_in_bus_4,a_ram_data_in_bus_3,a_ram_data_in_bus_2,a_ram_data_in_bus_1,a_ram_data_in_bus_0}),
	.address_a({wraddress_a_bus_7,wraddress_a_bus_6,wraddress_a_bus_5,wraddress_a_bus_4,wraddress_a_bus_3,wraddress_a_bus_2,wraddress_a_bus_1,wraddress_a_bus_0}),
	.address_b({rdaddress_a_bus_7,rdaddress_a_bus_6,rdaddress_a_bus_5,rdaddress_a_bus_4,rdaddress_a_bus_3,rdaddress_a_bus_2,rdaddress_a_bus_1,rdaddress_a_bus_0}),
	.clock0(clk));

endmodule

module fft256_altsyncram_1 (
	q_b,
	clocken0,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[7:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_altsyncram_0ou3 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.clocken0(clocken0),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module fft256_altsyncram_0ou3 (
	q_b,
	clocken0,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[7:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 8;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 255;
defparam ram_block1a0.port_b_logical_ram_depth = 256;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.clk0_output_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "old";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 8;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock0";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 255;
defparam ram_block1a16.port_b_logical_ram_depth = 256;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 8;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 255;
defparam ram_block1a1.port_b_logical_ram_depth = 256;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.clk0_output_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "old";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 8;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock0";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 255;
defparam ram_block1a17.port_b_logical_ram_depth = 256;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 8;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 255;
defparam ram_block1a2.port_b_logical_ram_depth = 256;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.clk0_output_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "old";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 8;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock0";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 255;
defparam ram_block1a18.port_b_logical_ram_depth = 256;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 8;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 255;
defparam ram_block1a3.port_b_logical_ram_depth = 256;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.clk0_output_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "old";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 8;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock0";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 255;
defparam ram_block1a19.port_b_logical_ram_depth = 256;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 8;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 255;
defparam ram_block1a4.port_b_logical_ram_depth = 256;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.clk0_output_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "old";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 8;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock0";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 255;
defparam ram_block1a20.port_b_logical_ram_depth = 256;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 8;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 255;
defparam ram_block1a5.port_b_logical_ram_depth = 256;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.clk0_output_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "old";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 8;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock0";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 255;
defparam ram_block1a21.port_b_logical_ram_depth = 256;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 8;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 255;
defparam ram_block1a6.port_b_logical_ram_depth = 256;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.clk0_output_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "old";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 8;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "clock0";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 255;
defparam ram_block1a22.port_b_logical_ram_depth = 256;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 8;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 255;
defparam ram_block1a7.port_b_logical_ram_depth = 256;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.clk0_output_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "old";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 8;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "clock0";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 255;
defparam ram_block1a23.port_b_logical_ram_depth = 256;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 8;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 255;
defparam ram_block1a8.port_b_logical_ram_depth = 256;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.clk0_output_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "old";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 8;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 255;
defparam ram_block1a24.port_a_logical_ram_depth = 256;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 8;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "clock0";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 255;
defparam ram_block1a24.port_b_logical_ram_depth = 256;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 8;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 255;
defparam ram_block1a9.port_b_logical_ram_depth = 256;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.clk0_output_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "old";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 8;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 255;
defparam ram_block1a25.port_a_logical_ram_depth = 256;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 8;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "clock0";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 255;
defparam ram_block1a25.port_b_logical_ram_depth = 256;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 8;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 255;
defparam ram_block1a10.port_b_logical_ram_depth = 256;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.clk0_output_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "old";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 8;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 255;
defparam ram_block1a26.port_a_logical_ram_depth = 256;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 8;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "clock0";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 255;
defparam ram_block1a26.port_b_logical_ram_depth = 256;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 8;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 255;
defparam ram_block1a11.port_b_logical_ram_depth = 256;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.clk0_output_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "old";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 8;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 255;
defparam ram_block1a27.port_a_logical_ram_depth = 256;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 8;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "clock0";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 255;
defparam ram_block1a27.port_b_logical_ram_depth = 256;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 8;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 255;
defparam ram_block1a12.port_b_logical_ram_depth = 256;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.clk0_output_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "old";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 8;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 255;
defparam ram_block1a28.port_a_logical_ram_depth = 256;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 8;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "clock0";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 255;
defparam ram_block1a28.port_b_logical_ram_depth = 256;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 8;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 255;
defparam ram_block1a13.port_b_logical_ram_depth = 256;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.clk0_output_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "old";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 8;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 255;
defparam ram_block1a29.port_a_logical_ram_depth = 256;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 8;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "clock0";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 255;
defparam ram_block1a29.port_b_logical_ram_depth = 256;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 8;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 255;
defparam ram_block1a14.port_b_logical_ram_depth = 256;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.clk0_output_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "old";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 8;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 255;
defparam ram_block1a30.port_a_logical_ram_depth = 256;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 8;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "clock0";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 255;
defparam ram_block1a30.port_b_logical_ram_depth = 256;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 8;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 255;
defparam ram_block1a15.port_b_logical_ram_depth = 256;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.clk0_output_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1dp_ram_fft_121:\\gen_1_ram:gen_M4K:dat_A|asj_fft_data_ram_fft_121:dat_A|altsyncram:\\gen_M4K:altsyncram_component|altsyncram_0ou3:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "old";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 8;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 255;
defparam ram_block1a31.port_a_logical_ram_depth = 256;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 8;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "clock0";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 255;
defparam ram_block1a31.port_b_logical_ram_depth = 256;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";

endmodule

module fft256_asj_fft_1tdp_rom_fft_121 (
	q_a_0,
	q_b_0,
	q_a_1,
	q_b_1,
	q_a_2,
	q_b_2,
	q_a_3,
	q_b_3,
	q_a_4,
	q_b_4,
	q_a_5,
	q_b_5,
	q_a_6,
	q_b_6,
	q_a_7,
	q_b_7,
	q_a_8,
	q_b_8,
	q_a_9,
	q_b_9,
	q_a_10,
	q_b_10,
	q_a_11,
	q_b_11,
	q_a_12,
	q_b_12,
	q_a_13,
	q_b_13,
	q_a_14,
	q_b_14,
	q_a_15,
	q_b_15,
	twad_tempo_0,
	twad_tempe_1,
	twad_tempe_2,
	twad_tempe_3,
	twad_tempe_4,
	twad_tempe_5,
	twad_tempo_1,
	twad_tempo_2,
	twad_tempo_3,
	twad_tempo_4,
	twad_tempo_5,
	global_clock_enable,
	GND_port,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_b_0;
output 	q_a_1;
output 	q_b_1;
output 	q_a_2;
output 	q_b_2;
output 	q_a_3;
output 	q_b_3;
output 	q_a_4;
output 	q_b_4;
output 	q_a_5;
output 	q_b_5;
output 	q_a_6;
output 	q_b_6;
output 	q_a_7;
output 	q_b_7;
output 	q_a_8;
output 	q_b_8;
output 	q_a_9;
output 	q_b_9;
output 	q_a_10;
output 	q_b_10;
output 	q_a_11;
output 	q_b_11;
output 	q_a_12;
output 	q_b_12;
output 	q_a_13;
output 	q_b_13;
output 	q_a_14;
output 	q_b_14;
output 	q_a_15;
output 	q_b_15;
input 	twad_tempo_0;
input 	twad_tempe_1;
input 	twad_tempe_2;
input 	twad_tempe_3;
input 	twad_tempe_4;
input 	twad_tempe_5;
input 	twad_tempo_1;
input 	twad_tempo_2;
input 	twad_tempo_3;
input 	twad_tempo_4;
input 	twad_tempo_5;
input 	global_clock_enable;
input 	GND_port;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_asj_fft_twid_rom_tdp_fft_121 \gen_auto:sin_1n (
	.q_a({q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({twad_tempe_5,twad_tempe_4,twad_tempe_3,twad_tempe_2,twad_tempe_1,twad_tempo_0}),
	.address_b({twad_tempo_5,twad_tempo_4,twad_tempo_3,twad_tempo_2,twad_tempo_1,gnd}),
	.global_clock_enable(global_clock_enable),
	.GND_port(GND_port),
	.clock(clk));

endmodule

module fft256_asj_fft_twid_rom_tdp_fft_121 (
	q_a,
	q_b,
	address_a,
	address_b,
	global_clock_enable,
	GND_port,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_a;
output 	[15:0] q_b;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	global_clock_enable;
input 	GND_port;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_altsyncram_2 altsyncram_component(
	.q_a({q_a_unconnected_wire_31,q_a_unconnected_wire_30,q_a_unconnected_wire_29,q_a_unconnected_wire_28,q_a_unconnected_wire_27,q_a_unconnected_wire_26,q_a_unconnected_wire_25,q_a_unconnected_wire_24,q_a_unconnected_wire_23,q_a_unconnected_wire_22,q_a_unconnected_wire_21,
q_a_unconnected_wire_20,q_a_unconnected_wire_19,q_a_unconnected_wire_18,q_a_unconnected_wire_17,q_a_unconnected_wire_16,q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.q_b({q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,q_b_unconnected_wire_22,q_b_unconnected_wire_21,
q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],gnd}),
	.clocken0(global_clock_enable),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,GND_port,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.clock0(clock));

endmodule

module fft256_altsyncram_2 (
	q_a,
	q_b,
	address_a,
	address_b,
	clocken0,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
output 	[31:0] q_b;
input 	[7:0] address_a;
input 	[7:0] address_b;
input 	clocken0;
input 	[31:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_altsyncram_he72 auto_generated(
	.q_a({q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_a[0]}),
	.clocken0(clocken0),
	.data_a({data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15]}),
	.data_b({data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15],data_a[15]}),
	.clock0(clock0));

endmodule

module fft256_altsyncram_he72 (
	q_a,
	q_b,
	address_a,
	address_b,
	clocken0,
	data_a,
	data_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_a;
output 	[15:0] q_b;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clocken0;
input 	[15:0] data_a;
input 	[15:0] data_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "fft256_1n256sin.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1tdp_rom_fft_121:\\gen_se:gen_new:twrom|asj_fft_twid_rom_tdp_fft_121:\\gen_auto:sin_1n|altsyncram:altsyncram_component|altsyncram_he72:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "bidir_dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_in_clock = "clock0";
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.port_b_write_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = 64'h9BCB475E7C23CB20;

cycloneive_ram_block ram_block1a1(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "fft256_1n256sin.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1tdp_rom_fft_121:\\gen_se:gen_new:twrom|asj_fft_twid_rom_tdp_fft_121:\\gen_auto:sin_1n|altsyncram:altsyncram_component|altsyncram_he72:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "bidir_dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_in_clock = "clock0";
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.port_b_write_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = 64'h20821ACFBCF76EA8;

cycloneive_ram_block ram_block1a2(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "fft256_1n256sin.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1tdp_rom_fft_121:\\gen_se:gen_new:twrom|asj_fft_twid_rom_tdp_fft_121:\\gen_auto:sin_1n|altsyncram:altsyncram_component|altsyncram_he72:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "bidir_dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_in_clock = "clock0";
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.port_b_write_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = 64'hA634E9C44F7A6012;

cycloneive_ram_block ram_block1a3(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "fft256_1n256sin.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1tdp_rom_fft_121:\\gen_se:gen_new:twrom|asj_fft_twid_rom_tdp_fft_121:\\gen_auto:sin_1n|altsyncram:altsyncram_component|altsyncram_he72:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "bidir_dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_in_clock = "clock0";
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.port_b_write_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = 64'h4F7A0D682DCF577C;

cycloneive_ram_block ram_block1a4(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "fft256_1n256sin.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1tdp_rom_fft_121:\\gen_se:gen_new:twrom|asj_fft_twid_rom_tdp_fft_121:\\gen_auto:sin_1n|altsyncram:altsyncram_component|altsyncram_he72:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "bidir_dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_in_clock = "clock0";
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.port_b_write_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = 64'hC63068167FB7C500;

cycloneive_ram_block ram_block1a5(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "fft256_1n256sin.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1tdp_rom_fft_121:\\gen_se:gen_new:twrom|asj_fft_twid_rom_tdp_fft_121:\\gen_auto:sin_1n|altsyncram:altsyncram_component|altsyncram_he72:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "bidir_dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_in_clock = "clock0";
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.port_b_write_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = 64'hB0D253BA5E8539AA;

cycloneive_ram_block ram_block1a6(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "fft256_1n256sin.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1tdp_rom_fft_121:\\gen_se:gen_new:twrom|asj_fft_twid_rom_tdp_fft_121:\\gen_auto:sin_1n|altsyncram:altsyncram_component|altsyncram_he72:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "bidir_dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_in_clock = "clock0";
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.port_b_write_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = 64'hD0B33D7CC0D301CC;

cycloneive_ram_block ram_block1a7(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "fft256_1n256sin.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1tdp_rom_fft_121:\\gen_se:gen_new:twrom|asj_fft_twid_rom_tdp_fft_121:\\gen_auto:sin_1n|altsyncram:altsyncram_component|altsyncram_he72:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "bidir_dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_in_clock = "clock0";
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.port_b_write_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = 64'hE58C54FF6A4F01F0;

cycloneive_ram_block ram_block1a8(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "fft256_1n256sin.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1tdp_rom_fft_121:\\gen_se:gen_new:twrom|asj_fft_twid_rom_tdp_fft_121:\\gen_auto:sin_1n|altsyncram:altsyncram_component|altsyncram_he72:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "bidir_dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 6;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "clock0";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 63;
defparam ram_block1a8.port_a_logical_ram_depth = 64;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 6;
defparam ram_block1a8.port_b_data_in_clock = "clock0";
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 63;
defparam ram_block1a8.port_b_logical_ram_depth = 64;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.port_b_write_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = 64'hF92ACC00736A54AA;

cycloneive_ram_block ram_block1a9(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "fft256_1n256sin.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1tdp_rom_fft_121:\\gen_se:gen_new:twrom|asj_fft_twid_rom_tdp_fft_121:\\gen_auto:sin_1n|altsyncram:altsyncram_component|altsyncram_he72:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "bidir_dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 6;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "clock0";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 63;
defparam ram_block1a9.port_a_logical_ram_depth = 64;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 6;
defparam ram_block1a9.port_b_data_in_clock = "clock0";
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 63;
defparam ram_block1a9.port_b_logical_ram_depth = 64;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.port_b_write_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = 64'hFE3369552926CC66;

cycloneive_ram_block ram_block1a10(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "fft256_1n256sin.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1tdp_rom_fft_121:\\gen_se:gen_new:twrom|asj_fft_twid_rom_tdp_fft_121:\\gen_auto:sin_1n|altsyncram:altsyncram_component|altsyncram_he72:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "bidir_dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 6;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "clock0";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 63;
defparam ram_block1a10.port_a_logical_ram_depth = 64;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 6;
defparam ram_block1a10.port_b_data_in_clock = "clock0";
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 63;
defparam ram_block1a10.port_b_logical_ram_depth = 64;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.port_b_write_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = 64'hFFC38E664DB496B4;

cycloneive_ram_block ram_block1a11(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "fft256_1n256sin.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1tdp_rom_fft_121:\\gen_se:gen_new:twrom|asj_fft_twid_rom_tdp_fft_121:\\gen_auto:sin_1n|altsyncram:altsyncram_component|altsyncram_he72:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "bidir_dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 6;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "clock0";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 63;
defparam ram_block1a11.port_a_logical_ram_depth = 64;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 6;
defparam ram_block1a11.port_b_data_in_clock = "clock0";
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 63;
defparam ram_block1a11.port_b_logical_ram_depth = 64;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.port_b_write_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = 64'hFFFC0F878E38E738;

cycloneive_ram_block ram_block1a12(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "fft256_1n256sin.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1tdp_rom_fft_121:\\gen_se:gen_new:twrom|asj_fft_twid_rom_tdp_fft_121:\\gen_auto:sin_1n|altsyncram:altsyncram_component|altsyncram_he72:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "bidir_dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 6;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "clock0";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 63;
defparam ram_block1a12.port_a_logical_ram_depth = 64;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 6;
defparam ram_block1a12.port_b_data_in_clock = "clock0";
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 63;
defparam ram_block1a12.port_b_logical_ram_depth = 64;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.port_b_write_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = 64'hFFFFF007F03F07C0;

cycloneive_ram_block ram_block1a13(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "fft256_1n256sin.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1tdp_rom_fft_121:\\gen_se:gen_new:twrom|asj_fft_twid_rom_tdp_fft_121:\\gen_auto:sin_1n|altsyncram:altsyncram_component|altsyncram_he72:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "bidir_dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 6;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "clock0";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 63;
defparam ram_block1a13.port_a_logical_ram_depth = 64;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 6;
defparam ram_block1a13.port_b_data_in_clock = "clock0";
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 63;
defparam ram_block1a13.port_b_logical_ram_depth = 64;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.port_b_write_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = 64'hFFFFFFF8003FF800;

cycloneive_ram_block ram_block1a14(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "fft256_1n256sin.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1tdp_rom_fft_121:\\gen_se:gen_new:twrom|asj_fft_twid_rom_tdp_fft_121:\\gen_auto:sin_1n|altsyncram:altsyncram_component|altsyncram_he72:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "bidir_dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 6;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "clock0";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 63;
defparam ram_block1a14.port_a_logical_ram_depth = 64;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 6;
defparam ram_block1a14.port_b_data_in_clock = "clock0";
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 63;
defparam ram_block1a14.port_b_logical_ram_depth = 64;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.port_b_write_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init0 = 64'hFFFFFFFFFFC00000;

cycloneive_ram_block ram_block1a15(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "fft256_1n256sin.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|asj_fft_1tdp_rom_fft_121:\\gen_se:gen_new:twrom|asj_fft_twid_rom_tdp_fft_121:\\gen_auto:sin_1n|altsyncram:altsyncram_component|altsyncram_he72:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "bidir_dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 6;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "clock0";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 63;
defparam ram_block1a15.port_a_logical_ram_depth = 64;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 6;
defparam ram_block1a15.port_b_data_in_clock = "clock0";
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 63;
defparam ram_block1a15.port_b_logical_ram_depth = 64;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.port_b_write_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init0 = 64'h0000000000000000;

endmodule

module fft256_asj_fft_bfp_ctrl_fft_121 (
	rdy_for_next_block,
	global_clock_enable,
	blk_exp_0,
	blk_exp_1,
	blk_exp_2,
	blk_exp_3,
	blk_exp_4,
	blk_exp_5,
	sop_d,
	slb_i_0,
	Mux2,
	lut_out_0,
	tdl_arr_0,
	Mux1,
	lut_out_1,
	lut_out_2,
	lut_out_21,
	tdl_arr_9,
	slb_last_1,
	slb_last_0,
	slb_last_2,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	rdy_for_next_block;
input 	global_clock_enable;
output 	blk_exp_0;
output 	blk_exp_1;
output 	blk_exp_2;
output 	blk_exp_3;
output 	blk_exp_4;
output 	blk_exp_5;
input 	sop_d;
input 	slb_i_0;
input 	Mux2;
input 	lut_out_0;
output 	tdl_arr_0;
input 	Mux1;
input 	lut_out_1;
input 	lut_out_2;
input 	lut_out_21;
input 	tdl_arr_9;
output 	slb_last_1;
output 	slb_last_0;
output 	slb_last_2;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_so_crtl:gen_se_so:delay_next_pass|tdl_arr[12]~q ;
wire \blk_exp_acc[0]~6_combout ;
wire \blk_exp_acc[0]~8_combout ;
wire \blk_exp_acc[0]~9_combout ;
wire \blk_exp_acc[0]~10_combout ;
wire \blk_exp_acc[0]~q ;
wire \blk_exp~0_combout ;
wire \blk_exp[0]~1_combout ;
wire \blk_exp_acc[0]~7 ;
wire \blk_exp_acc[1]~11_combout ;
wire \blk_exp_acc[1]~q ;
wire \blk_exp~2_combout ;
wire \blk_exp_acc[1]~12 ;
wire \blk_exp_acc[2]~13_combout ;
wire \blk_exp_acc[2]~q ;
wire \blk_exp~3_combout ;
wire \blk_exp_acc[2]~14 ;
wire \blk_exp_acc[3]~15_combout ;
wire \blk_exp_acc[3]~q ;
wire \blk_exp~4_combout ;
wire \blk_exp_acc[3]~16 ;
wire \blk_exp_acc[4]~17_combout ;
wire \blk_exp_acc[4]~q ;
wire \blk_exp~5_combout ;
wire \blk_exp_acc[4]~18 ;
wire \blk_exp_acc[5]~19_combout ;
wire \blk_exp_acc[5]~q ;
wire \blk_exp~6_combout ;
wire \slb_last~0_combout ;
wire \slb_last[0]~1_combout ;
wire \slb_last[0]~2_combout ;
wire \slb_last~3_combout ;
wire \slb_last~4_combout ;


fft256_asj_fft_tdl_bit_fft_121 \gen_so_crtl:gen_se_so:delay_next_pass_2 (
	.global_clock_enable(global_clock_enable),
	.tdl_arr_0(tdl_arr_0),
	.data_in(tdl_arr_9),
	.clk(clk));

fft256_asj_fft_tdl_bit_rst_fft_121 \gen_so_crtl:gen_se_so:delay_next_pass (
	.global_clock_enable(global_clock_enable),
	.tdl_arr_12(\gen_so_crtl:gen_se_so:delay_next_pass|tdl_arr[12]~q ),
	.tdl_arr_9(tdl_arr_9),
	.clk(clk),
	.reset_n(reset_n));

dffeas \blk_exp[0] (
	.clk(clk),
	.d(\blk_exp~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_0),
	.prn(vcc));
defparam \blk_exp[0] .is_wysiwyg = "true";
defparam \blk_exp[0] .power_up = "low";

dffeas \blk_exp[1] (
	.clk(clk),
	.d(\blk_exp~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_1),
	.prn(vcc));
defparam \blk_exp[1] .is_wysiwyg = "true";
defparam \blk_exp[1] .power_up = "low";

dffeas \blk_exp[2] (
	.clk(clk),
	.d(\blk_exp~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_2),
	.prn(vcc));
defparam \blk_exp[2] .is_wysiwyg = "true";
defparam \blk_exp[2] .power_up = "low";

dffeas \blk_exp[3] (
	.clk(clk),
	.d(\blk_exp~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_3),
	.prn(vcc));
defparam \blk_exp[3] .is_wysiwyg = "true";
defparam \blk_exp[3] .power_up = "low";

dffeas \blk_exp[4] (
	.clk(clk),
	.d(\blk_exp~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_4),
	.prn(vcc));
defparam \blk_exp[4] .is_wysiwyg = "true";
defparam \blk_exp[4] .power_up = "low";

dffeas \blk_exp[5] (
	.clk(clk),
	.d(\blk_exp~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_5),
	.prn(vcc));
defparam \blk_exp[5] .is_wysiwyg = "true";
defparam \blk_exp[5] .power_up = "low";

dffeas \slb_last[1] (
	.clk(clk),
	.d(\slb_last~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_last[0]~2_combout ),
	.q(slb_last_1),
	.prn(vcc));
defparam \slb_last[1] .is_wysiwyg = "true";
defparam \slb_last[1] .power_up = "low";

dffeas \slb_last[0] (
	.clk(clk),
	.d(\slb_last~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_last[0]~2_combout ),
	.q(slb_last_0),
	.prn(vcc));
defparam \slb_last[0] .is_wysiwyg = "true";
defparam \slb_last[0] .power_up = "low";

dffeas \slb_last[2] (
	.clk(clk),
	.d(\slb_last~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_last[0]~2_combout ),
	.q(slb_last_2),
	.prn(vcc));
defparam \slb_last[2] .is_wysiwyg = "true";
defparam \slb_last[2] .power_up = "low";

cycloneive_lcell_comb \blk_exp_acc[0]~6 (
	.dataa(lut_out_0),
	.datab(\blk_exp_acc[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\blk_exp_acc[0]~6_combout ),
	.cout(\blk_exp_acc[0]~7 ));
defparam \blk_exp_acc[0]~6 .lut_mask = 16'h66EE;
defparam \blk_exp_acc[0]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp_acc[0]~8 (
	.dataa(reset_n),
	.datab(tdl_arr_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp_acc[0]~8_combout ),
	.cout());
defparam \blk_exp_acc[0]~8 .lut_mask = 16'h7777;
defparam \blk_exp_acc[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp_acc[0]~9 (
	.dataa(\gen_so_crtl:gen_se_so:delay_next_pass|tdl_arr[12]~q ),
	.datab(tdl_arr_0),
	.datac(rdy_for_next_block),
	.datad(sop_d),
	.cin(gnd),
	.combout(\blk_exp_acc[0]~9_combout ),
	.cout());
defparam \blk_exp_acc[0]~9 .lut_mask = 16'hBFFF;
defparam \blk_exp_acc[0]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp_acc[0]~10 (
	.dataa(global_clock_enable),
	.datab(reset_n),
	.datac(\blk_exp_acc[0]~9_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp_acc[0]~10_combout ),
	.cout());
defparam \blk_exp_acc[0]~10 .lut_mask = 16'hBFBF;
defparam \blk_exp_acc[0]~10 .sum_lutc_input = "datac";

dffeas \blk_exp_acc[0] (
	.clk(clk),
	.d(\blk_exp_acc[0]~6_combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[0]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[0]~q ),
	.prn(vcc));
defparam \blk_exp_acc[0] .is_wysiwyg = "true";
defparam \blk_exp_acc[0] .power_up = "low";

cycloneive_lcell_comb \blk_exp~0 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~0_combout ),
	.cout());
defparam \blk_exp~0 .lut_mask = 16'hEEEE;
defparam \blk_exp~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp[0]~1 (
	.dataa(sop_d),
	.datab(gnd),
	.datac(reset_n),
	.datad(global_clock_enable),
	.cin(gnd),
	.combout(\blk_exp[0]~1_combout ),
	.cout());
defparam \blk_exp[0]~1 .lut_mask = 16'hFFAF;
defparam \blk_exp[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp_acc[1]~11 (
	.dataa(lut_out_1),
	.datab(\blk_exp_acc[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\blk_exp_acc[0]~7 ),
	.combout(\blk_exp_acc[1]~11_combout ),
	.cout(\blk_exp_acc[1]~12 ));
defparam \blk_exp_acc[1]~11 .lut_mask = 16'h967F;
defparam \blk_exp_acc[1]~11 .sum_lutc_input = "cin";

dffeas \blk_exp_acc[1] (
	.clk(clk),
	.d(\blk_exp_acc[1]~11_combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[0]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[1]~q ),
	.prn(vcc));
defparam \blk_exp_acc[1] .is_wysiwyg = "true";
defparam \blk_exp_acc[1] .power_up = "low";

cycloneive_lcell_comb \blk_exp~2 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~2_combout ),
	.cout());
defparam \blk_exp~2 .lut_mask = 16'hEEEE;
defparam \blk_exp~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp_acc[2]~13 (
	.dataa(lut_out_21),
	.datab(\blk_exp_acc[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\blk_exp_acc[1]~12 ),
	.combout(\blk_exp_acc[2]~13_combout ),
	.cout(\blk_exp_acc[2]~14 ));
defparam \blk_exp_acc[2]~13 .lut_mask = 16'h96EF;
defparam \blk_exp_acc[2]~13 .sum_lutc_input = "cin";

dffeas \blk_exp_acc[2] (
	.clk(clk),
	.d(\blk_exp_acc[2]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[0]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[2]~q ),
	.prn(vcc));
defparam \blk_exp_acc[2] .is_wysiwyg = "true";
defparam \blk_exp_acc[2] .power_up = "low";

cycloneive_lcell_comb \blk_exp~3 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~3_combout ),
	.cout());
defparam \blk_exp~3 .lut_mask = 16'hEEEE;
defparam \blk_exp~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp_acc[3]~15 (
	.dataa(\blk_exp_acc[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\blk_exp_acc[2]~14 ),
	.combout(\blk_exp_acc[3]~15_combout ),
	.cout(\blk_exp_acc[3]~16 ));
defparam \blk_exp_acc[3]~15 .lut_mask = 16'h5A5F;
defparam \blk_exp_acc[3]~15 .sum_lutc_input = "cin";

dffeas \blk_exp_acc[3] (
	.clk(clk),
	.d(\blk_exp_acc[3]~15_combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[0]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[3]~q ),
	.prn(vcc));
defparam \blk_exp_acc[3] .is_wysiwyg = "true";
defparam \blk_exp_acc[3] .power_up = "low";

cycloneive_lcell_comb \blk_exp~4 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~4_combout ),
	.cout());
defparam \blk_exp~4 .lut_mask = 16'hEEEE;
defparam \blk_exp~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp_acc[4]~17 (
	.dataa(\blk_exp_acc[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\blk_exp_acc[3]~16 ),
	.combout(\blk_exp_acc[4]~17_combout ),
	.cout(\blk_exp_acc[4]~18 ));
defparam \blk_exp_acc[4]~17 .lut_mask = 16'h5AAF;
defparam \blk_exp_acc[4]~17 .sum_lutc_input = "cin";

dffeas \blk_exp_acc[4] (
	.clk(clk),
	.d(\blk_exp_acc[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[0]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[4]~q ),
	.prn(vcc));
defparam \blk_exp_acc[4] .is_wysiwyg = "true";
defparam \blk_exp_acc[4] .power_up = "low";

cycloneive_lcell_comb \blk_exp~5 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~5_combout ),
	.cout());
defparam \blk_exp~5 .lut_mask = 16'hEEEE;
defparam \blk_exp~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp_acc[5]~19 (
	.dataa(\blk_exp_acc[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\blk_exp_acc[4]~18 ),
	.combout(\blk_exp_acc[5]~19_combout ),
	.cout());
defparam \blk_exp_acc[5]~19 .lut_mask = 16'h5A5A;
defparam \blk_exp_acc[5]~19 .sum_lutc_input = "cin";

dffeas \blk_exp_acc[5] (
	.clk(clk),
	.d(\blk_exp_acc[5]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[0]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[5]~q ),
	.prn(vcc));
defparam \blk_exp_acc[5] .is_wysiwyg = "true";
defparam \blk_exp_acc[5] .power_up = "low";

cycloneive_lcell_comb \blk_exp~6 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~6_combout ),
	.cout());
defparam \blk_exp~6 .lut_mask = 16'hEEEE;
defparam \blk_exp~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \slb_last~0 (
	.dataa(reset_n),
	.datab(\gen_so_crtl:gen_se_so:delay_next_pass|tdl_arr[12]~q ),
	.datac(Mux1),
	.datad(sop_d),
	.cin(gnd),
	.combout(\slb_last~0_combout ),
	.cout());
defparam \slb_last~0 .lut_mask = 16'hFEFF;
defparam \slb_last~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \slb_last[0]~1 (
	.dataa(sop_d),
	.datab(tdl_arr_0),
	.datac(rdy_for_next_block),
	.datad(\gen_so_crtl:gen_se_so:delay_next_pass|tdl_arr[12]~q ),
	.cin(gnd),
	.combout(\slb_last[0]~1_combout ),
	.cout());
defparam \slb_last[0]~1 .lut_mask = 16'hEFFF;
defparam \slb_last[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \slb_last[0]~2 (
	.dataa(global_clock_enable),
	.datab(reset_n),
	.datac(\slb_last[0]~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\slb_last[0]~2_combout ),
	.cout());
defparam \slb_last[0]~2 .lut_mask = 16'hBFBF;
defparam \slb_last[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \slb_last~3 (
	.dataa(reset_n),
	.datab(Mux2),
	.datac(\gen_so_crtl:gen_se_so:delay_next_pass|tdl_arr[12]~q ),
	.datad(sop_d),
	.cin(gnd),
	.combout(\slb_last~3_combout ),
	.cout());
defparam \slb_last~3 .lut_mask = 16'hFEFF;
defparam \slb_last~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \slb_last~4 (
	.dataa(\gen_so_crtl:gen_se_so:delay_next_pass|tdl_arr[12]~q ),
	.datab(lut_out_2),
	.datac(sop_d),
	.datad(slb_i_0),
	.cin(gnd),
	.combout(\slb_last~4_combout ),
	.cout());
defparam \slb_last~4 .lut_mask = 16'hEFFF;
defparam \slb_last~4 .sum_lutc_input = "datac";

endmodule

module fft256_asj_fft_tdl_bit_fft_121 (
	global_clock_enable,
	tdl_arr_0,
	data_in,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_0;
input 	data_in;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \tdl_arr[0] (
	.clk(clk),
	.d(data_in),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_0),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

endmodule

module fft256_asj_fft_tdl_bit_rst_fft_121 (
	global_clock_enable,
	tdl_arr_12,
	tdl_arr_9,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_12;
input 	tdl_arr_9;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr~12_combout ;
wire \tdl_arr[0]~q ;
wire \tdl_arr~11_combout ;
wire \tdl_arr[1]~q ;
wire \tdl_arr~10_combout ;
wire \tdl_arr[2]~q ;
wire \tdl_arr~9_combout ;
wire \tdl_arr[3]~q ;
wire \tdl_arr~8_combout ;
wire \tdl_arr[4]~q ;
wire \tdl_arr~7_combout ;
wire \tdl_arr[5]~q ;
wire \tdl_arr~6_combout ;
wire \tdl_arr[6]~q ;
wire \tdl_arr~5_combout ;
wire \tdl_arr[7]~q ;
wire \tdl_arr~4_combout ;
wire \tdl_arr[8]~q ;
wire \tdl_arr~3_combout ;
wire \tdl_arr[9]~q ;
wire \tdl_arr~2_combout ;
wire \tdl_arr[10]~q ;
wire \tdl_arr~1_combout ;
wire \tdl_arr[11]~q ;
wire \tdl_arr~0_combout ;


dffeas \tdl_arr[12] (
	.clk(clk),
	.d(\tdl_arr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_12),
	.prn(vcc));
defparam \tdl_arr[12] .is_wysiwyg = "true";
defparam \tdl_arr[12] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~12 (
	.dataa(reset_n),
	.datab(tdl_arr_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~12_combout ),
	.cout());
defparam \tdl_arr~12 .lut_mask = 16'hEEEE;
defparam \tdl_arr~12 .sum_lutc_input = "datac";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(\tdl_arr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~11 (
	.dataa(reset_n),
	.datab(\tdl_arr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~11_combout ),
	.cout());
defparam \tdl_arr~11 .lut_mask = 16'hEEEE;
defparam \tdl_arr~11 .sum_lutc_input = "datac";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~10 (
	.dataa(reset_n),
	.datab(\tdl_arr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~10_combout ),
	.cout());
defparam \tdl_arr~10 .lut_mask = 16'hEEEE;
defparam \tdl_arr~10 .sum_lutc_input = "datac";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~9 (
	.dataa(reset_n),
	.datab(\tdl_arr[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~9_combout ),
	.cout());
defparam \tdl_arr~9 .lut_mask = 16'hEEEE;
defparam \tdl_arr~9 .sum_lutc_input = "datac";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~8 (
	.dataa(reset_n),
	.datab(\tdl_arr[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~8_combout ),
	.cout());
defparam \tdl_arr~8 .lut_mask = 16'hEEEE;
defparam \tdl_arr~8 .sum_lutc_input = "datac";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~7 (
	.dataa(reset_n),
	.datab(\tdl_arr[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~7_combout ),
	.cout());
defparam \tdl_arr~7 .lut_mask = 16'hEEEE;
defparam \tdl_arr~7 .sum_lutc_input = "datac";

dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5]~q ),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~6 (
	.dataa(reset_n),
	.datab(\tdl_arr[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~6_combout ),
	.cout());
defparam \tdl_arr~6 .lut_mask = 16'hEEEE;
defparam \tdl_arr~6 .sum_lutc_input = "datac";

dffeas \tdl_arr[6] (
	.clk(clk),
	.d(\tdl_arr~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[6]~q ),
	.prn(vcc));
defparam \tdl_arr[6] .is_wysiwyg = "true";
defparam \tdl_arr[6] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~5 (
	.dataa(reset_n),
	.datab(\tdl_arr[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~5_combout ),
	.cout());
defparam \tdl_arr~5 .lut_mask = 16'hEEEE;
defparam \tdl_arr~5 .sum_lutc_input = "datac";

dffeas \tdl_arr[7] (
	.clk(clk),
	.d(\tdl_arr~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[7]~q ),
	.prn(vcc));
defparam \tdl_arr[7] .is_wysiwyg = "true";
defparam \tdl_arr[7] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~4 (
	.dataa(reset_n),
	.datab(\tdl_arr[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~4_combout ),
	.cout());
defparam \tdl_arr~4 .lut_mask = 16'hEEEE;
defparam \tdl_arr~4 .sum_lutc_input = "datac";

dffeas \tdl_arr[8] (
	.clk(clk),
	.d(\tdl_arr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[8]~q ),
	.prn(vcc));
defparam \tdl_arr[8] .is_wysiwyg = "true";
defparam \tdl_arr[8] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~3 (
	.dataa(reset_n),
	.datab(\tdl_arr[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~3_combout ),
	.cout());
defparam \tdl_arr~3 .lut_mask = 16'hEEEE;
defparam \tdl_arr~3 .sum_lutc_input = "datac";

dffeas \tdl_arr[9] (
	.clk(clk),
	.d(\tdl_arr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[9]~q ),
	.prn(vcc));
defparam \tdl_arr[9] .is_wysiwyg = "true";
defparam \tdl_arr[9] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~2 (
	.dataa(reset_n),
	.datab(\tdl_arr[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~2_combout ),
	.cout());
defparam \tdl_arr~2 .lut_mask = 16'hEEEE;
defparam \tdl_arr~2 .sum_lutc_input = "datac";

dffeas \tdl_arr[10] (
	.clk(clk),
	.d(\tdl_arr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[10]~q ),
	.prn(vcc));
defparam \tdl_arr[10] .is_wysiwyg = "true";
defparam \tdl_arr[10] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~1 (
	.dataa(reset_n),
	.datab(\tdl_arr[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~1_combout ),
	.cout());
defparam \tdl_arr~1 .lut_mask = 16'hEEEE;
defparam \tdl_arr~1 .sum_lutc_input = "datac";

dffeas \tdl_arr[11] (
	.clk(clk),
	.d(\tdl_arr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[11]~q ),
	.prn(vcc));
defparam \tdl_arr[11] .is_wysiwyg = "true";
defparam \tdl_arr[11] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~0 (
	.dataa(reset_n),
	.datab(\tdl_arr[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~0_combout ),
	.cout());
defparam \tdl_arr~0 .lut_mask = 16'hEEEE;
defparam \tdl_arr~0 .sum_lutc_input = "datac";

endmodule

module fft256_asj_fft_dataadgen_fft_121 (
	k_count_wr_2,
	k_count_wr_0,
	k_count_wr_6,
	k_count_wr_3,
	k_count_wr_1,
	k_count_wr_7,
	k_count_wr_4,
	k_count_wr_5,
	global_clock_enable,
	rd_addr_a_0,
	rd_addr_a_1,
	rd_addr_a_2,
	rd_addr_a_3,
	rd_addr_a_4,
	rd_addr_a_5,
	rd_addr_a_6,
	rd_addr_a_7,
	p_tdl_0_18,
	p_tdl_1_18,
	p_tdl_2_18,
	clk)/* synthesis synthesis_greybox=1 */;
input 	k_count_wr_2;
input 	k_count_wr_0;
input 	k_count_wr_6;
input 	k_count_wr_3;
input 	k_count_wr_1;
input 	k_count_wr_7;
input 	k_count_wr_4;
input 	k_count_wr_5;
input 	global_clock_enable;
output 	rd_addr_a_0;
output 	rd_addr_a_1;
output 	rd_addr_a_2;
output 	rd_addr_a_3;
output 	rd_addr_a_4;
output 	rd_addr_a_5;
output 	rd_addr_a_6;
output 	rd_addr_a_7;
input 	p_tdl_0_18;
input 	p_tdl_1_18;
input 	p_tdl_2_18;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux7~0_combout ;
wire \Mux1~0_combout ;
wire \Mux7~1_combout ;
wire \Mux6~0_combout ;
wire \Mux6~1_combout ;
wire \Mux7~2_combout ;
wire \rd_addr_a[2]~0_combout ;
wire \Mux5~0_combout ;
wire \Mux5~1_combout ;
wire \Mux6~2_combout ;
wire \Mux4~0_combout ;
wire \Mux4~1_combout ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \rd_addr_a[5]~1_combout ;
wire \Mux3~2_combout ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \Mux2~2_combout ;
wire \Mux1~1_combout ;
wire \Mux1~2_combout ;
wire \Mux0~0_combout ;


dffeas \rd_addr_a[0] (
	.clk(clk),
	.d(\Mux7~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_a_0),
	.prn(vcc));
defparam \rd_addr_a[0] .is_wysiwyg = "true";
defparam \rd_addr_a[0] .power_up = "low";

dffeas \rd_addr_a[1] (
	.clk(clk),
	.d(\Mux6~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_a_1),
	.prn(vcc));
defparam \rd_addr_a[1] .is_wysiwyg = "true";
defparam \rd_addr_a[1] .power_up = "low";

dffeas \rd_addr_a[2] (
	.clk(clk),
	.d(\Mux5~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_a_2),
	.prn(vcc));
defparam \rd_addr_a[2] .is_wysiwyg = "true";
defparam \rd_addr_a[2] .power_up = "low";

dffeas \rd_addr_a[3] (
	.clk(clk),
	.d(\Mux4~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_a_3),
	.prn(vcc));
defparam \rd_addr_a[3] .is_wysiwyg = "true";
defparam \rd_addr_a[3] .power_up = "low";

dffeas \rd_addr_a[4] (
	.clk(clk),
	.d(\Mux3~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_a_4),
	.prn(vcc));
defparam \rd_addr_a[4] .is_wysiwyg = "true";
defparam \rd_addr_a[4] .power_up = "low";

dffeas \rd_addr_a[5] (
	.clk(clk),
	.d(\Mux2~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_a_5),
	.prn(vcc));
defparam \rd_addr_a[5] .is_wysiwyg = "true";
defparam \rd_addr_a[5] .power_up = "low";

dffeas \rd_addr_a[6] (
	.clk(clk),
	.d(\Mux1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_a_6),
	.prn(vcc));
defparam \rd_addr_a[6] .is_wysiwyg = "true";
defparam \rd_addr_a[6] .power_up = "low";

dffeas \rd_addr_a[7] (
	.clk(clk),
	.d(\Mux0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_a_7),
	.prn(vcc));
defparam \rd_addr_a[7] .is_wysiwyg = "true";
defparam \rd_addr_a[7] .power_up = "low";

cycloneive_lcell_comb \Mux7~0 (
	.dataa(k_count_wr_2),
	.datab(k_count_wr_0),
	.datac(p_tdl_0_18),
	.datad(p_tdl_1_18),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'hEFFE;
defparam \Mux7~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(p_tdl_0_18),
	.datad(p_tdl_1_18),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'h0FFF;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~1 (
	.dataa(\Mux7~0_combout ),
	.datab(k_count_wr_6),
	.datac(p_tdl_2_18),
	.datad(\Mux1~0_combout ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
defparam \Mux7~1 .lut_mask = 16'hEFFE;
defparam \Mux7~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~0 (
	.dataa(k_count_wr_3),
	.datab(k_count_wr_1),
	.datac(p_tdl_0_18),
	.datad(p_tdl_1_18),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'hEFFE;
defparam \Mux6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~1 (
	.dataa(\Mux6~0_combout ),
	.datab(k_count_wr_7),
	.datac(p_tdl_2_18),
	.datad(\Mux1~0_combout ),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
defparam \Mux6~1 .lut_mask = 16'hEFFE;
defparam \Mux6~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~2 (
	.dataa(k_count_wr_2),
	.datab(k_count_wr_4),
	.datac(gnd),
	.datad(p_tdl_2_18),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
defparam \Mux7~2 .lut_mask = 16'hAACC;
defparam \Mux7~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_addr_a[2]~0 (
	.dataa(p_tdl_2_18),
	.datab(gnd),
	.datac(p_tdl_0_18),
	.datad(p_tdl_1_18),
	.cin(gnd),
	.combout(\rd_addr_a[2]~0_combout ),
	.cout());
defparam \rd_addr_a[2]~0 .lut_mask = 16'hAFFA;
defparam \rd_addr_a[2]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~0 (
	.dataa(k_count_wr_0),
	.datab(\Mux7~2_combout ),
	.datac(p_tdl_1_18),
	.datad(\rd_addr_a[2]~0_combout ),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'hACFF;
defparam \Mux5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~1 (
	.dataa(\Mux5~0_combout ),
	.datab(k_count_wr_4),
	.datac(\rd_addr_a[2]~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
defparam \Mux5~1 .lut_mask = 16'hFEFE;
defparam \Mux5~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~2 (
	.dataa(k_count_wr_3),
	.datab(k_count_wr_5),
	.datac(gnd),
	.datad(p_tdl_2_18),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
defparam \Mux6~2 .lut_mask = 16'hAACC;
defparam \Mux6~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~0 (
	.dataa(k_count_wr_1),
	.datab(\Mux6~2_combout ),
	.datac(p_tdl_1_18),
	.datad(\rd_addr_a[2]~0_combout ),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'hACFF;
defparam \Mux4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~1 (
	.dataa(\Mux4~0_combout ),
	.datab(\rd_addr_a[2]~0_combout ),
	.datac(k_count_wr_5),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
defparam \Mux4~1 .lut_mask = 16'hFEFE;
defparam \Mux4~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~0 (
	.dataa(p_tdl_0_18),
	.datab(k_count_wr_0),
	.datac(p_tdl_1_18),
	.datad(k_count_wr_4),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hFFDE;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~1 (
	.dataa(k_count_wr_6),
	.datab(p_tdl_0_18),
	.datac(\Mux3~0_combout ),
	.datad(\Mux7~2_combout ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
defparam \Mux3~1 .lut_mask = 16'hFFBE;
defparam \Mux3~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_addr_a[5]~1 (
	.dataa(p_tdl_2_18),
	.datab(gnd),
	.datac(p_tdl_0_18),
	.datad(p_tdl_1_18),
	.cin(gnd),
	.combout(\rd_addr_a[5]~1_combout ),
	.cout());
defparam \rd_addr_a[5]~1 .lut_mask = 16'hA55A;
defparam \rd_addr_a[5]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~2 (
	.dataa(k_count_wr_2),
	.datab(\Mux3~1_combout ),
	.datac(gnd),
	.datad(\rd_addr_a[5]~1_combout ),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
defparam \Mux3~2 .lut_mask = 16'hAACC;
defparam \Mux3~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~0 (
	.dataa(p_tdl_0_18),
	.datab(k_count_wr_1),
	.datac(p_tdl_1_18),
	.datad(k_count_wr_5),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFFDE;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~1 (
	.dataa(k_count_wr_7),
	.datab(p_tdl_0_18),
	.datac(\Mux2~0_combout ),
	.datad(\Mux6~2_combout ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
defparam \Mux2~1 .lut_mask = 16'hFFBE;
defparam \Mux2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~2 (
	.dataa(k_count_wr_3),
	.datab(\Mux2~1_combout ),
	.datac(gnd),
	.datad(\rd_addr_a[5]~1_combout ),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
defparam \Mux2~2 .lut_mask = 16'hAACC;
defparam \Mux2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~1 (
	.dataa(gnd),
	.datab(p_tdl_1_18),
	.datac(p_tdl_0_18),
	.datad(p_tdl_2_18),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'h3FCF;
defparam \Mux1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~2 (
	.dataa(k_count_wr_6),
	.datab(k_count_wr_0),
	.datac(gnd),
	.datad(\Mux1~1_combout ),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
defparam \Mux1~2 .lut_mask = 16'hAACC;
defparam \Mux1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(k_count_wr_7),
	.datab(k_count_wr_1),
	.datac(gnd),
	.datad(\Mux1~1_combout ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hAACC;
defparam \Mux0~0 .sum_lutc_input = "datac";

endmodule

module fft256_asj_fft_dataadgen_fft_121_1 (
	global_clock_enable,
	rd_addr_a_0,
	rd_addr_a_1,
	rd_addr_a_2,
	rd_addr_a_3,
	rd_addr_a_4,
	rd_addr_a_5,
	rd_addr_a_6,
	rd_addr_a_7,
	p_2,
	p_0,
	p_1,
	rd_addr_a_01,
	k_count_2,
	k_count_0,
	k_count_6,
	k_count_3,
	k_count_1,
	k_count_7,
	k_count_4,
	k_count_5,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	rd_addr_a_0;
output 	rd_addr_a_1;
output 	rd_addr_a_2;
output 	rd_addr_a_3;
output 	rd_addr_a_4;
output 	rd_addr_a_5;
output 	rd_addr_a_6;
output 	rd_addr_a_7;
input 	p_2;
input 	p_0;
input 	p_1;
output 	rd_addr_a_01;
input 	k_count_2;
input 	k_count_0;
input 	k_count_6;
input 	k_count_3;
input 	k_count_1;
input 	k_count_7;
input 	k_count_4;
input 	k_count_5;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \Mux6~0_combout ;
wire \Mux6~1_combout ;
wire \Mux7~2_combout ;
wire \rd_addr_a[2]~1_combout ;
wire \Mux5~0_combout ;
wire \Mux5~1_combout ;
wire \Mux6~2_combout ;
wire \Mux4~0_combout ;
wire \Mux4~1_combout ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \rd_addr_a[4]~2_combout ;
wire \Mux3~2_combout ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \Mux2~2_combout ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \Mux0~0_combout ;


dffeas \rd_addr_a[0] (
	.clk(clk),
	.d(\Mux7~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_a_0),
	.prn(vcc));
defparam \rd_addr_a[0] .is_wysiwyg = "true";
defparam \rd_addr_a[0] .power_up = "low";

dffeas \rd_addr_a[1] (
	.clk(clk),
	.d(\Mux6~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_a_1),
	.prn(vcc));
defparam \rd_addr_a[1] .is_wysiwyg = "true";
defparam \rd_addr_a[1] .power_up = "low";

dffeas \rd_addr_a[2] (
	.clk(clk),
	.d(\Mux5~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_a_2),
	.prn(vcc));
defparam \rd_addr_a[2] .is_wysiwyg = "true";
defparam \rd_addr_a[2] .power_up = "low";

dffeas \rd_addr_a[3] (
	.clk(clk),
	.d(\Mux4~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_a_3),
	.prn(vcc));
defparam \rd_addr_a[3] .is_wysiwyg = "true";
defparam \rd_addr_a[3] .power_up = "low";

dffeas \rd_addr_a[4] (
	.clk(clk),
	.d(\Mux3~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_a_4),
	.prn(vcc));
defparam \rd_addr_a[4] .is_wysiwyg = "true";
defparam \rd_addr_a[4] .power_up = "low";

dffeas \rd_addr_a[5] (
	.clk(clk),
	.d(\Mux2~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_a_5),
	.prn(vcc));
defparam \rd_addr_a[5] .is_wysiwyg = "true";
defparam \rd_addr_a[5] .power_up = "low";

dffeas \rd_addr_a[6] (
	.clk(clk),
	.d(\Mux1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_a_6),
	.prn(vcc));
defparam \rd_addr_a[6] .is_wysiwyg = "true";
defparam \rd_addr_a[6] .power_up = "low";

dffeas \rd_addr_a[7] (
	.clk(clk),
	.d(\Mux0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_a_7),
	.prn(vcc));
defparam \rd_addr_a[7] .is_wysiwyg = "true";
defparam \rd_addr_a[7] .power_up = "low";

cycloneive_lcell_comb \rd_addr_a[0]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(rd_addr_a_01),
	.cout());
defparam \rd_addr_a[0]~0 .lut_mask = 16'h0FFF;
defparam \rd_addr_a[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~0 (
	.dataa(k_count_2),
	.datab(k_count_0),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'hEFFE;
defparam \Mux7~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~1 (
	.dataa(\Mux7~0_combout ),
	.datab(k_count_6),
	.datac(p_2),
	.datad(rd_addr_a_01),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
defparam \Mux7~1 .lut_mask = 16'hEFFE;
defparam \Mux7~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~0 (
	.dataa(k_count_3),
	.datab(k_count_1),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'hEFFE;
defparam \Mux6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~1 (
	.dataa(\Mux6~0_combout ),
	.datab(k_count_7),
	.datac(p_2),
	.datad(rd_addr_a_01),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
defparam \Mux6~1 .lut_mask = 16'hEFFE;
defparam \Mux6~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~2 (
	.dataa(k_count_2),
	.datab(k_count_4),
	.datac(gnd),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
defparam \Mux7~2 .lut_mask = 16'hAACC;
defparam \Mux7~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_addr_a[2]~1 (
	.dataa(p_2),
	.datab(gnd),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\rd_addr_a[2]~1_combout ),
	.cout());
defparam \rd_addr_a[2]~1 .lut_mask = 16'hAFFA;
defparam \rd_addr_a[2]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~0 (
	.dataa(k_count_0),
	.datab(\Mux7~2_combout ),
	.datac(p_1),
	.datad(\rd_addr_a[2]~1_combout ),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'hACFF;
defparam \Mux5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~1 (
	.dataa(\Mux5~0_combout ),
	.datab(k_count_4),
	.datac(\rd_addr_a[2]~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
defparam \Mux5~1 .lut_mask = 16'hFEFE;
defparam \Mux5~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~2 (
	.dataa(k_count_3),
	.datab(k_count_5),
	.datac(gnd),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
defparam \Mux6~2 .lut_mask = 16'hAACC;
defparam \Mux6~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~0 (
	.dataa(k_count_1),
	.datab(\Mux6~2_combout ),
	.datac(p_1),
	.datad(\rd_addr_a[2]~1_combout ),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'hACFF;
defparam \Mux4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~1 (
	.dataa(\Mux4~0_combout ),
	.datab(\rd_addr_a[2]~1_combout ),
	.datac(k_count_5),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
defparam \Mux4~1 .lut_mask = 16'hFEFE;
defparam \Mux4~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~0 (
	.dataa(p_0),
	.datab(k_count_0),
	.datac(p_1),
	.datad(k_count_4),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hFFDE;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~1 (
	.dataa(k_count_6),
	.datab(p_0),
	.datac(\Mux3~0_combout ),
	.datad(\Mux7~2_combout ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
defparam \Mux3~1 .lut_mask = 16'hFFBE;
defparam \Mux3~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_addr_a[4]~2 (
	.dataa(p_2),
	.datab(gnd),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\rd_addr_a[4]~2_combout ),
	.cout());
defparam \rd_addr_a[4]~2 .lut_mask = 16'hA55A;
defparam \rd_addr_a[4]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~2 (
	.dataa(k_count_2),
	.datab(\Mux3~1_combout ),
	.datac(gnd),
	.datad(\rd_addr_a[4]~2_combout ),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
defparam \Mux3~2 .lut_mask = 16'hAACC;
defparam \Mux3~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~0 (
	.dataa(p_1),
	.datab(k_count_7),
	.datac(p_0),
	.datad(k_count_5),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFFDE;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~1 (
	.dataa(k_count_1),
	.datab(p_1),
	.datac(\Mux2~0_combout ),
	.datad(\Mux6~2_combout ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
defparam \Mux2~1 .lut_mask = 16'hFFBE;
defparam \Mux2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~2 (
	.dataa(k_count_3),
	.datab(\Mux2~1_combout ),
	.datac(gnd),
	.datad(\rd_addr_a[4]~2_combout ),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
defparam \Mux2~2 .lut_mask = 16'hAACC;
defparam \Mux2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(gnd),
	.datab(p_1),
	.datac(p_0),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'h3FCF;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~1 (
	.dataa(k_count_6),
	.datab(k_count_0),
	.datac(gnd),
	.datad(\Mux1~0_combout ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hAACC;
defparam \Mux1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(k_count_7),
	.datab(k_count_1),
	.datac(gnd),
	.datad(\Mux1~0_combout ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hAACC;
defparam \Mux0~0 .sum_lutc_input = "datac";

endmodule

module fft256_asj_fft_dft_bfp_sgl_fft_121 (
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_31,
	twiddle_data_real_0,
	twiddle_data_real_15,
	twiddle_data_imag_1,
	twiddle_data_imag_2,
	twiddle_data_imag_3,
	twiddle_data_imag_4,
	twiddle_data_imag_5,
	twiddle_data_imag_6,
	twiddle_data_imag_7,
	twiddle_data_imag_8,
	twiddle_data_imag_9,
	twiddle_data_imag_10,
	twiddle_data_imag_11,
	twiddle_data_imag_12,
	twiddle_data_imag_13,
	twiddle_data_imag_14,
	twiddle_data_imag_15,
	source_valid_ctrl_sop,
	stall_reg,
	source_stall_int_d,
	global_clock_enable,
	slb_i_0,
	Mux2,
	lut_out_0,
	tdl_arr_0,
	Mux1,
	lut_out_1,
	lut_out_2,
	lut_out_21,
	real_out_0,
	real_out_1,
	real_out_2,
	real_out_3,
	real_out_4,
	real_out_5,
	real_out_6,
	real_out_7,
	real_out_8,
	real_out_9,
	real_out_10,
	real_out_11,
	real_out_12,
	real_out_13,
	real_out_14,
	real_out_15,
	tdl_arr_01,
	k_count_0,
	k_count_1,
	twiddle_data_real_1,
	twiddle_data_real_2,
	twiddle_data_real_3,
	twiddle_data_real_4,
	twiddle_data_real_5,
	twiddle_data_real_6,
	twiddle_data_real_7,
	twiddle_data_real_8,
	twiddle_data_real_9,
	twiddle_data_real_10,
	twiddle_data_real_11,
	twiddle_data_real_12,
	twiddle_data_real_13,
	twiddle_data_real_14,
	twiddle_data_imag_0,
	ram_data_out_0,
	ram_data_out_2,
	slb_last_1,
	ram_data_out_1,
	slb_last_0,
	slb_last_2,
	ram_data_out_14,
	ram_data_out_12,
	ram_data_out_13,
	ram_data_out_15,
	ram_data_out_11,
	ram_data_out_10,
	ram_data_out_9,
	ram_data_out_8,
	ram_data_out_7,
	ram_data_out_6,
	ram_data_out_5,
	ram_data_out_4,
	ram_data_out_3,
	ram_data_out_16,
	ram_data_out_18,
	ram_data_out_17,
	ram_data_out_28,
	ram_data_out_29,
	ram_data_out_30,
	ram_data_out_31,
	ram_data_out_27,
	ram_data_out_26,
	ram_data_out_25,
	ram_data_out_24,
	ram_data_out_23,
	ram_data_out_22,
	ram_data_out_21,
	ram_data_out_20,
	ram_data_out_19,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_31;
input 	twiddle_data_real_0;
input 	twiddle_data_real_15;
input 	twiddle_data_imag_1;
input 	twiddle_data_imag_2;
input 	twiddle_data_imag_3;
input 	twiddle_data_imag_4;
input 	twiddle_data_imag_5;
input 	twiddle_data_imag_6;
input 	twiddle_data_imag_7;
input 	twiddle_data_imag_8;
input 	twiddle_data_imag_9;
input 	twiddle_data_imag_10;
input 	twiddle_data_imag_11;
input 	twiddle_data_imag_12;
input 	twiddle_data_imag_13;
input 	twiddle_data_imag_14;
input 	twiddle_data_imag_15;
input 	source_valid_ctrl_sop;
input 	stall_reg;
input 	source_stall_int_d;
input 	global_clock_enable;
output 	slb_i_0;
output 	Mux2;
output 	lut_out_0;
input 	tdl_arr_0;
output 	Mux1;
output 	lut_out_1;
output 	lut_out_2;
output 	lut_out_21;
output 	real_out_0;
output 	real_out_1;
output 	real_out_2;
output 	real_out_3;
output 	real_out_4;
output 	real_out_5;
output 	real_out_6;
output 	real_out_7;
output 	real_out_8;
output 	real_out_9;
output 	real_out_10;
output 	real_out_11;
output 	real_out_12;
output 	real_out_13;
output 	real_out_14;
output 	real_out_15;
input 	tdl_arr_01;
input 	k_count_0;
input 	k_count_1;
input 	twiddle_data_real_1;
input 	twiddle_data_real_2;
input 	twiddle_data_real_3;
input 	twiddle_data_real_4;
input 	twiddle_data_real_5;
input 	twiddle_data_real_6;
input 	twiddle_data_real_7;
input 	twiddle_data_real_8;
input 	twiddle_data_real_9;
input 	twiddle_data_real_10;
input 	twiddle_data_real_11;
input 	twiddle_data_real_12;
input 	twiddle_data_real_13;
input 	twiddle_data_real_14;
input 	twiddle_data_imag_0;
input 	ram_data_out_0;
input 	ram_data_out_2;
input 	slb_last_1;
input 	ram_data_out_1;
input 	slb_last_0;
input 	slb_last_2;
input 	ram_data_out_14;
input 	ram_data_out_12;
input 	ram_data_out_13;
input 	ram_data_out_15;
input 	ram_data_out_11;
input 	ram_data_out_10;
input 	ram_data_out_9;
input 	ram_data_out_8;
input 	ram_data_out_7;
input 	ram_data_out_6;
input 	ram_data_out_5;
input 	ram_data_out_4;
input 	ram_data_out_3;
input 	ram_data_out_16;
input 	ram_data_out_18;
input 	ram_data_out_17;
input 	ram_data_out_28;
input 	ram_data_out_29;
input 	ram_data_out_30;
input 	ram_data_out_31;
input 	ram_data_out_27;
input 	ram_data_out_26;
input 	ram_data_out_25;
input 	ram_data_out_24;
input 	ram_data_out_23;
input 	ram_data_out_22;
input 	ram_data_out_21;
input 	ram_data_out_20;
input 	ram_data_out_19;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ;
wire \butterfly_st_imag[2]~q ;
wire \butterfly_st_imag[1]~q ;
wire \butterfly_st_imag[0]~q ;
wire \butterfly_st_imag[17]~q ;
wire \butterfly_st_imag[3]~q ;
wire \butterfly_st_imag[4]~q ;
wire \butterfly_st_imag[5]~q ;
wire \butterfly_st_imag[6]~q ;
wire \butterfly_st_imag[7]~q ;
wire \butterfly_st_imag[8]~q ;
wire \butterfly_st_imag[9]~q ;
wire \butterfly_st_imag[10]~q ;
wire \butterfly_st_imag[11]~q ;
wire \butterfly_st_imag[12]~q ;
wire \butterfly_st_imag[13]~q ;
wire \butterfly_st_imag[14]~q ;
wire \butterfly_st_imag[15]~q ;
wire \butterfly_st_imag[16]~q ;
wire \butterfly_st_real[2]~q ;
wire \butterfly_st_real[1]~q ;
wire \butterfly_st_real[0]~q ;
wire \butterfly_st_real[17]~q ;
wire \butterfly_st_real[3]~q ;
wire \butterfly_st_real[4]~q ;
wire \butterfly_st_real[5]~q ;
wire \butterfly_st_real[6]~q ;
wire \butterfly_st_real[7]~q ;
wire \butterfly_st_real[8]~q ;
wire \butterfly_st_real[9]~q ;
wire \butterfly_st_real[10]~q ;
wire \butterfly_st_real[11]~q ;
wire \butterfly_st_real[12]~q ;
wire \butterfly_st_real[13]~q ;
wire \butterfly_st_real[14]~q ;
wire \butterfly_st_real[15]~q ;
wire \butterfly_st_real[16]~q ;
wire \result_x2_x4_imag[2]~q ;
wire \result_x1_x3_imag[2]~q ;
wire \result_x2_x4_imag[1]~q ;
wire \result_x1_x3_imag[1]~q ;
wire \result_x2_x4_imag[0]~q ;
wire \result_x1_x3_imag[0]~q ;
wire \butterfly_st_imag[0]~19_cout ;
wire \butterfly_st_imag[0]~21 ;
wire \butterfly_st_imag[0]~20_combout ;
wire \butterfly_st_imag[1]~23 ;
wire \butterfly_st_imag[1]~22_combout ;
wire \butterfly_st_imag[2]~25 ;
wire \butterfly_st_imag[2]~24_combout ;
wire \result_x2_x4_imag[16]~q ;
wire \result_x1_x3_imag[16]~q ;
wire \result_x2_x4_imag[15]~q ;
wire \result_x1_x3_imag[15]~q ;
wire \result_x2_x4_imag[14]~q ;
wire \result_x1_x3_imag[14]~q ;
wire \result_x2_x4_imag[13]~q ;
wire \result_x1_x3_imag[13]~q ;
wire \result_x2_x4_imag[12]~q ;
wire \result_x1_x3_imag[12]~q ;
wire \result_x2_x4_imag[11]~q ;
wire \result_x1_x3_imag[11]~q ;
wire \result_x2_x4_imag[10]~q ;
wire \result_x1_x3_imag[10]~q ;
wire \result_x2_x4_imag[9]~q ;
wire \result_x1_x3_imag[9]~q ;
wire \result_x2_x4_imag[8]~q ;
wire \result_x1_x3_imag[8]~q ;
wire \result_x2_x4_imag[7]~q ;
wire \result_x1_x3_imag[7]~q ;
wire \result_x2_x4_imag[6]~q ;
wire \result_x1_x3_imag[6]~q ;
wire \result_x2_x4_imag[5]~q ;
wire \result_x1_x3_imag[5]~q ;
wire \result_x2_x4_imag[4]~q ;
wire \result_x1_x3_imag[4]~q ;
wire \result_x2_x4_imag[3]~q ;
wire \result_x1_x3_imag[3]~q ;
wire \butterfly_st_imag[3]~27 ;
wire \butterfly_st_imag[3]~26_combout ;
wire \butterfly_st_imag[4]~29 ;
wire \butterfly_st_imag[4]~28_combout ;
wire \butterfly_st_imag[5]~31 ;
wire \butterfly_st_imag[5]~30_combout ;
wire \butterfly_st_imag[6]~33 ;
wire \butterfly_st_imag[6]~32_combout ;
wire \butterfly_st_imag[7]~35 ;
wire \butterfly_st_imag[7]~34_combout ;
wire \butterfly_st_imag[8]~37 ;
wire \butterfly_st_imag[8]~36_combout ;
wire \butterfly_st_imag[9]~39 ;
wire \butterfly_st_imag[9]~38_combout ;
wire \butterfly_st_imag[10]~41 ;
wire \butterfly_st_imag[10]~40_combout ;
wire \butterfly_st_imag[11]~43 ;
wire \butterfly_st_imag[11]~42_combout ;
wire \butterfly_st_imag[12]~45 ;
wire \butterfly_st_imag[12]~44_combout ;
wire \butterfly_st_imag[13]~47 ;
wire \butterfly_st_imag[13]~46_combout ;
wire \butterfly_st_imag[14]~49 ;
wire \butterfly_st_imag[14]~48_combout ;
wire \butterfly_st_imag[15]~51 ;
wire \butterfly_st_imag[15]~50_combout ;
wire \butterfly_st_imag[16]~53 ;
wire \butterfly_st_imag[16]~52_combout ;
wire \butterfly_st_imag[17]~54_combout ;
wire \sr[0]~q ;
wire \result_x2_x4_real[2]~q ;
wire \result_x1_x3_real[2]~q ;
wire \result_x2_x4_real[1]~q ;
wire \result_x1_x3_real[1]~q ;
wire \result_x2_x4_real[0]~q ;
wire \result_x1_x3_real[0]~q ;
wire \butterfly_st_real[0]~19_cout ;
wire \butterfly_st_real[0]~21 ;
wire \butterfly_st_real[0]~20_combout ;
wire \butterfly_st_real[1]~23 ;
wire \butterfly_st_real[1]~22_combout ;
wire \butterfly_st_real[2]~25 ;
wire \butterfly_st_real[2]~24_combout ;
wire \result_x2_x4_real[16]~q ;
wire \result_x1_x3_real[16]~q ;
wire \result_x2_x4_real[15]~q ;
wire \result_x1_x3_real[15]~q ;
wire \result_x2_x4_real[14]~q ;
wire \result_x1_x3_real[14]~q ;
wire \result_x2_x4_real[13]~q ;
wire \result_x1_x3_real[13]~q ;
wire \result_x2_x4_real[12]~q ;
wire \result_x1_x3_real[12]~q ;
wire \result_x2_x4_real[11]~q ;
wire \result_x1_x3_real[11]~q ;
wire \result_x2_x4_real[10]~q ;
wire \result_x1_x3_real[10]~q ;
wire \result_x2_x4_real[9]~q ;
wire \result_x1_x3_real[9]~q ;
wire \result_x2_x4_real[8]~q ;
wire \result_x1_x3_real[8]~q ;
wire \result_x2_x4_real[7]~q ;
wire \result_x1_x3_real[7]~q ;
wire \result_x2_x4_real[6]~q ;
wire \result_x1_x3_real[6]~q ;
wire \result_x2_x4_real[5]~q ;
wire \result_x1_x3_real[5]~q ;
wire \result_x2_x4_real[4]~q ;
wire \result_x1_x3_real[4]~q ;
wire \result_x2_x4_real[3]~q ;
wire \result_x1_x3_real[3]~q ;
wire \butterfly_st_real[3]~27 ;
wire \butterfly_st_real[3]~26_combout ;
wire \butterfly_st_real[4]~29 ;
wire \butterfly_st_real[4]~28_combout ;
wire \butterfly_st_real[5]~31 ;
wire \butterfly_st_real[5]~30_combout ;
wire \butterfly_st_real[6]~33 ;
wire \butterfly_st_real[6]~32_combout ;
wire \butterfly_st_real[7]~35 ;
wire \butterfly_st_real[7]~34_combout ;
wire \butterfly_st_real[8]~37 ;
wire \butterfly_st_real[8]~36_combout ;
wire \butterfly_st_real[9]~39 ;
wire \butterfly_st_real[9]~38_combout ;
wire \butterfly_st_real[10]~41 ;
wire \butterfly_st_real[10]~40_combout ;
wire \butterfly_st_real[11]~43 ;
wire \butterfly_st_real[11]~42_combout ;
wire \butterfly_st_real[12]~45 ;
wire \butterfly_st_real[12]~44_combout ;
wire \butterfly_st_real[13]~47 ;
wire \butterfly_st_real[13]~46_combout ;
wire \butterfly_st_real[14]~49 ;
wire \butterfly_st_real[14]~48_combout ;
wire \butterfly_st_real[15]~51 ;
wire \butterfly_st_real[15]~50_combout ;
wire \butterfly_st_real[16]~53 ;
wire \butterfly_st_real[16]~52_combout ;
wire \butterfly_st_real[17]~54_combout ;
wire \result_x2_x4_imag[0]~18_cout ;
wire \result_x2_x4_imag[0]~20 ;
wire \result_x2_x4_imag[0]~19_combout ;
wire \result_x2_x4_imag[1]~22 ;
wire \result_x2_x4_imag[1]~21_combout ;
wire \result_x2_x4_imag[2]~24 ;
wire \result_x2_x4_imag[2]~23_combout ;
wire \result_x1_x3_imag[0]~18_cout ;
wire \result_x1_x3_imag[0]~20 ;
wire \result_x1_x3_imag[0]~19_combout ;
wire \result_x1_x3_imag[1]~22 ;
wire \result_x1_x3_imag[1]~21_combout ;
wire \result_x1_x3_imag[2]~24 ;
wire \result_x1_x3_imag[2]~23_combout ;
wire \result_x2_x4_imag[3]~26 ;
wire \result_x2_x4_imag[3]~25_combout ;
wire \result_x2_x4_imag[4]~28 ;
wire \result_x2_x4_imag[4]~27_combout ;
wire \result_x2_x4_imag[5]~30 ;
wire \result_x2_x4_imag[5]~29_combout ;
wire \result_x2_x4_imag[6]~32 ;
wire \result_x2_x4_imag[6]~31_combout ;
wire \result_x2_x4_imag[7]~34 ;
wire \result_x2_x4_imag[7]~33_combout ;
wire \result_x2_x4_imag[8]~36 ;
wire \result_x2_x4_imag[8]~35_combout ;
wire \result_x2_x4_imag[9]~38 ;
wire \result_x2_x4_imag[9]~37_combout ;
wire \result_x2_x4_imag[10]~40 ;
wire \result_x2_x4_imag[10]~39_combout ;
wire \result_x2_x4_imag[11]~42 ;
wire \result_x2_x4_imag[11]~41_combout ;
wire \result_x2_x4_imag[12]~44 ;
wire \result_x2_x4_imag[12]~43_combout ;
wire \result_x2_x4_imag[13]~46 ;
wire \result_x2_x4_imag[13]~45_combout ;
wire \result_x2_x4_imag[14]~48 ;
wire \result_x2_x4_imag[14]~47_combout ;
wire \result_x2_x4_imag[15]~50 ;
wire \result_x2_x4_imag[15]~49_combout ;
wire \result_x2_x4_imag[16]~51_combout ;
wire \result_x1_x3_imag[3]~26 ;
wire \result_x1_x3_imag[3]~25_combout ;
wire \result_x1_x3_imag[4]~28 ;
wire \result_x1_x3_imag[4]~27_combout ;
wire \result_x1_x3_imag[5]~30 ;
wire \result_x1_x3_imag[5]~29_combout ;
wire \result_x1_x3_imag[6]~32 ;
wire \result_x1_x3_imag[6]~31_combout ;
wire \result_x1_x3_imag[7]~34 ;
wire \result_x1_x3_imag[7]~33_combout ;
wire \result_x1_x3_imag[8]~36 ;
wire \result_x1_x3_imag[8]~35_combout ;
wire \result_x1_x3_imag[9]~38 ;
wire \result_x1_x3_imag[9]~37_combout ;
wire \result_x1_x3_imag[10]~40 ;
wire \result_x1_x3_imag[10]~39_combout ;
wire \result_x1_x3_imag[11]~42 ;
wire \result_x1_x3_imag[11]~41_combout ;
wire \result_x1_x3_imag[12]~44 ;
wire \result_x1_x3_imag[12]~43_combout ;
wire \result_x1_x3_imag[13]~46 ;
wire \result_x1_x3_imag[13]~45_combout ;
wire \result_x1_x3_imag[14]~48 ;
wire \result_x1_x3_imag[14]~47_combout ;
wire \result_x1_x3_imag[15]~50 ;
wire \result_x1_x3_imag[15]~49_combout ;
wire \result_x1_x3_imag[16]~51_combout ;
wire \result_x2_x4_real[0]~18_cout ;
wire \result_x2_x4_real[0]~20 ;
wire \result_x2_x4_real[0]~19_combout ;
wire \result_x2_x4_real[1]~22 ;
wire \result_x2_x4_real[1]~21_combout ;
wire \result_x2_x4_real[2]~24 ;
wire \result_x2_x4_real[2]~23_combout ;
wire \result_x1_x3_real[0]~18_cout ;
wire \result_x1_x3_real[0]~20 ;
wire \result_x1_x3_real[0]~19_combout ;
wire \result_x1_x3_real[1]~22 ;
wire \result_x1_x3_real[1]~21_combout ;
wire \result_x1_x3_real[2]~24 ;
wire \result_x1_x3_real[2]~23_combout ;
wire \result_x2_x4_real[3]~26 ;
wire \result_x2_x4_real[3]~25_combout ;
wire \result_x2_x4_real[4]~28 ;
wire \result_x2_x4_real[4]~27_combout ;
wire \result_x2_x4_real[5]~30 ;
wire \result_x2_x4_real[5]~29_combout ;
wire \result_x2_x4_real[6]~32 ;
wire \result_x2_x4_real[6]~31_combout ;
wire \result_x2_x4_real[7]~34 ;
wire \result_x2_x4_real[7]~33_combout ;
wire \result_x2_x4_real[8]~36 ;
wire \result_x2_x4_real[8]~35_combout ;
wire \result_x2_x4_real[9]~38 ;
wire \result_x2_x4_real[9]~37_combout ;
wire \result_x2_x4_real[10]~40 ;
wire \result_x2_x4_real[10]~39_combout ;
wire \result_x2_x4_real[11]~42 ;
wire \result_x2_x4_real[11]~41_combout ;
wire \result_x2_x4_real[12]~44 ;
wire \result_x2_x4_real[12]~43_combout ;
wire \result_x2_x4_real[13]~46 ;
wire \result_x2_x4_real[13]~45_combout ;
wire \result_x2_x4_real[14]~48 ;
wire \result_x2_x4_real[14]~47_combout ;
wire \result_x2_x4_real[15]~50 ;
wire \result_x2_x4_real[15]~49_combout ;
wire \result_x2_x4_real[16]~51_combout ;
wire \result_x1_x3_real[3]~26 ;
wire \result_x1_x3_real[3]~25_combout ;
wire \result_x1_x3_real[4]~28 ;
wire \result_x1_x3_real[4]~27_combout ;
wire \result_x1_x3_real[5]~30 ;
wire \result_x1_x3_real[5]~29_combout ;
wire \result_x1_x3_real[6]~32 ;
wire \result_x1_x3_real[6]~31_combout ;
wire \result_x1_x3_real[7]~34 ;
wire \result_x1_x3_real[7]~33_combout ;
wire \result_x1_x3_real[8]~36 ;
wire \result_x1_x3_real[8]~35_combout ;
wire \result_x1_x3_real[9]~38 ;
wire \result_x1_x3_real[9]~37_combout ;
wire \result_x1_x3_real[10]~40 ;
wire \result_x1_x3_real[10]~39_combout ;
wire \result_x1_x3_real[11]~42 ;
wire \result_x1_x3_real[11]~41_combout ;
wire \result_x1_x3_real[12]~44 ;
wire \result_x1_x3_real[12]~43_combout ;
wire \result_x1_x3_real[13]~46 ;
wire \result_x1_x3_real[13]~45_combout ;
wire \result_x1_x3_real[14]~48 ;
wire \result_x1_x3_real[14]~47_combout ;
wire \result_x1_x3_real[15]~50 ;
wire \result_x1_x3_real[15]~49_combout ;
wire \result_x1_x3_real[16]~51_combout ;
wire \bfp_scale|i_array_out[0][2]~q ;
wire \bfp_scale|i_array_out[0][13]~q ;
wire \bfp_scale|i_array_out[0][12]~q ;
wire \bfp_scale|i_array_out[0][11]~q ;
wire \bfp_scale|i_array_out[0][10]~q ;
wire \bfp_scale|i_array_out[0][9]~q ;
wire \bfp_scale|i_array_out[0][8]~q ;
wire \bfp_scale|i_array_out[0][7]~q ;
wire \bfp_scale|i_array_out[0][6]~q ;
wire \bfp_scale|i_array_out[0][5]~q ;
wire \bfp_scale|i_array_out[0][4]~q ;
wire \bfp_scale|i_array_out[0][3]~q ;
wire \bfp_scale|r_array_out[0][2]~q ;
wire \bfp_scale|r_array_out[0][13]~q ;
wire \bfp_scale|r_array_out[0][12]~q ;
wire \bfp_scale|r_array_out[0][11]~q ;
wire \bfp_scale|r_array_out[0][10]~q ;
wire \bfp_scale|r_array_out[0][9]~q ;
wire \bfp_scale|r_array_out[0][8]~q ;
wire \bfp_scale|r_array_out[0][7]~q ;
wire \bfp_scale|r_array_out[0][6]~q ;
wire \bfp_scale|r_array_out[0][5]~q ;
wire \bfp_scale|r_array_out[0][4]~q ;
wire \bfp_scale|r_array_out[0][3]~q ;
wire \si[0]~q ;
wire \Add10~1_combout ;
wire \Add10~2_combout ;
wire \Add10~3_combout ;
wire \Add10~4_combout ;
wire \Add10~5_combout ;
wire \Add10~6_combout ;
wire \Add10~7_combout ;
wire \Add10~8_combout ;
wire \Add10~9_combout ;
wire \Add10~10_combout ;
wire \Add10~11_combout ;
wire \Add10~12_combout ;
wire \Add10~13_combout ;
wire \Add10~14_combout ;
wire \Add10~15_combout ;
wire \Add10~16_combout ;
wire \Add10~17_combout ;
wire \Add4~1_combout ;
wire \Add4~2_combout ;
wire \Add4~3_combout ;
wire \Add4~4_combout ;
wire \Add4~5_combout ;
wire \Add4~6_combout ;
wire \Add4~7_combout ;
wire \Add4~8_combout ;
wire \Add4~9_combout ;
wire \Add4~10_combout ;
wire \Add4~11_combout ;
wire \Add4~12_combout ;
wire \Add4~13_combout ;
wire \Add4~14_combout ;
wire \Add4~15_combout ;
wire \Add4~16_combout ;
wire \Add4~17_combout ;
wire \sel_arr[9][1]~q ;
wire \si~0_combout ;
wire \si[1]~q ;
wire \x_4_imag_held[2]~q ;
wire \Add8~1_combout ;
wire \x_2_imag_held[2]~q ;
wire \x_4_imag_held[1]~q ;
wire \Add8~2_combout ;
wire \x_2_imag_held[1]~q ;
wire \x_4_imag_held[0]~q ;
wire \Add8~3_combout ;
wire \x_2_imag_held[0]~q ;
wire \x_3_imag_held[2]~q ;
wire \Add6~1_combout ;
wire \x_1_imag_held[2]~q ;
wire \x_3_imag_held[1]~q ;
wire \Add6~2_combout ;
wire \x_1_imag_held[1]~q ;
wire \x_3_imag_held[0]~q ;
wire \Add6~3_combout ;
wire \x_1_imag_held[0]~q ;
wire \x_4_imag_held[15]~q ;
wire \Add8~4_combout ;
wire \x_2_imag_held[15]~q ;
wire \x_4_imag_held[14]~q ;
wire \Add8~5_combout ;
wire \x_2_imag_held[14]~q ;
wire \x_4_imag_held[13]~q ;
wire \Add8~6_combout ;
wire \x_2_imag_held[13]~q ;
wire \x_4_imag_held[12]~q ;
wire \Add8~7_combout ;
wire \x_2_imag_held[12]~q ;
wire \x_4_imag_held[11]~q ;
wire \Add8~8_combout ;
wire \x_2_imag_held[11]~q ;
wire \x_4_imag_held[10]~q ;
wire \Add8~9_combout ;
wire \x_2_imag_held[10]~q ;
wire \x_4_imag_held[9]~q ;
wire \Add8~10_combout ;
wire \x_2_imag_held[9]~q ;
wire \x_4_imag_held[8]~q ;
wire \Add8~11_combout ;
wire \x_2_imag_held[8]~q ;
wire \x_4_imag_held[7]~q ;
wire \Add8~12_combout ;
wire \x_2_imag_held[7]~q ;
wire \x_4_imag_held[6]~q ;
wire \Add8~13_combout ;
wire \x_2_imag_held[6]~q ;
wire \x_4_imag_held[5]~q ;
wire \Add8~14_combout ;
wire \x_2_imag_held[5]~q ;
wire \x_4_imag_held[4]~q ;
wire \Add8~15_combout ;
wire \x_2_imag_held[4]~q ;
wire \x_4_imag_held[3]~q ;
wire \Add8~16_combout ;
wire \x_2_imag_held[3]~q ;
wire \x_3_imag_held[15]~q ;
wire \Add6~4_combout ;
wire \x_1_imag_held[15]~q ;
wire \x_3_imag_held[14]~q ;
wire \Add6~5_combout ;
wire \x_1_imag_held[14]~q ;
wire \x_3_imag_held[13]~q ;
wire \Add6~6_combout ;
wire \x_1_imag_held[13]~q ;
wire \x_3_imag_held[12]~q ;
wire \Add6~7_combout ;
wire \x_1_imag_held[12]~q ;
wire \x_3_imag_held[11]~q ;
wire \Add6~8_combout ;
wire \x_1_imag_held[11]~q ;
wire \x_3_imag_held[10]~q ;
wire \Add6~9_combout ;
wire \x_1_imag_held[10]~q ;
wire \x_3_imag_held[9]~q ;
wire \Add6~10_combout ;
wire \x_1_imag_held[9]~q ;
wire \x_3_imag_held[8]~q ;
wire \Add6~11_combout ;
wire \x_1_imag_held[8]~q ;
wire \x_3_imag_held[7]~q ;
wire \Add6~12_combout ;
wire \x_1_imag_held[7]~q ;
wire \x_3_imag_held[6]~q ;
wire \Add6~13_combout ;
wire \x_1_imag_held[6]~q ;
wire \x_3_imag_held[5]~q ;
wire \Add6~14_combout ;
wire \x_1_imag_held[5]~q ;
wire \x_3_imag_held[4]~q ;
wire \Add6~15_combout ;
wire \x_1_imag_held[4]~q ;
wire \x_3_imag_held[3]~q ;
wire \Add6~16_combout ;
wire \x_1_imag_held[3]~q ;
wire \sel_arr[9][0]~q ;
wire \Mux264~0_combout ;
wire \x_4_real_held[2]~q ;
wire \Add2~1_combout ;
wire \x_2_real_held[2]~q ;
wire \x_4_real_held[1]~q ;
wire \Add2~2_combout ;
wire \x_2_real_held[1]~q ;
wire \x_4_real_held[0]~q ;
wire \Add2~3_combout ;
wire \x_2_real_held[0]~q ;
wire \x_3_real_held[2]~q ;
wire \Add0~1_combout ;
wire \x_1_real_held[2]~q ;
wire \x_3_real_held[1]~q ;
wire \Add0~2_combout ;
wire \x_1_real_held[1]~q ;
wire \x_3_real_held[0]~q ;
wire \Add0~3_combout ;
wire \x_1_real_held[0]~q ;
wire \x_4_real_held[15]~q ;
wire \Add2~4_combout ;
wire \x_2_real_held[15]~q ;
wire \x_4_real_held[14]~q ;
wire \Add2~5_combout ;
wire \x_2_real_held[14]~q ;
wire \x_4_real_held[13]~q ;
wire \Add2~6_combout ;
wire \x_2_real_held[13]~q ;
wire \x_4_real_held[12]~q ;
wire \Add2~7_combout ;
wire \x_2_real_held[12]~q ;
wire \x_4_real_held[11]~q ;
wire \Add2~8_combout ;
wire \x_2_real_held[11]~q ;
wire \x_4_real_held[10]~q ;
wire \Add2~9_combout ;
wire \x_2_real_held[10]~q ;
wire \x_4_real_held[9]~q ;
wire \Add2~10_combout ;
wire \x_2_real_held[9]~q ;
wire \x_4_real_held[8]~q ;
wire \Add2~11_combout ;
wire \x_2_real_held[8]~q ;
wire \x_4_real_held[7]~q ;
wire \Add2~12_combout ;
wire \x_2_real_held[7]~q ;
wire \x_4_real_held[6]~q ;
wire \Add2~13_combout ;
wire \x_2_real_held[6]~q ;
wire \x_4_real_held[5]~q ;
wire \Add2~14_combout ;
wire \x_2_real_held[5]~q ;
wire \x_4_real_held[4]~q ;
wire \Add2~15_combout ;
wire \x_2_real_held[4]~q ;
wire \x_4_real_held[3]~q ;
wire \Add2~16_combout ;
wire \x_2_real_held[3]~q ;
wire \x_3_real_held[15]~q ;
wire \Add0~4_combout ;
wire \x_1_real_held[15]~q ;
wire \x_3_real_held[14]~q ;
wire \Add0~5_combout ;
wire \x_1_real_held[14]~q ;
wire \x_3_real_held[13]~q ;
wire \Add0~6_combout ;
wire \x_1_real_held[13]~q ;
wire \x_3_real_held[12]~q ;
wire \Add0~7_combout ;
wire \x_1_real_held[12]~q ;
wire \x_3_real_held[11]~q ;
wire \Add0~8_combout ;
wire \x_1_real_held[11]~q ;
wire \x_3_real_held[10]~q ;
wire \Add0~9_combout ;
wire \x_1_real_held[10]~q ;
wire \x_3_real_held[9]~q ;
wire \Add0~10_combout ;
wire \x_1_real_held[9]~q ;
wire \x_3_real_held[8]~q ;
wire \Add0~11_combout ;
wire \x_1_real_held[8]~q ;
wire \x_3_real_held[7]~q ;
wire \Add0~12_combout ;
wire \x_1_real_held[7]~q ;
wire \x_3_real_held[6]~q ;
wire \Add0~13_combout ;
wire \x_1_real_held[6]~q ;
wire \x_3_real_held[5]~q ;
wire \Add0~14_combout ;
wire \x_1_real_held[5]~q ;
wire \x_3_real_held[4]~q ;
wire \Add0~15_combout ;
wire \x_1_real_held[4]~q ;
wire \x_3_real_held[3]~q ;
wire \Add0~16_combout ;
wire \x_1_real_held[3]~q ;
wire \sel_arr[8][1]~q ;
wire \sel_arr~0_combout ;
wire \si~1_combout ;
wire \butterfly_st1[3][1][2]~q ;
wire \Mux261~0_combout ;
wire \butterfly_st1[1][1][2]~q ;
wire \Mux227~0_combout ;
wire \butterfly_st1[3][1][1]~q ;
wire \Mux262~0_combout ;
wire \butterfly_st1[1][1][1]~q ;
wire \Mux228~0_combout ;
wire \butterfly_st1[3][1][0]~q ;
wire \Mux263~0_combout ;
wire \butterfly_st1[1][1][0]~q ;
wire \Mux229~0_combout ;
wire \butterfly_st1[2][1][2]~q ;
wire \x_3_imag_held[0]~0_combout ;
wire \butterfly_st1[0][1][2]~q ;
wire \butterfly_st1[2][1][1]~q ;
wire \butterfly_st1[0][1][1]~q ;
wire \butterfly_st1[2][1][0]~q ;
wire \butterfly_st1[0][1][0]~q ;
wire \butterfly_st1[3][1][15]~q ;
wire \Mux248~0_combout ;
wire \butterfly_st1[1][1][15]~q ;
wire \Mux214~0_combout ;
wire \butterfly_st1[3][1][14]~q ;
wire \Mux249~0_combout ;
wire \butterfly_st1[1][1][14]~q ;
wire \Mux215~0_combout ;
wire \butterfly_st1[3][1][13]~q ;
wire \Mux250~0_combout ;
wire \butterfly_st1[1][1][13]~q ;
wire \Mux216~0_combout ;
wire \butterfly_st1[3][1][12]~q ;
wire \Mux251~0_combout ;
wire \butterfly_st1[1][1][12]~q ;
wire \Mux217~0_combout ;
wire \butterfly_st1[3][1][11]~q ;
wire \Mux252~0_combout ;
wire \butterfly_st1[1][1][11]~q ;
wire \Mux218~0_combout ;
wire \butterfly_st1[3][1][10]~q ;
wire \Mux253~0_combout ;
wire \butterfly_st1[1][1][10]~q ;
wire \Mux219~0_combout ;
wire \butterfly_st1[3][1][9]~q ;
wire \Mux254~0_combout ;
wire \butterfly_st1[1][1][9]~q ;
wire \Mux220~0_combout ;
wire \butterfly_st1[3][1][8]~q ;
wire \Mux255~0_combout ;
wire \butterfly_st1[1][1][8]~q ;
wire \Mux221~0_combout ;
wire \butterfly_st1[3][1][7]~q ;
wire \Mux256~0_combout ;
wire \butterfly_st1[1][1][7]~q ;
wire \Mux222~0_combout ;
wire \butterfly_st1[3][1][6]~q ;
wire \Mux257~0_combout ;
wire \butterfly_st1[1][1][6]~q ;
wire \Mux223~0_combout ;
wire \butterfly_st1[3][1][5]~q ;
wire \Mux258~0_combout ;
wire \butterfly_st1[1][1][5]~q ;
wire \Mux224~0_combout ;
wire \butterfly_st1[3][1][4]~q ;
wire \Mux259~0_combout ;
wire \butterfly_st1[1][1][4]~q ;
wire \Mux225~0_combout ;
wire \butterfly_st1[3][1][3]~q ;
wire \Mux260~0_combout ;
wire \butterfly_st1[1][1][3]~q ;
wire \Mux226~0_combout ;
wire \butterfly_st1[2][1][15]~q ;
wire \butterfly_st1[0][1][15]~q ;
wire \butterfly_st1[2][1][14]~q ;
wire \butterfly_st1[0][1][14]~q ;
wire \butterfly_st1[2][1][13]~q ;
wire \butterfly_st1[0][1][13]~q ;
wire \butterfly_st1[2][1][12]~q ;
wire \butterfly_st1[0][1][12]~q ;
wire \butterfly_st1[2][1][11]~q ;
wire \butterfly_st1[0][1][11]~q ;
wire \butterfly_st1[2][1][10]~q ;
wire \butterfly_st1[0][1][10]~q ;
wire \butterfly_st1[2][1][9]~q ;
wire \butterfly_st1[0][1][9]~q ;
wire \butterfly_st1[2][1][8]~q ;
wire \butterfly_st1[0][1][8]~q ;
wire \butterfly_st1[2][1][7]~q ;
wire \butterfly_st1[0][1][7]~q ;
wire \butterfly_st1[2][1][6]~q ;
wire \butterfly_st1[0][1][6]~q ;
wire \butterfly_st1[2][1][5]~q ;
wire \butterfly_st1[0][1][5]~q ;
wire \butterfly_st1[2][1][4]~q ;
wire \butterfly_st1[0][1][4]~q ;
wire \butterfly_st1[2][1][3]~q ;
wire \butterfly_st1[0][1][3]~q ;
wire \sel_arr[8][0]~q ;
wire \sel_arr~1_combout ;
wire \butterfly_st1[3][0][2]~q ;
wire \Mux193~0_combout ;
wire \butterfly_st1[1][0][2]~q ;
wire \Mux159~0_combout ;
wire \butterfly_st1[3][0][1]~q ;
wire \Mux194~0_combout ;
wire \butterfly_st1[1][0][1]~q ;
wire \Mux160~0_combout ;
wire \butterfly_st1[3][0][0]~q ;
wire \Mux195~0_combout ;
wire \butterfly_st1[1][0][0]~q ;
wire \Mux161~0_combout ;
wire \butterfly_st1[2][0][2]~q ;
wire \butterfly_st1[0][0][2]~q ;
wire \butterfly_st1[2][0][1]~q ;
wire \butterfly_st1[0][0][1]~q ;
wire \butterfly_st1[2][0][0]~q ;
wire \butterfly_st1[0][0][0]~q ;
wire \butterfly_st1[3][0][15]~q ;
wire \Mux180~0_combout ;
wire \butterfly_st1[1][0][15]~q ;
wire \Mux146~0_combout ;
wire \butterfly_st1[3][0][14]~q ;
wire \Mux181~0_combout ;
wire \butterfly_st1[1][0][14]~q ;
wire \Mux147~0_combout ;
wire \butterfly_st1[3][0][13]~q ;
wire \Mux182~0_combout ;
wire \butterfly_st1[1][0][13]~q ;
wire \Mux148~0_combout ;
wire \butterfly_st1[3][0][12]~q ;
wire \Mux183~0_combout ;
wire \butterfly_st1[1][0][12]~q ;
wire \Mux149~0_combout ;
wire \butterfly_st1[3][0][11]~q ;
wire \Mux184~0_combout ;
wire \butterfly_st1[1][0][11]~q ;
wire \Mux150~0_combout ;
wire \butterfly_st1[3][0][10]~q ;
wire \Mux185~0_combout ;
wire \butterfly_st1[1][0][10]~q ;
wire \Mux151~0_combout ;
wire \butterfly_st1[3][0][9]~q ;
wire \Mux186~0_combout ;
wire \butterfly_st1[1][0][9]~q ;
wire \Mux152~0_combout ;
wire \butterfly_st1[3][0][8]~q ;
wire \Mux187~0_combout ;
wire \butterfly_st1[1][0][8]~q ;
wire \Mux153~0_combout ;
wire \butterfly_st1[3][0][7]~q ;
wire \Mux188~0_combout ;
wire \butterfly_st1[1][0][7]~q ;
wire \Mux154~0_combout ;
wire \butterfly_st1[3][0][6]~q ;
wire \Mux189~0_combout ;
wire \butterfly_st1[1][0][6]~q ;
wire \Mux155~0_combout ;
wire \butterfly_st1[3][0][5]~q ;
wire \Mux190~0_combout ;
wire \butterfly_st1[1][0][5]~q ;
wire \Mux156~0_combout ;
wire \butterfly_st1[3][0][4]~q ;
wire \Mux191~0_combout ;
wire \butterfly_st1[1][0][4]~q ;
wire \Mux157~0_combout ;
wire \butterfly_st1[3][0][3]~q ;
wire \Mux192~0_combout ;
wire \butterfly_st1[1][0][3]~q ;
wire \Mux158~0_combout ;
wire \butterfly_st1[2][0][15]~q ;
wire \butterfly_st1[0][0][15]~q ;
wire \butterfly_st1[2][0][14]~q ;
wire \butterfly_st1[0][0][14]~q ;
wire \butterfly_st1[2][0][13]~q ;
wire \butterfly_st1[0][0][13]~q ;
wire \butterfly_st1[2][0][12]~q ;
wire \butterfly_st1[0][0][12]~q ;
wire \butterfly_st1[2][0][11]~q ;
wire \butterfly_st1[0][0][11]~q ;
wire \butterfly_st1[2][0][10]~q ;
wire \butterfly_st1[0][0][10]~q ;
wire \butterfly_st1[2][0][9]~q ;
wire \butterfly_st1[0][0][9]~q ;
wire \butterfly_st1[2][0][8]~q ;
wire \butterfly_st1[0][0][8]~q ;
wire \butterfly_st1[2][0][7]~q ;
wire \butterfly_st1[0][0][7]~q ;
wire \butterfly_st1[2][0][6]~q ;
wire \butterfly_st1[0][0][6]~q ;
wire \butterfly_st1[2][0][5]~q ;
wire \butterfly_st1[0][0][5]~q ;
wire \butterfly_st1[2][0][4]~q ;
wire \butterfly_st1[0][0][4]~q ;
wire \butterfly_st1[2][0][3]~q ;
wire \butterfly_st1[0][0][3]~q ;
wire \sel_arr[7][1]~q ;
wire \sel_arr~2_combout ;
wire \butterfly_st1~0_combout ;
wire \sel_arr[5][0]~q ;
wire \sel_arr[5][1]~q ;
wire \butterfly_st1[3][1][0]~0_combout ;
wire \butterfly_st1[1][1][0]~0_combout ;
wire \bfp_scale|i_array_out[0][1]~q ;
wire \butterfly_st1~1_combout ;
wire \bfp_scale|i_array_out[0][0]~q ;
wire \butterfly_st1~2_combout ;
wire \butterfly_st1[2][1][0]~0_combout ;
wire \butterfly_st1[0][1][0]~0_combout ;
wire \bfp_scale|i_array_out[0][15]~q ;
wire \butterfly_st1~3_combout ;
wire \bfp_scale|i_array_out[0][14]~q ;
wire \butterfly_st1~4_combout ;
wire \butterfly_st1~5_combout ;
wire \butterfly_st1~6_combout ;
wire \butterfly_st1~7_combout ;
wire \butterfly_st1~8_combout ;
wire \butterfly_st1~9_combout ;
wire \butterfly_st1~10_combout ;
wire \butterfly_st1~11_combout ;
wire \butterfly_st1~12_combout ;
wire \butterfly_st1~13_combout ;
wire \butterfly_st1~14_combout ;
wire \butterfly_st1~15_combout ;
wire \sel_arr[7][0]~q ;
wire \sel_arr~3_combout ;
wire \butterfly_st1~16_combout ;
wire \bfp_scale|r_array_out[0][1]~q ;
wire \butterfly_st1~17_combout ;
wire \bfp_scale|r_array_out[0][0]~q ;
wire \butterfly_st1~18_combout ;
wire \bfp_scale|r_array_out[0][15]~q ;
wire \butterfly_st1~19_combout ;
wire \bfp_scale|r_array_out[0][14]~q ;
wire \butterfly_st1~20_combout ;
wire \butterfly_st1~21_combout ;
wire \butterfly_st1~22_combout ;
wire \butterfly_st1~23_combout ;
wire \butterfly_st1~24_combout ;
wire \butterfly_st1~25_combout ;
wire \butterfly_st1~26_combout ;
wire \butterfly_st1~27_combout ;
wire \butterfly_st1~28_combout ;
wire \butterfly_st1~29_combout ;
wire \butterfly_st1~30_combout ;
wire \butterfly_st1~31_combout ;
wire \sel_arr[6][1]~q ;
wire \sel_arr~4_combout ;
wire \sel_arr[4][0]~q ;
wire \sel_arr~5_combout ;
wire \sel_arr[4][1]~q ;
wire \sel_arr~6_combout ;
wire \sel_arr[6][0]~q ;
wire \sel_arr~7_combout ;
wire \sel_arr~8_combout ;
wire \sel_arr[3][0]~q ;
wire \sel_arr~9_combout ;
wire \sel_arr[3][1]~q ;
wire \sel_arr~10_combout ;
wire \sel_arr~11_combout ;
wire \sel_arr[2][0]~q ;
wire \sel_arr~12_combout ;
wire \sel_arr[2][1]~q ;
wire \sel_arr~13_combout ;
wire \sel_arr[1][0]~q ;
wire \sel_arr~14_combout ;
wire \sel_arr[1][1]~q ;
wire \sel_arr~15_combout ;
wire \sel_arr[0][0]~q ;
wire \sel_arr~16_combout ;
wire \sel_arr[0][1]~q ;
wire \sel_arr~17_combout ;
wire \sel_arr~18_combout ;
wire \sel_arr~19_combout ;


fft256_asj_fft_cmult_can_fft_121 \gen_da0:gen_canonic:cm1 (
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_2(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_12(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_15(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_161(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_171(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ),
	.twiddle_data_real_0(twiddle_data_real_0),
	.twiddle_data_real_15(twiddle_data_real_15),
	.pipeline_dffe_210(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_32(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_101(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_111(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_121(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_131(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_141(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_151(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_162(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_172(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ),
	.twiddle_data_imag_1(twiddle_data_imag_1),
	.twiddle_data_imag_2(twiddle_data_imag_2),
	.twiddle_data_imag_3(twiddle_data_imag_3),
	.twiddle_data_imag_4(twiddle_data_imag_4),
	.twiddle_data_imag_5(twiddle_data_imag_5),
	.twiddle_data_imag_6(twiddle_data_imag_6),
	.twiddle_data_imag_7(twiddle_data_imag_7),
	.twiddle_data_imag_8(twiddle_data_imag_8),
	.twiddle_data_imag_9(twiddle_data_imag_9),
	.twiddle_data_imag_10(twiddle_data_imag_10),
	.twiddle_data_imag_11(twiddle_data_imag_11),
	.twiddle_data_imag_12(twiddle_data_imag_12),
	.twiddle_data_imag_13(twiddle_data_imag_13),
	.twiddle_data_imag_14(twiddle_data_imag_14),
	.twiddle_data_imag_15(twiddle_data_imag_15),
	.global_clock_enable(global_clock_enable),
	.real_out_0(real_out_0),
	.real_out_1(real_out_1),
	.real_out_2(real_out_2),
	.real_out_3(real_out_3),
	.real_out_4(real_out_4),
	.real_out_5(real_out_5),
	.real_out_6(real_out_6),
	.real_out_7(real_out_7),
	.real_out_8(real_out_8),
	.real_out_9(real_out_9),
	.real_out_10(real_out_10),
	.real_out_11(real_out_11),
	.real_out_12(real_out_12),
	.real_out_13(real_out_13),
	.real_out_14(real_out_14),
	.real_out_15(real_out_15),
	.twiddle_data_real_1(twiddle_data_real_1),
	.twiddle_data_real_2(twiddle_data_real_2),
	.twiddle_data_real_3(twiddle_data_real_3),
	.twiddle_data_real_4(twiddle_data_real_4),
	.twiddle_data_real_5(twiddle_data_real_5),
	.twiddle_data_real_6(twiddle_data_real_6),
	.twiddle_data_real_7(twiddle_data_real_7),
	.twiddle_data_real_8(twiddle_data_real_8),
	.twiddle_data_real_9(twiddle_data_real_9),
	.twiddle_data_real_10(twiddle_data_real_10),
	.twiddle_data_real_11(twiddle_data_real_11),
	.twiddle_data_real_12(twiddle_data_real_12),
	.twiddle_data_real_13(twiddle_data_real_13),
	.twiddle_data_real_14(twiddle_data_real_14),
	.twiddle_data_imag_0(twiddle_data_imag_0),
	.clk(clk),
	.reset(reset));

fft256_asj_fft_bfp_i_fft_121 bfp_scale(
	.i_array_out_2_0(\bfp_scale|i_array_out[0][2]~q ),
	.i_array_out_13_0(\bfp_scale|i_array_out[0][13]~q ),
	.i_array_out_12_0(\bfp_scale|i_array_out[0][12]~q ),
	.i_array_out_11_0(\bfp_scale|i_array_out[0][11]~q ),
	.i_array_out_10_0(\bfp_scale|i_array_out[0][10]~q ),
	.i_array_out_9_0(\bfp_scale|i_array_out[0][9]~q ),
	.i_array_out_8_0(\bfp_scale|i_array_out[0][8]~q ),
	.i_array_out_7_0(\bfp_scale|i_array_out[0][7]~q ),
	.i_array_out_6_0(\bfp_scale|i_array_out[0][6]~q ),
	.i_array_out_5_0(\bfp_scale|i_array_out[0][5]~q ),
	.i_array_out_4_0(\bfp_scale|i_array_out[0][4]~q ),
	.i_array_out_3_0(\bfp_scale|i_array_out[0][3]~q ),
	.r_array_out_2_0(\bfp_scale|r_array_out[0][2]~q ),
	.r_array_out_13_0(\bfp_scale|r_array_out[0][13]~q ),
	.r_array_out_12_0(\bfp_scale|r_array_out[0][12]~q ),
	.r_array_out_11_0(\bfp_scale|r_array_out[0][11]~q ),
	.r_array_out_10_0(\bfp_scale|r_array_out[0][10]~q ),
	.r_array_out_9_0(\bfp_scale|r_array_out[0][9]~q ),
	.r_array_out_8_0(\bfp_scale|r_array_out[0][8]~q ),
	.r_array_out_7_0(\bfp_scale|r_array_out[0][7]~q ),
	.r_array_out_6_0(\bfp_scale|r_array_out[0][6]~q ),
	.r_array_out_5_0(\bfp_scale|r_array_out[0][5]~q ),
	.r_array_out_4_0(\bfp_scale|r_array_out[0][4]~q ),
	.r_array_out_3_0(\bfp_scale|r_array_out[0][3]~q ),
	.global_clock_enable(global_clock_enable),
	.i_array_out_1_0(\bfp_scale|i_array_out[0][1]~q ),
	.i_array_out_0_0(\bfp_scale|i_array_out[0][0]~q ),
	.i_array_out_15_0(\bfp_scale|i_array_out[0][15]~q ),
	.i_array_out_14_0(\bfp_scale|i_array_out[0][14]~q ),
	.r_array_out_1_0(\bfp_scale|r_array_out[0][1]~q ),
	.r_array_out_0_0(\bfp_scale|r_array_out[0][0]~q ),
	.r_array_out_15_0(\bfp_scale|r_array_out[0][15]~q ),
	.r_array_out_14_0(\bfp_scale|r_array_out[0][14]~q ),
	.ram_data_out_0(ram_data_out_0),
	.ram_data_out_2(ram_data_out_2),
	.slb_last_1(slb_last_1),
	.ram_data_out_1(ram_data_out_1),
	.slb_last_0(slb_last_0),
	.slb_last_2(slb_last_2),
	.ram_data_out_14(ram_data_out_14),
	.ram_data_out_12(ram_data_out_12),
	.ram_data_out_13(ram_data_out_13),
	.ram_data_out_15(ram_data_out_15),
	.ram_data_out_11(ram_data_out_11),
	.ram_data_out_10(ram_data_out_10),
	.ram_data_out_9(ram_data_out_9),
	.ram_data_out_8(ram_data_out_8),
	.ram_data_out_7(ram_data_out_7),
	.ram_data_out_6(ram_data_out_6),
	.ram_data_out_5(ram_data_out_5),
	.ram_data_out_4(ram_data_out_4),
	.ram_data_out_3(ram_data_out_3),
	.ram_data_out_16(ram_data_out_16),
	.ram_data_out_18(ram_data_out_18),
	.ram_data_out_17(ram_data_out_17),
	.ram_data_out_28(ram_data_out_28),
	.ram_data_out_29(ram_data_out_29),
	.ram_data_out_30(ram_data_out_30),
	.ram_data_out_31(ram_data_out_31),
	.ram_data_out_27(ram_data_out_27),
	.ram_data_out_26(ram_data_out_26),
	.ram_data_out_25(ram_data_out_25),
	.ram_data_out_24(ram_data_out_24),
	.ram_data_out_23(ram_data_out_23),
	.ram_data_out_22(ram_data_out_22),
	.ram_data_out_21(ram_data_out_21),
	.ram_data_out_20(ram_data_out_20),
	.ram_data_out_19(ram_data_out_19),
	.clk(clk));

fft256_asj_fft_bfp_o_fft_121 bfp_detect(
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_31(pipeline_dffe_31),
	.source_valid_ctrl_sop(source_valid_ctrl_sop),
	.stall_reg(stall_reg),
	.source_stall_int_d(source_stall_int_d),
	.global_clock_enable(global_clock_enable),
	.slb_i_0(slb_i_0),
	.Mux2(Mux2),
	.lut_out_0(lut_out_0),
	.tdl_arr_0(tdl_arr_0),
	.Mux1(Mux1),
	.lut_out_1(lut_out_1),
	.lut_out_2(lut_out_2),
	.lut_out_21(lut_out_21),
	.real_out_11(real_out_11),
	.real_out_12(real_out_12),
	.real_out_13(real_out_13),
	.real_out_14(real_out_14),
	.real_out_15(real_out_15),
	.tdl_arr_01(tdl_arr_01),
	.clk(clk),
	.reset_n(reset));

fft256_asj_fft_pround_fft_121_3 \gen_full_rnd:u1 (
	.pipeline_dffe_2(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_12(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_15(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_16(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ),
	.butterfly_st_imag_2(\butterfly_st_imag[2]~q ),
	.butterfly_st_imag_1(\butterfly_st_imag[1]~q ),
	.butterfly_st_imag_0(\butterfly_st_imag[0]~q ),
	.butterfly_st_imag_17(\butterfly_st_imag[17]~q ),
	.butterfly_st_imag_3(\butterfly_st_imag[3]~q ),
	.butterfly_st_imag_4(\butterfly_st_imag[4]~q ),
	.butterfly_st_imag_5(\butterfly_st_imag[5]~q ),
	.butterfly_st_imag_6(\butterfly_st_imag[6]~q ),
	.butterfly_st_imag_7(\butterfly_st_imag[7]~q ),
	.butterfly_st_imag_8(\butterfly_st_imag[8]~q ),
	.butterfly_st_imag_9(\butterfly_st_imag[9]~q ),
	.butterfly_st_imag_10(\butterfly_st_imag[10]~q ),
	.butterfly_st_imag_11(\butterfly_st_imag[11]~q ),
	.butterfly_st_imag_12(\butterfly_st_imag[12]~q ),
	.butterfly_st_imag_13(\butterfly_st_imag[13]~q ),
	.butterfly_st_imag_14(\butterfly_st_imag[14]~q ),
	.butterfly_st_imag_15(\butterfly_st_imag[15]~q ),
	.butterfly_st_imag_16(\butterfly_st_imag[16]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fft256_asj_fft_pround_fft_121_2 \gen_full_rnd:u0 (
	.pipeline_dffe_2(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_12(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_15(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_16(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ),
	.butterfly_st_real_2(\butterfly_st_real[2]~q ),
	.butterfly_st_real_1(\butterfly_st_real[1]~q ),
	.butterfly_st_real_0(\butterfly_st_real[0]~q ),
	.butterfly_st_real_17(\butterfly_st_real[17]~q ),
	.butterfly_st_real_3(\butterfly_st_real[3]~q ),
	.butterfly_st_real_4(\butterfly_st_real[4]~q ),
	.butterfly_st_real_5(\butterfly_st_real[5]~q ),
	.butterfly_st_real_6(\butterfly_st_real[6]~q ),
	.butterfly_st_real_7(\butterfly_st_real[7]~q ),
	.butterfly_st_real_8(\butterfly_st_real[8]~q ),
	.butterfly_st_real_9(\butterfly_st_real[9]~q ),
	.butterfly_st_real_10(\butterfly_st_real[10]~q ),
	.butterfly_st_real_11(\butterfly_st_real[11]~q ),
	.butterfly_st_real_12(\butterfly_st_real[12]~q ),
	.butterfly_st_real_13(\butterfly_st_real[13]~q ),
	.butterfly_st_real_14(\butterfly_st_real[14]~q ),
	.butterfly_st_real_15(\butterfly_st_real[15]~q ),
	.butterfly_st_real_16(\butterfly_st_real[16]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

dffeas \butterfly_st_imag[2] (
	.clk(clk),
	.d(\butterfly_st_imag[2]~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[2]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[2] .is_wysiwyg = "true";
defparam \butterfly_st_imag[2] .power_up = "low";

dffeas \butterfly_st_imag[1] (
	.clk(clk),
	.d(\butterfly_st_imag[1]~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[1]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[1] .is_wysiwyg = "true";
defparam \butterfly_st_imag[1] .power_up = "low";

dffeas \butterfly_st_imag[0] (
	.clk(clk),
	.d(\butterfly_st_imag[0]~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[0]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[0] .is_wysiwyg = "true";
defparam \butterfly_st_imag[0] .power_up = "low";

dffeas \butterfly_st_imag[17] (
	.clk(clk),
	.d(\butterfly_st_imag[17]~54_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[17]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[17] .is_wysiwyg = "true";
defparam \butterfly_st_imag[17] .power_up = "low";

dffeas \butterfly_st_imag[3] (
	.clk(clk),
	.d(\butterfly_st_imag[3]~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[3]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[3] .is_wysiwyg = "true";
defparam \butterfly_st_imag[3] .power_up = "low";

dffeas \butterfly_st_imag[4] (
	.clk(clk),
	.d(\butterfly_st_imag[4]~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[4]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[4] .is_wysiwyg = "true";
defparam \butterfly_st_imag[4] .power_up = "low";

dffeas \butterfly_st_imag[5] (
	.clk(clk),
	.d(\butterfly_st_imag[5]~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[5]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[5] .is_wysiwyg = "true";
defparam \butterfly_st_imag[5] .power_up = "low";

dffeas \butterfly_st_imag[6] (
	.clk(clk),
	.d(\butterfly_st_imag[6]~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[6]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[6] .is_wysiwyg = "true";
defparam \butterfly_st_imag[6] .power_up = "low";

dffeas \butterfly_st_imag[7] (
	.clk(clk),
	.d(\butterfly_st_imag[7]~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[7]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[7] .is_wysiwyg = "true";
defparam \butterfly_st_imag[7] .power_up = "low";

dffeas \butterfly_st_imag[8] (
	.clk(clk),
	.d(\butterfly_st_imag[8]~36_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[8]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[8] .is_wysiwyg = "true";
defparam \butterfly_st_imag[8] .power_up = "low";

dffeas \butterfly_st_imag[9] (
	.clk(clk),
	.d(\butterfly_st_imag[9]~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[9]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[9] .is_wysiwyg = "true";
defparam \butterfly_st_imag[9] .power_up = "low";

dffeas \butterfly_st_imag[10] (
	.clk(clk),
	.d(\butterfly_st_imag[10]~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[10]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[10] .is_wysiwyg = "true";
defparam \butterfly_st_imag[10] .power_up = "low";

dffeas \butterfly_st_imag[11] (
	.clk(clk),
	.d(\butterfly_st_imag[11]~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[11]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[11] .is_wysiwyg = "true";
defparam \butterfly_st_imag[11] .power_up = "low";

dffeas \butterfly_st_imag[12] (
	.clk(clk),
	.d(\butterfly_st_imag[12]~44_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[12]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[12] .is_wysiwyg = "true";
defparam \butterfly_st_imag[12] .power_up = "low";

dffeas \butterfly_st_imag[13] (
	.clk(clk),
	.d(\butterfly_st_imag[13]~46_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[13]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[13] .is_wysiwyg = "true";
defparam \butterfly_st_imag[13] .power_up = "low";

dffeas \butterfly_st_imag[14] (
	.clk(clk),
	.d(\butterfly_st_imag[14]~48_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[14]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[14] .is_wysiwyg = "true";
defparam \butterfly_st_imag[14] .power_up = "low";

dffeas \butterfly_st_imag[15] (
	.clk(clk),
	.d(\butterfly_st_imag[15]~50_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[15]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[15] .is_wysiwyg = "true";
defparam \butterfly_st_imag[15] .power_up = "low";

dffeas \butterfly_st_imag[16] (
	.clk(clk),
	.d(\butterfly_st_imag[16]~52_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_imag[16]~q ),
	.prn(vcc));
defparam \butterfly_st_imag[16] .is_wysiwyg = "true";
defparam \butterfly_st_imag[16] .power_up = "low";

dffeas \butterfly_st_real[2] (
	.clk(clk),
	.d(\butterfly_st_real[2]~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[2]~q ),
	.prn(vcc));
defparam \butterfly_st_real[2] .is_wysiwyg = "true";
defparam \butterfly_st_real[2] .power_up = "low";

dffeas \butterfly_st_real[1] (
	.clk(clk),
	.d(\butterfly_st_real[1]~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[1]~q ),
	.prn(vcc));
defparam \butterfly_st_real[1] .is_wysiwyg = "true";
defparam \butterfly_st_real[1] .power_up = "low";

dffeas \butterfly_st_real[0] (
	.clk(clk),
	.d(\butterfly_st_real[0]~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[0]~q ),
	.prn(vcc));
defparam \butterfly_st_real[0] .is_wysiwyg = "true";
defparam \butterfly_st_real[0] .power_up = "low";

dffeas \butterfly_st_real[17] (
	.clk(clk),
	.d(\butterfly_st_real[17]~54_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[17]~q ),
	.prn(vcc));
defparam \butterfly_st_real[17] .is_wysiwyg = "true";
defparam \butterfly_st_real[17] .power_up = "low";

dffeas \butterfly_st_real[3] (
	.clk(clk),
	.d(\butterfly_st_real[3]~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[3]~q ),
	.prn(vcc));
defparam \butterfly_st_real[3] .is_wysiwyg = "true";
defparam \butterfly_st_real[3] .power_up = "low";

dffeas \butterfly_st_real[4] (
	.clk(clk),
	.d(\butterfly_st_real[4]~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[4]~q ),
	.prn(vcc));
defparam \butterfly_st_real[4] .is_wysiwyg = "true";
defparam \butterfly_st_real[4] .power_up = "low";

dffeas \butterfly_st_real[5] (
	.clk(clk),
	.d(\butterfly_st_real[5]~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[5]~q ),
	.prn(vcc));
defparam \butterfly_st_real[5] .is_wysiwyg = "true";
defparam \butterfly_st_real[5] .power_up = "low";

dffeas \butterfly_st_real[6] (
	.clk(clk),
	.d(\butterfly_st_real[6]~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[6]~q ),
	.prn(vcc));
defparam \butterfly_st_real[6] .is_wysiwyg = "true";
defparam \butterfly_st_real[6] .power_up = "low";

dffeas \butterfly_st_real[7] (
	.clk(clk),
	.d(\butterfly_st_real[7]~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[7]~q ),
	.prn(vcc));
defparam \butterfly_st_real[7] .is_wysiwyg = "true";
defparam \butterfly_st_real[7] .power_up = "low";

dffeas \butterfly_st_real[8] (
	.clk(clk),
	.d(\butterfly_st_real[8]~36_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[8]~q ),
	.prn(vcc));
defparam \butterfly_st_real[8] .is_wysiwyg = "true";
defparam \butterfly_st_real[8] .power_up = "low";

dffeas \butterfly_st_real[9] (
	.clk(clk),
	.d(\butterfly_st_real[9]~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[9]~q ),
	.prn(vcc));
defparam \butterfly_st_real[9] .is_wysiwyg = "true";
defparam \butterfly_st_real[9] .power_up = "low";

dffeas \butterfly_st_real[10] (
	.clk(clk),
	.d(\butterfly_st_real[10]~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[10]~q ),
	.prn(vcc));
defparam \butterfly_st_real[10] .is_wysiwyg = "true";
defparam \butterfly_st_real[10] .power_up = "low";

dffeas \butterfly_st_real[11] (
	.clk(clk),
	.d(\butterfly_st_real[11]~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[11]~q ),
	.prn(vcc));
defparam \butterfly_st_real[11] .is_wysiwyg = "true";
defparam \butterfly_st_real[11] .power_up = "low";

dffeas \butterfly_st_real[12] (
	.clk(clk),
	.d(\butterfly_st_real[12]~44_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[12]~q ),
	.prn(vcc));
defparam \butterfly_st_real[12] .is_wysiwyg = "true";
defparam \butterfly_st_real[12] .power_up = "low";

dffeas \butterfly_st_real[13] (
	.clk(clk),
	.d(\butterfly_st_real[13]~46_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[13]~q ),
	.prn(vcc));
defparam \butterfly_st_real[13] .is_wysiwyg = "true";
defparam \butterfly_st_real[13] .power_up = "low";

dffeas \butterfly_st_real[14] (
	.clk(clk),
	.d(\butterfly_st_real[14]~48_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[14]~q ),
	.prn(vcc));
defparam \butterfly_st_real[14] .is_wysiwyg = "true";
defparam \butterfly_st_real[14] .power_up = "low";

dffeas \butterfly_st_real[15] (
	.clk(clk),
	.d(\butterfly_st_real[15]~50_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[15]~q ),
	.prn(vcc));
defparam \butterfly_st_real[15] .is_wysiwyg = "true";
defparam \butterfly_st_real[15] .power_up = "low";

dffeas \butterfly_st_real[16] (
	.clk(clk),
	.d(\butterfly_st_real[16]~52_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st_real[16]~q ),
	.prn(vcc));
defparam \butterfly_st_real[16] .is_wysiwyg = "true";
defparam \butterfly_st_real[16] .power_up = "low";

dffeas \result_x2_x4_imag[2] (
	.clk(clk),
	.d(\result_x2_x4_imag[2]~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_imag[2]~q ),
	.prn(vcc));
defparam \result_x2_x4_imag[2] .is_wysiwyg = "true";
defparam \result_x2_x4_imag[2] .power_up = "low";

dffeas \result_x1_x3_imag[2] (
	.clk(clk),
	.d(\result_x1_x3_imag[2]~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_imag[2]~q ),
	.prn(vcc));
defparam \result_x1_x3_imag[2] .is_wysiwyg = "true";
defparam \result_x1_x3_imag[2] .power_up = "low";

dffeas \result_x2_x4_imag[1] (
	.clk(clk),
	.d(\result_x2_x4_imag[1]~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_imag[1]~q ),
	.prn(vcc));
defparam \result_x2_x4_imag[1] .is_wysiwyg = "true";
defparam \result_x2_x4_imag[1] .power_up = "low";

dffeas \result_x1_x3_imag[1] (
	.clk(clk),
	.d(\result_x1_x3_imag[1]~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_imag[1]~q ),
	.prn(vcc));
defparam \result_x1_x3_imag[1] .is_wysiwyg = "true";
defparam \result_x1_x3_imag[1] .power_up = "low";

dffeas \result_x2_x4_imag[0] (
	.clk(clk),
	.d(\result_x2_x4_imag[0]~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_imag[0]~q ),
	.prn(vcc));
defparam \result_x2_x4_imag[0] .is_wysiwyg = "true";
defparam \result_x2_x4_imag[0] .power_up = "low";

dffeas \result_x1_x3_imag[0] (
	.clk(clk),
	.d(\result_x1_x3_imag[0]~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_imag[0]~q ),
	.prn(vcc));
defparam \result_x1_x3_imag[0] .is_wysiwyg = "true";
defparam \result_x1_x3_imag[0] .power_up = "low";

cycloneive_lcell_comb \butterfly_st_imag[0]~19 (
	.dataa(\si[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\butterfly_st_imag[0]~19_cout ));
defparam \butterfly_st_imag[0]~19 .lut_mask = 16'h0055;
defparam \butterfly_st_imag[0]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st_imag[0]~20 (
	.dataa(\Add10~3_combout ),
	.datab(\result_x1_x3_imag[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_imag[0]~19_cout ),
	.combout(\butterfly_st_imag[0]~20_combout ),
	.cout(\butterfly_st_imag[0]~21 ));
defparam \butterfly_st_imag[0]~20 .lut_mask = 16'h96BF;
defparam \butterfly_st_imag[0]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_imag[1]~22 (
	.dataa(\Add10~2_combout ),
	.datab(\result_x1_x3_imag[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_imag[0]~21 ),
	.combout(\butterfly_st_imag[1]~22_combout ),
	.cout(\butterfly_st_imag[1]~23 ));
defparam \butterfly_st_imag[1]~22 .lut_mask = 16'h96DF;
defparam \butterfly_st_imag[1]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_imag[2]~24 (
	.dataa(\Add10~1_combout ),
	.datab(\result_x1_x3_imag[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_imag[1]~23 ),
	.combout(\butterfly_st_imag[2]~24_combout ),
	.cout(\butterfly_st_imag[2]~25 ));
defparam \butterfly_st_imag[2]~24 .lut_mask = 16'h96BF;
defparam \butterfly_st_imag[2]~24 .sum_lutc_input = "cin";

dffeas \result_x2_x4_imag[16] (
	.clk(clk),
	.d(\result_x2_x4_imag[16]~51_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_imag[16]~q ),
	.prn(vcc));
defparam \result_x2_x4_imag[16] .is_wysiwyg = "true";
defparam \result_x2_x4_imag[16] .power_up = "low";

dffeas \result_x1_x3_imag[16] (
	.clk(clk),
	.d(\result_x1_x3_imag[16]~51_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_imag[16]~q ),
	.prn(vcc));
defparam \result_x1_x3_imag[16] .is_wysiwyg = "true";
defparam \result_x1_x3_imag[16] .power_up = "low";

dffeas \result_x2_x4_imag[15] (
	.clk(clk),
	.d(\result_x2_x4_imag[15]~49_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_imag[15]~q ),
	.prn(vcc));
defparam \result_x2_x4_imag[15] .is_wysiwyg = "true";
defparam \result_x2_x4_imag[15] .power_up = "low";

dffeas \result_x1_x3_imag[15] (
	.clk(clk),
	.d(\result_x1_x3_imag[15]~49_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_imag[15]~q ),
	.prn(vcc));
defparam \result_x1_x3_imag[15] .is_wysiwyg = "true";
defparam \result_x1_x3_imag[15] .power_up = "low";

dffeas \result_x2_x4_imag[14] (
	.clk(clk),
	.d(\result_x2_x4_imag[14]~47_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_imag[14]~q ),
	.prn(vcc));
defparam \result_x2_x4_imag[14] .is_wysiwyg = "true";
defparam \result_x2_x4_imag[14] .power_up = "low";

dffeas \result_x1_x3_imag[14] (
	.clk(clk),
	.d(\result_x1_x3_imag[14]~47_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_imag[14]~q ),
	.prn(vcc));
defparam \result_x1_x3_imag[14] .is_wysiwyg = "true";
defparam \result_x1_x3_imag[14] .power_up = "low";

dffeas \result_x2_x4_imag[13] (
	.clk(clk),
	.d(\result_x2_x4_imag[13]~45_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_imag[13]~q ),
	.prn(vcc));
defparam \result_x2_x4_imag[13] .is_wysiwyg = "true";
defparam \result_x2_x4_imag[13] .power_up = "low";

dffeas \result_x1_x3_imag[13] (
	.clk(clk),
	.d(\result_x1_x3_imag[13]~45_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_imag[13]~q ),
	.prn(vcc));
defparam \result_x1_x3_imag[13] .is_wysiwyg = "true";
defparam \result_x1_x3_imag[13] .power_up = "low";

dffeas \result_x2_x4_imag[12] (
	.clk(clk),
	.d(\result_x2_x4_imag[12]~43_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_imag[12]~q ),
	.prn(vcc));
defparam \result_x2_x4_imag[12] .is_wysiwyg = "true";
defparam \result_x2_x4_imag[12] .power_up = "low";

dffeas \result_x1_x3_imag[12] (
	.clk(clk),
	.d(\result_x1_x3_imag[12]~43_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_imag[12]~q ),
	.prn(vcc));
defparam \result_x1_x3_imag[12] .is_wysiwyg = "true";
defparam \result_x1_x3_imag[12] .power_up = "low";

dffeas \result_x2_x4_imag[11] (
	.clk(clk),
	.d(\result_x2_x4_imag[11]~41_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_imag[11]~q ),
	.prn(vcc));
defparam \result_x2_x4_imag[11] .is_wysiwyg = "true";
defparam \result_x2_x4_imag[11] .power_up = "low";

dffeas \result_x1_x3_imag[11] (
	.clk(clk),
	.d(\result_x1_x3_imag[11]~41_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_imag[11]~q ),
	.prn(vcc));
defparam \result_x1_x3_imag[11] .is_wysiwyg = "true";
defparam \result_x1_x3_imag[11] .power_up = "low";

dffeas \result_x2_x4_imag[10] (
	.clk(clk),
	.d(\result_x2_x4_imag[10]~39_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_imag[10]~q ),
	.prn(vcc));
defparam \result_x2_x4_imag[10] .is_wysiwyg = "true";
defparam \result_x2_x4_imag[10] .power_up = "low";

dffeas \result_x1_x3_imag[10] (
	.clk(clk),
	.d(\result_x1_x3_imag[10]~39_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_imag[10]~q ),
	.prn(vcc));
defparam \result_x1_x3_imag[10] .is_wysiwyg = "true";
defparam \result_x1_x3_imag[10] .power_up = "low";

dffeas \result_x2_x4_imag[9] (
	.clk(clk),
	.d(\result_x2_x4_imag[9]~37_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_imag[9]~q ),
	.prn(vcc));
defparam \result_x2_x4_imag[9] .is_wysiwyg = "true";
defparam \result_x2_x4_imag[9] .power_up = "low";

dffeas \result_x1_x3_imag[9] (
	.clk(clk),
	.d(\result_x1_x3_imag[9]~37_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_imag[9]~q ),
	.prn(vcc));
defparam \result_x1_x3_imag[9] .is_wysiwyg = "true";
defparam \result_x1_x3_imag[9] .power_up = "low";

dffeas \result_x2_x4_imag[8] (
	.clk(clk),
	.d(\result_x2_x4_imag[8]~35_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_imag[8]~q ),
	.prn(vcc));
defparam \result_x2_x4_imag[8] .is_wysiwyg = "true";
defparam \result_x2_x4_imag[8] .power_up = "low";

dffeas \result_x1_x3_imag[8] (
	.clk(clk),
	.d(\result_x1_x3_imag[8]~35_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_imag[8]~q ),
	.prn(vcc));
defparam \result_x1_x3_imag[8] .is_wysiwyg = "true";
defparam \result_x1_x3_imag[8] .power_up = "low";

dffeas \result_x2_x4_imag[7] (
	.clk(clk),
	.d(\result_x2_x4_imag[7]~33_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_imag[7]~q ),
	.prn(vcc));
defparam \result_x2_x4_imag[7] .is_wysiwyg = "true";
defparam \result_x2_x4_imag[7] .power_up = "low";

dffeas \result_x1_x3_imag[7] (
	.clk(clk),
	.d(\result_x1_x3_imag[7]~33_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_imag[7]~q ),
	.prn(vcc));
defparam \result_x1_x3_imag[7] .is_wysiwyg = "true";
defparam \result_x1_x3_imag[7] .power_up = "low";

dffeas \result_x2_x4_imag[6] (
	.clk(clk),
	.d(\result_x2_x4_imag[6]~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_imag[6]~q ),
	.prn(vcc));
defparam \result_x2_x4_imag[6] .is_wysiwyg = "true";
defparam \result_x2_x4_imag[6] .power_up = "low";

dffeas \result_x1_x3_imag[6] (
	.clk(clk),
	.d(\result_x1_x3_imag[6]~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_imag[6]~q ),
	.prn(vcc));
defparam \result_x1_x3_imag[6] .is_wysiwyg = "true";
defparam \result_x1_x3_imag[6] .power_up = "low";

dffeas \result_x2_x4_imag[5] (
	.clk(clk),
	.d(\result_x2_x4_imag[5]~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_imag[5]~q ),
	.prn(vcc));
defparam \result_x2_x4_imag[5] .is_wysiwyg = "true";
defparam \result_x2_x4_imag[5] .power_up = "low";

dffeas \result_x1_x3_imag[5] (
	.clk(clk),
	.d(\result_x1_x3_imag[5]~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_imag[5]~q ),
	.prn(vcc));
defparam \result_x1_x3_imag[5] .is_wysiwyg = "true";
defparam \result_x1_x3_imag[5] .power_up = "low";

dffeas \result_x2_x4_imag[4] (
	.clk(clk),
	.d(\result_x2_x4_imag[4]~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_imag[4]~q ),
	.prn(vcc));
defparam \result_x2_x4_imag[4] .is_wysiwyg = "true";
defparam \result_x2_x4_imag[4] .power_up = "low";

dffeas \result_x1_x3_imag[4] (
	.clk(clk),
	.d(\result_x1_x3_imag[4]~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_imag[4]~q ),
	.prn(vcc));
defparam \result_x1_x3_imag[4] .is_wysiwyg = "true";
defparam \result_x1_x3_imag[4] .power_up = "low";

dffeas \result_x2_x4_imag[3] (
	.clk(clk),
	.d(\result_x2_x4_imag[3]~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_imag[3]~q ),
	.prn(vcc));
defparam \result_x2_x4_imag[3] .is_wysiwyg = "true";
defparam \result_x2_x4_imag[3] .power_up = "low";

dffeas \result_x1_x3_imag[3] (
	.clk(clk),
	.d(\result_x1_x3_imag[3]~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_imag[3]~q ),
	.prn(vcc));
defparam \result_x1_x3_imag[3] .is_wysiwyg = "true";
defparam \result_x1_x3_imag[3] .power_up = "low";

cycloneive_lcell_comb \butterfly_st_imag[3]~26 (
	.dataa(\Add10~17_combout ),
	.datab(\result_x1_x3_imag[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_imag[2]~25 ),
	.combout(\butterfly_st_imag[3]~26_combout ),
	.cout(\butterfly_st_imag[3]~27 ));
defparam \butterfly_st_imag[3]~26 .lut_mask = 16'h96DF;
defparam \butterfly_st_imag[3]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_imag[4]~28 (
	.dataa(\Add10~16_combout ),
	.datab(\result_x1_x3_imag[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_imag[3]~27 ),
	.combout(\butterfly_st_imag[4]~28_combout ),
	.cout(\butterfly_st_imag[4]~29 ));
defparam \butterfly_st_imag[4]~28 .lut_mask = 16'h96BF;
defparam \butterfly_st_imag[4]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_imag[5]~30 (
	.dataa(\Add10~15_combout ),
	.datab(\result_x1_x3_imag[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_imag[4]~29 ),
	.combout(\butterfly_st_imag[5]~30_combout ),
	.cout(\butterfly_st_imag[5]~31 ));
defparam \butterfly_st_imag[5]~30 .lut_mask = 16'h96DF;
defparam \butterfly_st_imag[5]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_imag[6]~32 (
	.dataa(\Add10~14_combout ),
	.datab(\result_x1_x3_imag[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_imag[5]~31 ),
	.combout(\butterfly_st_imag[6]~32_combout ),
	.cout(\butterfly_st_imag[6]~33 ));
defparam \butterfly_st_imag[6]~32 .lut_mask = 16'h96BF;
defparam \butterfly_st_imag[6]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_imag[7]~34 (
	.dataa(\Add10~13_combout ),
	.datab(\result_x1_x3_imag[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_imag[6]~33 ),
	.combout(\butterfly_st_imag[7]~34_combout ),
	.cout(\butterfly_st_imag[7]~35 ));
defparam \butterfly_st_imag[7]~34 .lut_mask = 16'h96DF;
defparam \butterfly_st_imag[7]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_imag[8]~36 (
	.dataa(\Add10~12_combout ),
	.datab(\result_x1_x3_imag[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_imag[7]~35 ),
	.combout(\butterfly_st_imag[8]~36_combout ),
	.cout(\butterfly_st_imag[8]~37 ));
defparam \butterfly_st_imag[8]~36 .lut_mask = 16'h96BF;
defparam \butterfly_st_imag[8]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_imag[9]~38 (
	.dataa(\Add10~11_combout ),
	.datab(\result_x1_x3_imag[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_imag[8]~37 ),
	.combout(\butterfly_st_imag[9]~38_combout ),
	.cout(\butterfly_st_imag[9]~39 ));
defparam \butterfly_st_imag[9]~38 .lut_mask = 16'h96DF;
defparam \butterfly_st_imag[9]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_imag[10]~40 (
	.dataa(\Add10~10_combout ),
	.datab(\result_x1_x3_imag[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_imag[9]~39 ),
	.combout(\butterfly_st_imag[10]~40_combout ),
	.cout(\butterfly_st_imag[10]~41 ));
defparam \butterfly_st_imag[10]~40 .lut_mask = 16'h96BF;
defparam \butterfly_st_imag[10]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_imag[11]~42 (
	.dataa(\Add10~9_combout ),
	.datab(\result_x1_x3_imag[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_imag[10]~41 ),
	.combout(\butterfly_st_imag[11]~42_combout ),
	.cout(\butterfly_st_imag[11]~43 ));
defparam \butterfly_st_imag[11]~42 .lut_mask = 16'h96DF;
defparam \butterfly_st_imag[11]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_imag[12]~44 (
	.dataa(\Add10~8_combout ),
	.datab(\result_x1_x3_imag[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_imag[11]~43 ),
	.combout(\butterfly_st_imag[12]~44_combout ),
	.cout(\butterfly_st_imag[12]~45 ));
defparam \butterfly_st_imag[12]~44 .lut_mask = 16'h96BF;
defparam \butterfly_st_imag[12]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_imag[13]~46 (
	.dataa(\Add10~7_combout ),
	.datab(\result_x1_x3_imag[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_imag[12]~45 ),
	.combout(\butterfly_st_imag[13]~46_combout ),
	.cout(\butterfly_st_imag[13]~47 ));
defparam \butterfly_st_imag[13]~46 .lut_mask = 16'h96DF;
defparam \butterfly_st_imag[13]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_imag[14]~48 (
	.dataa(\Add10~6_combout ),
	.datab(\result_x1_x3_imag[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_imag[13]~47 ),
	.combout(\butterfly_st_imag[14]~48_combout ),
	.cout(\butterfly_st_imag[14]~49 ));
defparam \butterfly_st_imag[14]~48 .lut_mask = 16'h96BF;
defparam \butterfly_st_imag[14]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_imag[15]~50 (
	.dataa(\Add10~5_combout ),
	.datab(\result_x1_x3_imag[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_imag[14]~49 ),
	.combout(\butterfly_st_imag[15]~50_combout ),
	.cout(\butterfly_st_imag[15]~51 ));
defparam \butterfly_st_imag[15]~50 .lut_mask = 16'h96DF;
defparam \butterfly_st_imag[15]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_imag[16]~52 (
	.dataa(\Add10~4_combout ),
	.datab(\result_x1_x3_imag[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_imag[15]~51 ),
	.combout(\butterfly_st_imag[16]~52_combout ),
	.cout(\butterfly_st_imag[16]~53 ));
defparam \butterfly_st_imag[16]~52 .lut_mask = 16'h96BF;
defparam \butterfly_st_imag[16]~52 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_imag[17]~54 (
	.dataa(\Add10~4_combout ),
	.datab(\result_x1_x3_imag[16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st_imag[16]~53 ),
	.combout(\butterfly_st_imag[17]~54_combout ),
	.cout());
defparam \butterfly_st_imag[17]~54 .lut_mask = 16'h9696;
defparam \butterfly_st_imag[17]~54 .sum_lutc_input = "cin";

dffeas \sr[0] (
	.clk(clk),
	.d(\Mux264~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sr[0]~q ),
	.prn(vcc));
defparam \sr[0] .is_wysiwyg = "true";
defparam \sr[0] .power_up = "low";

dffeas \result_x2_x4_real[2] (
	.clk(clk),
	.d(\result_x2_x4_real[2]~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_real[2]~q ),
	.prn(vcc));
defparam \result_x2_x4_real[2] .is_wysiwyg = "true";
defparam \result_x2_x4_real[2] .power_up = "low";

dffeas \result_x1_x3_real[2] (
	.clk(clk),
	.d(\result_x1_x3_real[2]~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_real[2]~q ),
	.prn(vcc));
defparam \result_x1_x3_real[2] .is_wysiwyg = "true";
defparam \result_x1_x3_real[2] .power_up = "low";

dffeas \result_x2_x4_real[1] (
	.clk(clk),
	.d(\result_x2_x4_real[1]~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_real[1]~q ),
	.prn(vcc));
defparam \result_x2_x4_real[1] .is_wysiwyg = "true";
defparam \result_x2_x4_real[1] .power_up = "low";

dffeas \result_x1_x3_real[1] (
	.clk(clk),
	.d(\result_x1_x3_real[1]~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_real[1]~q ),
	.prn(vcc));
defparam \result_x1_x3_real[1] .is_wysiwyg = "true";
defparam \result_x1_x3_real[1] .power_up = "low";

dffeas \result_x2_x4_real[0] (
	.clk(clk),
	.d(\result_x2_x4_real[0]~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_real[0]~q ),
	.prn(vcc));
defparam \result_x2_x4_real[0] .is_wysiwyg = "true";
defparam \result_x2_x4_real[0] .power_up = "low";

dffeas \result_x1_x3_real[0] (
	.clk(clk),
	.d(\result_x1_x3_real[0]~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_real[0]~q ),
	.prn(vcc));
defparam \result_x1_x3_real[0] .is_wysiwyg = "true";
defparam \result_x1_x3_real[0] .power_up = "low";

cycloneive_lcell_comb \butterfly_st_real[0]~19 (
	.dataa(\sr[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\butterfly_st_real[0]~19_cout ));
defparam \butterfly_st_real[0]~19 .lut_mask = 16'h0055;
defparam \butterfly_st_real[0]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st_real[0]~20 (
	.dataa(\Add4~3_combout ),
	.datab(\result_x1_x3_real[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_real[0]~19_cout ),
	.combout(\butterfly_st_real[0]~20_combout ),
	.cout(\butterfly_st_real[0]~21 ));
defparam \butterfly_st_real[0]~20 .lut_mask = 16'h96BF;
defparam \butterfly_st_real[0]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_real[1]~22 (
	.dataa(\Add4~2_combout ),
	.datab(\result_x1_x3_real[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_real[0]~21 ),
	.combout(\butterfly_st_real[1]~22_combout ),
	.cout(\butterfly_st_real[1]~23 ));
defparam \butterfly_st_real[1]~22 .lut_mask = 16'h96DF;
defparam \butterfly_st_real[1]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_real[2]~24 (
	.dataa(\Add4~1_combout ),
	.datab(\result_x1_x3_real[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_real[1]~23 ),
	.combout(\butterfly_st_real[2]~24_combout ),
	.cout(\butterfly_st_real[2]~25 ));
defparam \butterfly_st_real[2]~24 .lut_mask = 16'h96BF;
defparam \butterfly_st_real[2]~24 .sum_lutc_input = "cin";

dffeas \result_x2_x4_real[16] (
	.clk(clk),
	.d(\result_x2_x4_real[16]~51_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_real[16]~q ),
	.prn(vcc));
defparam \result_x2_x4_real[16] .is_wysiwyg = "true";
defparam \result_x2_x4_real[16] .power_up = "low";

dffeas \result_x1_x3_real[16] (
	.clk(clk),
	.d(\result_x1_x3_real[16]~51_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_real[16]~q ),
	.prn(vcc));
defparam \result_x1_x3_real[16] .is_wysiwyg = "true";
defparam \result_x1_x3_real[16] .power_up = "low";

dffeas \result_x2_x4_real[15] (
	.clk(clk),
	.d(\result_x2_x4_real[15]~49_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_real[15]~q ),
	.prn(vcc));
defparam \result_x2_x4_real[15] .is_wysiwyg = "true";
defparam \result_x2_x4_real[15] .power_up = "low";

dffeas \result_x1_x3_real[15] (
	.clk(clk),
	.d(\result_x1_x3_real[15]~49_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_real[15]~q ),
	.prn(vcc));
defparam \result_x1_x3_real[15] .is_wysiwyg = "true";
defparam \result_x1_x3_real[15] .power_up = "low";

dffeas \result_x2_x4_real[14] (
	.clk(clk),
	.d(\result_x2_x4_real[14]~47_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_real[14]~q ),
	.prn(vcc));
defparam \result_x2_x4_real[14] .is_wysiwyg = "true";
defparam \result_x2_x4_real[14] .power_up = "low";

dffeas \result_x1_x3_real[14] (
	.clk(clk),
	.d(\result_x1_x3_real[14]~47_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_real[14]~q ),
	.prn(vcc));
defparam \result_x1_x3_real[14] .is_wysiwyg = "true";
defparam \result_x1_x3_real[14] .power_up = "low";

dffeas \result_x2_x4_real[13] (
	.clk(clk),
	.d(\result_x2_x4_real[13]~45_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_real[13]~q ),
	.prn(vcc));
defparam \result_x2_x4_real[13] .is_wysiwyg = "true";
defparam \result_x2_x4_real[13] .power_up = "low";

dffeas \result_x1_x3_real[13] (
	.clk(clk),
	.d(\result_x1_x3_real[13]~45_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_real[13]~q ),
	.prn(vcc));
defparam \result_x1_x3_real[13] .is_wysiwyg = "true";
defparam \result_x1_x3_real[13] .power_up = "low";

dffeas \result_x2_x4_real[12] (
	.clk(clk),
	.d(\result_x2_x4_real[12]~43_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_real[12]~q ),
	.prn(vcc));
defparam \result_x2_x4_real[12] .is_wysiwyg = "true";
defparam \result_x2_x4_real[12] .power_up = "low";

dffeas \result_x1_x3_real[12] (
	.clk(clk),
	.d(\result_x1_x3_real[12]~43_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_real[12]~q ),
	.prn(vcc));
defparam \result_x1_x3_real[12] .is_wysiwyg = "true";
defparam \result_x1_x3_real[12] .power_up = "low";

dffeas \result_x2_x4_real[11] (
	.clk(clk),
	.d(\result_x2_x4_real[11]~41_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_real[11]~q ),
	.prn(vcc));
defparam \result_x2_x4_real[11] .is_wysiwyg = "true";
defparam \result_x2_x4_real[11] .power_up = "low";

dffeas \result_x1_x3_real[11] (
	.clk(clk),
	.d(\result_x1_x3_real[11]~41_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_real[11]~q ),
	.prn(vcc));
defparam \result_x1_x3_real[11] .is_wysiwyg = "true";
defparam \result_x1_x3_real[11] .power_up = "low";

dffeas \result_x2_x4_real[10] (
	.clk(clk),
	.d(\result_x2_x4_real[10]~39_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_real[10]~q ),
	.prn(vcc));
defparam \result_x2_x4_real[10] .is_wysiwyg = "true";
defparam \result_x2_x4_real[10] .power_up = "low";

dffeas \result_x1_x3_real[10] (
	.clk(clk),
	.d(\result_x1_x3_real[10]~39_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_real[10]~q ),
	.prn(vcc));
defparam \result_x1_x3_real[10] .is_wysiwyg = "true";
defparam \result_x1_x3_real[10] .power_up = "low";

dffeas \result_x2_x4_real[9] (
	.clk(clk),
	.d(\result_x2_x4_real[9]~37_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_real[9]~q ),
	.prn(vcc));
defparam \result_x2_x4_real[9] .is_wysiwyg = "true";
defparam \result_x2_x4_real[9] .power_up = "low";

dffeas \result_x1_x3_real[9] (
	.clk(clk),
	.d(\result_x1_x3_real[9]~37_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_real[9]~q ),
	.prn(vcc));
defparam \result_x1_x3_real[9] .is_wysiwyg = "true";
defparam \result_x1_x3_real[9] .power_up = "low";

dffeas \result_x2_x4_real[8] (
	.clk(clk),
	.d(\result_x2_x4_real[8]~35_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_real[8]~q ),
	.prn(vcc));
defparam \result_x2_x4_real[8] .is_wysiwyg = "true";
defparam \result_x2_x4_real[8] .power_up = "low";

dffeas \result_x1_x3_real[8] (
	.clk(clk),
	.d(\result_x1_x3_real[8]~35_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_real[8]~q ),
	.prn(vcc));
defparam \result_x1_x3_real[8] .is_wysiwyg = "true";
defparam \result_x1_x3_real[8] .power_up = "low";

dffeas \result_x2_x4_real[7] (
	.clk(clk),
	.d(\result_x2_x4_real[7]~33_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_real[7]~q ),
	.prn(vcc));
defparam \result_x2_x4_real[7] .is_wysiwyg = "true";
defparam \result_x2_x4_real[7] .power_up = "low";

dffeas \result_x1_x3_real[7] (
	.clk(clk),
	.d(\result_x1_x3_real[7]~33_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_real[7]~q ),
	.prn(vcc));
defparam \result_x1_x3_real[7] .is_wysiwyg = "true";
defparam \result_x1_x3_real[7] .power_up = "low";

dffeas \result_x2_x4_real[6] (
	.clk(clk),
	.d(\result_x2_x4_real[6]~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_real[6]~q ),
	.prn(vcc));
defparam \result_x2_x4_real[6] .is_wysiwyg = "true";
defparam \result_x2_x4_real[6] .power_up = "low";

dffeas \result_x1_x3_real[6] (
	.clk(clk),
	.d(\result_x1_x3_real[6]~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_real[6]~q ),
	.prn(vcc));
defparam \result_x1_x3_real[6] .is_wysiwyg = "true";
defparam \result_x1_x3_real[6] .power_up = "low";

dffeas \result_x2_x4_real[5] (
	.clk(clk),
	.d(\result_x2_x4_real[5]~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_real[5]~q ),
	.prn(vcc));
defparam \result_x2_x4_real[5] .is_wysiwyg = "true";
defparam \result_x2_x4_real[5] .power_up = "low";

dffeas \result_x1_x3_real[5] (
	.clk(clk),
	.d(\result_x1_x3_real[5]~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_real[5]~q ),
	.prn(vcc));
defparam \result_x1_x3_real[5] .is_wysiwyg = "true";
defparam \result_x1_x3_real[5] .power_up = "low";

dffeas \result_x2_x4_real[4] (
	.clk(clk),
	.d(\result_x2_x4_real[4]~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_real[4]~q ),
	.prn(vcc));
defparam \result_x2_x4_real[4] .is_wysiwyg = "true";
defparam \result_x2_x4_real[4] .power_up = "low";

dffeas \result_x1_x3_real[4] (
	.clk(clk),
	.d(\result_x1_x3_real[4]~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_real[4]~q ),
	.prn(vcc));
defparam \result_x1_x3_real[4] .is_wysiwyg = "true";
defparam \result_x1_x3_real[4] .power_up = "low";

dffeas \result_x2_x4_real[3] (
	.clk(clk),
	.d(\result_x2_x4_real[3]~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x2_x4_real[3]~q ),
	.prn(vcc));
defparam \result_x2_x4_real[3] .is_wysiwyg = "true";
defparam \result_x2_x4_real[3] .power_up = "low";

dffeas \result_x1_x3_real[3] (
	.clk(clk),
	.d(\result_x1_x3_real[3]~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_x1_x3_real[3]~q ),
	.prn(vcc));
defparam \result_x1_x3_real[3] .is_wysiwyg = "true";
defparam \result_x1_x3_real[3] .power_up = "low";

cycloneive_lcell_comb \butterfly_st_real[3]~26 (
	.dataa(\Add4~17_combout ),
	.datab(\result_x1_x3_real[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_real[2]~25 ),
	.combout(\butterfly_st_real[3]~26_combout ),
	.cout(\butterfly_st_real[3]~27 ));
defparam \butterfly_st_real[3]~26 .lut_mask = 16'h96DF;
defparam \butterfly_st_real[3]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_real[4]~28 (
	.dataa(\Add4~16_combout ),
	.datab(\result_x1_x3_real[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_real[3]~27 ),
	.combout(\butterfly_st_real[4]~28_combout ),
	.cout(\butterfly_st_real[4]~29 ));
defparam \butterfly_st_real[4]~28 .lut_mask = 16'h96BF;
defparam \butterfly_st_real[4]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_real[5]~30 (
	.dataa(\Add4~15_combout ),
	.datab(\result_x1_x3_real[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_real[4]~29 ),
	.combout(\butterfly_st_real[5]~30_combout ),
	.cout(\butterfly_st_real[5]~31 ));
defparam \butterfly_st_real[5]~30 .lut_mask = 16'h96DF;
defparam \butterfly_st_real[5]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_real[6]~32 (
	.dataa(\Add4~14_combout ),
	.datab(\result_x1_x3_real[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_real[5]~31 ),
	.combout(\butterfly_st_real[6]~32_combout ),
	.cout(\butterfly_st_real[6]~33 ));
defparam \butterfly_st_real[6]~32 .lut_mask = 16'h96BF;
defparam \butterfly_st_real[6]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_real[7]~34 (
	.dataa(\Add4~13_combout ),
	.datab(\result_x1_x3_real[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_real[6]~33 ),
	.combout(\butterfly_st_real[7]~34_combout ),
	.cout(\butterfly_st_real[7]~35 ));
defparam \butterfly_st_real[7]~34 .lut_mask = 16'h96DF;
defparam \butterfly_st_real[7]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_real[8]~36 (
	.dataa(\Add4~12_combout ),
	.datab(\result_x1_x3_real[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_real[7]~35 ),
	.combout(\butterfly_st_real[8]~36_combout ),
	.cout(\butterfly_st_real[8]~37 ));
defparam \butterfly_st_real[8]~36 .lut_mask = 16'h96BF;
defparam \butterfly_st_real[8]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_real[9]~38 (
	.dataa(\Add4~11_combout ),
	.datab(\result_x1_x3_real[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_real[8]~37 ),
	.combout(\butterfly_st_real[9]~38_combout ),
	.cout(\butterfly_st_real[9]~39 ));
defparam \butterfly_st_real[9]~38 .lut_mask = 16'h96DF;
defparam \butterfly_st_real[9]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_real[10]~40 (
	.dataa(\Add4~10_combout ),
	.datab(\result_x1_x3_real[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_real[9]~39 ),
	.combout(\butterfly_st_real[10]~40_combout ),
	.cout(\butterfly_st_real[10]~41 ));
defparam \butterfly_st_real[10]~40 .lut_mask = 16'h96BF;
defparam \butterfly_st_real[10]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_real[11]~42 (
	.dataa(\Add4~9_combout ),
	.datab(\result_x1_x3_real[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_real[10]~41 ),
	.combout(\butterfly_st_real[11]~42_combout ),
	.cout(\butterfly_st_real[11]~43 ));
defparam \butterfly_st_real[11]~42 .lut_mask = 16'h96DF;
defparam \butterfly_st_real[11]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_real[12]~44 (
	.dataa(\Add4~8_combout ),
	.datab(\result_x1_x3_real[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_real[11]~43 ),
	.combout(\butterfly_st_real[12]~44_combout ),
	.cout(\butterfly_st_real[12]~45 ));
defparam \butterfly_st_real[12]~44 .lut_mask = 16'h96BF;
defparam \butterfly_st_real[12]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_real[13]~46 (
	.dataa(\Add4~7_combout ),
	.datab(\result_x1_x3_real[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_real[12]~45 ),
	.combout(\butterfly_st_real[13]~46_combout ),
	.cout(\butterfly_st_real[13]~47 ));
defparam \butterfly_st_real[13]~46 .lut_mask = 16'h96DF;
defparam \butterfly_st_real[13]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_real[14]~48 (
	.dataa(\Add4~6_combout ),
	.datab(\result_x1_x3_real[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_real[13]~47 ),
	.combout(\butterfly_st_real[14]~48_combout ),
	.cout(\butterfly_st_real[14]~49 ));
defparam \butterfly_st_real[14]~48 .lut_mask = 16'h96BF;
defparam \butterfly_st_real[14]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_real[15]~50 (
	.dataa(\Add4~5_combout ),
	.datab(\result_x1_x3_real[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_real[14]~49 ),
	.combout(\butterfly_st_real[15]~50_combout ),
	.cout(\butterfly_st_real[15]~51 ));
defparam \butterfly_st_real[15]~50 .lut_mask = 16'h96DF;
defparam \butterfly_st_real[15]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_real[16]~52 (
	.dataa(\Add4~4_combout ),
	.datab(\result_x1_x3_real[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st_real[15]~51 ),
	.combout(\butterfly_st_real[16]~52_combout ),
	.cout(\butterfly_st_real[16]~53 ));
defparam \butterfly_st_real[16]~52 .lut_mask = 16'h96BF;
defparam \butterfly_st_real[16]~52 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st_real[17]~54 (
	.dataa(\Add4~4_combout ),
	.datab(\result_x1_x3_real[16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st_real[16]~53 ),
	.combout(\butterfly_st_real[17]~54_combout ),
	.cout());
defparam \butterfly_st_real[17]~54 .lut_mask = 16'h9696;
defparam \butterfly_st_real[17]~54 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_imag[0]~18 (
	.dataa(\si[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\result_x2_x4_imag[0]~18_cout ));
defparam \result_x2_x4_imag[0]~18 .lut_mask = 16'h0055;
defparam \result_x2_x4_imag[0]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \result_x2_x4_imag[0]~19 (
	.dataa(\Add8~3_combout ),
	.datab(\x_2_imag_held[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_imag[0]~18_cout ),
	.combout(\result_x2_x4_imag[0]~19_combout ),
	.cout(\result_x2_x4_imag[0]~20 ));
defparam \result_x2_x4_imag[0]~19 .lut_mask = 16'h96BF;
defparam \result_x2_x4_imag[0]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_imag[1]~21 (
	.dataa(\Add8~2_combout ),
	.datab(\x_2_imag_held[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_imag[0]~20 ),
	.combout(\result_x2_x4_imag[1]~21_combout ),
	.cout(\result_x2_x4_imag[1]~22 ));
defparam \result_x2_x4_imag[1]~21 .lut_mask = 16'h96DF;
defparam \result_x2_x4_imag[1]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_imag[2]~23 (
	.dataa(\Add8~1_combout ),
	.datab(\x_2_imag_held[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_imag[1]~22 ),
	.combout(\result_x2_x4_imag[2]~23_combout ),
	.cout(\result_x2_x4_imag[2]~24 ));
defparam \result_x2_x4_imag[2]~23 .lut_mask = 16'h96BF;
defparam \result_x2_x4_imag[2]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_imag[0]~18 (
	.dataa(\si[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\result_x1_x3_imag[0]~18_cout ));
defparam \result_x1_x3_imag[0]~18 .lut_mask = 16'h0055;
defparam \result_x1_x3_imag[0]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \result_x1_x3_imag[0]~19 (
	.dataa(\Add6~3_combout ),
	.datab(\x_1_imag_held[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_imag[0]~18_cout ),
	.combout(\result_x1_x3_imag[0]~19_combout ),
	.cout(\result_x1_x3_imag[0]~20 ));
defparam \result_x1_x3_imag[0]~19 .lut_mask = 16'h96BF;
defparam \result_x1_x3_imag[0]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_imag[1]~21 (
	.dataa(\Add6~2_combout ),
	.datab(\x_1_imag_held[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_imag[0]~20 ),
	.combout(\result_x1_x3_imag[1]~21_combout ),
	.cout(\result_x1_x3_imag[1]~22 ));
defparam \result_x1_x3_imag[1]~21 .lut_mask = 16'h96DF;
defparam \result_x1_x3_imag[1]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_imag[2]~23 (
	.dataa(\Add6~1_combout ),
	.datab(\x_1_imag_held[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_imag[1]~22 ),
	.combout(\result_x1_x3_imag[2]~23_combout ),
	.cout(\result_x1_x3_imag[2]~24 ));
defparam \result_x1_x3_imag[2]~23 .lut_mask = 16'h96BF;
defparam \result_x1_x3_imag[2]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_imag[3]~25 (
	.dataa(\Add8~16_combout ),
	.datab(\x_2_imag_held[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_imag[2]~24 ),
	.combout(\result_x2_x4_imag[3]~25_combout ),
	.cout(\result_x2_x4_imag[3]~26 ));
defparam \result_x2_x4_imag[3]~25 .lut_mask = 16'h96DF;
defparam \result_x2_x4_imag[3]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_imag[4]~27 (
	.dataa(\Add8~15_combout ),
	.datab(\x_2_imag_held[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_imag[3]~26 ),
	.combout(\result_x2_x4_imag[4]~27_combout ),
	.cout(\result_x2_x4_imag[4]~28 ));
defparam \result_x2_x4_imag[4]~27 .lut_mask = 16'h96BF;
defparam \result_x2_x4_imag[4]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_imag[5]~29 (
	.dataa(\Add8~14_combout ),
	.datab(\x_2_imag_held[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_imag[4]~28 ),
	.combout(\result_x2_x4_imag[5]~29_combout ),
	.cout(\result_x2_x4_imag[5]~30 ));
defparam \result_x2_x4_imag[5]~29 .lut_mask = 16'h96DF;
defparam \result_x2_x4_imag[5]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_imag[6]~31 (
	.dataa(\Add8~13_combout ),
	.datab(\x_2_imag_held[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_imag[5]~30 ),
	.combout(\result_x2_x4_imag[6]~31_combout ),
	.cout(\result_x2_x4_imag[6]~32 ));
defparam \result_x2_x4_imag[6]~31 .lut_mask = 16'h96BF;
defparam \result_x2_x4_imag[6]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_imag[7]~33 (
	.dataa(\Add8~12_combout ),
	.datab(\x_2_imag_held[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_imag[6]~32 ),
	.combout(\result_x2_x4_imag[7]~33_combout ),
	.cout(\result_x2_x4_imag[7]~34 ));
defparam \result_x2_x4_imag[7]~33 .lut_mask = 16'h96DF;
defparam \result_x2_x4_imag[7]~33 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_imag[8]~35 (
	.dataa(\Add8~11_combout ),
	.datab(\x_2_imag_held[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_imag[7]~34 ),
	.combout(\result_x2_x4_imag[8]~35_combout ),
	.cout(\result_x2_x4_imag[8]~36 ));
defparam \result_x2_x4_imag[8]~35 .lut_mask = 16'h96BF;
defparam \result_x2_x4_imag[8]~35 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_imag[9]~37 (
	.dataa(\Add8~10_combout ),
	.datab(\x_2_imag_held[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_imag[8]~36 ),
	.combout(\result_x2_x4_imag[9]~37_combout ),
	.cout(\result_x2_x4_imag[9]~38 ));
defparam \result_x2_x4_imag[9]~37 .lut_mask = 16'h96DF;
defparam \result_x2_x4_imag[9]~37 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_imag[10]~39 (
	.dataa(\Add8~9_combout ),
	.datab(\x_2_imag_held[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_imag[9]~38 ),
	.combout(\result_x2_x4_imag[10]~39_combout ),
	.cout(\result_x2_x4_imag[10]~40 ));
defparam \result_x2_x4_imag[10]~39 .lut_mask = 16'h96BF;
defparam \result_x2_x4_imag[10]~39 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_imag[11]~41 (
	.dataa(\Add8~8_combout ),
	.datab(\x_2_imag_held[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_imag[10]~40 ),
	.combout(\result_x2_x4_imag[11]~41_combout ),
	.cout(\result_x2_x4_imag[11]~42 ));
defparam \result_x2_x4_imag[11]~41 .lut_mask = 16'h96DF;
defparam \result_x2_x4_imag[11]~41 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_imag[12]~43 (
	.dataa(\Add8~7_combout ),
	.datab(\x_2_imag_held[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_imag[11]~42 ),
	.combout(\result_x2_x4_imag[12]~43_combout ),
	.cout(\result_x2_x4_imag[12]~44 ));
defparam \result_x2_x4_imag[12]~43 .lut_mask = 16'h96BF;
defparam \result_x2_x4_imag[12]~43 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_imag[13]~45 (
	.dataa(\Add8~6_combout ),
	.datab(\x_2_imag_held[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_imag[12]~44 ),
	.combout(\result_x2_x4_imag[13]~45_combout ),
	.cout(\result_x2_x4_imag[13]~46 ));
defparam \result_x2_x4_imag[13]~45 .lut_mask = 16'h96DF;
defparam \result_x2_x4_imag[13]~45 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_imag[14]~47 (
	.dataa(\Add8~5_combout ),
	.datab(\x_2_imag_held[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_imag[13]~46 ),
	.combout(\result_x2_x4_imag[14]~47_combout ),
	.cout(\result_x2_x4_imag[14]~48 ));
defparam \result_x2_x4_imag[14]~47 .lut_mask = 16'h96BF;
defparam \result_x2_x4_imag[14]~47 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_imag[15]~49 (
	.dataa(\Add8~4_combout ),
	.datab(\x_2_imag_held[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_imag[14]~48 ),
	.combout(\result_x2_x4_imag[15]~49_combout ),
	.cout(\result_x2_x4_imag[15]~50 ));
defparam \result_x2_x4_imag[15]~49 .lut_mask = 16'h96DF;
defparam \result_x2_x4_imag[15]~49 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_imag[16]~51 (
	.dataa(\Add8~4_combout ),
	.datab(\x_2_imag_held[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\result_x2_x4_imag[15]~50 ),
	.combout(\result_x2_x4_imag[16]~51_combout ),
	.cout());
defparam \result_x2_x4_imag[16]~51 .lut_mask = 16'h9696;
defparam \result_x2_x4_imag[16]~51 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_imag[3]~25 (
	.dataa(\Add6~16_combout ),
	.datab(\x_1_imag_held[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_imag[2]~24 ),
	.combout(\result_x1_x3_imag[3]~25_combout ),
	.cout(\result_x1_x3_imag[3]~26 ));
defparam \result_x1_x3_imag[3]~25 .lut_mask = 16'h96DF;
defparam \result_x1_x3_imag[3]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_imag[4]~27 (
	.dataa(\Add6~15_combout ),
	.datab(\x_1_imag_held[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_imag[3]~26 ),
	.combout(\result_x1_x3_imag[4]~27_combout ),
	.cout(\result_x1_x3_imag[4]~28 ));
defparam \result_x1_x3_imag[4]~27 .lut_mask = 16'h96BF;
defparam \result_x1_x3_imag[4]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_imag[5]~29 (
	.dataa(\Add6~14_combout ),
	.datab(\x_1_imag_held[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_imag[4]~28 ),
	.combout(\result_x1_x3_imag[5]~29_combout ),
	.cout(\result_x1_x3_imag[5]~30 ));
defparam \result_x1_x3_imag[5]~29 .lut_mask = 16'h96DF;
defparam \result_x1_x3_imag[5]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_imag[6]~31 (
	.dataa(\Add6~13_combout ),
	.datab(\x_1_imag_held[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_imag[5]~30 ),
	.combout(\result_x1_x3_imag[6]~31_combout ),
	.cout(\result_x1_x3_imag[6]~32 ));
defparam \result_x1_x3_imag[6]~31 .lut_mask = 16'h96BF;
defparam \result_x1_x3_imag[6]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_imag[7]~33 (
	.dataa(\Add6~12_combout ),
	.datab(\x_1_imag_held[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_imag[6]~32 ),
	.combout(\result_x1_x3_imag[7]~33_combout ),
	.cout(\result_x1_x3_imag[7]~34 ));
defparam \result_x1_x3_imag[7]~33 .lut_mask = 16'h96DF;
defparam \result_x1_x3_imag[7]~33 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_imag[8]~35 (
	.dataa(\Add6~11_combout ),
	.datab(\x_1_imag_held[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_imag[7]~34 ),
	.combout(\result_x1_x3_imag[8]~35_combout ),
	.cout(\result_x1_x3_imag[8]~36 ));
defparam \result_x1_x3_imag[8]~35 .lut_mask = 16'h96BF;
defparam \result_x1_x3_imag[8]~35 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_imag[9]~37 (
	.dataa(\Add6~10_combout ),
	.datab(\x_1_imag_held[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_imag[8]~36 ),
	.combout(\result_x1_x3_imag[9]~37_combout ),
	.cout(\result_x1_x3_imag[9]~38 ));
defparam \result_x1_x3_imag[9]~37 .lut_mask = 16'h96DF;
defparam \result_x1_x3_imag[9]~37 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_imag[10]~39 (
	.dataa(\Add6~9_combout ),
	.datab(\x_1_imag_held[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_imag[9]~38 ),
	.combout(\result_x1_x3_imag[10]~39_combout ),
	.cout(\result_x1_x3_imag[10]~40 ));
defparam \result_x1_x3_imag[10]~39 .lut_mask = 16'h96BF;
defparam \result_x1_x3_imag[10]~39 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_imag[11]~41 (
	.dataa(\Add6~8_combout ),
	.datab(\x_1_imag_held[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_imag[10]~40 ),
	.combout(\result_x1_x3_imag[11]~41_combout ),
	.cout(\result_x1_x3_imag[11]~42 ));
defparam \result_x1_x3_imag[11]~41 .lut_mask = 16'h96DF;
defparam \result_x1_x3_imag[11]~41 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_imag[12]~43 (
	.dataa(\Add6~7_combout ),
	.datab(\x_1_imag_held[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_imag[11]~42 ),
	.combout(\result_x1_x3_imag[12]~43_combout ),
	.cout(\result_x1_x3_imag[12]~44 ));
defparam \result_x1_x3_imag[12]~43 .lut_mask = 16'h96BF;
defparam \result_x1_x3_imag[12]~43 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_imag[13]~45 (
	.dataa(\Add6~6_combout ),
	.datab(\x_1_imag_held[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_imag[12]~44 ),
	.combout(\result_x1_x3_imag[13]~45_combout ),
	.cout(\result_x1_x3_imag[13]~46 ));
defparam \result_x1_x3_imag[13]~45 .lut_mask = 16'h96DF;
defparam \result_x1_x3_imag[13]~45 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_imag[14]~47 (
	.dataa(\Add6~5_combout ),
	.datab(\x_1_imag_held[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_imag[13]~46 ),
	.combout(\result_x1_x3_imag[14]~47_combout ),
	.cout(\result_x1_x3_imag[14]~48 ));
defparam \result_x1_x3_imag[14]~47 .lut_mask = 16'h96BF;
defparam \result_x1_x3_imag[14]~47 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_imag[15]~49 (
	.dataa(\Add6~4_combout ),
	.datab(\x_1_imag_held[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_imag[14]~48 ),
	.combout(\result_x1_x3_imag[15]~49_combout ),
	.cout(\result_x1_x3_imag[15]~50 ));
defparam \result_x1_x3_imag[15]~49 .lut_mask = 16'h96DF;
defparam \result_x1_x3_imag[15]~49 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_imag[16]~51 (
	.dataa(\Add6~4_combout ),
	.datab(\x_1_imag_held[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\result_x1_x3_imag[15]~50 ),
	.combout(\result_x1_x3_imag[16]~51_combout ),
	.cout());
defparam \result_x1_x3_imag[16]~51 .lut_mask = 16'h9696;
defparam \result_x1_x3_imag[16]~51 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_real[0]~18 (
	.dataa(\si[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\result_x2_x4_real[0]~18_cout ));
defparam \result_x2_x4_real[0]~18 .lut_mask = 16'h0055;
defparam \result_x2_x4_real[0]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \result_x2_x4_real[0]~19 (
	.dataa(\Add2~3_combout ),
	.datab(\x_2_real_held[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_real[0]~18_cout ),
	.combout(\result_x2_x4_real[0]~19_combout ),
	.cout(\result_x2_x4_real[0]~20 ));
defparam \result_x2_x4_real[0]~19 .lut_mask = 16'h96BF;
defparam \result_x2_x4_real[0]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_real[1]~21 (
	.dataa(\Add2~2_combout ),
	.datab(\x_2_real_held[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_real[0]~20 ),
	.combout(\result_x2_x4_real[1]~21_combout ),
	.cout(\result_x2_x4_real[1]~22 ));
defparam \result_x2_x4_real[1]~21 .lut_mask = 16'h96DF;
defparam \result_x2_x4_real[1]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_real[2]~23 (
	.dataa(\Add2~1_combout ),
	.datab(\x_2_real_held[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_real[1]~22 ),
	.combout(\result_x2_x4_real[2]~23_combout ),
	.cout(\result_x2_x4_real[2]~24 ));
defparam \result_x2_x4_real[2]~23 .lut_mask = 16'h96BF;
defparam \result_x2_x4_real[2]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_real[0]~18 (
	.dataa(\si[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\result_x1_x3_real[0]~18_cout ));
defparam \result_x1_x3_real[0]~18 .lut_mask = 16'h0055;
defparam \result_x1_x3_real[0]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \result_x1_x3_real[0]~19 (
	.dataa(\Add0~3_combout ),
	.datab(\x_1_real_held[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_real[0]~18_cout ),
	.combout(\result_x1_x3_real[0]~19_combout ),
	.cout(\result_x1_x3_real[0]~20 ));
defparam \result_x1_x3_real[0]~19 .lut_mask = 16'h96BF;
defparam \result_x1_x3_real[0]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_real[1]~21 (
	.dataa(\Add0~2_combout ),
	.datab(\x_1_real_held[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_real[0]~20 ),
	.combout(\result_x1_x3_real[1]~21_combout ),
	.cout(\result_x1_x3_real[1]~22 ));
defparam \result_x1_x3_real[1]~21 .lut_mask = 16'h96DF;
defparam \result_x1_x3_real[1]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_real[2]~23 (
	.dataa(\Add0~1_combout ),
	.datab(\x_1_real_held[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_real[1]~22 ),
	.combout(\result_x1_x3_real[2]~23_combout ),
	.cout(\result_x1_x3_real[2]~24 ));
defparam \result_x1_x3_real[2]~23 .lut_mask = 16'h96BF;
defparam \result_x1_x3_real[2]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_real[3]~25 (
	.dataa(\Add2~16_combout ),
	.datab(\x_2_real_held[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_real[2]~24 ),
	.combout(\result_x2_x4_real[3]~25_combout ),
	.cout(\result_x2_x4_real[3]~26 ));
defparam \result_x2_x4_real[3]~25 .lut_mask = 16'h96DF;
defparam \result_x2_x4_real[3]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_real[4]~27 (
	.dataa(\Add2~15_combout ),
	.datab(\x_2_real_held[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_real[3]~26 ),
	.combout(\result_x2_x4_real[4]~27_combout ),
	.cout(\result_x2_x4_real[4]~28 ));
defparam \result_x2_x4_real[4]~27 .lut_mask = 16'h96BF;
defparam \result_x2_x4_real[4]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_real[5]~29 (
	.dataa(\Add2~14_combout ),
	.datab(\x_2_real_held[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_real[4]~28 ),
	.combout(\result_x2_x4_real[5]~29_combout ),
	.cout(\result_x2_x4_real[5]~30 ));
defparam \result_x2_x4_real[5]~29 .lut_mask = 16'h96DF;
defparam \result_x2_x4_real[5]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_real[6]~31 (
	.dataa(\Add2~13_combout ),
	.datab(\x_2_real_held[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_real[5]~30 ),
	.combout(\result_x2_x4_real[6]~31_combout ),
	.cout(\result_x2_x4_real[6]~32 ));
defparam \result_x2_x4_real[6]~31 .lut_mask = 16'h96BF;
defparam \result_x2_x4_real[6]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_real[7]~33 (
	.dataa(\Add2~12_combout ),
	.datab(\x_2_real_held[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_real[6]~32 ),
	.combout(\result_x2_x4_real[7]~33_combout ),
	.cout(\result_x2_x4_real[7]~34 ));
defparam \result_x2_x4_real[7]~33 .lut_mask = 16'h96DF;
defparam \result_x2_x4_real[7]~33 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_real[8]~35 (
	.dataa(\Add2~11_combout ),
	.datab(\x_2_real_held[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_real[7]~34 ),
	.combout(\result_x2_x4_real[8]~35_combout ),
	.cout(\result_x2_x4_real[8]~36 ));
defparam \result_x2_x4_real[8]~35 .lut_mask = 16'h96BF;
defparam \result_x2_x4_real[8]~35 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_real[9]~37 (
	.dataa(\Add2~10_combout ),
	.datab(\x_2_real_held[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_real[8]~36 ),
	.combout(\result_x2_x4_real[9]~37_combout ),
	.cout(\result_x2_x4_real[9]~38 ));
defparam \result_x2_x4_real[9]~37 .lut_mask = 16'h96DF;
defparam \result_x2_x4_real[9]~37 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_real[10]~39 (
	.dataa(\Add2~9_combout ),
	.datab(\x_2_real_held[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_real[9]~38 ),
	.combout(\result_x2_x4_real[10]~39_combout ),
	.cout(\result_x2_x4_real[10]~40 ));
defparam \result_x2_x4_real[10]~39 .lut_mask = 16'h96BF;
defparam \result_x2_x4_real[10]~39 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_real[11]~41 (
	.dataa(\Add2~8_combout ),
	.datab(\x_2_real_held[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_real[10]~40 ),
	.combout(\result_x2_x4_real[11]~41_combout ),
	.cout(\result_x2_x4_real[11]~42 ));
defparam \result_x2_x4_real[11]~41 .lut_mask = 16'h96DF;
defparam \result_x2_x4_real[11]~41 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_real[12]~43 (
	.dataa(\Add2~7_combout ),
	.datab(\x_2_real_held[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_real[11]~42 ),
	.combout(\result_x2_x4_real[12]~43_combout ),
	.cout(\result_x2_x4_real[12]~44 ));
defparam \result_x2_x4_real[12]~43 .lut_mask = 16'h96BF;
defparam \result_x2_x4_real[12]~43 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_real[13]~45 (
	.dataa(\Add2~6_combout ),
	.datab(\x_2_real_held[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_real[12]~44 ),
	.combout(\result_x2_x4_real[13]~45_combout ),
	.cout(\result_x2_x4_real[13]~46 ));
defparam \result_x2_x4_real[13]~45 .lut_mask = 16'h96DF;
defparam \result_x2_x4_real[13]~45 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_real[14]~47 (
	.dataa(\Add2~5_combout ),
	.datab(\x_2_real_held[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_real[13]~46 ),
	.combout(\result_x2_x4_real[14]~47_combout ),
	.cout(\result_x2_x4_real[14]~48 ));
defparam \result_x2_x4_real[14]~47 .lut_mask = 16'h96BF;
defparam \result_x2_x4_real[14]~47 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_real[15]~49 (
	.dataa(\Add2~4_combout ),
	.datab(\x_2_real_held[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x2_x4_real[14]~48 ),
	.combout(\result_x2_x4_real[15]~49_combout ),
	.cout(\result_x2_x4_real[15]~50 ));
defparam \result_x2_x4_real[15]~49 .lut_mask = 16'h96DF;
defparam \result_x2_x4_real[15]~49 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x2_x4_real[16]~51 (
	.dataa(\Add2~4_combout ),
	.datab(\x_2_real_held[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\result_x2_x4_real[15]~50 ),
	.combout(\result_x2_x4_real[16]~51_combout ),
	.cout());
defparam \result_x2_x4_real[16]~51 .lut_mask = 16'h9696;
defparam \result_x2_x4_real[16]~51 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_real[3]~25 (
	.dataa(\Add0~16_combout ),
	.datab(\x_1_real_held[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_real[2]~24 ),
	.combout(\result_x1_x3_real[3]~25_combout ),
	.cout(\result_x1_x3_real[3]~26 ));
defparam \result_x1_x3_real[3]~25 .lut_mask = 16'h96DF;
defparam \result_x1_x3_real[3]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_real[4]~27 (
	.dataa(\Add0~15_combout ),
	.datab(\x_1_real_held[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_real[3]~26 ),
	.combout(\result_x1_x3_real[4]~27_combout ),
	.cout(\result_x1_x3_real[4]~28 ));
defparam \result_x1_x3_real[4]~27 .lut_mask = 16'h96BF;
defparam \result_x1_x3_real[4]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_real[5]~29 (
	.dataa(\Add0~14_combout ),
	.datab(\x_1_real_held[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_real[4]~28 ),
	.combout(\result_x1_x3_real[5]~29_combout ),
	.cout(\result_x1_x3_real[5]~30 ));
defparam \result_x1_x3_real[5]~29 .lut_mask = 16'h96DF;
defparam \result_x1_x3_real[5]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_real[6]~31 (
	.dataa(\Add0~13_combout ),
	.datab(\x_1_real_held[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_real[5]~30 ),
	.combout(\result_x1_x3_real[6]~31_combout ),
	.cout(\result_x1_x3_real[6]~32 ));
defparam \result_x1_x3_real[6]~31 .lut_mask = 16'h96BF;
defparam \result_x1_x3_real[6]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_real[7]~33 (
	.dataa(\Add0~12_combout ),
	.datab(\x_1_real_held[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_real[6]~32 ),
	.combout(\result_x1_x3_real[7]~33_combout ),
	.cout(\result_x1_x3_real[7]~34 ));
defparam \result_x1_x3_real[7]~33 .lut_mask = 16'h96DF;
defparam \result_x1_x3_real[7]~33 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_real[8]~35 (
	.dataa(\Add0~11_combout ),
	.datab(\x_1_real_held[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_real[7]~34 ),
	.combout(\result_x1_x3_real[8]~35_combout ),
	.cout(\result_x1_x3_real[8]~36 ));
defparam \result_x1_x3_real[8]~35 .lut_mask = 16'h96BF;
defparam \result_x1_x3_real[8]~35 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_real[9]~37 (
	.dataa(\Add0~10_combout ),
	.datab(\x_1_real_held[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_real[8]~36 ),
	.combout(\result_x1_x3_real[9]~37_combout ),
	.cout(\result_x1_x3_real[9]~38 ));
defparam \result_x1_x3_real[9]~37 .lut_mask = 16'h96DF;
defparam \result_x1_x3_real[9]~37 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_real[10]~39 (
	.dataa(\Add0~9_combout ),
	.datab(\x_1_real_held[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_real[9]~38 ),
	.combout(\result_x1_x3_real[10]~39_combout ),
	.cout(\result_x1_x3_real[10]~40 ));
defparam \result_x1_x3_real[10]~39 .lut_mask = 16'h96BF;
defparam \result_x1_x3_real[10]~39 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_real[11]~41 (
	.dataa(\Add0~8_combout ),
	.datab(\x_1_real_held[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_real[10]~40 ),
	.combout(\result_x1_x3_real[11]~41_combout ),
	.cout(\result_x1_x3_real[11]~42 ));
defparam \result_x1_x3_real[11]~41 .lut_mask = 16'h96DF;
defparam \result_x1_x3_real[11]~41 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_real[12]~43 (
	.dataa(\Add0~7_combout ),
	.datab(\x_1_real_held[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_real[11]~42 ),
	.combout(\result_x1_x3_real[12]~43_combout ),
	.cout(\result_x1_x3_real[12]~44 ));
defparam \result_x1_x3_real[12]~43 .lut_mask = 16'h96BF;
defparam \result_x1_x3_real[12]~43 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_real[13]~45 (
	.dataa(\Add0~6_combout ),
	.datab(\x_1_real_held[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_real[12]~44 ),
	.combout(\result_x1_x3_real[13]~45_combout ),
	.cout(\result_x1_x3_real[13]~46 ));
defparam \result_x1_x3_real[13]~45 .lut_mask = 16'h96DF;
defparam \result_x1_x3_real[13]~45 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_real[14]~47 (
	.dataa(\Add0~5_combout ),
	.datab(\x_1_real_held[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_real[13]~46 ),
	.combout(\result_x1_x3_real[14]~47_combout ),
	.cout(\result_x1_x3_real[14]~48 ));
defparam \result_x1_x3_real[14]~47 .lut_mask = 16'h96BF;
defparam \result_x1_x3_real[14]~47 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_real[15]~49 (
	.dataa(\Add0~4_combout ),
	.datab(\x_1_real_held[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_x1_x3_real[14]~48 ),
	.combout(\result_x1_x3_real[15]~49_combout ),
	.cout(\result_x1_x3_real[15]~50 ));
defparam \result_x1_x3_real[15]~49 .lut_mask = 16'h96DF;
defparam \result_x1_x3_real[15]~49 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_x1_x3_real[16]~51 (
	.dataa(\Add0~4_combout ),
	.datab(\x_1_real_held[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\result_x1_x3_real[15]~50 ),
	.combout(\result_x1_x3_real[16]~51_combout ),
	.cout());
defparam \result_x1_x3_real[16]~51 .lut_mask = 16'h9696;
defparam \result_x1_x3_real[16]~51 .sum_lutc_input = "cin";

dffeas \si[0] (
	.clk(clk),
	.d(\si~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\si[0]~q ),
	.prn(vcc));
defparam \si[0] .is_wysiwyg = "true";
defparam \si[0] .power_up = "low";

cycloneive_lcell_comb \Add10~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[0]~q ),
	.datad(\result_x2_x4_imag[2]~q ),
	.cin(gnd),
	.combout(\Add10~1_combout ),
	.cout());
defparam \Add10~1 .lut_mask = 16'h0FF0;
defparam \Add10~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add10~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[0]~q ),
	.datad(\result_x2_x4_imag[1]~q ),
	.cin(gnd),
	.combout(\Add10~2_combout ),
	.cout());
defparam \Add10~2 .lut_mask = 16'h0FF0;
defparam \Add10~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add10~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[0]~q ),
	.datad(\result_x2_x4_imag[0]~q ),
	.cin(gnd),
	.combout(\Add10~3_combout ),
	.cout());
defparam \Add10~3 .lut_mask = 16'h0FF0;
defparam \Add10~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add10~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[0]~q ),
	.datad(\result_x2_x4_imag[16]~q ),
	.cin(gnd),
	.combout(\Add10~4_combout ),
	.cout());
defparam \Add10~4 .lut_mask = 16'h0FF0;
defparam \Add10~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add10~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[0]~q ),
	.datad(\result_x2_x4_imag[15]~q ),
	.cin(gnd),
	.combout(\Add10~5_combout ),
	.cout());
defparam \Add10~5 .lut_mask = 16'h0FF0;
defparam \Add10~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add10~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[0]~q ),
	.datad(\result_x2_x4_imag[14]~q ),
	.cin(gnd),
	.combout(\Add10~6_combout ),
	.cout());
defparam \Add10~6 .lut_mask = 16'h0FF0;
defparam \Add10~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add10~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[0]~q ),
	.datad(\result_x2_x4_imag[13]~q ),
	.cin(gnd),
	.combout(\Add10~7_combout ),
	.cout());
defparam \Add10~7 .lut_mask = 16'h0FF0;
defparam \Add10~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add10~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[0]~q ),
	.datad(\result_x2_x4_imag[12]~q ),
	.cin(gnd),
	.combout(\Add10~8_combout ),
	.cout());
defparam \Add10~8 .lut_mask = 16'h0FF0;
defparam \Add10~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add10~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[0]~q ),
	.datad(\result_x2_x4_imag[11]~q ),
	.cin(gnd),
	.combout(\Add10~9_combout ),
	.cout());
defparam \Add10~9 .lut_mask = 16'h0FF0;
defparam \Add10~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add10~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[0]~q ),
	.datad(\result_x2_x4_imag[10]~q ),
	.cin(gnd),
	.combout(\Add10~10_combout ),
	.cout());
defparam \Add10~10 .lut_mask = 16'h0FF0;
defparam \Add10~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add10~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[0]~q ),
	.datad(\result_x2_x4_imag[9]~q ),
	.cin(gnd),
	.combout(\Add10~11_combout ),
	.cout());
defparam \Add10~11 .lut_mask = 16'h0FF0;
defparam \Add10~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add10~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[0]~q ),
	.datad(\result_x2_x4_imag[8]~q ),
	.cin(gnd),
	.combout(\Add10~12_combout ),
	.cout());
defparam \Add10~12 .lut_mask = 16'h0FF0;
defparam \Add10~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add10~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[0]~q ),
	.datad(\result_x2_x4_imag[7]~q ),
	.cin(gnd),
	.combout(\Add10~13_combout ),
	.cout());
defparam \Add10~13 .lut_mask = 16'h0FF0;
defparam \Add10~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add10~14 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[0]~q ),
	.datad(\result_x2_x4_imag[6]~q ),
	.cin(gnd),
	.combout(\Add10~14_combout ),
	.cout());
defparam \Add10~14 .lut_mask = 16'h0FF0;
defparam \Add10~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add10~15 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[0]~q ),
	.datad(\result_x2_x4_imag[5]~q ),
	.cin(gnd),
	.combout(\Add10~15_combout ),
	.cout());
defparam \Add10~15 .lut_mask = 16'h0FF0;
defparam \Add10~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add10~16 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[0]~q ),
	.datad(\result_x2_x4_imag[4]~q ),
	.cin(gnd),
	.combout(\Add10~16_combout ),
	.cout());
defparam \Add10~16 .lut_mask = 16'h0FF0;
defparam \Add10~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add10~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[0]~q ),
	.datad(\result_x2_x4_imag[3]~q ),
	.cin(gnd),
	.combout(\Add10~17_combout ),
	.cout());
defparam \Add10~17 .lut_mask = 16'h0FF0;
defparam \Add10~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sr[0]~q ),
	.datad(\result_x2_x4_real[2]~q ),
	.cin(gnd),
	.combout(\Add4~1_combout ),
	.cout());
defparam \Add4~1 .lut_mask = 16'h0FF0;
defparam \Add4~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add4~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sr[0]~q ),
	.datad(\result_x2_x4_real[1]~q ),
	.cin(gnd),
	.combout(\Add4~2_combout ),
	.cout());
defparam \Add4~2 .lut_mask = 16'h0FF0;
defparam \Add4~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add4~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sr[0]~q ),
	.datad(\result_x2_x4_real[0]~q ),
	.cin(gnd),
	.combout(\Add4~3_combout ),
	.cout());
defparam \Add4~3 .lut_mask = 16'h0FF0;
defparam \Add4~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add4~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sr[0]~q ),
	.datad(\result_x2_x4_real[16]~q ),
	.cin(gnd),
	.combout(\Add4~4_combout ),
	.cout());
defparam \Add4~4 .lut_mask = 16'h0FF0;
defparam \Add4~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add4~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sr[0]~q ),
	.datad(\result_x2_x4_real[15]~q ),
	.cin(gnd),
	.combout(\Add4~5_combout ),
	.cout());
defparam \Add4~5 .lut_mask = 16'h0FF0;
defparam \Add4~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add4~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sr[0]~q ),
	.datad(\result_x2_x4_real[14]~q ),
	.cin(gnd),
	.combout(\Add4~6_combout ),
	.cout());
defparam \Add4~6 .lut_mask = 16'h0FF0;
defparam \Add4~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add4~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sr[0]~q ),
	.datad(\result_x2_x4_real[13]~q ),
	.cin(gnd),
	.combout(\Add4~7_combout ),
	.cout());
defparam \Add4~7 .lut_mask = 16'h0FF0;
defparam \Add4~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add4~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sr[0]~q ),
	.datad(\result_x2_x4_real[12]~q ),
	.cin(gnd),
	.combout(\Add4~8_combout ),
	.cout());
defparam \Add4~8 .lut_mask = 16'h0FF0;
defparam \Add4~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sr[0]~q ),
	.datad(\result_x2_x4_real[11]~q ),
	.cin(gnd),
	.combout(\Add4~9_combout ),
	.cout());
defparam \Add4~9 .lut_mask = 16'h0FF0;
defparam \Add4~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add4~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sr[0]~q ),
	.datad(\result_x2_x4_real[10]~q ),
	.cin(gnd),
	.combout(\Add4~10_combout ),
	.cout());
defparam \Add4~10 .lut_mask = 16'h0FF0;
defparam \Add4~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add4~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sr[0]~q ),
	.datad(\result_x2_x4_real[9]~q ),
	.cin(gnd),
	.combout(\Add4~11_combout ),
	.cout());
defparam \Add4~11 .lut_mask = 16'h0FF0;
defparam \Add4~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add4~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sr[0]~q ),
	.datad(\result_x2_x4_real[8]~q ),
	.cin(gnd),
	.combout(\Add4~12_combout ),
	.cout());
defparam \Add4~12 .lut_mask = 16'h0FF0;
defparam \Add4~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add4~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sr[0]~q ),
	.datad(\result_x2_x4_real[7]~q ),
	.cin(gnd),
	.combout(\Add4~13_combout ),
	.cout());
defparam \Add4~13 .lut_mask = 16'h0FF0;
defparam \Add4~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add4~14 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sr[0]~q ),
	.datad(\result_x2_x4_real[6]~q ),
	.cin(gnd),
	.combout(\Add4~14_combout ),
	.cout());
defparam \Add4~14 .lut_mask = 16'h0FF0;
defparam \Add4~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add4~15 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sr[0]~q ),
	.datad(\result_x2_x4_real[5]~q ),
	.cin(gnd),
	.combout(\Add4~15_combout ),
	.cout());
defparam \Add4~15 .lut_mask = 16'h0FF0;
defparam \Add4~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add4~16 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sr[0]~q ),
	.datad(\result_x2_x4_real[4]~q ),
	.cin(gnd),
	.combout(\Add4~16_combout ),
	.cout());
defparam \Add4~16 .lut_mask = 16'h0FF0;
defparam \Add4~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add4~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sr[0]~q ),
	.datad(\result_x2_x4_real[3]~q ),
	.cin(gnd),
	.combout(\Add4~17_combout ),
	.cout());
defparam \Add4~17 .lut_mask = 16'h0FF0;
defparam \Add4~17 .sum_lutc_input = "datac";

dffeas \sel_arr[9][1] (
	.clk(clk),
	.d(\sel_arr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[9][1]~q ),
	.prn(vcc));
defparam \sel_arr[9][1] .is_wysiwyg = "true";
defparam \sel_arr[9][1] .power_up = "low";

cycloneive_lcell_comb \si~0 (
	.dataa(\sel_arr[9][1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset),
	.cin(gnd),
	.combout(\si~0_combout ),
	.cout());
defparam \si~0 .lut_mask = 16'hFF55;
defparam \si~0 .sum_lutc_input = "datac";

dffeas \si[1] (
	.clk(clk),
	.d(\si~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\si[1]~q ),
	.prn(vcc));
defparam \si[1] .is_wysiwyg = "true";
defparam \si[1] .power_up = "low";

dffeas \x_4_imag_held[2] (
	.clk(clk),
	.d(\Mux261~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_imag_held[2]~q ),
	.prn(vcc));
defparam \x_4_imag_held[2] .is_wysiwyg = "true";
defparam \x_4_imag_held[2] .power_up = "low";

cycloneive_lcell_comb \Add8~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_imag_held[2]~q ),
	.cin(gnd),
	.combout(\Add8~1_combout ),
	.cout());
defparam \Add8~1 .lut_mask = 16'h0FF0;
defparam \Add8~1 .sum_lutc_input = "datac";

dffeas \x_2_imag_held[2] (
	.clk(clk),
	.d(\Mux227~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_imag_held[2]~q ),
	.prn(vcc));
defparam \x_2_imag_held[2] .is_wysiwyg = "true";
defparam \x_2_imag_held[2] .power_up = "low";

dffeas \x_4_imag_held[1] (
	.clk(clk),
	.d(\Mux262~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_imag_held[1]~q ),
	.prn(vcc));
defparam \x_4_imag_held[1] .is_wysiwyg = "true";
defparam \x_4_imag_held[1] .power_up = "low";

cycloneive_lcell_comb \Add8~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_imag_held[1]~q ),
	.cin(gnd),
	.combout(\Add8~2_combout ),
	.cout());
defparam \Add8~2 .lut_mask = 16'h0FF0;
defparam \Add8~2 .sum_lutc_input = "datac";

dffeas \x_2_imag_held[1] (
	.clk(clk),
	.d(\Mux228~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_imag_held[1]~q ),
	.prn(vcc));
defparam \x_2_imag_held[1] .is_wysiwyg = "true";
defparam \x_2_imag_held[1] .power_up = "low";

dffeas \x_4_imag_held[0] (
	.clk(clk),
	.d(\Mux263~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_imag_held[0]~q ),
	.prn(vcc));
defparam \x_4_imag_held[0] .is_wysiwyg = "true";
defparam \x_4_imag_held[0] .power_up = "low";

cycloneive_lcell_comb \Add8~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_imag_held[0]~q ),
	.cin(gnd),
	.combout(\Add8~3_combout ),
	.cout());
defparam \Add8~3 .lut_mask = 16'h0FF0;
defparam \Add8~3 .sum_lutc_input = "datac";

dffeas \x_2_imag_held[0] (
	.clk(clk),
	.d(\Mux229~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_imag_held[0]~q ),
	.prn(vcc));
defparam \x_2_imag_held[0] .is_wysiwyg = "true";
defparam \x_2_imag_held[0] .power_up = "low";

dffeas \x_3_imag_held[2] (
	.clk(clk),
	.d(\butterfly_st1[2][1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_imag_held[2]~q ),
	.prn(vcc));
defparam \x_3_imag_held[2] .is_wysiwyg = "true";
defparam \x_3_imag_held[2] .power_up = "low";

cycloneive_lcell_comb \Add6~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_imag_held[2]~q ),
	.cin(gnd),
	.combout(\Add6~1_combout ),
	.cout());
defparam \Add6~1 .lut_mask = 16'h0FF0;
defparam \Add6~1 .sum_lutc_input = "datac";

dffeas \x_1_imag_held[2] (
	.clk(clk),
	.d(\butterfly_st1[0][1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_imag_held[2]~q ),
	.prn(vcc));
defparam \x_1_imag_held[2] .is_wysiwyg = "true";
defparam \x_1_imag_held[2] .power_up = "low";

dffeas \x_3_imag_held[1] (
	.clk(clk),
	.d(\butterfly_st1[2][1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_imag_held[1]~q ),
	.prn(vcc));
defparam \x_3_imag_held[1] .is_wysiwyg = "true";
defparam \x_3_imag_held[1] .power_up = "low";

cycloneive_lcell_comb \Add6~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_imag_held[1]~q ),
	.cin(gnd),
	.combout(\Add6~2_combout ),
	.cout());
defparam \Add6~2 .lut_mask = 16'h0FF0;
defparam \Add6~2 .sum_lutc_input = "datac";

dffeas \x_1_imag_held[1] (
	.clk(clk),
	.d(\butterfly_st1[0][1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_imag_held[1]~q ),
	.prn(vcc));
defparam \x_1_imag_held[1] .is_wysiwyg = "true";
defparam \x_1_imag_held[1] .power_up = "low";

dffeas \x_3_imag_held[0] (
	.clk(clk),
	.d(\butterfly_st1[2][1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_imag_held[0]~q ),
	.prn(vcc));
defparam \x_3_imag_held[0] .is_wysiwyg = "true";
defparam \x_3_imag_held[0] .power_up = "low";

cycloneive_lcell_comb \Add6~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_imag_held[0]~q ),
	.cin(gnd),
	.combout(\Add6~3_combout ),
	.cout());
defparam \Add6~3 .lut_mask = 16'h0FF0;
defparam \Add6~3 .sum_lutc_input = "datac";

dffeas \x_1_imag_held[0] (
	.clk(clk),
	.d(\butterfly_st1[0][1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_imag_held[0]~q ),
	.prn(vcc));
defparam \x_1_imag_held[0] .is_wysiwyg = "true";
defparam \x_1_imag_held[0] .power_up = "low";

dffeas \x_4_imag_held[15] (
	.clk(clk),
	.d(\Mux248~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_imag_held[15]~q ),
	.prn(vcc));
defparam \x_4_imag_held[15] .is_wysiwyg = "true";
defparam \x_4_imag_held[15] .power_up = "low";

cycloneive_lcell_comb \Add8~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_imag_held[15]~q ),
	.cin(gnd),
	.combout(\Add8~4_combout ),
	.cout());
defparam \Add8~4 .lut_mask = 16'h0FF0;
defparam \Add8~4 .sum_lutc_input = "datac";

dffeas \x_2_imag_held[15] (
	.clk(clk),
	.d(\Mux214~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_imag_held[15]~q ),
	.prn(vcc));
defparam \x_2_imag_held[15] .is_wysiwyg = "true";
defparam \x_2_imag_held[15] .power_up = "low";

dffeas \x_4_imag_held[14] (
	.clk(clk),
	.d(\Mux249~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_imag_held[14]~q ),
	.prn(vcc));
defparam \x_4_imag_held[14] .is_wysiwyg = "true";
defparam \x_4_imag_held[14] .power_up = "low";

cycloneive_lcell_comb \Add8~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_imag_held[14]~q ),
	.cin(gnd),
	.combout(\Add8~5_combout ),
	.cout());
defparam \Add8~5 .lut_mask = 16'h0FF0;
defparam \Add8~5 .sum_lutc_input = "datac";

dffeas \x_2_imag_held[14] (
	.clk(clk),
	.d(\Mux215~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_imag_held[14]~q ),
	.prn(vcc));
defparam \x_2_imag_held[14] .is_wysiwyg = "true";
defparam \x_2_imag_held[14] .power_up = "low";

dffeas \x_4_imag_held[13] (
	.clk(clk),
	.d(\Mux250~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_imag_held[13]~q ),
	.prn(vcc));
defparam \x_4_imag_held[13] .is_wysiwyg = "true";
defparam \x_4_imag_held[13] .power_up = "low";

cycloneive_lcell_comb \Add8~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_imag_held[13]~q ),
	.cin(gnd),
	.combout(\Add8~6_combout ),
	.cout());
defparam \Add8~6 .lut_mask = 16'h0FF0;
defparam \Add8~6 .sum_lutc_input = "datac";

dffeas \x_2_imag_held[13] (
	.clk(clk),
	.d(\Mux216~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_imag_held[13]~q ),
	.prn(vcc));
defparam \x_2_imag_held[13] .is_wysiwyg = "true";
defparam \x_2_imag_held[13] .power_up = "low";

dffeas \x_4_imag_held[12] (
	.clk(clk),
	.d(\Mux251~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_imag_held[12]~q ),
	.prn(vcc));
defparam \x_4_imag_held[12] .is_wysiwyg = "true";
defparam \x_4_imag_held[12] .power_up = "low";

cycloneive_lcell_comb \Add8~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_imag_held[12]~q ),
	.cin(gnd),
	.combout(\Add8~7_combout ),
	.cout());
defparam \Add8~7 .lut_mask = 16'h0FF0;
defparam \Add8~7 .sum_lutc_input = "datac";

dffeas \x_2_imag_held[12] (
	.clk(clk),
	.d(\Mux217~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_imag_held[12]~q ),
	.prn(vcc));
defparam \x_2_imag_held[12] .is_wysiwyg = "true";
defparam \x_2_imag_held[12] .power_up = "low";

dffeas \x_4_imag_held[11] (
	.clk(clk),
	.d(\Mux252~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_imag_held[11]~q ),
	.prn(vcc));
defparam \x_4_imag_held[11] .is_wysiwyg = "true";
defparam \x_4_imag_held[11] .power_up = "low";

cycloneive_lcell_comb \Add8~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_imag_held[11]~q ),
	.cin(gnd),
	.combout(\Add8~8_combout ),
	.cout());
defparam \Add8~8 .lut_mask = 16'h0FF0;
defparam \Add8~8 .sum_lutc_input = "datac";

dffeas \x_2_imag_held[11] (
	.clk(clk),
	.d(\Mux218~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_imag_held[11]~q ),
	.prn(vcc));
defparam \x_2_imag_held[11] .is_wysiwyg = "true";
defparam \x_2_imag_held[11] .power_up = "low";

dffeas \x_4_imag_held[10] (
	.clk(clk),
	.d(\Mux253~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_imag_held[10]~q ),
	.prn(vcc));
defparam \x_4_imag_held[10] .is_wysiwyg = "true";
defparam \x_4_imag_held[10] .power_up = "low";

cycloneive_lcell_comb \Add8~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_imag_held[10]~q ),
	.cin(gnd),
	.combout(\Add8~9_combout ),
	.cout());
defparam \Add8~9 .lut_mask = 16'h0FF0;
defparam \Add8~9 .sum_lutc_input = "datac";

dffeas \x_2_imag_held[10] (
	.clk(clk),
	.d(\Mux219~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_imag_held[10]~q ),
	.prn(vcc));
defparam \x_2_imag_held[10] .is_wysiwyg = "true";
defparam \x_2_imag_held[10] .power_up = "low";

dffeas \x_4_imag_held[9] (
	.clk(clk),
	.d(\Mux254~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_imag_held[9]~q ),
	.prn(vcc));
defparam \x_4_imag_held[9] .is_wysiwyg = "true";
defparam \x_4_imag_held[9] .power_up = "low";

cycloneive_lcell_comb \Add8~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_imag_held[9]~q ),
	.cin(gnd),
	.combout(\Add8~10_combout ),
	.cout());
defparam \Add8~10 .lut_mask = 16'h0FF0;
defparam \Add8~10 .sum_lutc_input = "datac";

dffeas \x_2_imag_held[9] (
	.clk(clk),
	.d(\Mux220~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_imag_held[9]~q ),
	.prn(vcc));
defparam \x_2_imag_held[9] .is_wysiwyg = "true";
defparam \x_2_imag_held[9] .power_up = "low";

dffeas \x_4_imag_held[8] (
	.clk(clk),
	.d(\Mux255~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_imag_held[8]~q ),
	.prn(vcc));
defparam \x_4_imag_held[8] .is_wysiwyg = "true";
defparam \x_4_imag_held[8] .power_up = "low";

cycloneive_lcell_comb \Add8~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_imag_held[8]~q ),
	.cin(gnd),
	.combout(\Add8~11_combout ),
	.cout());
defparam \Add8~11 .lut_mask = 16'h0FF0;
defparam \Add8~11 .sum_lutc_input = "datac";

dffeas \x_2_imag_held[8] (
	.clk(clk),
	.d(\Mux221~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_imag_held[8]~q ),
	.prn(vcc));
defparam \x_2_imag_held[8] .is_wysiwyg = "true";
defparam \x_2_imag_held[8] .power_up = "low";

dffeas \x_4_imag_held[7] (
	.clk(clk),
	.d(\Mux256~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_imag_held[7]~q ),
	.prn(vcc));
defparam \x_4_imag_held[7] .is_wysiwyg = "true";
defparam \x_4_imag_held[7] .power_up = "low";

cycloneive_lcell_comb \Add8~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_imag_held[7]~q ),
	.cin(gnd),
	.combout(\Add8~12_combout ),
	.cout());
defparam \Add8~12 .lut_mask = 16'h0FF0;
defparam \Add8~12 .sum_lutc_input = "datac";

dffeas \x_2_imag_held[7] (
	.clk(clk),
	.d(\Mux222~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_imag_held[7]~q ),
	.prn(vcc));
defparam \x_2_imag_held[7] .is_wysiwyg = "true";
defparam \x_2_imag_held[7] .power_up = "low";

dffeas \x_4_imag_held[6] (
	.clk(clk),
	.d(\Mux257~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_imag_held[6]~q ),
	.prn(vcc));
defparam \x_4_imag_held[6] .is_wysiwyg = "true";
defparam \x_4_imag_held[6] .power_up = "low";

cycloneive_lcell_comb \Add8~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_imag_held[6]~q ),
	.cin(gnd),
	.combout(\Add8~13_combout ),
	.cout());
defparam \Add8~13 .lut_mask = 16'h0FF0;
defparam \Add8~13 .sum_lutc_input = "datac";

dffeas \x_2_imag_held[6] (
	.clk(clk),
	.d(\Mux223~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_imag_held[6]~q ),
	.prn(vcc));
defparam \x_2_imag_held[6] .is_wysiwyg = "true";
defparam \x_2_imag_held[6] .power_up = "low";

dffeas \x_4_imag_held[5] (
	.clk(clk),
	.d(\Mux258~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_imag_held[5]~q ),
	.prn(vcc));
defparam \x_4_imag_held[5] .is_wysiwyg = "true";
defparam \x_4_imag_held[5] .power_up = "low";

cycloneive_lcell_comb \Add8~14 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_imag_held[5]~q ),
	.cin(gnd),
	.combout(\Add8~14_combout ),
	.cout());
defparam \Add8~14 .lut_mask = 16'h0FF0;
defparam \Add8~14 .sum_lutc_input = "datac";

dffeas \x_2_imag_held[5] (
	.clk(clk),
	.d(\Mux224~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_imag_held[5]~q ),
	.prn(vcc));
defparam \x_2_imag_held[5] .is_wysiwyg = "true";
defparam \x_2_imag_held[5] .power_up = "low";

dffeas \x_4_imag_held[4] (
	.clk(clk),
	.d(\Mux259~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_imag_held[4]~q ),
	.prn(vcc));
defparam \x_4_imag_held[4] .is_wysiwyg = "true";
defparam \x_4_imag_held[4] .power_up = "low";

cycloneive_lcell_comb \Add8~15 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_imag_held[4]~q ),
	.cin(gnd),
	.combout(\Add8~15_combout ),
	.cout());
defparam \Add8~15 .lut_mask = 16'h0FF0;
defparam \Add8~15 .sum_lutc_input = "datac";

dffeas \x_2_imag_held[4] (
	.clk(clk),
	.d(\Mux225~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_imag_held[4]~q ),
	.prn(vcc));
defparam \x_2_imag_held[4] .is_wysiwyg = "true";
defparam \x_2_imag_held[4] .power_up = "low";

dffeas \x_4_imag_held[3] (
	.clk(clk),
	.d(\Mux260~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_imag_held[3]~q ),
	.prn(vcc));
defparam \x_4_imag_held[3] .is_wysiwyg = "true";
defparam \x_4_imag_held[3] .power_up = "low";

cycloneive_lcell_comb \Add8~16 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_imag_held[3]~q ),
	.cin(gnd),
	.combout(\Add8~16_combout ),
	.cout());
defparam \Add8~16 .lut_mask = 16'h0FF0;
defparam \Add8~16 .sum_lutc_input = "datac";

dffeas \x_2_imag_held[3] (
	.clk(clk),
	.d(\Mux226~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_imag_held[3]~q ),
	.prn(vcc));
defparam \x_2_imag_held[3] .is_wysiwyg = "true";
defparam \x_2_imag_held[3] .power_up = "low";

dffeas \x_3_imag_held[15] (
	.clk(clk),
	.d(\butterfly_st1[2][1][15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_imag_held[15]~q ),
	.prn(vcc));
defparam \x_3_imag_held[15] .is_wysiwyg = "true";
defparam \x_3_imag_held[15] .power_up = "low";

cycloneive_lcell_comb \Add6~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_imag_held[15]~q ),
	.cin(gnd),
	.combout(\Add6~4_combout ),
	.cout());
defparam \Add6~4 .lut_mask = 16'h0FF0;
defparam \Add6~4 .sum_lutc_input = "datac";

dffeas \x_1_imag_held[15] (
	.clk(clk),
	.d(\butterfly_st1[0][1][15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_imag_held[15]~q ),
	.prn(vcc));
defparam \x_1_imag_held[15] .is_wysiwyg = "true";
defparam \x_1_imag_held[15] .power_up = "low";

dffeas \x_3_imag_held[14] (
	.clk(clk),
	.d(\butterfly_st1[2][1][14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_imag_held[14]~q ),
	.prn(vcc));
defparam \x_3_imag_held[14] .is_wysiwyg = "true";
defparam \x_3_imag_held[14] .power_up = "low";

cycloneive_lcell_comb \Add6~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_imag_held[14]~q ),
	.cin(gnd),
	.combout(\Add6~5_combout ),
	.cout());
defparam \Add6~5 .lut_mask = 16'h0FF0;
defparam \Add6~5 .sum_lutc_input = "datac";

dffeas \x_1_imag_held[14] (
	.clk(clk),
	.d(\butterfly_st1[0][1][14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_imag_held[14]~q ),
	.prn(vcc));
defparam \x_1_imag_held[14] .is_wysiwyg = "true";
defparam \x_1_imag_held[14] .power_up = "low";

dffeas \x_3_imag_held[13] (
	.clk(clk),
	.d(\butterfly_st1[2][1][13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_imag_held[13]~q ),
	.prn(vcc));
defparam \x_3_imag_held[13] .is_wysiwyg = "true";
defparam \x_3_imag_held[13] .power_up = "low";

cycloneive_lcell_comb \Add6~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_imag_held[13]~q ),
	.cin(gnd),
	.combout(\Add6~6_combout ),
	.cout());
defparam \Add6~6 .lut_mask = 16'h0FF0;
defparam \Add6~6 .sum_lutc_input = "datac";

dffeas \x_1_imag_held[13] (
	.clk(clk),
	.d(\butterfly_st1[0][1][13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_imag_held[13]~q ),
	.prn(vcc));
defparam \x_1_imag_held[13] .is_wysiwyg = "true";
defparam \x_1_imag_held[13] .power_up = "low";

dffeas \x_3_imag_held[12] (
	.clk(clk),
	.d(\butterfly_st1[2][1][12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_imag_held[12]~q ),
	.prn(vcc));
defparam \x_3_imag_held[12] .is_wysiwyg = "true";
defparam \x_3_imag_held[12] .power_up = "low";

cycloneive_lcell_comb \Add6~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_imag_held[12]~q ),
	.cin(gnd),
	.combout(\Add6~7_combout ),
	.cout());
defparam \Add6~7 .lut_mask = 16'h0FF0;
defparam \Add6~7 .sum_lutc_input = "datac";

dffeas \x_1_imag_held[12] (
	.clk(clk),
	.d(\butterfly_st1[0][1][12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_imag_held[12]~q ),
	.prn(vcc));
defparam \x_1_imag_held[12] .is_wysiwyg = "true";
defparam \x_1_imag_held[12] .power_up = "low";

dffeas \x_3_imag_held[11] (
	.clk(clk),
	.d(\butterfly_st1[2][1][11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_imag_held[11]~q ),
	.prn(vcc));
defparam \x_3_imag_held[11] .is_wysiwyg = "true";
defparam \x_3_imag_held[11] .power_up = "low";

cycloneive_lcell_comb \Add6~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_imag_held[11]~q ),
	.cin(gnd),
	.combout(\Add6~8_combout ),
	.cout());
defparam \Add6~8 .lut_mask = 16'h0FF0;
defparam \Add6~8 .sum_lutc_input = "datac";

dffeas \x_1_imag_held[11] (
	.clk(clk),
	.d(\butterfly_st1[0][1][11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_imag_held[11]~q ),
	.prn(vcc));
defparam \x_1_imag_held[11] .is_wysiwyg = "true";
defparam \x_1_imag_held[11] .power_up = "low";

dffeas \x_3_imag_held[10] (
	.clk(clk),
	.d(\butterfly_st1[2][1][10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_imag_held[10]~q ),
	.prn(vcc));
defparam \x_3_imag_held[10] .is_wysiwyg = "true";
defparam \x_3_imag_held[10] .power_up = "low";

cycloneive_lcell_comb \Add6~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_imag_held[10]~q ),
	.cin(gnd),
	.combout(\Add6~9_combout ),
	.cout());
defparam \Add6~9 .lut_mask = 16'h0FF0;
defparam \Add6~9 .sum_lutc_input = "datac";

dffeas \x_1_imag_held[10] (
	.clk(clk),
	.d(\butterfly_st1[0][1][10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_imag_held[10]~q ),
	.prn(vcc));
defparam \x_1_imag_held[10] .is_wysiwyg = "true";
defparam \x_1_imag_held[10] .power_up = "low";

dffeas \x_3_imag_held[9] (
	.clk(clk),
	.d(\butterfly_st1[2][1][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_imag_held[9]~q ),
	.prn(vcc));
defparam \x_3_imag_held[9] .is_wysiwyg = "true";
defparam \x_3_imag_held[9] .power_up = "low";

cycloneive_lcell_comb \Add6~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_imag_held[9]~q ),
	.cin(gnd),
	.combout(\Add6~10_combout ),
	.cout());
defparam \Add6~10 .lut_mask = 16'h0FF0;
defparam \Add6~10 .sum_lutc_input = "datac";

dffeas \x_1_imag_held[9] (
	.clk(clk),
	.d(\butterfly_st1[0][1][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_imag_held[9]~q ),
	.prn(vcc));
defparam \x_1_imag_held[9] .is_wysiwyg = "true";
defparam \x_1_imag_held[9] .power_up = "low";

dffeas \x_3_imag_held[8] (
	.clk(clk),
	.d(\butterfly_st1[2][1][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_imag_held[8]~q ),
	.prn(vcc));
defparam \x_3_imag_held[8] .is_wysiwyg = "true";
defparam \x_3_imag_held[8] .power_up = "low";

cycloneive_lcell_comb \Add6~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_imag_held[8]~q ),
	.cin(gnd),
	.combout(\Add6~11_combout ),
	.cout());
defparam \Add6~11 .lut_mask = 16'h0FF0;
defparam \Add6~11 .sum_lutc_input = "datac";

dffeas \x_1_imag_held[8] (
	.clk(clk),
	.d(\butterfly_st1[0][1][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_imag_held[8]~q ),
	.prn(vcc));
defparam \x_1_imag_held[8] .is_wysiwyg = "true";
defparam \x_1_imag_held[8] .power_up = "low";

dffeas \x_3_imag_held[7] (
	.clk(clk),
	.d(\butterfly_st1[2][1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_imag_held[7]~q ),
	.prn(vcc));
defparam \x_3_imag_held[7] .is_wysiwyg = "true";
defparam \x_3_imag_held[7] .power_up = "low";

cycloneive_lcell_comb \Add6~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_imag_held[7]~q ),
	.cin(gnd),
	.combout(\Add6~12_combout ),
	.cout());
defparam \Add6~12 .lut_mask = 16'h0FF0;
defparam \Add6~12 .sum_lutc_input = "datac";

dffeas \x_1_imag_held[7] (
	.clk(clk),
	.d(\butterfly_st1[0][1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_imag_held[7]~q ),
	.prn(vcc));
defparam \x_1_imag_held[7] .is_wysiwyg = "true";
defparam \x_1_imag_held[7] .power_up = "low";

dffeas \x_3_imag_held[6] (
	.clk(clk),
	.d(\butterfly_st1[2][1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_imag_held[6]~q ),
	.prn(vcc));
defparam \x_3_imag_held[6] .is_wysiwyg = "true";
defparam \x_3_imag_held[6] .power_up = "low";

cycloneive_lcell_comb \Add6~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_imag_held[6]~q ),
	.cin(gnd),
	.combout(\Add6~13_combout ),
	.cout());
defparam \Add6~13 .lut_mask = 16'h0FF0;
defparam \Add6~13 .sum_lutc_input = "datac";

dffeas \x_1_imag_held[6] (
	.clk(clk),
	.d(\butterfly_st1[0][1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_imag_held[6]~q ),
	.prn(vcc));
defparam \x_1_imag_held[6] .is_wysiwyg = "true";
defparam \x_1_imag_held[6] .power_up = "low";

dffeas \x_3_imag_held[5] (
	.clk(clk),
	.d(\butterfly_st1[2][1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_imag_held[5]~q ),
	.prn(vcc));
defparam \x_3_imag_held[5] .is_wysiwyg = "true";
defparam \x_3_imag_held[5] .power_up = "low";

cycloneive_lcell_comb \Add6~14 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_imag_held[5]~q ),
	.cin(gnd),
	.combout(\Add6~14_combout ),
	.cout());
defparam \Add6~14 .lut_mask = 16'h0FF0;
defparam \Add6~14 .sum_lutc_input = "datac";

dffeas \x_1_imag_held[5] (
	.clk(clk),
	.d(\butterfly_st1[0][1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_imag_held[5]~q ),
	.prn(vcc));
defparam \x_1_imag_held[5] .is_wysiwyg = "true";
defparam \x_1_imag_held[5] .power_up = "low";

dffeas \x_3_imag_held[4] (
	.clk(clk),
	.d(\butterfly_st1[2][1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_imag_held[4]~q ),
	.prn(vcc));
defparam \x_3_imag_held[4] .is_wysiwyg = "true";
defparam \x_3_imag_held[4] .power_up = "low";

cycloneive_lcell_comb \Add6~15 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_imag_held[4]~q ),
	.cin(gnd),
	.combout(\Add6~15_combout ),
	.cout());
defparam \Add6~15 .lut_mask = 16'h0FF0;
defparam \Add6~15 .sum_lutc_input = "datac";

dffeas \x_1_imag_held[4] (
	.clk(clk),
	.d(\butterfly_st1[0][1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_imag_held[4]~q ),
	.prn(vcc));
defparam \x_1_imag_held[4] .is_wysiwyg = "true";
defparam \x_1_imag_held[4] .power_up = "low";

dffeas \x_3_imag_held[3] (
	.clk(clk),
	.d(\butterfly_st1[2][1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_imag_held[3]~q ),
	.prn(vcc));
defparam \x_3_imag_held[3] .is_wysiwyg = "true";
defparam \x_3_imag_held[3] .power_up = "low";

cycloneive_lcell_comb \Add6~16 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_imag_held[3]~q ),
	.cin(gnd),
	.combout(\Add6~16_combout ),
	.cout());
defparam \Add6~16 .lut_mask = 16'h0FF0;
defparam \Add6~16 .sum_lutc_input = "datac";

dffeas \x_1_imag_held[3] (
	.clk(clk),
	.d(\butterfly_st1[0][1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_imag_held[3]~q ),
	.prn(vcc));
defparam \x_1_imag_held[3] .is_wysiwyg = "true";
defparam \x_1_imag_held[3] .power_up = "low";

dffeas \sel_arr[9][0] (
	.clk(clk),
	.d(\sel_arr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[9][0]~q ),
	.prn(vcc));
defparam \sel_arr[9][0] .is_wysiwyg = "true";
defparam \sel_arr[9][0] .power_up = "low";

cycloneive_lcell_comb \Mux264~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux264~0_combout ),
	.cout());
defparam \Mux264~0 .lut_mask = 16'h0FF0;
defparam \Mux264~0 .sum_lutc_input = "datac";

dffeas \x_4_real_held[2] (
	.clk(clk),
	.d(\Mux193~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_real_held[2]~q ),
	.prn(vcc));
defparam \x_4_real_held[2] .is_wysiwyg = "true";
defparam \x_4_real_held[2] .power_up = "low";

cycloneive_lcell_comb \Add2~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_real_held[2]~q ),
	.cin(gnd),
	.combout(\Add2~1_combout ),
	.cout());
defparam \Add2~1 .lut_mask = 16'h0FF0;
defparam \Add2~1 .sum_lutc_input = "datac";

dffeas \x_2_real_held[2] (
	.clk(clk),
	.d(\Mux159~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_real_held[2]~q ),
	.prn(vcc));
defparam \x_2_real_held[2] .is_wysiwyg = "true";
defparam \x_2_real_held[2] .power_up = "low";

dffeas \x_4_real_held[1] (
	.clk(clk),
	.d(\Mux194~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_real_held[1]~q ),
	.prn(vcc));
defparam \x_4_real_held[1] .is_wysiwyg = "true";
defparam \x_4_real_held[1] .power_up = "low";

cycloneive_lcell_comb \Add2~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_real_held[1]~q ),
	.cin(gnd),
	.combout(\Add2~2_combout ),
	.cout());
defparam \Add2~2 .lut_mask = 16'h0FF0;
defparam \Add2~2 .sum_lutc_input = "datac";

dffeas \x_2_real_held[1] (
	.clk(clk),
	.d(\Mux160~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_real_held[1]~q ),
	.prn(vcc));
defparam \x_2_real_held[1] .is_wysiwyg = "true";
defparam \x_2_real_held[1] .power_up = "low";

dffeas \x_4_real_held[0] (
	.clk(clk),
	.d(\Mux195~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_real_held[0]~q ),
	.prn(vcc));
defparam \x_4_real_held[0] .is_wysiwyg = "true";
defparam \x_4_real_held[0] .power_up = "low";

cycloneive_lcell_comb \Add2~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_real_held[0]~q ),
	.cin(gnd),
	.combout(\Add2~3_combout ),
	.cout());
defparam \Add2~3 .lut_mask = 16'h0FF0;
defparam \Add2~3 .sum_lutc_input = "datac";

dffeas \x_2_real_held[0] (
	.clk(clk),
	.d(\Mux161~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_real_held[0]~q ),
	.prn(vcc));
defparam \x_2_real_held[0] .is_wysiwyg = "true";
defparam \x_2_real_held[0] .power_up = "low";

dffeas \x_3_real_held[2] (
	.clk(clk),
	.d(\butterfly_st1[2][0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_real_held[2]~q ),
	.prn(vcc));
defparam \x_3_real_held[2] .is_wysiwyg = "true";
defparam \x_3_real_held[2] .power_up = "low";

cycloneive_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_real_held[2]~q ),
	.cin(gnd),
	.combout(\Add0~1_combout ),
	.cout());
defparam \Add0~1 .lut_mask = 16'h0FF0;
defparam \Add0~1 .sum_lutc_input = "datac";

dffeas \x_1_real_held[2] (
	.clk(clk),
	.d(\butterfly_st1[0][0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_real_held[2]~q ),
	.prn(vcc));
defparam \x_1_real_held[2] .is_wysiwyg = "true";
defparam \x_1_real_held[2] .power_up = "low";

dffeas \x_3_real_held[1] (
	.clk(clk),
	.d(\butterfly_st1[2][0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_real_held[1]~q ),
	.prn(vcc));
defparam \x_3_real_held[1] .is_wysiwyg = "true";
defparam \x_3_real_held[1] .power_up = "low";

cycloneive_lcell_comb \Add0~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_real_held[1]~q ),
	.cin(gnd),
	.combout(\Add0~2_combout ),
	.cout());
defparam \Add0~2 .lut_mask = 16'h0FF0;
defparam \Add0~2 .sum_lutc_input = "datac";

dffeas \x_1_real_held[1] (
	.clk(clk),
	.d(\butterfly_st1[0][0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_real_held[1]~q ),
	.prn(vcc));
defparam \x_1_real_held[1] .is_wysiwyg = "true";
defparam \x_1_real_held[1] .power_up = "low";

dffeas \x_3_real_held[0] (
	.clk(clk),
	.d(\butterfly_st1[2][0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_real_held[0]~q ),
	.prn(vcc));
defparam \x_3_real_held[0] .is_wysiwyg = "true";
defparam \x_3_real_held[0] .power_up = "low";

cycloneive_lcell_comb \Add0~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_real_held[0]~q ),
	.cin(gnd),
	.combout(\Add0~3_combout ),
	.cout());
defparam \Add0~3 .lut_mask = 16'h0FF0;
defparam \Add0~3 .sum_lutc_input = "datac";

dffeas \x_1_real_held[0] (
	.clk(clk),
	.d(\butterfly_st1[0][0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_real_held[0]~q ),
	.prn(vcc));
defparam \x_1_real_held[0] .is_wysiwyg = "true";
defparam \x_1_real_held[0] .power_up = "low";

dffeas \x_4_real_held[15] (
	.clk(clk),
	.d(\Mux180~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_real_held[15]~q ),
	.prn(vcc));
defparam \x_4_real_held[15] .is_wysiwyg = "true";
defparam \x_4_real_held[15] .power_up = "low";

cycloneive_lcell_comb \Add2~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_real_held[15]~q ),
	.cin(gnd),
	.combout(\Add2~4_combout ),
	.cout());
defparam \Add2~4 .lut_mask = 16'h0FF0;
defparam \Add2~4 .sum_lutc_input = "datac";

dffeas \x_2_real_held[15] (
	.clk(clk),
	.d(\Mux146~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_real_held[15]~q ),
	.prn(vcc));
defparam \x_2_real_held[15] .is_wysiwyg = "true";
defparam \x_2_real_held[15] .power_up = "low";

dffeas \x_4_real_held[14] (
	.clk(clk),
	.d(\Mux181~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_real_held[14]~q ),
	.prn(vcc));
defparam \x_4_real_held[14] .is_wysiwyg = "true";
defparam \x_4_real_held[14] .power_up = "low";

cycloneive_lcell_comb \Add2~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_real_held[14]~q ),
	.cin(gnd),
	.combout(\Add2~5_combout ),
	.cout());
defparam \Add2~5 .lut_mask = 16'h0FF0;
defparam \Add2~5 .sum_lutc_input = "datac";

dffeas \x_2_real_held[14] (
	.clk(clk),
	.d(\Mux147~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_real_held[14]~q ),
	.prn(vcc));
defparam \x_2_real_held[14] .is_wysiwyg = "true";
defparam \x_2_real_held[14] .power_up = "low";

dffeas \x_4_real_held[13] (
	.clk(clk),
	.d(\Mux182~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_real_held[13]~q ),
	.prn(vcc));
defparam \x_4_real_held[13] .is_wysiwyg = "true";
defparam \x_4_real_held[13] .power_up = "low";

cycloneive_lcell_comb \Add2~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_real_held[13]~q ),
	.cin(gnd),
	.combout(\Add2~6_combout ),
	.cout());
defparam \Add2~6 .lut_mask = 16'h0FF0;
defparam \Add2~6 .sum_lutc_input = "datac";

dffeas \x_2_real_held[13] (
	.clk(clk),
	.d(\Mux148~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_real_held[13]~q ),
	.prn(vcc));
defparam \x_2_real_held[13] .is_wysiwyg = "true";
defparam \x_2_real_held[13] .power_up = "low";

dffeas \x_4_real_held[12] (
	.clk(clk),
	.d(\Mux183~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_real_held[12]~q ),
	.prn(vcc));
defparam \x_4_real_held[12] .is_wysiwyg = "true";
defparam \x_4_real_held[12] .power_up = "low";

cycloneive_lcell_comb \Add2~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_real_held[12]~q ),
	.cin(gnd),
	.combout(\Add2~7_combout ),
	.cout());
defparam \Add2~7 .lut_mask = 16'h0FF0;
defparam \Add2~7 .sum_lutc_input = "datac";

dffeas \x_2_real_held[12] (
	.clk(clk),
	.d(\Mux149~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_real_held[12]~q ),
	.prn(vcc));
defparam \x_2_real_held[12] .is_wysiwyg = "true";
defparam \x_2_real_held[12] .power_up = "low";

dffeas \x_4_real_held[11] (
	.clk(clk),
	.d(\Mux184~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_real_held[11]~q ),
	.prn(vcc));
defparam \x_4_real_held[11] .is_wysiwyg = "true";
defparam \x_4_real_held[11] .power_up = "low";

cycloneive_lcell_comb \Add2~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_real_held[11]~q ),
	.cin(gnd),
	.combout(\Add2~8_combout ),
	.cout());
defparam \Add2~8 .lut_mask = 16'h0FF0;
defparam \Add2~8 .sum_lutc_input = "datac";

dffeas \x_2_real_held[11] (
	.clk(clk),
	.d(\Mux150~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_real_held[11]~q ),
	.prn(vcc));
defparam \x_2_real_held[11] .is_wysiwyg = "true";
defparam \x_2_real_held[11] .power_up = "low";

dffeas \x_4_real_held[10] (
	.clk(clk),
	.d(\Mux185~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_real_held[10]~q ),
	.prn(vcc));
defparam \x_4_real_held[10] .is_wysiwyg = "true";
defparam \x_4_real_held[10] .power_up = "low";

cycloneive_lcell_comb \Add2~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_real_held[10]~q ),
	.cin(gnd),
	.combout(\Add2~9_combout ),
	.cout());
defparam \Add2~9 .lut_mask = 16'h0FF0;
defparam \Add2~9 .sum_lutc_input = "datac";

dffeas \x_2_real_held[10] (
	.clk(clk),
	.d(\Mux151~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_real_held[10]~q ),
	.prn(vcc));
defparam \x_2_real_held[10] .is_wysiwyg = "true";
defparam \x_2_real_held[10] .power_up = "low";

dffeas \x_4_real_held[9] (
	.clk(clk),
	.d(\Mux186~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_real_held[9]~q ),
	.prn(vcc));
defparam \x_4_real_held[9] .is_wysiwyg = "true";
defparam \x_4_real_held[9] .power_up = "low";

cycloneive_lcell_comb \Add2~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_real_held[9]~q ),
	.cin(gnd),
	.combout(\Add2~10_combout ),
	.cout());
defparam \Add2~10 .lut_mask = 16'h0FF0;
defparam \Add2~10 .sum_lutc_input = "datac";

dffeas \x_2_real_held[9] (
	.clk(clk),
	.d(\Mux152~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_real_held[9]~q ),
	.prn(vcc));
defparam \x_2_real_held[9] .is_wysiwyg = "true";
defparam \x_2_real_held[9] .power_up = "low";

dffeas \x_4_real_held[8] (
	.clk(clk),
	.d(\Mux187~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_real_held[8]~q ),
	.prn(vcc));
defparam \x_4_real_held[8] .is_wysiwyg = "true";
defparam \x_4_real_held[8] .power_up = "low";

cycloneive_lcell_comb \Add2~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_real_held[8]~q ),
	.cin(gnd),
	.combout(\Add2~11_combout ),
	.cout());
defparam \Add2~11 .lut_mask = 16'h0FF0;
defparam \Add2~11 .sum_lutc_input = "datac";

dffeas \x_2_real_held[8] (
	.clk(clk),
	.d(\Mux153~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_real_held[8]~q ),
	.prn(vcc));
defparam \x_2_real_held[8] .is_wysiwyg = "true";
defparam \x_2_real_held[8] .power_up = "low";

dffeas \x_4_real_held[7] (
	.clk(clk),
	.d(\Mux188~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_real_held[7]~q ),
	.prn(vcc));
defparam \x_4_real_held[7] .is_wysiwyg = "true";
defparam \x_4_real_held[7] .power_up = "low";

cycloneive_lcell_comb \Add2~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_real_held[7]~q ),
	.cin(gnd),
	.combout(\Add2~12_combout ),
	.cout());
defparam \Add2~12 .lut_mask = 16'h0FF0;
defparam \Add2~12 .sum_lutc_input = "datac";

dffeas \x_2_real_held[7] (
	.clk(clk),
	.d(\Mux154~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_real_held[7]~q ),
	.prn(vcc));
defparam \x_2_real_held[7] .is_wysiwyg = "true";
defparam \x_2_real_held[7] .power_up = "low";

dffeas \x_4_real_held[6] (
	.clk(clk),
	.d(\Mux189~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_real_held[6]~q ),
	.prn(vcc));
defparam \x_4_real_held[6] .is_wysiwyg = "true";
defparam \x_4_real_held[6] .power_up = "low";

cycloneive_lcell_comb \Add2~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_real_held[6]~q ),
	.cin(gnd),
	.combout(\Add2~13_combout ),
	.cout());
defparam \Add2~13 .lut_mask = 16'h0FF0;
defparam \Add2~13 .sum_lutc_input = "datac";

dffeas \x_2_real_held[6] (
	.clk(clk),
	.d(\Mux155~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_real_held[6]~q ),
	.prn(vcc));
defparam \x_2_real_held[6] .is_wysiwyg = "true";
defparam \x_2_real_held[6] .power_up = "low";

dffeas \x_4_real_held[5] (
	.clk(clk),
	.d(\Mux190~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_real_held[5]~q ),
	.prn(vcc));
defparam \x_4_real_held[5] .is_wysiwyg = "true";
defparam \x_4_real_held[5] .power_up = "low";

cycloneive_lcell_comb \Add2~14 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_real_held[5]~q ),
	.cin(gnd),
	.combout(\Add2~14_combout ),
	.cout());
defparam \Add2~14 .lut_mask = 16'h0FF0;
defparam \Add2~14 .sum_lutc_input = "datac";

dffeas \x_2_real_held[5] (
	.clk(clk),
	.d(\Mux156~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_real_held[5]~q ),
	.prn(vcc));
defparam \x_2_real_held[5] .is_wysiwyg = "true";
defparam \x_2_real_held[5] .power_up = "low";

dffeas \x_4_real_held[4] (
	.clk(clk),
	.d(\Mux191~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_real_held[4]~q ),
	.prn(vcc));
defparam \x_4_real_held[4] .is_wysiwyg = "true";
defparam \x_4_real_held[4] .power_up = "low";

cycloneive_lcell_comb \Add2~15 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_real_held[4]~q ),
	.cin(gnd),
	.combout(\Add2~15_combout ),
	.cout());
defparam \Add2~15 .lut_mask = 16'h0FF0;
defparam \Add2~15 .sum_lutc_input = "datac";

dffeas \x_2_real_held[4] (
	.clk(clk),
	.d(\Mux157~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_real_held[4]~q ),
	.prn(vcc));
defparam \x_2_real_held[4] .is_wysiwyg = "true";
defparam \x_2_real_held[4] .power_up = "low";

dffeas \x_4_real_held[3] (
	.clk(clk),
	.d(\Mux192~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_4_real_held[3]~q ),
	.prn(vcc));
defparam \x_4_real_held[3] .is_wysiwyg = "true";
defparam \x_4_real_held[3] .power_up = "low";

cycloneive_lcell_comb \Add2~16 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_4_real_held[3]~q ),
	.cin(gnd),
	.combout(\Add2~16_combout ),
	.cout());
defparam \Add2~16 .lut_mask = 16'h0FF0;
defparam \Add2~16 .sum_lutc_input = "datac";

dffeas \x_2_real_held[3] (
	.clk(clk),
	.d(\Mux158~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\x_2_real_held[3]~q ),
	.prn(vcc));
defparam \x_2_real_held[3] .is_wysiwyg = "true";
defparam \x_2_real_held[3] .power_up = "low";

dffeas \x_3_real_held[15] (
	.clk(clk),
	.d(\butterfly_st1[2][0][15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_real_held[15]~q ),
	.prn(vcc));
defparam \x_3_real_held[15] .is_wysiwyg = "true";
defparam \x_3_real_held[15] .power_up = "low";

cycloneive_lcell_comb \Add0~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_real_held[15]~q ),
	.cin(gnd),
	.combout(\Add0~4_combout ),
	.cout());
defparam \Add0~4 .lut_mask = 16'h0FF0;
defparam \Add0~4 .sum_lutc_input = "datac";

dffeas \x_1_real_held[15] (
	.clk(clk),
	.d(\butterfly_st1[0][0][15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_real_held[15]~q ),
	.prn(vcc));
defparam \x_1_real_held[15] .is_wysiwyg = "true";
defparam \x_1_real_held[15] .power_up = "low";

dffeas \x_3_real_held[14] (
	.clk(clk),
	.d(\butterfly_st1[2][0][14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_real_held[14]~q ),
	.prn(vcc));
defparam \x_3_real_held[14] .is_wysiwyg = "true";
defparam \x_3_real_held[14] .power_up = "low";

cycloneive_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_real_held[14]~q ),
	.cin(gnd),
	.combout(\Add0~5_combout ),
	.cout());
defparam \Add0~5 .lut_mask = 16'h0FF0;
defparam \Add0~5 .sum_lutc_input = "datac";

dffeas \x_1_real_held[14] (
	.clk(clk),
	.d(\butterfly_st1[0][0][14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_real_held[14]~q ),
	.prn(vcc));
defparam \x_1_real_held[14] .is_wysiwyg = "true";
defparam \x_1_real_held[14] .power_up = "low";

dffeas \x_3_real_held[13] (
	.clk(clk),
	.d(\butterfly_st1[2][0][13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_real_held[13]~q ),
	.prn(vcc));
defparam \x_3_real_held[13] .is_wysiwyg = "true";
defparam \x_3_real_held[13] .power_up = "low";

cycloneive_lcell_comb \Add0~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_real_held[13]~q ),
	.cin(gnd),
	.combout(\Add0~6_combout ),
	.cout());
defparam \Add0~6 .lut_mask = 16'h0FF0;
defparam \Add0~6 .sum_lutc_input = "datac";

dffeas \x_1_real_held[13] (
	.clk(clk),
	.d(\butterfly_st1[0][0][13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_real_held[13]~q ),
	.prn(vcc));
defparam \x_1_real_held[13] .is_wysiwyg = "true";
defparam \x_1_real_held[13] .power_up = "low";

dffeas \x_3_real_held[12] (
	.clk(clk),
	.d(\butterfly_st1[2][0][12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_real_held[12]~q ),
	.prn(vcc));
defparam \x_3_real_held[12] .is_wysiwyg = "true";
defparam \x_3_real_held[12] .power_up = "low";

cycloneive_lcell_comb \Add0~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_real_held[12]~q ),
	.cin(gnd),
	.combout(\Add0~7_combout ),
	.cout());
defparam \Add0~7 .lut_mask = 16'h0FF0;
defparam \Add0~7 .sum_lutc_input = "datac";

dffeas \x_1_real_held[12] (
	.clk(clk),
	.d(\butterfly_st1[0][0][12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_real_held[12]~q ),
	.prn(vcc));
defparam \x_1_real_held[12] .is_wysiwyg = "true";
defparam \x_1_real_held[12] .power_up = "low";

dffeas \x_3_real_held[11] (
	.clk(clk),
	.d(\butterfly_st1[2][0][11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_real_held[11]~q ),
	.prn(vcc));
defparam \x_3_real_held[11] .is_wysiwyg = "true";
defparam \x_3_real_held[11] .power_up = "low";

cycloneive_lcell_comb \Add0~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_real_held[11]~q ),
	.cin(gnd),
	.combout(\Add0~8_combout ),
	.cout());
defparam \Add0~8 .lut_mask = 16'h0FF0;
defparam \Add0~8 .sum_lutc_input = "datac";

dffeas \x_1_real_held[11] (
	.clk(clk),
	.d(\butterfly_st1[0][0][11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_real_held[11]~q ),
	.prn(vcc));
defparam \x_1_real_held[11] .is_wysiwyg = "true";
defparam \x_1_real_held[11] .power_up = "low";

dffeas \x_3_real_held[10] (
	.clk(clk),
	.d(\butterfly_st1[2][0][10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_real_held[10]~q ),
	.prn(vcc));
defparam \x_3_real_held[10] .is_wysiwyg = "true";
defparam \x_3_real_held[10] .power_up = "low";

cycloneive_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_real_held[10]~q ),
	.cin(gnd),
	.combout(\Add0~9_combout ),
	.cout());
defparam \Add0~9 .lut_mask = 16'h0FF0;
defparam \Add0~9 .sum_lutc_input = "datac";

dffeas \x_1_real_held[10] (
	.clk(clk),
	.d(\butterfly_st1[0][0][10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_real_held[10]~q ),
	.prn(vcc));
defparam \x_1_real_held[10] .is_wysiwyg = "true";
defparam \x_1_real_held[10] .power_up = "low";

dffeas \x_3_real_held[9] (
	.clk(clk),
	.d(\butterfly_st1[2][0][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_real_held[9]~q ),
	.prn(vcc));
defparam \x_3_real_held[9] .is_wysiwyg = "true";
defparam \x_3_real_held[9] .power_up = "low";

cycloneive_lcell_comb \Add0~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_real_held[9]~q ),
	.cin(gnd),
	.combout(\Add0~10_combout ),
	.cout());
defparam \Add0~10 .lut_mask = 16'h0FF0;
defparam \Add0~10 .sum_lutc_input = "datac";

dffeas \x_1_real_held[9] (
	.clk(clk),
	.d(\butterfly_st1[0][0][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_real_held[9]~q ),
	.prn(vcc));
defparam \x_1_real_held[9] .is_wysiwyg = "true";
defparam \x_1_real_held[9] .power_up = "low";

dffeas \x_3_real_held[8] (
	.clk(clk),
	.d(\butterfly_st1[2][0][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_real_held[8]~q ),
	.prn(vcc));
defparam \x_3_real_held[8] .is_wysiwyg = "true";
defparam \x_3_real_held[8] .power_up = "low";

cycloneive_lcell_comb \Add0~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_real_held[8]~q ),
	.cin(gnd),
	.combout(\Add0~11_combout ),
	.cout());
defparam \Add0~11 .lut_mask = 16'h0FF0;
defparam \Add0~11 .sum_lutc_input = "datac";

dffeas \x_1_real_held[8] (
	.clk(clk),
	.d(\butterfly_st1[0][0][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_real_held[8]~q ),
	.prn(vcc));
defparam \x_1_real_held[8] .is_wysiwyg = "true";
defparam \x_1_real_held[8] .power_up = "low";

dffeas \x_3_real_held[7] (
	.clk(clk),
	.d(\butterfly_st1[2][0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_real_held[7]~q ),
	.prn(vcc));
defparam \x_3_real_held[7] .is_wysiwyg = "true";
defparam \x_3_real_held[7] .power_up = "low";

cycloneive_lcell_comb \Add0~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_real_held[7]~q ),
	.cin(gnd),
	.combout(\Add0~12_combout ),
	.cout());
defparam \Add0~12 .lut_mask = 16'h0FF0;
defparam \Add0~12 .sum_lutc_input = "datac";

dffeas \x_1_real_held[7] (
	.clk(clk),
	.d(\butterfly_st1[0][0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_real_held[7]~q ),
	.prn(vcc));
defparam \x_1_real_held[7] .is_wysiwyg = "true";
defparam \x_1_real_held[7] .power_up = "low";

dffeas \x_3_real_held[6] (
	.clk(clk),
	.d(\butterfly_st1[2][0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_real_held[6]~q ),
	.prn(vcc));
defparam \x_3_real_held[6] .is_wysiwyg = "true";
defparam \x_3_real_held[6] .power_up = "low";

cycloneive_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_real_held[6]~q ),
	.cin(gnd),
	.combout(\Add0~13_combout ),
	.cout());
defparam \Add0~13 .lut_mask = 16'h0FF0;
defparam \Add0~13 .sum_lutc_input = "datac";

dffeas \x_1_real_held[6] (
	.clk(clk),
	.d(\butterfly_st1[0][0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_real_held[6]~q ),
	.prn(vcc));
defparam \x_1_real_held[6] .is_wysiwyg = "true";
defparam \x_1_real_held[6] .power_up = "low";

dffeas \x_3_real_held[5] (
	.clk(clk),
	.d(\butterfly_st1[2][0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_real_held[5]~q ),
	.prn(vcc));
defparam \x_3_real_held[5] .is_wysiwyg = "true";
defparam \x_3_real_held[5] .power_up = "low";

cycloneive_lcell_comb \Add0~14 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_real_held[5]~q ),
	.cin(gnd),
	.combout(\Add0~14_combout ),
	.cout());
defparam \Add0~14 .lut_mask = 16'h0FF0;
defparam \Add0~14 .sum_lutc_input = "datac";

dffeas \x_1_real_held[5] (
	.clk(clk),
	.d(\butterfly_st1[0][0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_real_held[5]~q ),
	.prn(vcc));
defparam \x_1_real_held[5] .is_wysiwyg = "true";
defparam \x_1_real_held[5] .power_up = "low";

dffeas \x_3_real_held[4] (
	.clk(clk),
	.d(\butterfly_st1[2][0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_real_held[4]~q ),
	.prn(vcc));
defparam \x_3_real_held[4] .is_wysiwyg = "true";
defparam \x_3_real_held[4] .power_up = "low";

cycloneive_lcell_comb \Add0~15 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_real_held[4]~q ),
	.cin(gnd),
	.combout(\Add0~15_combout ),
	.cout());
defparam \Add0~15 .lut_mask = 16'h0FF0;
defparam \Add0~15 .sum_lutc_input = "datac";

dffeas \x_1_real_held[4] (
	.clk(clk),
	.d(\butterfly_st1[0][0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_real_held[4]~q ),
	.prn(vcc));
defparam \x_1_real_held[4] .is_wysiwyg = "true";
defparam \x_1_real_held[4] .power_up = "low";

dffeas \x_3_real_held[3] (
	.clk(clk),
	.d(\butterfly_st1[2][0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_3_real_held[3]~q ),
	.prn(vcc));
defparam \x_3_real_held[3] .is_wysiwyg = "true";
defparam \x_3_real_held[3] .power_up = "low";

cycloneive_lcell_comb \Add0~16 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\si[1]~q ),
	.datad(\x_3_real_held[3]~q ),
	.cin(gnd),
	.combout(\Add0~16_combout ),
	.cout());
defparam \Add0~16 .lut_mask = 16'h0FF0;
defparam \Add0~16 .sum_lutc_input = "datac";

dffeas \x_1_real_held[3] (
	.clk(clk),
	.d(\butterfly_st1[0][0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\x_3_imag_held[0]~0_combout ),
	.q(\x_1_real_held[3]~q ),
	.prn(vcc));
defparam \x_1_real_held[3] .is_wysiwyg = "true";
defparam \x_1_real_held[3] .power_up = "low";

dffeas \sel_arr[8][1] (
	.clk(clk),
	.d(\sel_arr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[8][1]~q ),
	.prn(vcc));
defparam \sel_arr[8][1] .is_wysiwyg = "true";
defparam \sel_arr[8][1] .power_up = "low";

cycloneive_lcell_comb \sel_arr~0 (
	.dataa(reset),
	.datab(\sel_arr[8][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~0_combout ),
	.cout());
defparam \sel_arr~0 .lut_mask = 16'hEEEE;
defparam \sel_arr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \si~1 (
	.dataa(\sel_arr[9][0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset),
	.cin(gnd),
	.combout(\si~1_combout ),
	.cout());
defparam \si~1 .lut_mask = 16'hFF55;
defparam \si~1 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][1][2] (
	.clk(clk),
	.d(\butterfly_st1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][2] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][2] .power_up = "low";

cycloneive_lcell_comb \Mux261~0 (
	.dataa(\x_4_real_held[2]~q ),
	.datab(\butterfly_st1[3][1][2]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux261~0_combout ),
	.cout());
defparam \Mux261~0 .lut_mask = 16'hEFFE;
defparam \Mux261~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][1][2] (
	.clk(clk),
	.d(\butterfly_st1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][2] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][2] .power_up = "low";

cycloneive_lcell_comb \Mux227~0 (
	.dataa(\x_2_real_held[2]~q ),
	.datab(\butterfly_st1[1][1][2]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux227~0_combout ),
	.cout());
defparam \Mux227~0 .lut_mask = 16'hEFFE;
defparam \Mux227~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][1][1] (
	.clk(clk),
	.d(\butterfly_st1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][1] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][1] .power_up = "low";

cycloneive_lcell_comb \Mux262~0 (
	.dataa(\x_4_real_held[1]~q ),
	.datab(\butterfly_st1[3][1][1]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux262~0_combout ),
	.cout());
defparam \Mux262~0 .lut_mask = 16'hEFFE;
defparam \Mux262~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][1][1] (
	.clk(clk),
	.d(\butterfly_st1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][1] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][1] .power_up = "low";

cycloneive_lcell_comb \Mux228~0 (
	.dataa(\x_2_real_held[1]~q ),
	.datab(\butterfly_st1[1][1][1]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux228~0_combout ),
	.cout());
defparam \Mux228~0 .lut_mask = 16'hEFFE;
defparam \Mux228~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][1][0] (
	.clk(clk),
	.d(\butterfly_st1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][0] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][0] .power_up = "low";

cycloneive_lcell_comb \Mux263~0 (
	.dataa(\x_4_real_held[0]~q ),
	.datab(\butterfly_st1[3][1][0]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux263~0_combout ),
	.cout());
defparam \Mux263~0 .lut_mask = 16'hEFFE;
defparam \Mux263~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][1][0] (
	.clk(clk),
	.d(\butterfly_st1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][0] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][0] .power_up = "low";

cycloneive_lcell_comb \Mux229~0 (
	.dataa(\x_2_real_held[0]~q ),
	.datab(\butterfly_st1[1][1][0]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux229~0_combout ),
	.cout());
defparam \Mux229~0 .lut_mask = 16'hEFFE;
defparam \Mux229~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[2][1][2] (
	.clk(clk),
	.d(\butterfly_st1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][2] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][2] .power_up = "low";

cycloneive_lcell_comb \x_3_imag_held[0]~0 (
	.dataa(global_clock_enable),
	.datab(\sel_arr[9][1]~q ),
	.datac(\sel_arr[9][0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\x_3_imag_held[0]~0_combout ),
	.cout());
defparam \x_3_imag_held[0]~0 .lut_mask = 16'hBFBF;
defparam \x_3_imag_held[0]~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[0][1][2] (
	.clk(clk),
	.d(\butterfly_st1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][2] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][2] .power_up = "low";

dffeas \butterfly_st1[2][1][1] (
	.clk(clk),
	.d(\butterfly_st1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][1] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][1] .power_up = "low";

dffeas \butterfly_st1[0][1][1] (
	.clk(clk),
	.d(\butterfly_st1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][1] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][1] .power_up = "low";

dffeas \butterfly_st1[2][1][0] (
	.clk(clk),
	.d(\butterfly_st1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][0] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][0] .power_up = "low";

dffeas \butterfly_st1[0][1][0] (
	.clk(clk),
	.d(\butterfly_st1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][0] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][0] .power_up = "low";

dffeas \butterfly_st1[3][1][15] (
	.clk(clk),
	.d(\butterfly_st1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][1][15]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][15] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][15] .power_up = "low";

cycloneive_lcell_comb \Mux248~0 (
	.dataa(\x_4_real_held[15]~q ),
	.datab(\butterfly_st1[3][1][15]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux248~0_combout ),
	.cout());
defparam \Mux248~0 .lut_mask = 16'hEFFE;
defparam \Mux248~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][1][15] (
	.clk(clk),
	.d(\butterfly_st1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][1][15]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][15] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][15] .power_up = "low";

cycloneive_lcell_comb \Mux214~0 (
	.dataa(\x_2_real_held[15]~q ),
	.datab(\butterfly_st1[1][1][15]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux214~0_combout ),
	.cout());
defparam \Mux214~0 .lut_mask = 16'hEFFE;
defparam \Mux214~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][1][14] (
	.clk(clk),
	.d(\butterfly_st1~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][1][14]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][14] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][14] .power_up = "low";

cycloneive_lcell_comb \Mux249~0 (
	.dataa(\x_4_real_held[14]~q ),
	.datab(\butterfly_st1[3][1][14]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux249~0_combout ),
	.cout());
defparam \Mux249~0 .lut_mask = 16'hEFFE;
defparam \Mux249~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][1][14] (
	.clk(clk),
	.d(\butterfly_st1~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][1][14]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][14] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][14] .power_up = "low";

cycloneive_lcell_comb \Mux215~0 (
	.dataa(\x_2_real_held[14]~q ),
	.datab(\butterfly_st1[1][1][14]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux215~0_combout ),
	.cout());
defparam \Mux215~0 .lut_mask = 16'hEFFE;
defparam \Mux215~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][1][13] (
	.clk(clk),
	.d(\butterfly_st1~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][1][13]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][13] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][13] .power_up = "low";

cycloneive_lcell_comb \Mux250~0 (
	.dataa(\x_4_real_held[13]~q ),
	.datab(\butterfly_st1[3][1][13]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux250~0_combout ),
	.cout());
defparam \Mux250~0 .lut_mask = 16'hEFFE;
defparam \Mux250~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][1][13] (
	.clk(clk),
	.d(\butterfly_st1~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][1][13]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][13] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][13] .power_up = "low";

cycloneive_lcell_comb \Mux216~0 (
	.dataa(\x_2_real_held[13]~q ),
	.datab(\butterfly_st1[1][1][13]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux216~0_combout ),
	.cout());
defparam \Mux216~0 .lut_mask = 16'hEFFE;
defparam \Mux216~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][1][12] (
	.clk(clk),
	.d(\butterfly_st1~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][1][12]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][12] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][12] .power_up = "low";

cycloneive_lcell_comb \Mux251~0 (
	.dataa(\x_4_real_held[12]~q ),
	.datab(\butterfly_st1[3][1][12]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux251~0_combout ),
	.cout());
defparam \Mux251~0 .lut_mask = 16'hEFFE;
defparam \Mux251~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][1][12] (
	.clk(clk),
	.d(\butterfly_st1~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][1][12]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][12] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][12] .power_up = "low";

cycloneive_lcell_comb \Mux217~0 (
	.dataa(\x_2_real_held[12]~q ),
	.datab(\butterfly_st1[1][1][12]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux217~0_combout ),
	.cout());
defparam \Mux217~0 .lut_mask = 16'hEFFE;
defparam \Mux217~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][1][11] (
	.clk(clk),
	.d(\butterfly_st1~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][1][11]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][11] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][11] .power_up = "low";

cycloneive_lcell_comb \Mux252~0 (
	.dataa(\x_4_real_held[11]~q ),
	.datab(\butterfly_st1[3][1][11]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux252~0_combout ),
	.cout());
defparam \Mux252~0 .lut_mask = 16'hEFFE;
defparam \Mux252~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][1][11] (
	.clk(clk),
	.d(\butterfly_st1~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][1][11]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][11] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][11] .power_up = "low";

cycloneive_lcell_comb \Mux218~0 (
	.dataa(\x_2_real_held[11]~q ),
	.datab(\butterfly_st1[1][1][11]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux218~0_combout ),
	.cout());
defparam \Mux218~0 .lut_mask = 16'hEFFE;
defparam \Mux218~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][1][10] (
	.clk(clk),
	.d(\butterfly_st1~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][1][10]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][10] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][10] .power_up = "low";

cycloneive_lcell_comb \Mux253~0 (
	.dataa(\x_4_real_held[10]~q ),
	.datab(\butterfly_st1[3][1][10]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux253~0_combout ),
	.cout());
defparam \Mux253~0 .lut_mask = 16'hEFFE;
defparam \Mux253~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][1][10] (
	.clk(clk),
	.d(\butterfly_st1~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][1][10]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][10] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][10] .power_up = "low";

cycloneive_lcell_comb \Mux219~0 (
	.dataa(\x_2_real_held[10]~q ),
	.datab(\butterfly_st1[1][1][10]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux219~0_combout ),
	.cout());
defparam \Mux219~0 .lut_mask = 16'hEFFE;
defparam \Mux219~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][1][9] (
	.clk(clk),
	.d(\butterfly_st1~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][9] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][9] .power_up = "low";

cycloneive_lcell_comb \Mux254~0 (
	.dataa(\x_4_real_held[9]~q ),
	.datab(\butterfly_st1[3][1][9]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux254~0_combout ),
	.cout());
defparam \Mux254~0 .lut_mask = 16'hEFFE;
defparam \Mux254~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][1][9] (
	.clk(clk),
	.d(\butterfly_st1~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][9] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][9] .power_up = "low";

cycloneive_lcell_comb \Mux220~0 (
	.dataa(\x_2_real_held[9]~q ),
	.datab(\butterfly_st1[1][1][9]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux220~0_combout ),
	.cout());
defparam \Mux220~0 .lut_mask = 16'hEFFE;
defparam \Mux220~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][1][8] (
	.clk(clk),
	.d(\butterfly_st1~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][8] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][8] .power_up = "low";

cycloneive_lcell_comb \Mux255~0 (
	.dataa(\x_4_real_held[8]~q ),
	.datab(\butterfly_st1[3][1][8]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux255~0_combout ),
	.cout());
defparam \Mux255~0 .lut_mask = 16'hEFFE;
defparam \Mux255~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][1][8] (
	.clk(clk),
	.d(\butterfly_st1~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][8] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][8] .power_up = "low";

cycloneive_lcell_comb \Mux221~0 (
	.dataa(\x_2_real_held[8]~q ),
	.datab(\butterfly_st1[1][1][8]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux221~0_combout ),
	.cout());
defparam \Mux221~0 .lut_mask = 16'hEFFE;
defparam \Mux221~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][1][7] (
	.clk(clk),
	.d(\butterfly_st1~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][7] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][7] .power_up = "low";

cycloneive_lcell_comb \Mux256~0 (
	.dataa(\x_4_real_held[7]~q ),
	.datab(\butterfly_st1[3][1][7]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux256~0_combout ),
	.cout());
defparam \Mux256~0 .lut_mask = 16'hEFFE;
defparam \Mux256~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][1][7] (
	.clk(clk),
	.d(\butterfly_st1~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][7] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][7] .power_up = "low";

cycloneive_lcell_comb \Mux222~0 (
	.dataa(\x_2_real_held[7]~q ),
	.datab(\butterfly_st1[1][1][7]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux222~0_combout ),
	.cout());
defparam \Mux222~0 .lut_mask = 16'hEFFE;
defparam \Mux222~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][1][6] (
	.clk(clk),
	.d(\butterfly_st1~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][6] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][6] .power_up = "low";

cycloneive_lcell_comb \Mux257~0 (
	.dataa(\x_4_real_held[6]~q ),
	.datab(\butterfly_st1[3][1][6]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux257~0_combout ),
	.cout());
defparam \Mux257~0 .lut_mask = 16'hEFFE;
defparam \Mux257~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][1][6] (
	.clk(clk),
	.d(\butterfly_st1~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][6] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][6] .power_up = "low";

cycloneive_lcell_comb \Mux223~0 (
	.dataa(\x_2_real_held[6]~q ),
	.datab(\butterfly_st1[1][1][6]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux223~0_combout ),
	.cout());
defparam \Mux223~0 .lut_mask = 16'hEFFE;
defparam \Mux223~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][1][5] (
	.clk(clk),
	.d(\butterfly_st1~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][5] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][5] .power_up = "low";

cycloneive_lcell_comb \Mux258~0 (
	.dataa(\x_4_real_held[5]~q ),
	.datab(\butterfly_st1[3][1][5]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux258~0_combout ),
	.cout());
defparam \Mux258~0 .lut_mask = 16'hEFFE;
defparam \Mux258~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][1][5] (
	.clk(clk),
	.d(\butterfly_st1~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][5] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][5] .power_up = "low";

cycloneive_lcell_comb \Mux224~0 (
	.dataa(\x_2_real_held[5]~q ),
	.datab(\butterfly_st1[1][1][5]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux224~0_combout ),
	.cout());
defparam \Mux224~0 .lut_mask = 16'hEFFE;
defparam \Mux224~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][1][4] (
	.clk(clk),
	.d(\butterfly_st1~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][4] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][4] .power_up = "low";

cycloneive_lcell_comb \Mux259~0 (
	.dataa(\x_4_real_held[4]~q ),
	.datab(\butterfly_st1[3][1][4]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux259~0_combout ),
	.cout());
defparam \Mux259~0 .lut_mask = 16'hEFFE;
defparam \Mux259~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][1][4] (
	.clk(clk),
	.d(\butterfly_st1~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][4] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][4] .power_up = "low";

cycloneive_lcell_comb \Mux225~0 (
	.dataa(\x_2_real_held[4]~q ),
	.datab(\butterfly_st1[1][1][4]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux225~0_combout ),
	.cout());
defparam \Mux225~0 .lut_mask = 16'hEFFE;
defparam \Mux225~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][1][3] (
	.clk(clk),
	.d(\butterfly_st1~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][3] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][3] .power_up = "low";

cycloneive_lcell_comb \Mux260~0 (
	.dataa(\x_4_real_held[3]~q ),
	.datab(\butterfly_st1[3][1][3]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux260~0_combout ),
	.cout());
defparam \Mux260~0 .lut_mask = 16'hEFFE;
defparam \Mux260~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][1][3] (
	.clk(clk),
	.d(\butterfly_st1~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][3] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][3] .power_up = "low";

cycloneive_lcell_comb \Mux226~0 (
	.dataa(\x_2_real_held[3]~q ),
	.datab(\butterfly_st1[1][1][3]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux226~0_combout ),
	.cout());
defparam \Mux226~0 .lut_mask = 16'hEFFE;
defparam \Mux226~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[2][1][15] (
	.clk(clk),
	.d(\butterfly_st1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][1][15]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][15] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][15] .power_up = "low";

dffeas \butterfly_st1[0][1][15] (
	.clk(clk),
	.d(\butterfly_st1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][1][15]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][15] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][15] .power_up = "low";

dffeas \butterfly_st1[2][1][14] (
	.clk(clk),
	.d(\butterfly_st1~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][1][14]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][14] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][14] .power_up = "low";

dffeas \butterfly_st1[0][1][14] (
	.clk(clk),
	.d(\butterfly_st1~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][1][14]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][14] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][14] .power_up = "low";

dffeas \butterfly_st1[2][1][13] (
	.clk(clk),
	.d(\butterfly_st1~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][1][13]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][13] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][13] .power_up = "low";

dffeas \butterfly_st1[0][1][13] (
	.clk(clk),
	.d(\butterfly_st1~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][1][13]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][13] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][13] .power_up = "low";

dffeas \butterfly_st1[2][1][12] (
	.clk(clk),
	.d(\butterfly_st1~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][1][12]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][12] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][12] .power_up = "low";

dffeas \butterfly_st1[0][1][12] (
	.clk(clk),
	.d(\butterfly_st1~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][1][12]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][12] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][12] .power_up = "low";

dffeas \butterfly_st1[2][1][11] (
	.clk(clk),
	.d(\butterfly_st1~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][1][11]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][11] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][11] .power_up = "low";

dffeas \butterfly_st1[0][1][11] (
	.clk(clk),
	.d(\butterfly_st1~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][1][11]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][11] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][11] .power_up = "low";

dffeas \butterfly_st1[2][1][10] (
	.clk(clk),
	.d(\butterfly_st1~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][1][10]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][10] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][10] .power_up = "low";

dffeas \butterfly_st1[0][1][10] (
	.clk(clk),
	.d(\butterfly_st1~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][1][10]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][10] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][10] .power_up = "low";

dffeas \butterfly_st1[2][1][9] (
	.clk(clk),
	.d(\butterfly_st1~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][9] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][9] .power_up = "low";

dffeas \butterfly_st1[0][1][9] (
	.clk(clk),
	.d(\butterfly_st1~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][9] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][9] .power_up = "low";

dffeas \butterfly_st1[2][1][8] (
	.clk(clk),
	.d(\butterfly_st1~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][8] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][8] .power_up = "low";

dffeas \butterfly_st1[0][1][8] (
	.clk(clk),
	.d(\butterfly_st1~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][8] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][8] .power_up = "low";

dffeas \butterfly_st1[2][1][7] (
	.clk(clk),
	.d(\butterfly_st1~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][7] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][7] .power_up = "low";

dffeas \butterfly_st1[0][1][7] (
	.clk(clk),
	.d(\butterfly_st1~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][7] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][7] .power_up = "low";

dffeas \butterfly_st1[2][1][6] (
	.clk(clk),
	.d(\butterfly_st1~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][6] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][6] .power_up = "low";

dffeas \butterfly_st1[0][1][6] (
	.clk(clk),
	.d(\butterfly_st1~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][6] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][6] .power_up = "low";

dffeas \butterfly_st1[2][1][5] (
	.clk(clk),
	.d(\butterfly_st1~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][5] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][5] .power_up = "low";

dffeas \butterfly_st1[0][1][5] (
	.clk(clk),
	.d(\butterfly_st1~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][5] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][5] .power_up = "low";

dffeas \butterfly_st1[2][1][4] (
	.clk(clk),
	.d(\butterfly_st1~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][4] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][4] .power_up = "low";

dffeas \butterfly_st1[0][1][4] (
	.clk(clk),
	.d(\butterfly_st1~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][4] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][4] .power_up = "low";

dffeas \butterfly_st1[2][1][3] (
	.clk(clk),
	.d(\butterfly_st1~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][3] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][3] .power_up = "low";

dffeas \butterfly_st1[0][1][3] (
	.clk(clk),
	.d(\butterfly_st1~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][3] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][3] .power_up = "low";

dffeas \sel_arr[8][0] (
	.clk(clk),
	.d(\sel_arr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[8][0]~q ),
	.prn(vcc));
defparam \sel_arr[8][0] .is_wysiwyg = "true";
defparam \sel_arr[8][0] .power_up = "low";

cycloneive_lcell_comb \sel_arr~1 (
	.dataa(reset),
	.datab(\sel_arr[8][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~1_combout ),
	.cout());
defparam \sel_arr~1 .lut_mask = 16'hEEEE;
defparam \sel_arr~1 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][0][2] (
	.clk(clk),
	.d(\butterfly_st1~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][2] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][2] .power_up = "low";

cycloneive_lcell_comb \Mux193~0 (
	.dataa(\x_4_imag_held[2]~q ),
	.datab(\butterfly_st1[3][0][2]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux193~0_combout ),
	.cout());
defparam \Mux193~0 .lut_mask = 16'hEFFE;
defparam \Mux193~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][0][2] (
	.clk(clk),
	.d(\butterfly_st1~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][2] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][2] .power_up = "low";

cycloneive_lcell_comb \Mux159~0 (
	.dataa(\x_2_imag_held[2]~q ),
	.datab(\butterfly_st1[1][0][2]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux159~0_combout ),
	.cout());
defparam \Mux159~0 .lut_mask = 16'hEFFE;
defparam \Mux159~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][0][1] (
	.clk(clk),
	.d(\butterfly_st1~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][1] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][1] .power_up = "low";

cycloneive_lcell_comb \Mux194~0 (
	.dataa(\x_4_imag_held[1]~q ),
	.datab(\butterfly_st1[3][0][1]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux194~0_combout ),
	.cout());
defparam \Mux194~0 .lut_mask = 16'hEFFE;
defparam \Mux194~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][0][1] (
	.clk(clk),
	.d(\butterfly_st1~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][1] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][1] .power_up = "low";

cycloneive_lcell_comb \Mux160~0 (
	.dataa(\x_2_imag_held[1]~q ),
	.datab(\butterfly_st1[1][0][1]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux160~0_combout ),
	.cout());
defparam \Mux160~0 .lut_mask = 16'hEFFE;
defparam \Mux160~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][0][0] (
	.clk(clk),
	.d(\butterfly_st1~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][0] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][0] .power_up = "low";

cycloneive_lcell_comb \Mux195~0 (
	.dataa(\x_4_imag_held[0]~q ),
	.datab(\butterfly_st1[3][0][0]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux195~0_combout ),
	.cout());
defparam \Mux195~0 .lut_mask = 16'hEFFE;
defparam \Mux195~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][0][0] (
	.clk(clk),
	.d(\butterfly_st1~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][0] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][0] .power_up = "low";

cycloneive_lcell_comb \Mux161~0 (
	.dataa(\x_2_imag_held[0]~q ),
	.datab(\butterfly_st1[1][0][0]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux161~0_combout ),
	.cout());
defparam \Mux161~0 .lut_mask = 16'hEFFE;
defparam \Mux161~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[2][0][2] (
	.clk(clk),
	.d(\butterfly_st1~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][2] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][2] .power_up = "low";

dffeas \butterfly_st1[0][0][2] (
	.clk(clk),
	.d(\butterfly_st1~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][2] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][2] .power_up = "low";

dffeas \butterfly_st1[2][0][1] (
	.clk(clk),
	.d(\butterfly_st1~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][1] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][1] .power_up = "low";

dffeas \butterfly_st1[0][0][1] (
	.clk(clk),
	.d(\butterfly_st1~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][1] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][1] .power_up = "low";

dffeas \butterfly_st1[2][0][0] (
	.clk(clk),
	.d(\butterfly_st1~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][0] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][0] .power_up = "low";

dffeas \butterfly_st1[0][0][0] (
	.clk(clk),
	.d(\butterfly_st1~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][0] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][0] .power_up = "low";

dffeas \butterfly_st1[3][0][15] (
	.clk(clk),
	.d(\butterfly_st1~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][0][15]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][15] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][15] .power_up = "low";

cycloneive_lcell_comb \Mux180~0 (
	.dataa(\x_4_imag_held[15]~q ),
	.datab(\butterfly_st1[3][0][15]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux180~0_combout ),
	.cout());
defparam \Mux180~0 .lut_mask = 16'hEFFE;
defparam \Mux180~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][0][15] (
	.clk(clk),
	.d(\butterfly_st1~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][0][15]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][15] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][15] .power_up = "low";

cycloneive_lcell_comb \Mux146~0 (
	.dataa(\x_2_imag_held[15]~q ),
	.datab(\butterfly_st1[1][0][15]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux146~0_combout ),
	.cout());
defparam \Mux146~0 .lut_mask = 16'hEFFE;
defparam \Mux146~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][0][14] (
	.clk(clk),
	.d(\butterfly_st1~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][0][14]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][14] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][14] .power_up = "low";

cycloneive_lcell_comb \Mux181~0 (
	.dataa(\x_4_imag_held[14]~q ),
	.datab(\butterfly_st1[3][0][14]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux181~0_combout ),
	.cout());
defparam \Mux181~0 .lut_mask = 16'hEFFE;
defparam \Mux181~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][0][14] (
	.clk(clk),
	.d(\butterfly_st1~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][0][14]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][14] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][14] .power_up = "low";

cycloneive_lcell_comb \Mux147~0 (
	.dataa(\x_2_imag_held[14]~q ),
	.datab(\butterfly_st1[1][0][14]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux147~0_combout ),
	.cout());
defparam \Mux147~0 .lut_mask = 16'hEFFE;
defparam \Mux147~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][0][13] (
	.clk(clk),
	.d(\butterfly_st1~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][0][13]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][13] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][13] .power_up = "low";

cycloneive_lcell_comb \Mux182~0 (
	.dataa(\x_4_imag_held[13]~q ),
	.datab(\butterfly_st1[3][0][13]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux182~0_combout ),
	.cout());
defparam \Mux182~0 .lut_mask = 16'hEFFE;
defparam \Mux182~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][0][13] (
	.clk(clk),
	.d(\butterfly_st1~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][0][13]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][13] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][13] .power_up = "low";

cycloneive_lcell_comb \Mux148~0 (
	.dataa(\x_2_imag_held[13]~q ),
	.datab(\butterfly_st1[1][0][13]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux148~0_combout ),
	.cout());
defparam \Mux148~0 .lut_mask = 16'hEFFE;
defparam \Mux148~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][0][12] (
	.clk(clk),
	.d(\butterfly_st1~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][0][12]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][12] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][12] .power_up = "low";

cycloneive_lcell_comb \Mux183~0 (
	.dataa(\x_4_imag_held[12]~q ),
	.datab(\butterfly_st1[3][0][12]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux183~0_combout ),
	.cout());
defparam \Mux183~0 .lut_mask = 16'hEFFE;
defparam \Mux183~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][0][12] (
	.clk(clk),
	.d(\butterfly_st1~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][0][12]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][12] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][12] .power_up = "low";

cycloneive_lcell_comb \Mux149~0 (
	.dataa(\x_2_imag_held[12]~q ),
	.datab(\butterfly_st1[1][0][12]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux149~0_combout ),
	.cout());
defparam \Mux149~0 .lut_mask = 16'hEFFE;
defparam \Mux149~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][0][11] (
	.clk(clk),
	.d(\butterfly_st1~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][0][11]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][11] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][11] .power_up = "low";

cycloneive_lcell_comb \Mux184~0 (
	.dataa(\x_4_imag_held[11]~q ),
	.datab(\butterfly_st1[3][0][11]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux184~0_combout ),
	.cout());
defparam \Mux184~0 .lut_mask = 16'hEFFE;
defparam \Mux184~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][0][11] (
	.clk(clk),
	.d(\butterfly_st1~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][0][11]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][11] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][11] .power_up = "low";

cycloneive_lcell_comb \Mux150~0 (
	.dataa(\x_2_imag_held[11]~q ),
	.datab(\butterfly_st1[1][0][11]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux150~0_combout ),
	.cout());
defparam \Mux150~0 .lut_mask = 16'hEFFE;
defparam \Mux150~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][0][10] (
	.clk(clk),
	.d(\butterfly_st1~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][0][10]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][10] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][10] .power_up = "low";

cycloneive_lcell_comb \Mux185~0 (
	.dataa(\x_4_imag_held[10]~q ),
	.datab(\butterfly_st1[3][0][10]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux185~0_combout ),
	.cout());
defparam \Mux185~0 .lut_mask = 16'hEFFE;
defparam \Mux185~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][0][10] (
	.clk(clk),
	.d(\butterfly_st1~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][0][10]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][10] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][10] .power_up = "low";

cycloneive_lcell_comb \Mux151~0 (
	.dataa(\x_2_imag_held[10]~q ),
	.datab(\butterfly_st1[1][0][10]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux151~0_combout ),
	.cout());
defparam \Mux151~0 .lut_mask = 16'hEFFE;
defparam \Mux151~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][0][9] (
	.clk(clk),
	.d(\butterfly_st1~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][9] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][9] .power_up = "low";

cycloneive_lcell_comb \Mux186~0 (
	.dataa(\x_4_imag_held[9]~q ),
	.datab(\butterfly_st1[3][0][9]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux186~0_combout ),
	.cout());
defparam \Mux186~0 .lut_mask = 16'hEFFE;
defparam \Mux186~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][0][9] (
	.clk(clk),
	.d(\butterfly_st1~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][9] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][9] .power_up = "low";

cycloneive_lcell_comb \Mux152~0 (
	.dataa(\x_2_imag_held[9]~q ),
	.datab(\butterfly_st1[1][0][9]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux152~0_combout ),
	.cout());
defparam \Mux152~0 .lut_mask = 16'hEFFE;
defparam \Mux152~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][0][8] (
	.clk(clk),
	.d(\butterfly_st1~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][8] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][8] .power_up = "low";

cycloneive_lcell_comb \Mux187~0 (
	.dataa(\x_4_imag_held[8]~q ),
	.datab(\butterfly_st1[3][0][8]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux187~0_combout ),
	.cout());
defparam \Mux187~0 .lut_mask = 16'hEFFE;
defparam \Mux187~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][0][8] (
	.clk(clk),
	.d(\butterfly_st1~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][8] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][8] .power_up = "low";

cycloneive_lcell_comb \Mux153~0 (
	.dataa(\x_2_imag_held[8]~q ),
	.datab(\butterfly_st1[1][0][8]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux153~0_combout ),
	.cout());
defparam \Mux153~0 .lut_mask = 16'hEFFE;
defparam \Mux153~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][0][7] (
	.clk(clk),
	.d(\butterfly_st1~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][7] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][7] .power_up = "low";

cycloneive_lcell_comb \Mux188~0 (
	.dataa(\x_4_imag_held[7]~q ),
	.datab(\butterfly_st1[3][0][7]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux188~0_combout ),
	.cout());
defparam \Mux188~0 .lut_mask = 16'hEFFE;
defparam \Mux188~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][0][7] (
	.clk(clk),
	.d(\butterfly_st1~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][7] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][7] .power_up = "low";

cycloneive_lcell_comb \Mux154~0 (
	.dataa(\x_2_imag_held[7]~q ),
	.datab(\butterfly_st1[1][0][7]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux154~0_combout ),
	.cout());
defparam \Mux154~0 .lut_mask = 16'hEFFE;
defparam \Mux154~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][0][6] (
	.clk(clk),
	.d(\butterfly_st1~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][6] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][6] .power_up = "low";

cycloneive_lcell_comb \Mux189~0 (
	.dataa(\x_4_imag_held[6]~q ),
	.datab(\butterfly_st1[3][0][6]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux189~0_combout ),
	.cout());
defparam \Mux189~0 .lut_mask = 16'hEFFE;
defparam \Mux189~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][0][6] (
	.clk(clk),
	.d(\butterfly_st1~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][6] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][6] .power_up = "low";

cycloneive_lcell_comb \Mux155~0 (
	.dataa(\x_2_imag_held[6]~q ),
	.datab(\butterfly_st1[1][0][6]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux155~0_combout ),
	.cout());
defparam \Mux155~0 .lut_mask = 16'hEFFE;
defparam \Mux155~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][0][5] (
	.clk(clk),
	.d(\butterfly_st1~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][5] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][5] .power_up = "low";

cycloneive_lcell_comb \Mux190~0 (
	.dataa(\x_4_imag_held[5]~q ),
	.datab(\butterfly_st1[3][0][5]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux190~0_combout ),
	.cout());
defparam \Mux190~0 .lut_mask = 16'hEFFE;
defparam \Mux190~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][0][5] (
	.clk(clk),
	.d(\butterfly_st1~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][5] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][5] .power_up = "low";

cycloneive_lcell_comb \Mux156~0 (
	.dataa(\x_2_imag_held[5]~q ),
	.datab(\butterfly_st1[1][0][5]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux156~0_combout ),
	.cout());
defparam \Mux156~0 .lut_mask = 16'hEFFE;
defparam \Mux156~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][0][4] (
	.clk(clk),
	.d(\butterfly_st1~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][4] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][4] .power_up = "low";

cycloneive_lcell_comb \Mux191~0 (
	.dataa(\x_4_imag_held[4]~q ),
	.datab(\butterfly_st1[3][0][4]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux191~0_combout ),
	.cout());
defparam \Mux191~0 .lut_mask = 16'hEFFE;
defparam \Mux191~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][0][4] (
	.clk(clk),
	.d(\butterfly_st1~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][4] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][4] .power_up = "low";

cycloneive_lcell_comb \Mux157~0 (
	.dataa(\x_2_imag_held[4]~q ),
	.datab(\butterfly_st1[1][0][4]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux157~0_combout ),
	.cout());
defparam \Mux157~0 .lut_mask = 16'hEFFE;
defparam \Mux157~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[3][0][3] (
	.clk(clk),
	.d(\butterfly_st1~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[3][1][0]~0_combout ),
	.q(\butterfly_st1[3][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][3] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][3] .power_up = "low";

cycloneive_lcell_comb \Mux192~0 (
	.dataa(\x_4_imag_held[3]~q ),
	.datab(\butterfly_st1[3][0][3]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux192~0_combout ),
	.cout());
defparam \Mux192~0 .lut_mask = 16'hEFFE;
defparam \Mux192~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[1][0][3] (
	.clk(clk),
	.d(\butterfly_st1~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[1][1][0]~0_combout ),
	.q(\butterfly_st1[1][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][3] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][3] .power_up = "low";

cycloneive_lcell_comb \Mux158~0 (
	.dataa(\x_2_imag_held[3]~q ),
	.datab(\butterfly_st1[1][0][3]~q ),
	.datac(\sel_arr[9][1]~q ),
	.datad(\sel_arr[9][0]~q ),
	.cin(gnd),
	.combout(\Mux158~0_combout ),
	.cout());
defparam \Mux158~0 .lut_mask = 16'hEFFE;
defparam \Mux158~0 .sum_lutc_input = "datac";

dffeas \butterfly_st1[2][0][15] (
	.clk(clk),
	.d(\butterfly_st1~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][0][15]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][15] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][15] .power_up = "low";

dffeas \butterfly_st1[0][0][15] (
	.clk(clk),
	.d(\butterfly_st1~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][0][15]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][15] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][15] .power_up = "low";

dffeas \butterfly_st1[2][0][14] (
	.clk(clk),
	.d(\butterfly_st1~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][0][14]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][14] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][14] .power_up = "low";

dffeas \butterfly_st1[0][0][14] (
	.clk(clk),
	.d(\butterfly_st1~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][0][14]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][14] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][14] .power_up = "low";

dffeas \butterfly_st1[2][0][13] (
	.clk(clk),
	.d(\butterfly_st1~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][0][13]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][13] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][13] .power_up = "low";

dffeas \butterfly_st1[0][0][13] (
	.clk(clk),
	.d(\butterfly_st1~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][0][13]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][13] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][13] .power_up = "low";

dffeas \butterfly_st1[2][0][12] (
	.clk(clk),
	.d(\butterfly_st1~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][0][12]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][12] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][12] .power_up = "low";

dffeas \butterfly_st1[0][0][12] (
	.clk(clk),
	.d(\butterfly_st1~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][0][12]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][12] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][12] .power_up = "low";

dffeas \butterfly_st1[2][0][11] (
	.clk(clk),
	.d(\butterfly_st1~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][0][11]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][11] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][11] .power_up = "low";

dffeas \butterfly_st1[0][0][11] (
	.clk(clk),
	.d(\butterfly_st1~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][0][11]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][11] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][11] .power_up = "low";

dffeas \butterfly_st1[2][0][10] (
	.clk(clk),
	.d(\butterfly_st1~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][0][10]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][10] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][10] .power_up = "low";

dffeas \butterfly_st1[0][0][10] (
	.clk(clk),
	.d(\butterfly_st1~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][0][10]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][10] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][10] .power_up = "low";

dffeas \butterfly_st1[2][0][9] (
	.clk(clk),
	.d(\butterfly_st1~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][9] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][9] .power_up = "low";

dffeas \butterfly_st1[0][0][9] (
	.clk(clk),
	.d(\butterfly_st1~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][9] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][9] .power_up = "low";

dffeas \butterfly_st1[2][0][8] (
	.clk(clk),
	.d(\butterfly_st1~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][8] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][8] .power_up = "low";

dffeas \butterfly_st1[0][0][8] (
	.clk(clk),
	.d(\butterfly_st1~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][8] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][8] .power_up = "low";

dffeas \butterfly_st1[2][0][7] (
	.clk(clk),
	.d(\butterfly_st1~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][7] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][7] .power_up = "low";

dffeas \butterfly_st1[0][0][7] (
	.clk(clk),
	.d(\butterfly_st1~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][7] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][7] .power_up = "low";

dffeas \butterfly_st1[2][0][6] (
	.clk(clk),
	.d(\butterfly_st1~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][6] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][6] .power_up = "low";

dffeas \butterfly_st1[0][0][6] (
	.clk(clk),
	.d(\butterfly_st1~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][6] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][6] .power_up = "low";

dffeas \butterfly_st1[2][0][5] (
	.clk(clk),
	.d(\butterfly_st1~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][5] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][5] .power_up = "low";

dffeas \butterfly_st1[0][0][5] (
	.clk(clk),
	.d(\butterfly_st1~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][5] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][5] .power_up = "low";

dffeas \butterfly_st1[2][0][4] (
	.clk(clk),
	.d(\butterfly_st1~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][4] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][4] .power_up = "low";

dffeas \butterfly_st1[0][0][4] (
	.clk(clk),
	.d(\butterfly_st1~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][4] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][4] .power_up = "low";

dffeas \butterfly_st1[2][0][3] (
	.clk(clk),
	.d(\butterfly_st1~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[2][1][0]~0_combout ),
	.q(\butterfly_st1[2][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][3] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][3] .power_up = "low";

dffeas \butterfly_st1[0][0][3] (
	.clk(clk),
	.d(\butterfly_st1~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\butterfly_st1[0][1][0]~0_combout ),
	.q(\butterfly_st1[0][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][3] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][3] .power_up = "low";

dffeas \sel_arr[7][1] (
	.clk(clk),
	.d(\sel_arr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[7][1]~q ),
	.prn(vcc));
defparam \sel_arr[7][1] .is_wysiwyg = "true";
defparam \sel_arr[7][1] .power_up = "low";

cycloneive_lcell_comb \sel_arr~2 (
	.dataa(reset),
	.datab(\sel_arr[7][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~2_combout ),
	.cout());
defparam \sel_arr~2 .lut_mask = 16'hEEEE;
defparam \sel_arr~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~0 (
	.dataa(reset),
	.datab(\bfp_scale|i_array_out[0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~0_combout ),
	.cout());
defparam \butterfly_st1~0 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~0 .sum_lutc_input = "datac";

dffeas \sel_arr[5][0] (
	.clk(clk),
	.d(\sel_arr~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[5][0]~q ),
	.prn(vcc));
defparam \sel_arr[5][0] .is_wysiwyg = "true";
defparam \sel_arr[5][0] .power_up = "low";

dffeas \sel_arr[5][1] (
	.clk(clk),
	.d(\sel_arr~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[5][1]~q ),
	.prn(vcc));
defparam \sel_arr[5][1] .is_wysiwyg = "true";
defparam \sel_arr[5][1] .power_up = "low";

cycloneive_lcell_comb \butterfly_st1[3][1][0]~0 (
	.dataa(\sel_arr[5][0]~q ),
	.datab(\sel_arr[5][1]~q ),
	.datac(reset),
	.datad(global_clock_enable),
	.cin(gnd),
	.combout(\butterfly_st1[3][1][0]~0_combout ),
	.cout());
defparam \butterfly_st1[3][1][0]~0 .lut_mask = 16'hFFEF;
defparam \butterfly_st1[3][1][0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1[1][1][0]~0 (
	.dataa(\sel_arr[5][0]~q ),
	.datab(\sel_arr[5][1]~q ),
	.datac(reset),
	.datad(global_clock_enable),
	.cin(gnd),
	.combout(\butterfly_st1[1][1][0]~0_combout ),
	.cout());
defparam \butterfly_st1[1][1][0]~0 .lut_mask = 16'hFFBF;
defparam \butterfly_st1[1][1][0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~1 (
	.dataa(reset),
	.datab(\bfp_scale|i_array_out[0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~1_combout ),
	.cout());
defparam \butterfly_st1~1 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~2 (
	.dataa(reset),
	.datab(\bfp_scale|i_array_out[0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~2_combout ),
	.cout());
defparam \butterfly_st1~2 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1[2][1][0]~0 (
	.dataa(\sel_arr[5][1]~q ),
	.datab(\sel_arr[5][0]~q ),
	.datac(reset),
	.datad(global_clock_enable),
	.cin(gnd),
	.combout(\butterfly_st1[2][1][0]~0_combout ),
	.cout());
defparam \butterfly_st1[2][1][0]~0 .lut_mask = 16'hFFBF;
defparam \butterfly_st1[2][1][0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1[0][1][0]~0 (
	.dataa(global_clock_enable),
	.datab(reset),
	.datac(\sel_arr[5][0]~q ),
	.datad(\sel_arr[5][1]~q ),
	.cin(gnd),
	.combout(\butterfly_st1[0][1][0]~0_combout ),
	.cout());
defparam \butterfly_st1[0][1][0]~0 .lut_mask = 16'hBFFF;
defparam \butterfly_st1[0][1][0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~3 (
	.dataa(reset),
	.datab(\bfp_scale|i_array_out[0][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~3_combout ),
	.cout());
defparam \butterfly_st1~3 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~4 (
	.dataa(reset),
	.datab(\bfp_scale|i_array_out[0][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~4_combout ),
	.cout());
defparam \butterfly_st1~4 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~5 (
	.dataa(reset),
	.datab(\bfp_scale|i_array_out[0][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~5_combout ),
	.cout());
defparam \butterfly_st1~5 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~6 (
	.dataa(reset),
	.datab(\bfp_scale|i_array_out[0][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~6_combout ),
	.cout());
defparam \butterfly_st1~6 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~7 (
	.dataa(reset),
	.datab(\bfp_scale|i_array_out[0][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~7_combout ),
	.cout());
defparam \butterfly_st1~7 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~8 (
	.dataa(reset),
	.datab(\bfp_scale|i_array_out[0][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~8_combout ),
	.cout());
defparam \butterfly_st1~8 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~9 (
	.dataa(reset),
	.datab(\bfp_scale|i_array_out[0][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~9_combout ),
	.cout());
defparam \butterfly_st1~9 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~10 (
	.dataa(reset),
	.datab(\bfp_scale|i_array_out[0][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~10_combout ),
	.cout());
defparam \butterfly_st1~10 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~11 (
	.dataa(reset),
	.datab(\bfp_scale|i_array_out[0][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~11_combout ),
	.cout());
defparam \butterfly_st1~11 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~12 (
	.dataa(reset),
	.datab(\bfp_scale|i_array_out[0][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~12_combout ),
	.cout());
defparam \butterfly_st1~12 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~13 (
	.dataa(reset),
	.datab(\bfp_scale|i_array_out[0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~13_combout ),
	.cout());
defparam \butterfly_st1~13 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~14 (
	.dataa(reset),
	.datab(\bfp_scale|i_array_out[0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~14_combout ),
	.cout());
defparam \butterfly_st1~14 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~15 (
	.dataa(reset),
	.datab(\bfp_scale|i_array_out[0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~15_combout ),
	.cout());
defparam \butterfly_st1~15 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~15 .sum_lutc_input = "datac";

dffeas \sel_arr[7][0] (
	.clk(clk),
	.d(\sel_arr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[7][0]~q ),
	.prn(vcc));
defparam \sel_arr[7][0] .is_wysiwyg = "true";
defparam \sel_arr[7][0] .power_up = "low";

cycloneive_lcell_comb \sel_arr~3 (
	.dataa(reset),
	.datab(\sel_arr[7][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~3_combout ),
	.cout());
defparam \sel_arr~3 .lut_mask = 16'hEEEE;
defparam \sel_arr~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~16 (
	.dataa(reset),
	.datab(\bfp_scale|r_array_out[0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~16_combout ),
	.cout());
defparam \butterfly_st1~16 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~17 (
	.dataa(reset),
	.datab(\bfp_scale|r_array_out[0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~17_combout ),
	.cout());
defparam \butterfly_st1~17 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~18 (
	.dataa(reset),
	.datab(\bfp_scale|r_array_out[0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~18_combout ),
	.cout());
defparam \butterfly_st1~18 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~19 (
	.dataa(reset),
	.datab(\bfp_scale|r_array_out[0][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~19_combout ),
	.cout());
defparam \butterfly_st1~19 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~20 (
	.dataa(reset),
	.datab(\bfp_scale|r_array_out[0][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~20_combout ),
	.cout());
defparam \butterfly_st1~20 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~21 (
	.dataa(reset),
	.datab(\bfp_scale|r_array_out[0][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~21_combout ),
	.cout());
defparam \butterfly_st1~21 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~22 (
	.dataa(reset),
	.datab(\bfp_scale|r_array_out[0][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~22_combout ),
	.cout());
defparam \butterfly_st1~22 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~23 (
	.dataa(reset),
	.datab(\bfp_scale|r_array_out[0][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~23_combout ),
	.cout());
defparam \butterfly_st1~23 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~24 (
	.dataa(reset),
	.datab(\bfp_scale|r_array_out[0][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~24_combout ),
	.cout());
defparam \butterfly_st1~24 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~25 (
	.dataa(reset),
	.datab(\bfp_scale|r_array_out[0][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~25_combout ),
	.cout());
defparam \butterfly_st1~25 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~26 (
	.dataa(reset),
	.datab(\bfp_scale|r_array_out[0][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~26_combout ),
	.cout());
defparam \butterfly_st1~26 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~27 (
	.dataa(reset),
	.datab(\bfp_scale|r_array_out[0][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~27_combout ),
	.cout());
defparam \butterfly_st1~27 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~28 (
	.dataa(reset),
	.datab(\bfp_scale|r_array_out[0][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~28_combout ),
	.cout());
defparam \butterfly_st1~28 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~29 (
	.dataa(reset),
	.datab(\bfp_scale|r_array_out[0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~29_combout ),
	.cout());
defparam \butterfly_st1~29 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~30 (
	.dataa(reset),
	.datab(\bfp_scale|r_array_out[0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~30_combout ),
	.cout());
defparam \butterfly_st1~30 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1~31 (
	.dataa(reset),
	.datab(\bfp_scale|r_array_out[0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\butterfly_st1~31_combout ),
	.cout());
defparam \butterfly_st1~31 .lut_mask = 16'hEEEE;
defparam \butterfly_st1~31 .sum_lutc_input = "datac";

dffeas \sel_arr[6][1] (
	.clk(clk),
	.d(\sel_arr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[6][1]~q ),
	.prn(vcc));
defparam \sel_arr[6][1] .is_wysiwyg = "true";
defparam \sel_arr[6][1] .power_up = "low";

cycloneive_lcell_comb \sel_arr~4 (
	.dataa(reset),
	.datab(\sel_arr[6][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~4_combout ),
	.cout());
defparam \sel_arr~4 .lut_mask = 16'hEEEE;
defparam \sel_arr~4 .sum_lutc_input = "datac";

dffeas \sel_arr[4][0] (
	.clk(clk),
	.d(\sel_arr~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[4][0]~q ),
	.prn(vcc));
defparam \sel_arr[4][0] .is_wysiwyg = "true";
defparam \sel_arr[4][0] .power_up = "low";

cycloneive_lcell_comb \sel_arr~5 (
	.dataa(reset),
	.datab(\sel_arr[4][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~5_combout ),
	.cout());
defparam \sel_arr~5 .lut_mask = 16'hEEEE;
defparam \sel_arr~5 .sum_lutc_input = "datac";

dffeas \sel_arr[4][1] (
	.clk(clk),
	.d(\sel_arr~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[4][1]~q ),
	.prn(vcc));
defparam \sel_arr[4][1] .is_wysiwyg = "true";
defparam \sel_arr[4][1] .power_up = "low";

cycloneive_lcell_comb \sel_arr~6 (
	.dataa(reset),
	.datab(\sel_arr[4][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~6_combout ),
	.cout());
defparam \sel_arr~6 .lut_mask = 16'hEEEE;
defparam \sel_arr~6 .sum_lutc_input = "datac";

dffeas \sel_arr[6][0] (
	.clk(clk),
	.d(\sel_arr~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[6][0]~q ),
	.prn(vcc));
defparam \sel_arr[6][0] .is_wysiwyg = "true";
defparam \sel_arr[6][0] .power_up = "low";

cycloneive_lcell_comb \sel_arr~7 (
	.dataa(reset),
	.datab(\sel_arr[6][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~7_combout ),
	.cout());
defparam \sel_arr~7 .lut_mask = 16'hEEEE;
defparam \sel_arr~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sel_arr~8 (
	.dataa(reset),
	.datab(\sel_arr[5][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~8_combout ),
	.cout());
defparam \sel_arr~8 .lut_mask = 16'hEEEE;
defparam \sel_arr~8 .sum_lutc_input = "datac";

dffeas \sel_arr[3][0] (
	.clk(clk),
	.d(\sel_arr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[3][0]~q ),
	.prn(vcc));
defparam \sel_arr[3][0] .is_wysiwyg = "true";
defparam \sel_arr[3][0] .power_up = "low";

cycloneive_lcell_comb \sel_arr~9 (
	.dataa(reset),
	.datab(\sel_arr[3][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~9_combout ),
	.cout());
defparam \sel_arr~9 .lut_mask = 16'hEEEE;
defparam \sel_arr~9 .sum_lutc_input = "datac";

dffeas \sel_arr[3][1] (
	.clk(clk),
	.d(\sel_arr~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[3][1]~q ),
	.prn(vcc));
defparam \sel_arr[3][1] .is_wysiwyg = "true";
defparam \sel_arr[3][1] .power_up = "low";

cycloneive_lcell_comb \sel_arr~10 (
	.dataa(reset),
	.datab(\sel_arr[3][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~10_combout ),
	.cout());
defparam \sel_arr~10 .lut_mask = 16'hEEEE;
defparam \sel_arr~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sel_arr~11 (
	.dataa(reset),
	.datab(\sel_arr[5][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~11_combout ),
	.cout());
defparam \sel_arr~11 .lut_mask = 16'hEEEE;
defparam \sel_arr~11 .sum_lutc_input = "datac";

dffeas \sel_arr[2][0] (
	.clk(clk),
	.d(\sel_arr~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[2][0]~q ),
	.prn(vcc));
defparam \sel_arr[2][0] .is_wysiwyg = "true";
defparam \sel_arr[2][0] .power_up = "low";

cycloneive_lcell_comb \sel_arr~12 (
	.dataa(reset),
	.datab(\sel_arr[2][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~12_combout ),
	.cout());
defparam \sel_arr~12 .lut_mask = 16'hEEEE;
defparam \sel_arr~12 .sum_lutc_input = "datac";

dffeas \sel_arr[2][1] (
	.clk(clk),
	.d(\sel_arr~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[2][1]~q ),
	.prn(vcc));
defparam \sel_arr[2][1] .is_wysiwyg = "true";
defparam \sel_arr[2][1] .power_up = "low";

cycloneive_lcell_comb \sel_arr~13 (
	.dataa(reset),
	.datab(\sel_arr[2][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~13_combout ),
	.cout());
defparam \sel_arr~13 .lut_mask = 16'hEEEE;
defparam \sel_arr~13 .sum_lutc_input = "datac";

dffeas \sel_arr[1][0] (
	.clk(clk),
	.d(\sel_arr~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[1][0]~q ),
	.prn(vcc));
defparam \sel_arr[1][0] .is_wysiwyg = "true";
defparam \sel_arr[1][0] .power_up = "low";

cycloneive_lcell_comb \sel_arr~14 (
	.dataa(reset),
	.datab(\sel_arr[1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~14_combout ),
	.cout());
defparam \sel_arr~14 .lut_mask = 16'hEEEE;
defparam \sel_arr~14 .sum_lutc_input = "datac";

dffeas \sel_arr[1][1] (
	.clk(clk),
	.d(\sel_arr~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[1][1]~q ),
	.prn(vcc));
defparam \sel_arr[1][1] .is_wysiwyg = "true";
defparam \sel_arr[1][1] .power_up = "low";

cycloneive_lcell_comb \sel_arr~15 (
	.dataa(reset),
	.datab(\sel_arr[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~15_combout ),
	.cout());
defparam \sel_arr~15 .lut_mask = 16'hEEEE;
defparam \sel_arr~15 .sum_lutc_input = "datac";

dffeas \sel_arr[0][0] (
	.clk(clk),
	.d(\sel_arr~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[0][0]~q ),
	.prn(vcc));
defparam \sel_arr[0][0] .is_wysiwyg = "true";
defparam \sel_arr[0][0] .power_up = "low";

cycloneive_lcell_comb \sel_arr~16 (
	.dataa(reset),
	.datab(\sel_arr[0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~16_combout ),
	.cout());
defparam \sel_arr~16 .lut_mask = 16'hEEEE;
defparam \sel_arr~16 .sum_lutc_input = "datac";

dffeas \sel_arr[0][1] (
	.clk(clk),
	.d(\sel_arr~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sel_arr[0][1]~q ),
	.prn(vcc));
defparam \sel_arr[0][1] .is_wysiwyg = "true";
defparam \sel_arr[0][1] .power_up = "low";

cycloneive_lcell_comb \sel_arr~17 (
	.dataa(reset),
	.datab(\sel_arr[0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~17_combout ),
	.cout());
defparam \sel_arr~17 .lut_mask = 16'hEEEE;
defparam \sel_arr~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sel_arr~18 (
	.dataa(reset),
	.datab(k_count_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~18_combout ),
	.cout());
defparam \sel_arr~18 .lut_mask = 16'hEEEE;
defparam \sel_arr~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sel_arr~19 (
	.dataa(reset),
	.datab(k_count_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sel_arr~19_combout ),
	.cout());
defparam \sel_arr~19 .lut_mask = 16'hEEEE;
defparam \sel_arr~19 .sum_lutc_input = "datac";

endmodule

module fft256_asj_fft_bfp_i_fft_121 (
	i_array_out_2_0,
	i_array_out_13_0,
	i_array_out_12_0,
	i_array_out_11_0,
	i_array_out_10_0,
	i_array_out_9_0,
	i_array_out_8_0,
	i_array_out_7_0,
	i_array_out_6_0,
	i_array_out_5_0,
	i_array_out_4_0,
	i_array_out_3_0,
	r_array_out_2_0,
	r_array_out_13_0,
	r_array_out_12_0,
	r_array_out_11_0,
	r_array_out_10_0,
	r_array_out_9_0,
	r_array_out_8_0,
	r_array_out_7_0,
	r_array_out_6_0,
	r_array_out_5_0,
	r_array_out_4_0,
	r_array_out_3_0,
	global_clock_enable,
	i_array_out_1_0,
	i_array_out_0_0,
	i_array_out_15_0,
	i_array_out_14_0,
	r_array_out_1_0,
	r_array_out_0_0,
	r_array_out_15_0,
	r_array_out_14_0,
	ram_data_out_0,
	ram_data_out_2,
	slb_last_1,
	ram_data_out_1,
	slb_last_0,
	slb_last_2,
	ram_data_out_14,
	ram_data_out_12,
	ram_data_out_13,
	ram_data_out_15,
	ram_data_out_11,
	ram_data_out_10,
	ram_data_out_9,
	ram_data_out_8,
	ram_data_out_7,
	ram_data_out_6,
	ram_data_out_5,
	ram_data_out_4,
	ram_data_out_3,
	ram_data_out_16,
	ram_data_out_18,
	ram_data_out_17,
	ram_data_out_28,
	ram_data_out_29,
	ram_data_out_30,
	ram_data_out_31,
	ram_data_out_27,
	ram_data_out_26,
	ram_data_out_25,
	ram_data_out_24,
	ram_data_out_23,
	ram_data_out_22,
	ram_data_out_21,
	ram_data_out_20,
	ram_data_out_19,
	clk)/* synthesis synthesis_greybox=1 */;
output 	i_array_out_2_0;
output 	i_array_out_13_0;
output 	i_array_out_12_0;
output 	i_array_out_11_0;
output 	i_array_out_10_0;
output 	i_array_out_9_0;
output 	i_array_out_8_0;
output 	i_array_out_7_0;
output 	i_array_out_6_0;
output 	i_array_out_5_0;
output 	i_array_out_4_0;
output 	i_array_out_3_0;
output 	r_array_out_2_0;
output 	r_array_out_13_0;
output 	r_array_out_12_0;
output 	r_array_out_11_0;
output 	r_array_out_10_0;
output 	r_array_out_9_0;
output 	r_array_out_8_0;
output 	r_array_out_7_0;
output 	r_array_out_6_0;
output 	r_array_out_5_0;
output 	r_array_out_4_0;
output 	r_array_out_3_0;
input 	global_clock_enable;
output 	i_array_out_1_0;
output 	i_array_out_0_0;
output 	i_array_out_15_0;
output 	i_array_out_14_0;
output 	r_array_out_1_0;
output 	r_array_out_0_0;
output 	r_array_out_15_0;
output 	r_array_out_14_0;
input 	ram_data_out_0;
input 	ram_data_out_2;
input 	slb_last_1;
input 	ram_data_out_1;
input 	slb_last_0;
input 	slb_last_2;
input 	ram_data_out_14;
input 	ram_data_out_12;
input 	ram_data_out_13;
input 	ram_data_out_15;
input 	ram_data_out_11;
input 	ram_data_out_10;
input 	ram_data_out_9;
input 	ram_data_out_8;
input 	ram_data_out_7;
input 	ram_data_out_6;
input 	ram_data_out_5;
input 	ram_data_out_4;
input 	ram_data_out_3;
input 	ram_data_out_16;
input 	ram_data_out_18;
input 	ram_data_out_17;
input 	ram_data_out_28;
input 	ram_data_out_29;
input 	ram_data_out_30;
input 	ram_data_out_31;
input 	ram_data_out_27;
input 	ram_data_out_26;
input 	ram_data_out_25;
input 	ram_data_out_24;
input 	ram_data_out_23;
input 	ram_data_out_22;
input 	ram_data_out_21;
input 	ram_data_out_20;
input 	ram_data_out_19;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux28~0_combout ;
wire \Mux29~0_combout ;
wire \Mux18~0_combout ;
wire \Mux31~1_combout ;
wire \Mux18~1_combout ;
wire \Mux19~0_combout ;
wire \Mux31~2_combout ;
wire \Mux19~1_combout ;
wire \Mux20~0_combout ;
wire \Mux21~0_combout ;
wire \Mux20~1_combout ;
wire \Mux22~0_combout ;
wire \Mux21~1_combout ;
wire \Mux23~0_combout ;
wire \Mux22~1_combout ;
wire \Mux24~0_combout ;
wire \Mux23~1_combout ;
wire \Mux25~0_combout ;
wire \Mux24~1_combout ;
wire \Mux26~0_combout ;
wire \Mux25~1_combout ;
wire \Mux26~1_combout ;
wire \Mux26~2_combout ;
wire \Mux28~1_combout ;
wire \Mux27~0_combout ;
wire \Mux28~2_combout ;
wire \Mux12~0_combout ;
wire \Mux13~0_combout ;
wire \Mux2~0_combout ;
wire \Mux15~1_combout ;
wire \Mux2~1_combout ;
wire \Mux3~0_combout ;
wire \Mux15~2_combout ;
wire \Mux3~1_combout ;
wire \Mux4~0_combout ;
wire \Mux5~0_combout ;
wire \Mux4~1_combout ;
wire \Mux6~0_combout ;
wire \Mux5~1_combout ;
wire \Mux7~0_combout ;
wire \Mux6~1_combout ;
wire \Mux8~0_combout ;
wire \Mux7~1_combout ;
wire \Mux9~0_combout ;
wire \Mux8~1_combout ;
wire \Mux10~0_combout ;
wire \Mux9~1_combout ;
wire \Mux10~1_combout ;
wire \Mux10~2_combout ;
wire \Mux12~1_combout ;
wire \Mux11~0_combout ;
wire \Mux12~2_combout ;
wire \r_array_out[0][1]~0_combout ;
wire \Mux30~0_combout ;
wire \Mux31~0_combout ;
wire \r_array_out[0][15]~1_combout ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \Mux17~0_combout ;
wire \Mux17~1_combout ;
wire \Mux14~0_combout ;
wire \Mux15~0_combout ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;


dffeas \i_array_out[0][2] (
	.clk(clk),
	.d(\Mux29~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_2_0),
	.prn(vcc));
defparam \i_array_out[0][2] .is_wysiwyg = "true";
defparam \i_array_out[0][2] .power_up = "low";

dffeas \i_array_out[0][13] (
	.clk(clk),
	.d(\Mux18~1_combout ),
	.asdata(ram_data_out_9),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_13_0),
	.prn(vcc));
defparam \i_array_out[0][13] .is_wysiwyg = "true";
defparam \i_array_out[0][13] .power_up = "low";

dffeas \i_array_out[0][12] (
	.clk(clk),
	.d(\Mux19~1_combout ),
	.asdata(ram_data_out_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_12_0),
	.prn(vcc));
defparam \i_array_out[0][12] .is_wysiwyg = "true";
defparam \i_array_out[0][12] .power_up = "low";

dffeas \i_array_out[0][11] (
	.clk(clk),
	.d(\Mux20~1_combout ),
	.asdata(ram_data_out_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_11_0),
	.prn(vcc));
defparam \i_array_out[0][11] .is_wysiwyg = "true";
defparam \i_array_out[0][11] .power_up = "low";

dffeas \i_array_out[0][10] (
	.clk(clk),
	.d(\Mux21~1_combout ),
	.asdata(ram_data_out_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_10_0),
	.prn(vcc));
defparam \i_array_out[0][10] .is_wysiwyg = "true";
defparam \i_array_out[0][10] .power_up = "low";

dffeas \i_array_out[0][9] (
	.clk(clk),
	.d(\Mux22~1_combout ),
	.asdata(ram_data_out_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_9_0),
	.prn(vcc));
defparam \i_array_out[0][9] .is_wysiwyg = "true";
defparam \i_array_out[0][9] .power_up = "low";

dffeas \i_array_out[0][8] (
	.clk(clk),
	.d(\Mux23~1_combout ),
	.asdata(ram_data_out_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_8_0),
	.prn(vcc));
defparam \i_array_out[0][8] .is_wysiwyg = "true";
defparam \i_array_out[0][8] .power_up = "low";

dffeas \i_array_out[0][7] (
	.clk(clk),
	.d(\Mux24~1_combout ),
	.asdata(ram_data_out_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_7_0),
	.prn(vcc));
defparam \i_array_out[0][7] .is_wysiwyg = "true";
defparam \i_array_out[0][7] .power_up = "low";

dffeas \i_array_out[0][6] (
	.clk(clk),
	.d(\Mux25~1_combout ),
	.asdata(ram_data_out_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_6_0),
	.prn(vcc));
defparam \i_array_out[0][6] .is_wysiwyg = "true";
defparam \i_array_out[0][6] .power_up = "low";

dffeas \i_array_out[0][5] (
	.clk(clk),
	.d(\Mux26~2_combout ),
	.asdata(ram_data_out_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_5_0),
	.prn(vcc));
defparam \i_array_out[0][5] .is_wysiwyg = "true";
defparam \i_array_out[0][5] .power_up = "low";

dffeas \i_array_out[0][4] (
	.clk(clk),
	.d(\Mux27~0_combout ),
	.asdata(ram_data_out_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_4_0),
	.prn(vcc));
defparam \i_array_out[0][4] .is_wysiwyg = "true";
defparam \i_array_out[0][4] .power_up = "low";

dffeas \i_array_out[0][3] (
	.clk(clk),
	.d(\Mux28~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_3_0),
	.prn(vcc));
defparam \i_array_out[0][3] .is_wysiwyg = "true";
defparam \i_array_out[0][3] .power_up = "low";

dffeas \r_array_out[0][2] (
	.clk(clk),
	.d(\Mux13~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_2_0),
	.prn(vcc));
defparam \r_array_out[0][2] .is_wysiwyg = "true";
defparam \r_array_out[0][2] .power_up = "low";

dffeas \r_array_out[0][13] (
	.clk(clk),
	.d(\Mux2~1_combout ),
	.asdata(ram_data_out_25),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_13_0),
	.prn(vcc));
defparam \r_array_out[0][13] .is_wysiwyg = "true";
defparam \r_array_out[0][13] .power_up = "low";

dffeas \r_array_out[0][12] (
	.clk(clk),
	.d(\Mux3~1_combout ),
	.asdata(ram_data_out_24),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_12_0),
	.prn(vcc));
defparam \r_array_out[0][12] .is_wysiwyg = "true";
defparam \r_array_out[0][12] .power_up = "low";

dffeas \r_array_out[0][11] (
	.clk(clk),
	.d(\Mux4~1_combout ),
	.asdata(ram_data_out_23),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_11_0),
	.prn(vcc));
defparam \r_array_out[0][11] .is_wysiwyg = "true";
defparam \r_array_out[0][11] .power_up = "low";

dffeas \r_array_out[0][10] (
	.clk(clk),
	.d(\Mux5~1_combout ),
	.asdata(ram_data_out_22),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_10_0),
	.prn(vcc));
defparam \r_array_out[0][10] .is_wysiwyg = "true";
defparam \r_array_out[0][10] .power_up = "low";

dffeas \r_array_out[0][9] (
	.clk(clk),
	.d(\Mux6~1_combout ),
	.asdata(ram_data_out_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_9_0),
	.prn(vcc));
defparam \r_array_out[0][9] .is_wysiwyg = "true";
defparam \r_array_out[0][9] .power_up = "low";

dffeas \r_array_out[0][8] (
	.clk(clk),
	.d(\Mux7~1_combout ),
	.asdata(ram_data_out_20),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_8_0),
	.prn(vcc));
defparam \r_array_out[0][8] .is_wysiwyg = "true";
defparam \r_array_out[0][8] .power_up = "low";

dffeas \r_array_out[0][7] (
	.clk(clk),
	.d(\Mux8~1_combout ),
	.asdata(ram_data_out_19),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_7_0),
	.prn(vcc));
defparam \r_array_out[0][7] .is_wysiwyg = "true";
defparam \r_array_out[0][7] .power_up = "low";

dffeas \r_array_out[0][6] (
	.clk(clk),
	.d(\Mux9~1_combout ),
	.asdata(ram_data_out_18),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_6_0),
	.prn(vcc));
defparam \r_array_out[0][6] .is_wysiwyg = "true";
defparam \r_array_out[0][6] .power_up = "low";

dffeas \r_array_out[0][5] (
	.clk(clk),
	.d(\Mux10~2_combout ),
	.asdata(ram_data_out_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_5_0),
	.prn(vcc));
defparam \r_array_out[0][5] .is_wysiwyg = "true";
defparam \r_array_out[0][5] .power_up = "low";

dffeas \r_array_out[0][4] (
	.clk(clk),
	.d(\Mux11~0_combout ),
	.asdata(ram_data_out_16),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_4_0),
	.prn(vcc));
defparam \r_array_out[0][4] .is_wysiwyg = "true";
defparam \r_array_out[0][4] .power_up = "low";

dffeas \r_array_out[0][3] (
	.clk(clk),
	.d(\Mux12~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_3_0),
	.prn(vcc));
defparam \r_array_out[0][3] .is_wysiwyg = "true";
defparam \r_array_out[0][3] .power_up = "low";

dffeas \i_array_out[0][1] (
	.clk(clk),
	.d(\Mux30~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_1_0),
	.prn(vcc));
defparam \i_array_out[0][1] .is_wysiwyg = "true";
defparam \i_array_out[0][1] .power_up = "low";

dffeas \i_array_out[0][0] (
	.clk(clk),
	.d(\Mux31~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_0_0),
	.prn(vcc));
defparam \i_array_out[0][0] .is_wysiwyg = "true";
defparam \i_array_out[0][0] .power_up = "low";

dffeas \i_array_out[0][15] (
	.clk(clk),
	.d(\Mux16~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_15_0),
	.prn(vcc));
defparam \i_array_out[0][15] .is_wysiwyg = "true";
defparam \i_array_out[0][15] .power_up = "low";

dffeas \i_array_out[0][14] (
	.clk(clk),
	.d(\Mux17~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_14_0),
	.prn(vcc));
defparam \i_array_out[0][14] .is_wysiwyg = "true";
defparam \i_array_out[0][14] .power_up = "low";

dffeas \r_array_out[0][1] (
	.clk(clk),
	.d(\Mux14~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_1_0),
	.prn(vcc));
defparam \r_array_out[0][1] .is_wysiwyg = "true";
defparam \r_array_out[0][1] .power_up = "low";

dffeas \r_array_out[0][0] (
	.clk(clk),
	.d(\Mux15~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_0_0),
	.prn(vcc));
defparam \r_array_out[0][0] .is_wysiwyg = "true";
defparam \r_array_out[0][0] .power_up = "low";

dffeas \r_array_out[0][15] (
	.clk(clk),
	.d(\Mux0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_15_0),
	.prn(vcc));
defparam \r_array_out[0][15] .is_wysiwyg = "true";
defparam \r_array_out[0][15] .power_up = "low";

dffeas \r_array_out[0][14] (
	.clk(clk),
	.d(\Mux1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_14_0),
	.prn(vcc));
defparam \r_array_out[0][14] .is_wysiwyg = "true";
defparam \r_array_out[0][14] .power_up = "low";

cycloneive_lcell_comb \Mux28~0 (
	.dataa(ram_data_out_0),
	.datab(ram_data_out_2),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
defparam \Mux28~0 .lut_mask = 16'hAACC;
defparam \Mux28~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux29~0 (
	.dataa(\Mux28~0_combout ),
	.datab(ram_data_out_1),
	.datac(slb_last_0),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
defparam \Mux29~0 .lut_mask = 16'hACFF;
defparam \Mux29~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux18~0 (
	.dataa(slb_last_1),
	.datab(ram_data_out_10),
	.datac(ram_data_out_11),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
defparam \Mux18~0 .lut_mask = 16'hFAFC;
defparam \Mux18~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux31~1 (
	.dataa(ram_data_out_12),
	.datab(ram_data_out_13),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux31~1_combout ),
	.cout());
defparam \Mux31~1 .lut_mask = 16'hAACC;
defparam \Mux31~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux18~1 (
	.dataa(\Mux18~0_combout ),
	.datab(\Mux31~1_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
defparam \Mux18~1 .lut_mask = 16'hEEFF;
defparam \Mux18~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux19~0 (
	.dataa(slb_last_1),
	.datab(ram_data_out_9),
	.datac(ram_data_out_10),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
defparam \Mux19~0 .lut_mask = 16'hFAFC;
defparam \Mux19~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux31~2 (
	.dataa(ram_data_out_11),
	.datab(ram_data_out_12),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux31~2_combout ),
	.cout());
defparam \Mux31~2 .lut_mask = 16'hAACC;
defparam \Mux31~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux19~1 (
	.dataa(\Mux19~0_combout ),
	.datab(\Mux31~2_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux19~1_combout ),
	.cout());
defparam \Mux19~1 .lut_mask = 16'hEEFF;
defparam \Mux19~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux20~0 (
	.dataa(ram_data_out_9),
	.datab(ram_data_out_11),
	.datac(slb_last_1),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
defparam \Mux20~0 .lut_mask = 16'hACFF;
defparam \Mux20~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux21~0 (
	.dataa(ram_data_out_8),
	.datab(ram_data_out_10),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
defparam \Mux21~0 .lut_mask = 16'hAACC;
defparam \Mux21~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux20~1 (
	.dataa(\Mux20~0_combout ),
	.datab(slb_last_0),
	.datac(\Mux21~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
defparam \Mux20~1 .lut_mask = 16'hFEFE;
defparam \Mux20~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux22~0 (
	.dataa(ram_data_out_7),
	.datab(ram_data_out_9),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
defparam \Mux22~0 .lut_mask = 16'hAACC;
defparam \Mux22~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux21~1 (
	.dataa(\Mux22~0_combout ),
	.datab(\Mux21~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
defparam \Mux21~1 .lut_mask = 16'hAACC;
defparam \Mux21~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux23~0 (
	.dataa(ram_data_out_6),
	.datab(ram_data_out_8),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
defparam \Mux23~0 .lut_mask = 16'hAACC;
defparam \Mux23~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux22~1 (
	.dataa(\Mux23~0_combout ),
	.datab(\Mux22~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
defparam \Mux22~1 .lut_mask = 16'hAACC;
defparam \Mux22~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux24~0 (
	.dataa(ram_data_out_5),
	.datab(ram_data_out_7),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
defparam \Mux24~0 .lut_mask = 16'hAACC;
defparam \Mux24~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux23~1 (
	.dataa(\Mux24~0_combout ),
	.datab(\Mux23~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
defparam \Mux23~1 .lut_mask = 16'hAACC;
defparam \Mux23~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux25~0 (
	.dataa(ram_data_out_4),
	.datab(ram_data_out_6),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
defparam \Mux25~0 .lut_mask = 16'hAACC;
defparam \Mux25~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux24~1 (
	.dataa(\Mux25~0_combout ),
	.datab(\Mux24~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
defparam \Mux24~1 .lut_mask = 16'hAACC;
defparam \Mux24~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux26~0 (
	.dataa(ram_data_out_3),
	.datab(ram_data_out_5),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
defparam \Mux26~0 .lut_mask = 16'hAACC;
defparam \Mux26~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux25~1 (
	.dataa(\Mux26~0_combout ),
	.datab(\Mux25~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
defparam \Mux25~1 .lut_mask = 16'hAACC;
defparam \Mux25~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux26~1 (
	.dataa(ram_data_out_2),
	.datab(ram_data_out_4),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
defparam \Mux26~1 .lut_mask = 16'hAACC;
defparam \Mux26~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux26~2 (
	.dataa(\Mux26~1_combout ),
	.datab(\Mux26~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux26~2_combout ),
	.cout());
defparam \Mux26~2 .lut_mask = 16'hAACC;
defparam \Mux26~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux28~1 (
	.dataa(ram_data_out_1),
	.datab(ram_data_out_3),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
defparam \Mux28~1 .lut_mask = 16'hAACC;
defparam \Mux28~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux27~0 (
	.dataa(\Mux28~1_combout ),
	.datab(\Mux26~1_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
defparam \Mux27~0 .lut_mask = 16'hAACC;
defparam \Mux27~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux28~2 (
	.dataa(\Mux28~0_combout ),
	.datab(\Mux28~1_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux28~2_combout ),
	.cout());
defparam \Mux28~2 .lut_mask = 16'hAACC;
defparam \Mux28~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux12~0 (
	.dataa(ram_data_out_16),
	.datab(ram_data_out_18),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
defparam \Mux12~0 .lut_mask = 16'hAACC;
defparam \Mux12~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux13~0 (
	.dataa(\Mux12~0_combout ),
	.datab(ram_data_out_17),
	.datac(slb_last_0),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
defparam \Mux13~0 .lut_mask = 16'hACFF;
defparam \Mux13~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~0 (
	.dataa(slb_last_1),
	.datab(ram_data_out_26),
	.datac(ram_data_out_27),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFAFC;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux15~1 (
	.dataa(ram_data_out_28),
	.datab(ram_data_out_29),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
defparam \Mux15~1 .lut_mask = 16'hAACC;
defparam \Mux15~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~1 (
	.dataa(\Mux2~0_combout ),
	.datab(\Mux15~1_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
defparam \Mux2~1 .lut_mask = 16'hEEFF;
defparam \Mux2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~0 (
	.dataa(slb_last_1),
	.datab(ram_data_out_25),
	.datac(ram_data_out_26),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hFAFC;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux15~2 (
	.dataa(ram_data_out_27),
	.datab(ram_data_out_28),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux15~2_combout ),
	.cout());
defparam \Mux15~2 .lut_mask = 16'hAACC;
defparam \Mux15~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~1 (
	.dataa(\Mux3~0_combout ),
	.datab(\Mux15~2_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
defparam \Mux3~1 .lut_mask = 16'hEEFF;
defparam \Mux3~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~0 (
	.dataa(ram_data_out_25),
	.datab(ram_data_out_27),
	.datac(slb_last_1),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'hACFF;
defparam \Mux4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~0 (
	.dataa(ram_data_out_24),
	.datab(ram_data_out_26),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'hAACC;
defparam \Mux5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~1 (
	.dataa(\Mux4~0_combout ),
	.datab(slb_last_0),
	.datac(\Mux5~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
defparam \Mux4~1 .lut_mask = 16'hFEFE;
defparam \Mux4~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~0 (
	.dataa(ram_data_out_23),
	.datab(ram_data_out_25),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'hAACC;
defparam \Mux6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~1 (
	.dataa(\Mux6~0_combout ),
	.datab(\Mux5~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
defparam \Mux5~1 .lut_mask = 16'hAACC;
defparam \Mux5~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~0 (
	.dataa(ram_data_out_22),
	.datab(ram_data_out_24),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'hAACC;
defparam \Mux7~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~1 (
	.dataa(\Mux7~0_combout ),
	.datab(\Mux6~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
defparam \Mux6~1 .lut_mask = 16'hAACC;
defparam \Mux6~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux8~0 (
	.dataa(ram_data_out_21),
	.datab(ram_data_out_23),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
defparam \Mux8~0 .lut_mask = 16'hAACC;
defparam \Mux8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~1 (
	.dataa(\Mux8~0_combout ),
	.datab(\Mux7~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
defparam \Mux7~1 .lut_mask = 16'hAACC;
defparam \Mux7~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux9~0 (
	.dataa(ram_data_out_20),
	.datab(ram_data_out_22),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
defparam \Mux9~0 .lut_mask = 16'hAACC;
defparam \Mux9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux8~1 (
	.dataa(\Mux9~0_combout ),
	.datab(\Mux8~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
defparam \Mux8~1 .lut_mask = 16'hAACC;
defparam \Mux8~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~0 (
	.dataa(ram_data_out_19),
	.datab(ram_data_out_21),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
defparam \Mux10~0 .lut_mask = 16'hAACC;
defparam \Mux10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux9~1 (
	.dataa(\Mux10~0_combout ),
	.datab(\Mux9~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
defparam \Mux9~1 .lut_mask = 16'hAACC;
defparam \Mux9~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~1 (
	.dataa(ram_data_out_18),
	.datab(ram_data_out_20),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
defparam \Mux10~1 .lut_mask = 16'hAACC;
defparam \Mux10~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~2 (
	.dataa(\Mux10~1_combout ),
	.datab(\Mux10~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux10~2_combout ),
	.cout());
defparam \Mux10~2 .lut_mask = 16'hAACC;
defparam \Mux10~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux12~1 (
	.dataa(ram_data_out_17),
	.datab(ram_data_out_19),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
defparam \Mux12~1 .lut_mask = 16'hAACC;
defparam \Mux12~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux11~0 (
	.dataa(\Mux12~1_combout ),
	.datab(\Mux10~1_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
defparam \Mux11~0 .lut_mask = 16'hAACC;
defparam \Mux11~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux12~2 (
	.dataa(\Mux12~0_combout ),
	.datab(\Mux12~1_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux12~2_combout ),
	.cout());
defparam \Mux12~2 .lut_mask = 16'hAACC;
defparam \Mux12~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \r_array_out[0][1]~0 (
	.dataa(slb_last_1),
	.datab(slb_last_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\r_array_out[0][1]~0_combout ),
	.cout());
defparam \r_array_out[0][1]~0 .lut_mask = 16'hEEEE;
defparam \r_array_out[0][1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux30~0 (
	.dataa(ram_data_out_0),
	.datab(ram_data_out_1),
	.datac(slb_last_0),
	.datad(\r_array_out[0][1]~0_combout ),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
defparam \Mux30~0 .lut_mask = 16'hACFF;
defparam \Mux30~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux31~0 (
	.dataa(ram_data_out_0),
	.datab(slb_last_0),
	.datac(slb_last_1),
	.datad(slb_last_2),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
defparam \Mux31~0 .lut_mask = 16'hBFFF;
defparam \Mux31~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \r_array_out[0][15]~1 (
	.dataa(slb_last_2),
	.datab(slb_last_0),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\r_array_out[0][15]~1_combout ),
	.cout());
defparam \r_array_out[0][15]~1 .lut_mask = 16'hEEFF;
defparam \r_array_out[0][15]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~0 (
	.dataa(\r_array_out[0][15]~1_combout ),
	.datab(\Mux31~1_combout ),
	.datac(\r_array_out[0][1]~0_combout ),
	.datad(ram_data_out_15),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
defparam \Mux16~0 .lut_mask = 16'hFFDE;
defparam \Mux16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~1 (
	.dataa(ram_data_out_14),
	.datab(\r_array_out[0][15]~1_combout ),
	.datac(\Mux16~0_combout ),
	.datad(ram_data_out_11),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
defparam \Mux16~1 .lut_mask = 16'hFFBE;
defparam \Mux16~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux17~0 (
	.dataa(\r_array_out[0][15]~1_combout ),
	.datab(\Mux31~2_combout ),
	.datac(\r_array_out[0][1]~0_combout ),
	.datad(ram_data_out_14),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
defparam \Mux17~0 .lut_mask = 16'hFFDE;
defparam \Mux17~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux17~1 (
	.dataa(ram_data_out_13),
	.datab(\r_array_out[0][15]~1_combout ),
	.datac(\Mux17~0_combout ),
	.datad(ram_data_out_10),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
defparam \Mux17~1 .lut_mask = 16'hFFBE;
defparam \Mux17~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux14~0 (
	.dataa(ram_data_out_16),
	.datab(ram_data_out_17),
	.datac(slb_last_0),
	.datad(\r_array_out[0][1]~0_combout ),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
defparam \Mux14~0 .lut_mask = 16'hACFF;
defparam \Mux14~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux15~0 (
	.dataa(ram_data_out_16),
	.datab(slb_last_0),
	.datac(slb_last_1),
	.datad(slb_last_2),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
defparam \Mux15~0 .lut_mask = 16'hBFFF;
defparam \Mux15~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(\r_array_out[0][1]~0_combout ),
	.datab(ram_data_out_30),
	.datac(\r_array_out[0][15]~1_combout ),
	.datad(ram_data_out_31),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hFFDE;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~1 (
	.dataa(\Mux15~1_combout ),
	.datab(\r_array_out[0][1]~0_combout ),
	.datac(\Mux0~0_combout ),
	.datad(ram_data_out_27),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hFFBE;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(\r_array_out[0][15]~1_combout ),
	.datab(\Mux15~2_combout ),
	.datac(\r_array_out[0][1]~0_combout ),
	.datad(ram_data_out_30),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hFFDE;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~1 (
	.dataa(ram_data_out_29),
	.datab(\r_array_out[0][15]~1_combout ),
	.datac(\Mux1~0_combout ),
	.datad(ram_data_out_26),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hFFBE;
defparam \Mux1~1 .sum_lutc_input = "datac";

endmodule

module fft256_asj_fft_bfp_o_fft_121 (
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_31,
	source_valid_ctrl_sop,
	stall_reg,
	source_stall_int_d,
	global_clock_enable,
	slb_i_0,
	Mux2,
	lut_out_0,
	tdl_arr_0,
	Mux1,
	lut_out_1,
	lut_out_2,
	lut_out_21,
	real_out_11,
	real_out_12,
	real_out_13,
	real_out_14,
	real_out_15,
	tdl_arr_01,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	pipeline_dffe_27;
input 	pipeline_dffe_28;
input 	pipeline_dffe_29;
input 	pipeline_dffe_30;
input 	pipeline_dffe_31;
input 	source_valid_ctrl_sop;
input 	stall_reg;
input 	source_stall_int_d;
input 	global_clock_enable;
output 	slb_i_0;
output 	Mux2;
output 	lut_out_0;
input 	tdl_arr_0;
output 	Mux1;
output 	lut_out_1;
output 	lut_out_2;
output 	lut_out_21;
input 	real_out_11;
input 	real_out_12;
input 	real_out_13;
input 	real_out_14;
input 	real_out_15;
input 	tdl_arr_01;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \del_np_cnt[4]~q ;
wire \del_np_cnt[3]~12 ;
wire \del_np_cnt[4]~13_combout ;
wire \gen_blk_float:gen_1_input_bfp_o:delay_next_pass3|tdl_arr[2]~q ;
wire \gen_blk_float:gen_1_input_bfp_o:delay_next_pass|tdl_arr[8]~q ;
wire \del_np_cnt[0]~6 ;
wire \del_np_cnt[1]~8 ;
wire \del_np_cnt[2]~9_combout ;
wire \del_np_cnt[0]~5_combout ;
wire \del_np_cnt[0]~q ;
wire \del_np_cnt[1]~7_combout ;
wire \del_np_cnt[1]~q ;
wire \del_np_cnt[2]~10 ;
wire \del_np_cnt[3]~11_combout ;
wire \del_np_cnt[3]~q ;
wire \Equal1~0_combout ;
wire \Selector3~0_combout ;
wire \sdet.DISABLE~q ;
wire \delay_next_pass_counter~2_combout ;
wire \del_np_cnt[2]~q ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \sdet.ENABLE~q ;
wire \en_gain_lut_8_pts~q ;
wire \gain_lut_8pts~0_combout ;
wire \gain_lut_8pts~1_combout ;
wire \gain_lut_8pts[0]~q ;
wire \sdet.IDLE~0_combout ;
wire \sdet.IDLE~q ;
wire \Selector1~0_combout ;
wire \sdet.BLOCK_READY~q ;
wire \slb_i[3]~1_combout ;
wire \gain_lut_blk~0_combout ;
wire \gain_lut_blk[0]~q ;
wire \slb_i~0_combout ;
wire \slb_i[3]~2_combout ;
wire \gain_lut_8pts~2_combout ;
wire \gain_lut_8pts~3_combout ;
wire \gain_lut_8pts[1]~q ;
wire \gain_lut_blk~1_combout ;
wire \gain_lut_blk[1]~q ;
wire \slb_i~3_combout ;
wire \slb_i[1]~q ;
wire \gain_lut_8pts~4_combout ;
wire \gain_lut_8pts~5_combout ;
wire \gain_lut_8pts[2]~q ;
wire \gain_lut_blk~2_combout ;
wire \gain_lut_blk[2]~q ;
wire \slb_i~4_combout ;
wire \slb_i[2]~q ;
wire \gain_lut_8pts~6_combout ;
wire \gain_lut_8pts~7_combout ;
wire \gain_lut_8pts[3]~q ;
wire \gain_lut_blk~3_combout ;
wire \gain_lut_blk[3]~q ;
wire \slb_i~5_combout ;
wire \slb_i[3]~q ;


fft256_asj_fft_tdl_bit_fft_121_2 \gen_blk_float:gen_1_input_bfp_o:delay_next_pass3 (
	.global_clock_enable(global_clock_enable),
	.tdl_arr_2(\gen_blk_float:gen_1_input_bfp_o:delay_next_pass3|tdl_arr[2]~q ),
	.data_in(\gen_blk_float:gen_1_input_bfp_o:delay_next_pass|tdl_arr[8]~q ),
	.clk(clk));

fft256_asj_fft_tdl_bit_fft_121_1 \gen_blk_float:gen_1_input_bfp_o:delay_next_pass (
	.global_clock_enable(global_clock_enable),
	.tdl_arr_0(tdl_arr_0),
	.tdl_arr_8(\gen_blk_float:gen_1_input_bfp_o:delay_next_pass|tdl_arr[8]~q ),
	.clk(clk));

dffeas \del_np_cnt[4] (
	.clk(clk),
	.d(\del_np_cnt[4]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\delay_next_pass_counter~2_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_np_cnt[4]~q ),
	.prn(vcc));
defparam \del_np_cnt[4] .is_wysiwyg = "true";
defparam \del_np_cnt[4] .power_up = "low";

cycloneive_lcell_comb \del_np_cnt[3]~11 (
	.dataa(\del_np_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_np_cnt[2]~10 ),
	.combout(\del_np_cnt[3]~11_combout ),
	.cout(\del_np_cnt[3]~12 ));
defparam \del_np_cnt[3]~11 .lut_mask = 16'h5A5F;
defparam \del_np_cnt[3]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \del_np_cnt[4]~13 (
	.dataa(\del_np_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\del_np_cnt[3]~12 ),
	.combout(\del_np_cnt[4]~13_combout ),
	.cout());
defparam \del_np_cnt[4]~13 .lut_mask = 16'h5A5A;
defparam \del_np_cnt[4]~13 .sum_lutc_input = "cin";

dffeas \slb_i[0] (
	.clk(clk),
	.d(\slb_i~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_i[3]~2_combout ),
	.q(slb_i_0),
	.prn(vcc));
defparam \slb_i[0] .is_wysiwyg = "true";
defparam \slb_i[0] .power_up = "low";

cycloneive_lcell_comb \Mux2~0 (
	.dataa(slb_i_0),
	.datab(\slb_i[1]~q ),
	.datac(\slb_i[2]~q ),
	.datad(\slb_i[3]~q ),
	.cin(gnd),
	.combout(Mux2),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFBFF;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lut_out[0]~0 (
	.dataa(reset_n),
	.datab(Mux2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(lut_out_0),
	.cout());
defparam \lut_out[0]~0 .lut_mask = 16'hEEEE;
defparam \lut_out[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(slb_i_0),
	.datab(\slb_i[1]~q ),
	.datac(\slb_i[2]~q ),
	.datad(\slb_i[3]~q ),
	.cin(gnd),
	.combout(Mux1),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hEFFF;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lut_out[1]~1 (
	.dataa(reset_n),
	.datab(Mux1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(lut_out_1),
	.cout());
defparam \lut_out[1]~1 .lut_mask = 16'hEEEE;
defparam \lut_out[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lut_out[2]~2 (
	.dataa(reset_n),
	.datab(\slb_i[1]~q ),
	.datac(\slb_i[2]~q ),
	.datad(\slb_i[3]~q ),
	.cin(gnd),
	.combout(lut_out_2),
	.cout());
defparam \lut_out[2]~2 .lut_mask = 16'hBFFF;
defparam \lut_out[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lut_out[2]~3 (
	.dataa(lut_out_2),
	.datab(gnd),
	.datac(gnd),
	.datad(slb_i_0),
	.cin(gnd),
	.combout(lut_out_21),
	.cout());
defparam \lut_out[2]~3 .lut_mask = 16'hAAFF;
defparam \lut_out[2]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \del_np_cnt[0]~5 (
	.dataa(\del_np_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\del_np_cnt[0]~5_combout ),
	.cout(\del_np_cnt[0]~6 ));
defparam \del_np_cnt[0]~5 .lut_mask = 16'h55AA;
defparam \del_np_cnt[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \del_np_cnt[1]~7 (
	.dataa(\del_np_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_np_cnt[0]~6 ),
	.combout(\del_np_cnt[1]~7_combout ),
	.cout(\del_np_cnt[1]~8 ));
defparam \del_np_cnt[1]~7 .lut_mask = 16'h5A5F;
defparam \del_np_cnt[1]~7 .sum_lutc_input = "cin";

cycloneive_lcell_comb \del_np_cnt[2]~9 (
	.dataa(\del_np_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_np_cnt[1]~8 ),
	.combout(\del_np_cnt[2]~9_combout ),
	.cout(\del_np_cnt[2]~10 ));
defparam \del_np_cnt[2]~9 .lut_mask = 16'h5AAF;
defparam \del_np_cnt[2]~9 .sum_lutc_input = "cin";

dffeas \del_np_cnt[0] (
	.clk(clk),
	.d(\del_np_cnt[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\delay_next_pass_counter~2_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_np_cnt[0]~q ),
	.prn(vcc));
defparam \del_np_cnt[0] .is_wysiwyg = "true";
defparam \del_np_cnt[0] .power_up = "low";

dffeas \del_np_cnt[1] (
	.clk(clk),
	.d(\del_np_cnt[1]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\delay_next_pass_counter~2_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_np_cnt[1]~q ),
	.prn(vcc));
defparam \del_np_cnt[1] .is_wysiwyg = "true";
defparam \del_np_cnt[1] .power_up = "low";

dffeas \del_np_cnt[3] (
	.clk(clk),
	.d(\del_np_cnt[3]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\delay_next_pass_counter~2_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_np_cnt[3]~q ),
	.prn(vcc));
defparam \del_np_cnt[3] .is_wysiwyg = "true";
defparam \del_np_cnt[3] .power_up = "low";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(\Equal0~0_combout ),
	.datab(\del_np_cnt[0]~q ),
	.datac(\del_np_cnt[1]~q ),
	.datad(\del_np_cnt[3]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hFEFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~0 (
	.dataa(\gen_blk_float:gen_1_input_bfp_o:delay_next_pass|tdl_arr[8]~q ),
	.datab(\sdet.ENABLE~q ),
	.datac(\sdet.DISABLE~q ),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'hFEFF;
defparam \Selector3~0 .sum_lutc_input = "datac";

dffeas \sdet.DISABLE (
	.clk(clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdet.DISABLE~q ),
	.prn(vcc));
defparam \sdet.DISABLE .is_wysiwyg = "true";
defparam \sdet.DISABLE .power_up = "low";

cycloneive_lcell_comb \delay_next_pass_counter~2 (
	.dataa(\sdet.BLOCK_READY~q ),
	.datab(\sdet.DISABLE~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_next_pass_counter~2_combout ),
	.cout());
defparam \delay_next_pass_counter~2 .lut_mask = 16'h7777;
defparam \delay_next_pass_counter~2 .sum_lutc_input = "datac";

dffeas \del_np_cnt[2] (
	.clk(clk),
	.d(\del_np_cnt[2]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\delay_next_pass_counter~2_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_np_cnt[2]~q ),
	.prn(vcc));
defparam \del_np_cnt[2] .is_wysiwyg = "true";
defparam \del_np_cnt[2] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\del_np_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\del_np_cnt[2]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hAAFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\del_np_cnt[3]~q ),
	.datab(\Equal0~0_combout ),
	.datac(\del_np_cnt[0]~q ),
	.datad(\del_np_cnt[1]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hEFFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~0 (
	.dataa(\sdet.BLOCK_READY~q ),
	.datab(\Equal0~1_combout ),
	.datac(\sdet.DISABLE~q ),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hFFFE;
defparam \Selector2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~1 (
	.dataa(\sdet.ENABLE~q ),
	.datab(tdl_arr_01),
	.datac(\gen_blk_float:gen_1_input_bfp_o:delay_next_pass|tdl_arr[8]~q ),
	.datad(\Selector2~0_combout ),
	.cin(gnd),
	.combout(\Selector2~1_combout ),
	.cout());
defparam \Selector2~1 .lut_mask = 16'hFFBF;
defparam \Selector2~1 .sum_lutc_input = "datac";

dffeas \sdet.ENABLE (
	.clk(clk),
	.d(\Selector2~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdet.ENABLE~q ),
	.prn(vcc));
defparam \sdet.ENABLE .is_wysiwyg = "true";
defparam \sdet.ENABLE .power_up = "low";

dffeas en_gain_lut_8_pts(
	.clk(clk),
	.d(\sdet.ENABLE~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\en_gain_lut_8_pts~q ),
	.prn(vcc));
defparam en_gain_lut_8_pts.is_wysiwyg = "true";
defparam en_gain_lut_8_pts.power_up = "low";

cycloneive_lcell_comb \gain_lut_8pts~0 (
	.dataa(real_out_11),
	.datab(real_out_15),
	.datac(pipeline_dffe_27),
	.datad(pipeline_dffe_31),
	.cin(gnd),
	.combout(\gain_lut_8pts~0_combout ),
	.cout());
defparam \gain_lut_8pts~0 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~1 (
	.dataa(reset_n),
	.datab(\en_gain_lut_8_pts~q ),
	.datac(\gain_lut_8pts~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_8pts~1_combout ),
	.cout());
defparam \gain_lut_8pts~1 .lut_mask = 16'hFEFE;
defparam \gain_lut_8pts~1 .sum_lutc_input = "datac";

dffeas \gain_lut_8pts[0] (
	.clk(clk),
	.d(\gain_lut_8pts~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_8pts[0]~q ),
	.prn(vcc));
defparam \gain_lut_8pts[0] .is_wysiwyg = "true";
defparam \gain_lut_8pts[0] .power_up = "low";

cycloneive_lcell_comb \sdet.IDLE~0 (
	.dataa(tdl_arr_01),
	.datab(\sdet.ENABLE~q ),
	.datac(\gen_blk_float:gen_1_input_bfp_o:delay_next_pass|tdl_arr[8]~q ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\sdet.IDLE~0_combout ),
	.cout());
defparam \sdet.IDLE~0 .lut_mask = 16'hFFF7;
defparam \sdet.IDLE~0 .sum_lutc_input = "datac";

dffeas \sdet.IDLE (
	.clk(clk),
	.d(\sdet.IDLE~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdet.IDLE~q ),
	.prn(vcc));
defparam \sdet.IDLE .is_wysiwyg = "true";
defparam \sdet.IDLE .power_up = "low";

cycloneive_lcell_comb \Selector1~0 (
	.dataa(\sdet.BLOCK_READY~q ),
	.datab(gnd),
	.datac(\Equal0~1_combout ),
	.datad(\sdet.IDLE~q ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hAFFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

dffeas \sdet.BLOCK_READY (
	.clk(clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdet.BLOCK_READY~q ),
	.prn(vcc));
defparam \sdet.BLOCK_READY .is_wysiwyg = "true";
defparam \sdet.BLOCK_READY .power_up = "low";

cycloneive_lcell_comb \slb_i[3]~1 (
	.dataa(tdl_arr_01),
	.datab(\sdet.BLOCK_READY~q ),
	.datac(\gen_blk_float:gen_1_input_bfp_o:delay_next_pass3|tdl_arr[2]~q ),
	.datad(\sdet.IDLE~q ),
	.cin(gnd),
	.combout(\slb_i[3]~1_combout ),
	.cout());
defparam \slb_i[3]~1 .lut_mask = 16'hFEFF;
defparam \slb_i[3]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_blk~0 (
	.dataa(\gain_lut_blk[0]~q ),
	.datab(\gain_lut_8pts[0]~q ),
	.datac(gnd),
	.datad(\slb_i[3]~1_combout ),
	.cin(gnd),
	.combout(\gain_lut_blk~0_combout ),
	.cout());
defparam \gain_lut_blk~0 .lut_mask = 16'hEEFF;
defparam \gain_lut_blk~0 .sum_lutc_input = "datac";

dffeas \gain_lut_blk[0] (
	.clk(clk),
	.d(\gain_lut_blk~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_blk[0]~q ),
	.prn(vcc));
defparam \gain_lut_blk[0] .is_wysiwyg = "true";
defparam \gain_lut_blk[0] .power_up = "low";

cycloneive_lcell_comb \slb_i~0 (
	.dataa(\gain_lut_blk[0]~q ),
	.datab(\sdet.BLOCK_READY~q ),
	.datac(gnd),
	.datad(\sdet.IDLE~q ),
	.cin(gnd),
	.combout(\slb_i~0_combout ),
	.cout());
defparam \slb_i~0 .lut_mask = 16'hEEFF;
defparam \slb_i~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \slb_i[3]~2 (
	.dataa(\slb_i[3]~1_combout ),
	.datab(stall_reg),
	.datac(source_valid_ctrl_sop),
	.datad(source_stall_int_d),
	.cin(gnd),
	.combout(\slb_i[3]~2_combout ),
	.cout());
defparam \slb_i[3]~2 .lut_mask = 16'hACFF;
defparam \slb_i[3]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~2 (
	.dataa(real_out_12),
	.datab(real_out_15),
	.datac(pipeline_dffe_28),
	.datad(pipeline_dffe_31),
	.cin(gnd),
	.combout(\gain_lut_8pts~2_combout ),
	.cout());
defparam \gain_lut_8pts~2 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~3 (
	.dataa(reset_n),
	.datab(\en_gain_lut_8_pts~q ),
	.datac(\gain_lut_8pts~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_8pts~3_combout ),
	.cout());
defparam \gain_lut_8pts~3 .lut_mask = 16'hFEFE;
defparam \gain_lut_8pts~3 .sum_lutc_input = "datac";

dffeas \gain_lut_8pts[1] (
	.clk(clk),
	.d(\gain_lut_8pts~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_8pts[1]~q ),
	.prn(vcc));
defparam \gain_lut_8pts[1] .is_wysiwyg = "true";
defparam \gain_lut_8pts[1] .power_up = "low";

cycloneive_lcell_comb \gain_lut_blk~1 (
	.dataa(\gain_lut_blk[1]~q ),
	.datab(\gain_lut_8pts[1]~q ),
	.datac(gnd),
	.datad(\slb_i[3]~1_combout ),
	.cin(gnd),
	.combout(\gain_lut_blk~1_combout ),
	.cout());
defparam \gain_lut_blk~1 .lut_mask = 16'hEEFF;
defparam \gain_lut_blk~1 .sum_lutc_input = "datac";

dffeas \gain_lut_blk[1] (
	.clk(clk),
	.d(\gain_lut_blk~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_blk[1]~q ),
	.prn(vcc));
defparam \gain_lut_blk[1] .is_wysiwyg = "true";
defparam \gain_lut_blk[1] .power_up = "low";

cycloneive_lcell_comb \slb_i~3 (
	.dataa(\sdet.BLOCK_READY~q ),
	.datab(\gain_lut_blk[1]~q ),
	.datac(gnd),
	.datad(\sdet.IDLE~q ),
	.cin(gnd),
	.combout(\slb_i~3_combout ),
	.cout());
defparam \slb_i~3 .lut_mask = 16'hEEFF;
defparam \slb_i~3 .sum_lutc_input = "datac";

dffeas \slb_i[1] (
	.clk(clk),
	.d(\slb_i~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_i[3]~2_combout ),
	.q(\slb_i[1]~q ),
	.prn(vcc));
defparam \slb_i[1] .is_wysiwyg = "true";
defparam \slb_i[1] .power_up = "low";

cycloneive_lcell_comb \gain_lut_8pts~4 (
	.dataa(real_out_13),
	.datab(real_out_15),
	.datac(pipeline_dffe_29),
	.datad(pipeline_dffe_31),
	.cin(gnd),
	.combout(\gain_lut_8pts~4_combout ),
	.cout());
defparam \gain_lut_8pts~4 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~5 (
	.dataa(reset_n),
	.datab(\en_gain_lut_8_pts~q ),
	.datac(\gain_lut_8pts~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_8pts~5_combout ),
	.cout());
defparam \gain_lut_8pts~5 .lut_mask = 16'hFEFE;
defparam \gain_lut_8pts~5 .sum_lutc_input = "datac";

dffeas \gain_lut_8pts[2] (
	.clk(clk),
	.d(\gain_lut_8pts~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_8pts[2]~q ),
	.prn(vcc));
defparam \gain_lut_8pts[2] .is_wysiwyg = "true";
defparam \gain_lut_8pts[2] .power_up = "low";

cycloneive_lcell_comb \gain_lut_blk~2 (
	.dataa(\gain_lut_blk[2]~q ),
	.datab(\gain_lut_8pts[2]~q ),
	.datac(gnd),
	.datad(\slb_i[3]~1_combout ),
	.cin(gnd),
	.combout(\gain_lut_blk~2_combout ),
	.cout());
defparam \gain_lut_blk~2 .lut_mask = 16'hEEFF;
defparam \gain_lut_blk~2 .sum_lutc_input = "datac";

dffeas \gain_lut_blk[2] (
	.clk(clk),
	.d(\gain_lut_blk~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_blk[2]~q ),
	.prn(vcc));
defparam \gain_lut_blk[2] .is_wysiwyg = "true";
defparam \gain_lut_blk[2] .power_up = "low";

cycloneive_lcell_comb \slb_i~4 (
	.dataa(\sdet.BLOCK_READY~q ),
	.datab(\gain_lut_blk[2]~q ),
	.datac(gnd),
	.datad(\sdet.IDLE~q ),
	.cin(gnd),
	.combout(\slb_i~4_combout ),
	.cout());
defparam \slb_i~4 .lut_mask = 16'hEEFF;
defparam \slb_i~4 .sum_lutc_input = "datac";

dffeas \slb_i[2] (
	.clk(clk),
	.d(\slb_i~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_i[3]~2_combout ),
	.q(\slb_i[2]~q ),
	.prn(vcc));
defparam \slb_i[2] .is_wysiwyg = "true";
defparam \slb_i[2] .power_up = "low";

cycloneive_lcell_comb \gain_lut_8pts~6 (
	.dataa(real_out_14),
	.datab(real_out_15),
	.datac(pipeline_dffe_30),
	.datad(pipeline_dffe_31),
	.cin(gnd),
	.combout(\gain_lut_8pts~6_combout ),
	.cout());
defparam \gain_lut_8pts~6 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~7 (
	.dataa(reset_n),
	.datab(\en_gain_lut_8_pts~q ),
	.datac(\gain_lut_8pts~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_8pts~7_combout ),
	.cout());
defparam \gain_lut_8pts~7 .lut_mask = 16'hFEFE;
defparam \gain_lut_8pts~7 .sum_lutc_input = "datac";

dffeas \gain_lut_8pts[3] (
	.clk(clk),
	.d(\gain_lut_8pts~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_8pts[3]~q ),
	.prn(vcc));
defparam \gain_lut_8pts[3] .is_wysiwyg = "true";
defparam \gain_lut_8pts[3] .power_up = "low";

cycloneive_lcell_comb \gain_lut_blk~3 (
	.dataa(\gain_lut_blk[3]~q ),
	.datab(\gain_lut_8pts[3]~q ),
	.datac(gnd),
	.datad(\slb_i[3]~1_combout ),
	.cin(gnd),
	.combout(\gain_lut_blk~3_combout ),
	.cout());
defparam \gain_lut_blk~3 .lut_mask = 16'hEEFF;
defparam \gain_lut_blk~3 .sum_lutc_input = "datac";

dffeas \gain_lut_blk[3] (
	.clk(clk),
	.d(\gain_lut_blk~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_blk[3]~q ),
	.prn(vcc));
defparam \gain_lut_blk[3] .is_wysiwyg = "true";
defparam \gain_lut_blk[3] .power_up = "low";

cycloneive_lcell_comb \slb_i~5 (
	.dataa(\sdet.BLOCK_READY~q ),
	.datab(\gain_lut_blk[3]~q ),
	.datac(gnd),
	.datad(\sdet.IDLE~q ),
	.cin(gnd),
	.combout(\slb_i~5_combout ),
	.cout());
defparam \slb_i~5 .lut_mask = 16'hEEFF;
defparam \slb_i~5 .sum_lutc_input = "datac";

dffeas \slb_i[3] (
	.clk(clk),
	.d(\slb_i~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_i[3]~2_combout ),
	.q(\slb_i[3]~q ),
	.prn(vcc));
defparam \slb_i[3] .is_wysiwyg = "true";
defparam \slb_i[3] .power_up = "low";

endmodule

module fft256_asj_fft_tdl_bit_fft_121_1 (
	global_clock_enable,
	tdl_arr_0,
	tdl_arr_8,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
input 	tdl_arr_0;
output 	tdl_arr_8;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[1]~q ;
wire \tdl_arr[2]~q ;
wire \tdl_arr[3]~q ;
wire \tdl_arr[4]~q ;
wire \tdl_arr[5]~q ;
wire \tdl_arr[6]~q ;
wire \tdl_arr[7]~q ;


dffeas \tdl_arr[8] (
	.clk(clk),
	.d(\tdl_arr[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_8),
	.prn(vcc));
defparam \tdl_arr[8] .is_wysiwyg = "true";
defparam \tdl_arr[8] .power_up = "low";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(tdl_arr_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5]~q ),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

dffeas \tdl_arr[6] (
	.clk(clk),
	.d(\tdl_arr[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[6]~q ),
	.prn(vcc));
defparam \tdl_arr[6] .is_wysiwyg = "true";
defparam \tdl_arr[6] .power_up = "low";

dffeas \tdl_arr[7] (
	.clk(clk),
	.d(\tdl_arr[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[7]~q ),
	.prn(vcc));
defparam \tdl_arr[7] .is_wysiwyg = "true";
defparam \tdl_arr[7] .power_up = "low";

endmodule

module fft256_asj_fft_tdl_bit_fft_121_2 (
	global_clock_enable,
	tdl_arr_2,
	data_in,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_2;
input 	data_in;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0]~q ;
wire \tdl_arr[1]~q ;


dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_2),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(data_in),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

endmodule

module fft256_asj_fft_cmult_can_fft_121 (
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_31,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_161,
	pipeline_dffe_171,
	twiddle_data_real_0,
	twiddle_data_real_15,
	pipeline_dffe_210,
	pipeline_dffe_32,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	pipeline_dffe_121,
	pipeline_dffe_131,
	pipeline_dffe_141,
	pipeline_dffe_151,
	pipeline_dffe_162,
	pipeline_dffe_172,
	twiddle_data_imag_1,
	twiddle_data_imag_2,
	twiddle_data_imag_3,
	twiddle_data_imag_4,
	twiddle_data_imag_5,
	twiddle_data_imag_6,
	twiddle_data_imag_7,
	twiddle_data_imag_8,
	twiddle_data_imag_9,
	twiddle_data_imag_10,
	twiddle_data_imag_11,
	twiddle_data_imag_12,
	twiddle_data_imag_13,
	twiddle_data_imag_14,
	twiddle_data_imag_15,
	global_clock_enable,
	real_out_0,
	real_out_1,
	real_out_2,
	real_out_3,
	real_out_4,
	real_out_5,
	real_out_6,
	real_out_7,
	real_out_8,
	real_out_9,
	real_out_10,
	real_out_11,
	real_out_12,
	real_out_13,
	real_out_14,
	real_out_15,
	twiddle_data_real_1,
	twiddle_data_real_2,
	twiddle_data_real_3,
	twiddle_data_real_4,
	twiddle_data_real_5,
	twiddle_data_real_6,
	twiddle_data_real_7,
	twiddle_data_real_8,
	twiddle_data_real_9,
	twiddle_data_real_10,
	twiddle_data_real_11,
	twiddle_data_real_12,
	twiddle_data_real_13,
	twiddle_data_real_14,
	twiddle_data_imag_0,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_31;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_12;
input 	pipeline_dffe_13;
input 	pipeline_dffe_14;
input 	pipeline_dffe_15;
input 	pipeline_dffe_161;
input 	pipeline_dffe_171;
input 	twiddle_data_real_0;
input 	twiddle_data_real_15;
input 	pipeline_dffe_210;
input 	pipeline_dffe_32;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	pipeline_dffe_121;
input 	pipeline_dffe_131;
input 	pipeline_dffe_141;
input 	pipeline_dffe_151;
input 	pipeline_dffe_162;
input 	pipeline_dffe_172;
input 	twiddle_data_imag_1;
input 	twiddle_data_imag_2;
input 	twiddle_data_imag_3;
input 	twiddle_data_imag_4;
input 	twiddle_data_imag_5;
input 	twiddle_data_imag_6;
input 	twiddle_data_imag_7;
input 	twiddle_data_imag_8;
input 	twiddle_data_imag_9;
input 	twiddle_data_imag_10;
input 	twiddle_data_imag_11;
input 	twiddle_data_imag_12;
input 	twiddle_data_imag_13;
input 	twiddle_data_imag_14;
input 	twiddle_data_imag_15;
input 	global_clock_enable;
output 	real_out_0;
output 	real_out_1;
output 	real_out_2;
output 	real_out_3;
output 	real_out_4;
output 	real_out_5;
output 	real_out_6;
output 	real_out_7;
output 	real_out_8;
output 	real_out_9;
output 	real_out_10;
output 	real_out_11;
output 	real_out_12;
output 	real_out_13;
output 	real_out_14;
output 	real_out_15;
input 	twiddle_data_real_1;
input 	twiddle_data_real_2;
input 	twiddle_data_real_3;
input 	twiddle_data_real_4;
input 	twiddle_data_real_5;
input 	twiddle_data_real_6;
input 	twiddle_data_real_7;
input 	twiddle_data_real_8;
input 	twiddle_data_real_9;
input 	twiddle_data_real_10;
input 	twiddle_data_real_11;
input 	twiddle_data_real_12;
input 	twiddle_data_real_13;
input 	twiddle_data_real_14;
input 	twiddle_data_imag_0;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ;
wire \result_imag_1[16]~q ;
wire \result_imag_1[15]~q ;
wire \result_imag_1[14]~q ;
wire \result_imag_1[13]~q ;
wire \result_imag_1[12]~q ;
wire \result_imag_1[11]~q ;
wire \result_imag_1[10]~q ;
wire \result_imag_1[9]~q ;
wire \result_imag_1[8]~q ;
wire \result_imag_1[7]~q ;
wire \result_imag_1[6]~q ;
wire \result_imag_1[5]~q ;
wire \result_imag_1[4]~q ;
wire \result_imag_1[3]~q ;
wire \result_imag_1[2]~q ;
wire \result_imag_1[1]~q ;
wire \result_imag_1[0]~q ;
wire \result_imag_1[31]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ;
wire \result_imag_1[17]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ;
wire \result_imag_1[18]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ;
wire \result_imag_1[19]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~q ;
wire \result_imag_1[20]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~q ;
wire \result_imag_1[21]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~q ;
wire \result_imag_1[22]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~q ;
wire \result_imag_1[23]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~q ;
wire \result_imag_1[24]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~q ;
wire \result_imag_1[25]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~q ;
wire \result_imag_1[26]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~q ;
wire \result_imag_1[27]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~q ;
wire \result_imag_1[28]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~q ;
wire \result_imag_1[29]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~q ;
wire \result_imag_1[30]~q ;
wire \gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~q ;
wire \result_real_1_tmp[16]~q ;
wire \result_real_1_tmp[15]~q ;
wire \result_real_1_tmp[14]~q ;
wire \result_real_1_tmp[13]~q ;
wire \result_real_1_tmp[12]~q ;
wire \result_real_1_tmp[11]~q ;
wire \result_real_1_tmp[10]~q ;
wire \result_real_1_tmp[9]~q ;
wire \result_real_1_tmp[8]~q ;
wire \result_real_1_tmp[7]~q ;
wire \result_real_1_tmp[6]~q ;
wire \result_real_1_tmp[5]~q ;
wire \result_real_1_tmp[4]~q ;
wire \result_real_1_tmp[3]~q ;
wire \result_real_1_tmp[2]~q ;
wire \result_real_1_tmp[1]~q ;
wire \result_real_1_tmp[0]~q ;
wire \result_real_1_tmp[31]~q ;
wire \addresult_ac_bd[16]~q ;
wire \addresult_ac_bd[15]~q ;
wire \addresult_ac_bd[14]~q ;
wire \addresult_ac_bd[13]~q ;
wire \addresult_ac_bd[12]~q ;
wire \addresult_ac_bd[11]~q ;
wire \addresult_ac_bd[10]~q ;
wire \addresult_ac_bd[9]~q ;
wire \addresult_ac_bd[8]~q ;
wire \addresult_ac_bd[7]~q ;
wire \addresult_ac_bd[6]~q ;
wire \addresult_ac_bd[5]~q ;
wire \addresult_ac_bd[4]~q ;
wire \addresult_ac_bd[3]~q ;
wire \addresult_ac_bd[2]~q ;
wire \addresult_ac_bd[1]~q ;
wire \addresult_ac_bd[0]~q ;
wire \result_imag_1[0]~33 ;
wire \result_imag_1[0]~32_combout ;
wire \result_imag_1[1]~35 ;
wire \result_imag_1[1]~34_combout ;
wire \result_imag_1[2]~37 ;
wire \result_imag_1[2]~36_combout ;
wire \result_imag_1[3]~39 ;
wire \result_imag_1[3]~38_combout ;
wire \result_imag_1[4]~41 ;
wire \result_imag_1[4]~40_combout ;
wire \result_imag_1[5]~43 ;
wire \result_imag_1[5]~42_combout ;
wire \result_imag_1[6]~45 ;
wire \result_imag_1[6]~44_combout ;
wire \result_imag_1[7]~47 ;
wire \result_imag_1[7]~46_combout ;
wire \result_imag_1[8]~49 ;
wire \result_imag_1[8]~48_combout ;
wire \result_imag_1[9]~51 ;
wire \result_imag_1[9]~50_combout ;
wire \result_imag_1[10]~53 ;
wire \result_imag_1[10]~52_combout ;
wire \result_imag_1[11]~55 ;
wire \result_imag_1[11]~54_combout ;
wire \result_imag_1[12]~57 ;
wire \result_imag_1[12]~56_combout ;
wire \result_imag_1[13]~59 ;
wire \result_imag_1[13]~58_combout ;
wire \result_imag_1[14]~61 ;
wire \result_imag_1[14]~60_combout ;
wire \result_imag_1[15]~63 ;
wire \result_imag_1[15]~62_combout ;
wire \result_imag_1[16]~65 ;
wire \result_imag_1[16]~64_combout ;
wire \addresult_ac_bd[31]~q ;
wire \addresult_ac_bd[30]~q ;
wire \addresult_ac_bd[29]~q ;
wire \addresult_ac_bd[28]~q ;
wire \addresult_ac_bd[27]~q ;
wire \addresult_ac_bd[26]~q ;
wire \addresult_ac_bd[25]~q ;
wire \addresult_ac_bd[24]~q ;
wire \addresult_ac_bd[23]~q ;
wire \addresult_ac_bd[22]~q ;
wire \addresult_ac_bd[21]~q ;
wire \addresult_ac_bd[20]~q ;
wire \addresult_ac_bd[19]~q ;
wire \addresult_ac_bd[18]~q ;
wire \addresult_ac_bd[17]~q ;
wire \result_imag_1[17]~67 ;
wire \result_imag_1[17]~66_combout ;
wire \result_imag_1[18]~69 ;
wire \result_imag_1[18]~68_combout ;
wire \result_imag_1[19]~71 ;
wire \result_imag_1[19]~70_combout ;
wire \result_imag_1[20]~73 ;
wire \result_imag_1[20]~72_combout ;
wire \result_imag_1[21]~75 ;
wire \result_imag_1[21]~74_combout ;
wire \result_imag_1[22]~77 ;
wire \result_imag_1[22]~76_combout ;
wire \result_imag_1[23]~79 ;
wire \result_imag_1[23]~78_combout ;
wire \result_imag_1[24]~81 ;
wire \result_imag_1[24]~80_combout ;
wire \result_imag_1[25]~83 ;
wire \result_imag_1[25]~82_combout ;
wire \result_imag_1[26]~85 ;
wire \result_imag_1[26]~84_combout ;
wire \result_imag_1[27]~87 ;
wire \result_imag_1[27]~86_combout ;
wire \result_imag_1[28]~89 ;
wire \result_imag_1[28]~88_combout ;
wire \result_imag_1[29]~91 ;
wire \result_imag_1[29]~90_combout ;
wire \result_imag_1[30]~93 ;
wire \result_imag_1[30]~92_combout ;
wire \result_imag_1[31]~94_combout ;
wire \result_real_1_tmp[17]~q ;
wire \result_real_1_tmp[18]~q ;
wire \result_real_1_tmp[19]~q ;
wire \result_real_1_tmp[20]~q ;
wire \result_real_1_tmp[21]~q ;
wire \result_real_1_tmp[22]~q ;
wire \result_real_1_tmp[23]~q ;
wire \result_real_1_tmp[24]~q ;
wire \result_real_1_tmp[25]~q ;
wire \result_real_1_tmp[26]~q ;
wire \result_real_1_tmp[27]~q ;
wire \result_real_1_tmp[28]~q ;
wire \result_real_1_tmp[29]~q ;
wire \result_real_1_tmp[30]~q ;
wire \result_real_1_tmp[0]~33 ;
wire \result_real_1_tmp[0]~32_combout ;
wire \result_real_1_tmp[1]~35 ;
wire \result_real_1_tmp[1]~34_combout ;
wire \result_real_1_tmp[2]~37 ;
wire \result_real_1_tmp[2]~36_combout ;
wire \result_real_1_tmp[3]~39 ;
wire \result_real_1_tmp[3]~38_combout ;
wire \result_real_1_tmp[4]~41 ;
wire \result_real_1_tmp[4]~40_combout ;
wire \result_real_1_tmp[5]~43 ;
wire \result_real_1_tmp[5]~42_combout ;
wire \result_real_1_tmp[6]~45 ;
wire \result_real_1_tmp[6]~44_combout ;
wire \result_real_1_tmp[7]~47 ;
wire \result_real_1_tmp[7]~46_combout ;
wire \result_real_1_tmp[8]~49 ;
wire \result_real_1_tmp[8]~48_combout ;
wire \result_real_1_tmp[9]~51 ;
wire \result_real_1_tmp[9]~50_combout ;
wire \result_real_1_tmp[10]~53 ;
wire \result_real_1_tmp[10]~52_combout ;
wire \result_real_1_tmp[11]~55 ;
wire \result_real_1_tmp[11]~54_combout ;
wire \result_real_1_tmp[12]~57 ;
wire \result_real_1_tmp[12]~56_combout ;
wire \result_real_1_tmp[13]~59 ;
wire \result_real_1_tmp[13]~58_combout ;
wire \result_real_1_tmp[14]~61 ;
wire \result_real_1_tmp[14]~60_combout ;
wire \result_real_1_tmp[15]~63 ;
wire \result_real_1_tmp[15]~62_combout ;
wire \result_real_1_tmp[16]~65 ;
wire \result_real_1_tmp[16]~64_combout ;
wire \result_real_1_tmp[17]~67 ;
wire \result_real_1_tmp[17]~66_combout ;
wire \result_real_1_tmp[18]~69 ;
wire \result_real_1_tmp[18]~68_combout ;
wire \result_real_1_tmp[19]~71 ;
wire \result_real_1_tmp[19]~70_combout ;
wire \result_real_1_tmp[20]~73 ;
wire \result_real_1_tmp[20]~72_combout ;
wire \result_real_1_tmp[21]~75 ;
wire \result_real_1_tmp[21]~74_combout ;
wire \result_real_1_tmp[22]~77 ;
wire \result_real_1_tmp[22]~76_combout ;
wire \result_real_1_tmp[23]~79 ;
wire \result_real_1_tmp[23]~78_combout ;
wire \result_real_1_tmp[24]~81 ;
wire \result_real_1_tmp[24]~80_combout ;
wire \result_real_1_tmp[25]~83 ;
wire \result_real_1_tmp[25]~82_combout ;
wire \result_real_1_tmp[26]~85 ;
wire \result_real_1_tmp[26]~84_combout ;
wire \result_real_1_tmp[27]~87 ;
wire \result_real_1_tmp[27]~86_combout ;
wire \result_real_1_tmp[28]~89 ;
wire \result_real_1_tmp[28]~88_combout ;
wire \result_real_1_tmp[29]~91 ;
wire \result_real_1_tmp[29]~90_combout ;
wire \result_real_1_tmp[30]~93 ;
wire \result_real_1_tmp[30]~92_combout ;
wire \result_real_1_tmp[31]~94_combout ;
wire \addresult_ac_bd[0]~33 ;
wire \addresult_ac_bd[0]~32_combout ;
wire \addresult_ac_bd[1]~35 ;
wire \addresult_ac_bd[1]~34_combout ;
wire \addresult_ac_bd[2]~37 ;
wire \addresult_ac_bd[2]~36_combout ;
wire \addresult_ac_bd[3]~39 ;
wire \addresult_ac_bd[3]~38_combout ;
wire \addresult_ac_bd[4]~41 ;
wire \addresult_ac_bd[4]~40_combout ;
wire \addresult_ac_bd[5]~43 ;
wire \addresult_ac_bd[5]~42_combout ;
wire \addresult_ac_bd[6]~45 ;
wire \addresult_ac_bd[6]~44_combout ;
wire \addresult_ac_bd[7]~47 ;
wire \addresult_ac_bd[7]~46_combout ;
wire \addresult_ac_bd[8]~49 ;
wire \addresult_ac_bd[8]~48_combout ;
wire \addresult_ac_bd[9]~51 ;
wire \addresult_ac_bd[9]~50_combout ;
wire \addresult_ac_bd[10]~53 ;
wire \addresult_ac_bd[10]~52_combout ;
wire \addresult_ac_bd[11]~55 ;
wire \addresult_ac_bd[11]~54_combout ;
wire \addresult_ac_bd[12]~57 ;
wire \addresult_ac_bd[12]~56_combout ;
wire \addresult_ac_bd[13]~59 ;
wire \addresult_ac_bd[13]~58_combout ;
wire \addresult_ac_bd[14]~61 ;
wire \addresult_ac_bd[14]~60_combout ;
wire \addresult_ac_bd[15]~63 ;
wire \addresult_ac_bd[15]~62_combout ;
wire \addresult_ac_bd[16]~65 ;
wire \addresult_ac_bd[16]~64_combout ;
wire \addresult_ac_bd[17]~67 ;
wire \addresult_ac_bd[17]~66_combout ;
wire \addresult_ac_bd[18]~69 ;
wire \addresult_ac_bd[18]~68_combout ;
wire \addresult_ac_bd[19]~71 ;
wire \addresult_ac_bd[19]~70_combout ;
wire \addresult_ac_bd[20]~73 ;
wire \addresult_ac_bd[20]~72_combout ;
wire \addresult_ac_bd[21]~75 ;
wire \addresult_ac_bd[21]~74_combout ;
wire \addresult_ac_bd[22]~77 ;
wire \addresult_ac_bd[22]~76_combout ;
wire \addresult_ac_bd[23]~79 ;
wire \addresult_ac_bd[23]~78_combout ;
wire \addresult_ac_bd[24]~81 ;
wire \addresult_ac_bd[24]~80_combout ;
wire \addresult_ac_bd[25]~83 ;
wire \addresult_ac_bd[25]~82_combout ;
wire \addresult_ac_bd[26]~85 ;
wire \addresult_ac_bd[26]~84_combout ;
wire \addresult_ac_bd[27]~87 ;
wire \addresult_ac_bd[27]~86_combout ;
wire \addresult_ac_bd[28]~89 ;
wire \addresult_ac_bd[28]~88_combout ;
wire \addresult_ac_bd[29]~91 ;
wire \addresult_ac_bd[29]~90_combout ;
wire \addresult_ac_bd[30]~93 ;
wire \addresult_ac_bd[30]~92_combout ;
wire \addresult_ac_bd[31]~94_combout ;
wire \addresult_a_b[0]~q ;
wire \addresult_a_b[1]~q ;
wire \addresult_a_b[2]~q ;
wire \addresult_a_b[3]~q ;
wire \addresult_a_b[4]~q ;
wire \addresult_a_b[5]~q ;
wire \addresult_a_b[6]~q ;
wire \addresult_a_b[7]~q ;
wire \addresult_a_b[8]~q ;
wire \addresult_a_b[9]~q ;
wire \addresult_a_b[10]~q ;
wire \addresult_a_b[11]~q ;
wire \addresult_a_b[12]~q ;
wire \addresult_a_b[13]~q ;
wire \addresult_a_b[14]~q ;
wire \addresult_a_b[15]~q ;
wire \addresult_a_b[16]~q ;
wire \addresult_c_d[0]~q ;
wire \addresult_c_d[1]~q ;
wire \addresult_c_d[2]~q ;
wire \addresult_c_d[3]~q ;
wire \addresult_c_d[4]~q ;
wire \addresult_c_d[5]~q ;
wire \addresult_c_d[6]~q ;
wire \addresult_c_d[7]~q ;
wire \addresult_c_d[8]~q ;
wire \addresult_c_d[9]~q ;
wire \addresult_c_d[10]~q ;
wire \addresult_c_d[11]~q ;
wire \addresult_c_d[12]~q ;
wire \addresult_c_d[13]~q ;
wire \addresult_c_d[14]~q ;
wire \addresult_c_d[15]~q ;
wire \addresult_c_d[16]~q ;
wire \addresult_a_b[0]~18 ;
wire \addresult_a_b[0]~17_combout ;
wire \addresult_a_b[1]~20 ;
wire \addresult_a_b[1]~19_combout ;
wire \addresult_a_b[2]~22 ;
wire \addresult_a_b[2]~21_combout ;
wire \addresult_a_b[3]~24 ;
wire \addresult_a_b[3]~23_combout ;
wire \addresult_a_b[4]~26 ;
wire \addresult_a_b[4]~25_combout ;
wire \addresult_a_b[5]~28 ;
wire \addresult_a_b[5]~27_combout ;
wire \addresult_a_b[6]~30 ;
wire \addresult_a_b[6]~29_combout ;
wire \addresult_a_b[7]~32 ;
wire \addresult_a_b[7]~31_combout ;
wire \addresult_a_b[8]~34 ;
wire \addresult_a_b[8]~33_combout ;
wire \addresult_a_b[9]~36 ;
wire \addresult_a_b[9]~35_combout ;
wire \addresult_a_b[10]~38 ;
wire \addresult_a_b[10]~37_combout ;
wire \addresult_a_b[11]~40 ;
wire \addresult_a_b[11]~39_combout ;
wire \addresult_a_b[12]~42 ;
wire \addresult_a_b[12]~41_combout ;
wire \addresult_a_b[13]~44 ;
wire \addresult_a_b[13]~43_combout ;
wire \addresult_a_b[14]~46 ;
wire \addresult_a_b[14]~45_combout ;
wire \addresult_a_b[15]~48 ;
wire \addresult_a_b[15]~47_combout ;
wire \addresult_a_b[16]~49_combout ;
wire \addresult_c_d[0]~18 ;
wire \addresult_c_d[0]~17_combout ;
wire \addresult_c_d[1]~20 ;
wire \addresult_c_d[1]~19_combout ;
wire \addresult_c_d[2]~22 ;
wire \addresult_c_d[2]~21_combout ;
wire \addresult_c_d[3]~24 ;
wire \addresult_c_d[3]~23_combout ;
wire \addresult_c_d[4]~26 ;
wire \addresult_c_d[4]~25_combout ;
wire \addresult_c_d[5]~28 ;
wire \addresult_c_d[5]~27_combout ;
wire \addresult_c_d[6]~30 ;
wire \addresult_c_d[6]~29_combout ;
wire \addresult_c_d[7]~32 ;
wire \addresult_c_d[7]~31_combout ;
wire \addresult_c_d[8]~34 ;
wire \addresult_c_d[8]~33_combout ;
wire \addresult_c_d[9]~36 ;
wire \addresult_c_d[9]~35_combout ;
wire \addresult_c_d[10]~38 ;
wire \addresult_c_d[10]~37_combout ;
wire \addresult_c_d[11]~40 ;
wire \addresult_c_d[11]~39_combout ;
wire \addresult_c_d[12]~42 ;
wire \addresult_c_d[12]~41_combout ;
wire \addresult_c_d[13]~44 ;
wire \addresult_c_d[13]~43_combout ;
wire \addresult_c_d[14]~46 ;
wire \addresult_c_d[14]~45_combout ;
wire \addresult_c_d[15]~48 ;
wire \addresult_c_d[15]~47_combout ;
wire \addresult_c_d[16]~49_combout ;
wire \result_a_b_c_d_se[16]~q ;
wire \result_a_b_c_d_se[15]~q ;
wire \result_a_b_c_d_se[14]~q ;
wire \result_a_b_c_d_se[13]~q ;
wire \result_a_b_c_d_se[12]~q ;
wire \result_a_b_c_d_se[11]~q ;
wire \result_a_b_c_d_se[10]~q ;
wire \result_a_b_c_d_se[9]~q ;
wire \result_a_b_c_d_se[8]~q ;
wire \result_a_b_c_d_se[7]~q ;
wire \result_a_b_c_d_se[6]~q ;
wire \result_a_b_c_d_se[5]~q ;
wire \result_a_b_c_d_se[4]~q ;
wire \result_a_b_c_d_se[3]~q ;
wire \result_a_b_c_d_se[2]~q ;
wire \result_a_b_c_d_se[1]~q ;
wire \result_a_b_c_d_se[0]~q ;
wire \result_a_b_c_d_se[31]~q ;
wire \result_a_b_c_d_se[30]~q ;
wire \result_a_b_c_d_se[29]~q ;
wire \result_a_b_c_d_se[28]~q ;
wire \result_a_b_c_d_se[27]~q ;
wire \result_a_b_c_d_se[26]~q ;
wire \result_a_b_c_d_se[25]~q ;
wire \result_a_b_c_d_se[24]~q ;
wire \result_a_b_c_d_se[23]~q ;
wire \result_a_b_c_d_se[22]~q ;
wire \result_a_b_c_d_se[21]~q ;
wire \result_a_b_c_d_se[20]~q ;
wire \result_a_b_c_d_se[19]~q ;
wire \result_a_b_c_d_se[18]~q ;
wire \result_a_b_c_d_se[17]~q ;
wire \result_a_c_se[16]~q ;
wire \result_b_d_se[16]~q ;
wire \result_a_c_se[15]~q ;
wire \result_b_d_se[15]~q ;
wire \result_a_c_se[14]~q ;
wire \result_b_d_se[14]~q ;
wire \result_a_c_se[13]~q ;
wire \result_b_d_se[13]~q ;
wire \result_a_c_se[12]~q ;
wire \result_b_d_se[12]~q ;
wire \result_a_c_se[11]~q ;
wire \result_b_d_se[11]~q ;
wire \result_a_c_se[10]~q ;
wire \result_b_d_se[10]~q ;
wire \result_a_c_se[9]~q ;
wire \result_b_d_se[9]~q ;
wire \result_a_c_se[8]~q ;
wire \result_b_d_se[8]~q ;
wire \result_a_c_se[7]~q ;
wire \result_b_d_se[7]~q ;
wire \result_a_c_se[6]~q ;
wire \result_b_d_se[6]~q ;
wire \result_a_c_se[5]~q ;
wire \result_b_d_se[5]~q ;
wire \result_a_c_se[4]~q ;
wire \result_b_d_se[4]~q ;
wire \result_a_c_se[3]~q ;
wire \result_b_d_se[3]~q ;
wire \result_a_c_se[2]~q ;
wire \result_b_d_se[2]~q ;
wire \result_a_c_se[1]~q ;
wire \result_b_d_se[1]~q ;
wire \result_a_c_se[0]~q ;
wire \result_b_d_se[0]~q ;
wire \result_a_c_se[31]~q ;
wire \result_b_d_se[31]~q ;
wire \result_a_c_se[30]~q ;
wire \result_b_d_se[30]~q ;
wire \result_a_c_se[29]~q ;
wire \result_b_d_se[29]~q ;
wire \result_a_c_se[28]~q ;
wire \result_b_d_se[28]~q ;
wire \result_a_c_se[27]~q ;
wire \result_b_d_se[27]~q ;
wire \result_a_c_se[26]~q ;
wire \result_b_d_se[26]~q ;
wire \result_a_c_se[25]~q ;
wire \result_b_d_se[25]~q ;
wire \result_a_c_se[24]~q ;
wire \result_b_d_se[24]~q ;
wire \result_a_c_se[23]~q ;
wire \result_b_d_se[23]~q ;
wire \result_a_c_se[22]~q ;
wire \result_b_d_se[22]~q ;
wire \result_a_c_se[21]~q ;
wire \result_b_d_se[21]~q ;
wire \result_a_c_se[20]~q ;
wire \result_b_d_se[20]~q ;
wire \result_a_c_se[19]~q ;
wire \result_b_d_se[19]~q ;
wire \result_a_c_se[18]~q ;
wire \result_b_d_se[18]~q ;
wire \result_a_c_se[17]~q ;
wire \result_b_d_se[17]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[16]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[15]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[14]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[13]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[12]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[11]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[10]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[9]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[8]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[7]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[6]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[5]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[4]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[3]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[2]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[1]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[0]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[31]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[30]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[29]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[28]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[27]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[26]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[25]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[24]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[23]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[22]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[21]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[20]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[19]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[18]~q ;
wire \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[17]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[16]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[16]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[15]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[15]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[14]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[14]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[13]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[13]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[12]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[12]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[11]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[11]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[10]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[10]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[9]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[9]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[8]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[8]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[7]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[7]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[6]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[6]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[5]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[5]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[4]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[4]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[3]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[3]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[2]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[2]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[1]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[1]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[0]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[0]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[31]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[31]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[30]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[30]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[29]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[29]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[28]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[28]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[27]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[27]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[26]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[26]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[25]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[25]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[24]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[24]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[23]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[23]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[22]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[22]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[21]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[21]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[20]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[20]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[19]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[19]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[18]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[18]~q ;
wire \gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[17]~q ;
wire \gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[17]~q ;


fft256_asj_fft_pround_fft_121_1 \gen_unsc:u1 (
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_31(pipeline_dffe_31),
	.result_imag_1_16(\result_imag_1[16]~q ),
	.result_imag_1_15(\result_imag_1[15]~q ),
	.result_imag_1_14(\result_imag_1[14]~q ),
	.result_imag_1_13(\result_imag_1[13]~q ),
	.result_imag_1_12(\result_imag_1[12]~q ),
	.result_imag_1_11(\result_imag_1[11]~q ),
	.result_imag_1_10(\result_imag_1[10]~q ),
	.result_imag_1_9(\result_imag_1[9]~q ),
	.result_imag_1_8(\result_imag_1[8]~q ),
	.result_imag_1_7(\result_imag_1[7]~q ),
	.result_imag_1_6(\result_imag_1[6]~q ),
	.result_imag_1_5(\result_imag_1[5]~q ),
	.result_imag_1_4(\result_imag_1[4]~q ),
	.result_imag_1_3(\result_imag_1[3]~q ),
	.result_imag_1_2(\result_imag_1[2]~q ),
	.result_imag_1_1(\result_imag_1[1]~q ),
	.result_imag_1_0(\result_imag_1[0]~q ),
	.result_imag_1_31(\result_imag_1[31]~q ),
	.result_imag_1_17(\result_imag_1[17]~q ),
	.result_imag_1_18(\result_imag_1[18]~q ),
	.result_imag_1_19(\result_imag_1[19]~q ),
	.result_imag_1_20(\result_imag_1[20]~q ),
	.result_imag_1_21(\result_imag_1[21]~q ),
	.result_imag_1_22(\result_imag_1[22]~q ),
	.result_imag_1_23(\result_imag_1[23]~q ),
	.result_imag_1_24(\result_imag_1[24]~q ),
	.result_imag_1_25(\result_imag_1[25]~q ),
	.result_imag_1_26(\result_imag_1[26]~q ),
	.result_imag_1_27(\result_imag_1[27]~q ),
	.result_imag_1_28(\result_imag_1[28]~q ),
	.result_imag_1_29(\result_imag_1[29]~q ),
	.result_imag_1_30(\result_imag_1[30]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fft256_asj_fft_pround_fft_121 \gen_unsc:u0 (
	.pipeline_dffe_16(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_18(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_19(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_20(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_21(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_22(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_23(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~q ),
	.pipeline_dffe_24(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~q ),
	.pipeline_dffe_25(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~q ),
	.pipeline_dffe_26(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~q ),
	.pipeline_dffe_27(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_28(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_29(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_30(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_31(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~q ),
	.result_real_1_tmp_16(\result_real_1_tmp[16]~q ),
	.result_real_1_tmp_15(\result_real_1_tmp[15]~q ),
	.result_real_1_tmp_14(\result_real_1_tmp[14]~q ),
	.result_real_1_tmp_13(\result_real_1_tmp[13]~q ),
	.result_real_1_tmp_12(\result_real_1_tmp[12]~q ),
	.result_real_1_tmp_11(\result_real_1_tmp[11]~q ),
	.result_real_1_tmp_10(\result_real_1_tmp[10]~q ),
	.result_real_1_tmp_9(\result_real_1_tmp[9]~q ),
	.result_real_1_tmp_8(\result_real_1_tmp[8]~q ),
	.result_real_1_tmp_7(\result_real_1_tmp[7]~q ),
	.result_real_1_tmp_6(\result_real_1_tmp[6]~q ),
	.result_real_1_tmp_5(\result_real_1_tmp[5]~q ),
	.result_real_1_tmp_4(\result_real_1_tmp[4]~q ),
	.result_real_1_tmp_3(\result_real_1_tmp[3]~q ),
	.result_real_1_tmp_2(\result_real_1_tmp[2]~q ),
	.result_real_1_tmp_1(\result_real_1_tmp[1]~q ),
	.result_real_1_tmp_0(\result_real_1_tmp[0]~q ),
	.result_real_1_tmp_31(\result_real_1_tmp[31]~q ),
	.result_real_1_tmp_17(\result_real_1_tmp[17]~q ),
	.result_real_1_tmp_18(\result_real_1_tmp[18]~q ),
	.result_real_1_tmp_19(\result_real_1_tmp[19]~q ),
	.result_real_1_tmp_20(\result_real_1_tmp[20]~q ),
	.result_real_1_tmp_21(\result_real_1_tmp[21]~q ),
	.result_real_1_tmp_22(\result_real_1_tmp[22]~q ),
	.result_real_1_tmp_23(\result_real_1_tmp[23]~q ),
	.result_real_1_tmp_24(\result_real_1_tmp[24]~q ),
	.result_real_1_tmp_25(\result_real_1_tmp[25]~q ),
	.result_real_1_tmp_26(\result_real_1_tmp[26]~q ),
	.result_real_1_tmp_27(\result_real_1_tmp[27]~q ),
	.result_real_1_tmp_28(\result_real_1_tmp[28]~q ),
	.result_real_1_tmp_29(\result_real_1_tmp[29]~q ),
	.result_real_1_tmp_30(\result_real_1_tmp[30]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fft256_LPM_MULT_1 \gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d (
	.dataa({\addresult_a_b[16]~q ,\addresult_a_b[15]~q ,\addresult_a_b[14]~q ,\addresult_a_b[13]~q ,\addresult_a_b[12]~q ,\addresult_a_b[11]~q ,\addresult_a_b[10]~q ,\addresult_a_b[9]~q ,\addresult_a_b[8]~q ,\addresult_a_b[7]~q ,\addresult_a_b[6]~q ,\addresult_a_b[5]~q ,
\addresult_a_b[4]~q ,\addresult_a_b[3]~q ,\addresult_a_b[2]~q ,\addresult_a_b[1]~q ,\addresult_a_b[0]~q }),
	.datab({\addresult_c_d[16]~q ,\addresult_c_d[15]~q ,\addresult_c_d[14]~q ,\addresult_c_d[13]~q ,\addresult_c_d[12]~q ,\addresult_c_d[11]~q ,\addresult_c_d[10]~q ,\addresult_c_d[9]~q ,\addresult_c_d[8]~q ,\addresult_c_d[7]~q ,\addresult_c_d[6]~q ,\addresult_c_d[5]~q ,
\addresult_c_d[4]~q ,\addresult_c_d[3]~q ,\addresult_c_d[2]~q ,\addresult_c_d[1]~q ,\addresult_c_d[0]~q }),
	.clken(global_clock_enable),
	.dffe3a_16(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[16]~q ),
	.dffe3a_15(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[15]~q ),
	.dffe3a_14(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[14]~q ),
	.dffe3a_13(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[13]~q ),
	.dffe3a_12(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[12]~q ),
	.dffe3a_11(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[11]~q ),
	.dffe3a_10(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[10]~q ),
	.dffe3a_9(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[9]~q ),
	.dffe3a_8(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[8]~q ),
	.dffe3a_7(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[7]~q ),
	.dffe3a_6(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[6]~q ),
	.dffe3a_5(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[5]~q ),
	.dffe3a_4(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[4]~q ),
	.dffe3a_3(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[3]~q ),
	.dffe3a_2(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[2]~q ),
	.dffe3a_1(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[1]~q ),
	.dffe3a_0(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[0]~q ),
	.dffe3a_31(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[31]~q ),
	.dffe3a_30(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[30]~q ),
	.dffe3a_29(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[29]~q ),
	.dffe3a_28(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[28]~q ),
	.dffe3a_27(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[27]~q ),
	.dffe3a_26(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[26]~q ),
	.dffe3a_25(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[25]~q ),
	.dffe3a_24(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[24]~q ),
	.dffe3a_23(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[23]~q ),
	.dffe3a_22(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[22]~q ),
	.dffe3a_21(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[21]~q ),
	.dffe3a_20(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[20]~q ),
	.dffe3a_19(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[19]~q ),
	.dffe3a_18(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[18]~q ),
	.dffe3a_17(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[17]~q ),
	.clock(clk));

fft256_LPM_MULT_3 \gen_ded_m1:gen_unext_m_bd:m_bd (
	.dataa({gnd,pipeline_dffe_172,pipeline_dffe_162,pipeline_dffe_151,pipeline_dffe_141,pipeline_dffe_131,pipeline_dffe_121,pipeline_dffe_111,pipeline_dffe_101,pipeline_dffe_91,pipeline_dffe_81,pipeline_dffe_71,pipeline_dffe_61,pipeline_dffe_51,pipeline_dffe_41,pipeline_dffe_32,
pipeline_dffe_210}),
	.datab({gnd,twiddle_data_imag_15,twiddle_data_imag_14,twiddle_data_imag_13,twiddle_data_imag_12,twiddle_data_imag_11,twiddle_data_imag_10,twiddle_data_imag_9,twiddle_data_imag_8,twiddle_data_imag_7,twiddle_data_imag_6,twiddle_data_imag_5,twiddle_data_imag_4,twiddle_data_imag_3,
twiddle_data_imag_2,twiddle_data_imag_1,twiddle_data_imag_0}),
	.clken(global_clock_enable),
	.dffe3a_16(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[16]~q ),
	.dffe3a_15(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[15]~q ),
	.dffe3a_14(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[14]~q ),
	.dffe3a_13(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[13]~q ),
	.dffe3a_12(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[12]~q ),
	.dffe3a_11(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[11]~q ),
	.dffe3a_10(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[10]~q ),
	.dffe3a_9(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[9]~q ),
	.dffe3a_8(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[8]~q ),
	.dffe3a_7(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[7]~q ),
	.dffe3a_6(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[6]~q ),
	.dffe3a_5(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[5]~q ),
	.dffe3a_4(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[4]~q ),
	.dffe3a_3(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[3]~q ),
	.dffe3a_2(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[2]~q ),
	.dffe3a_1(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[1]~q ),
	.dffe3a_0(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[0]~q ),
	.dffe3a_31(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[31]~q ),
	.dffe3a_30(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[30]~q ),
	.dffe3a_29(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[29]~q ),
	.dffe3a_28(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[28]~q ),
	.dffe3a_27(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[27]~q ),
	.dffe3a_26(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[26]~q ),
	.dffe3a_25(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[25]~q ),
	.dffe3a_24(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[24]~q ),
	.dffe3a_23(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[23]~q ),
	.dffe3a_22(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[22]~q ),
	.dffe3a_21(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[21]~q ),
	.dffe3a_20(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[20]~q ),
	.dffe3a_19(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[19]~q ),
	.dffe3a_18(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[18]~q ),
	.dffe3a_17(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[17]~q ),
	.clock(clk));

fft256_LPM_MULT_2 \gen_ded_m1:gen_unext_m_ac:m_ac (
	.dataa({gnd,pipeline_dffe_171,pipeline_dffe_161,pipeline_dffe_15,pipeline_dffe_14,pipeline_dffe_13,pipeline_dffe_12,pipeline_dffe_11,pipeline_dffe_10,pipeline_dffe_9,pipeline_dffe_8,pipeline_dffe_7,pipeline_dffe_6,pipeline_dffe_5,pipeline_dffe_4,pipeline_dffe_3,pipeline_dffe_2}),
	.datab({gnd,twiddle_data_real_15,twiddle_data_real_14,twiddle_data_real_13,twiddle_data_real_12,twiddle_data_real_11,twiddle_data_real_10,twiddle_data_real_9,twiddle_data_real_8,twiddle_data_real_7,twiddle_data_real_6,twiddle_data_real_5,twiddle_data_real_4,twiddle_data_real_3,
twiddle_data_real_2,twiddle_data_real_1,twiddle_data_real_0}),
	.clken(global_clock_enable),
	.dffe3a_16(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[16]~q ),
	.dffe3a_15(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[15]~q ),
	.dffe3a_14(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[14]~q ),
	.dffe3a_13(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[13]~q ),
	.dffe3a_12(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[12]~q ),
	.dffe3a_11(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[11]~q ),
	.dffe3a_10(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[10]~q ),
	.dffe3a_9(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[9]~q ),
	.dffe3a_8(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[8]~q ),
	.dffe3a_7(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[7]~q ),
	.dffe3a_6(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[6]~q ),
	.dffe3a_5(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[5]~q ),
	.dffe3a_4(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[4]~q ),
	.dffe3a_3(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[3]~q ),
	.dffe3a_2(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[2]~q ),
	.dffe3a_1(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[1]~q ),
	.dffe3a_0(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[0]~q ),
	.dffe3a_31(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[31]~q ),
	.dffe3a_30(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[30]~q ),
	.dffe3a_29(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[29]~q ),
	.dffe3a_28(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[28]~q ),
	.dffe3a_27(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[27]~q ),
	.dffe3a_26(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[26]~q ),
	.dffe3a_25(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[25]~q ),
	.dffe3a_24(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[24]~q ),
	.dffe3a_23(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[23]~q ),
	.dffe3a_22(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[22]~q ),
	.dffe3a_21(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[21]~q ),
	.dffe3a_20(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[20]~q ),
	.dffe3a_19(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[19]~q ),
	.dffe3a_18(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[18]~q ),
	.dffe3a_17(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[17]~q ),
	.clock(clk));

dffeas \result_imag_1[16] (
	.clk(clk),
	.d(\result_imag_1[16]~64_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[16]~q ),
	.prn(vcc));
defparam \result_imag_1[16] .is_wysiwyg = "true";
defparam \result_imag_1[16] .power_up = "low";

dffeas \result_imag_1[15] (
	.clk(clk),
	.d(\result_imag_1[15]~62_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[15]~q ),
	.prn(vcc));
defparam \result_imag_1[15] .is_wysiwyg = "true";
defparam \result_imag_1[15] .power_up = "low";

dffeas \result_imag_1[14] (
	.clk(clk),
	.d(\result_imag_1[14]~60_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[14]~q ),
	.prn(vcc));
defparam \result_imag_1[14] .is_wysiwyg = "true";
defparam \result_imag_1[14] .power_up = "low";

dffeas \result_imag_1[13] (
	.clk(clk),
	.d(\result_imag_1[13]~58_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[13]~q ),
	.prn(vcc));
defparam \result_imag_1[13] .is_wysiwyg = "true";
defparam \result_imag_1[13] .power_up = "low";

dffeas \result_imag_1[12] (
	.clk(clk),
	.d(\result_imag_1[12]~56_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[12]~q ),
	.prn(vcc));
defparam \result_imag_1[12] .is_wysiwyg = "true";
defparam \result_imag_1[12] .power_up = "low";

dffeas \result_imag_1[11] (
	.clk(clk),
	.d(\result_imag_1[11]~54_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[11]~q ),
	.prn(vcc));
defparam \result_imag_1[11] .is_wysiwyg = "true";
defparam \result_imag_1[11] .power_up = "low";

dffeas \result_imag_1[10] (
	.clk(clk),
	.d(\result_imag_1[10]~52_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[10]~q ),
	.prn(vcc));
defparam \result_imag_1[10] .is_wysiwyg = "true";
defparam \result_imag_1[10] .power_up = "low";

dffeas \result_imag_1[9] (
	.clk(clk),
	.d(\result_imag_1[9]~50_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[9]~q ),
	.prn(vcc));
defparam \result_imag_1[9] .is_wysiwyg = "true";
defparam \result_imag_1[9] .power_up = "low";

dffeas \result_imag_1[8] (
	.clk(clk),
	.d(\result_imag_1[8]~48_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[8]~q ),
	.prn(vcc));
defparam \result_imag_1[8] .is_wysiwyg = "true";
defparam \result_imag_1[8] .power_up = "low";

dffeas \result_imag_1[7] (
	.clk(clk),
	.d(\result_imag_1[7]~46_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[7]~q ),
	.prn(vcc));
defparam \result_imag_1[7] .is_wysiwyg = "true";
defparam \result_imag_1[7] .power_up = "low";

dffeas \result_imag_1[6] (
	.clk(clk),
	.d(\result_imag_1[6]~44_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[6]~q ),
	.prn(vcc));
defparam \result_imag_1[6] .is_wysiwyg = "true";
defparam \result_imag_1[6] .power_up = "low";

dffeas \result_imag_1[5] (
	.clk(clk),
	.d(\result_imag_1[5]~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[5]~q ),
	.prn(vcc));
defparam \result_imag_1[5] .is_wysiwyg = "true";
defparam \result_imag_1[5] .power_up = "low";

dffeas \result_imag_1[4] (
	.clk(clk),
	.d(\result_imag_1[4]~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[4]~q ),
	.prn(vcc));
defparam \result_imag_1[4] .is_wysiwyg = "true";
defparam \result_imag_1[4] .power_up = "low";

dffeas \result_imag_1[3] (
	.clk(clk),
	.d(\result_imag_1[3]~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[3]~q ),
	.prn(vcc));
defparam \result_imag_1[3] .is_wysiwyg = "true";
defparam \result_imag_1[3] .power_up = "low";

dffeas \result_imag_1[2] (
	.clk(clk),
	.d(\result_imag_1[2]~36_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[2]~q ),
	.prn(vcc));
defparam \result_imag_1[2] .is_wysiwyg = "true";
defparam \result_imag_1[2] .power_up = "low";

dffeas \result_imag_1[1] (
	.clk(clk),
	.d(\result_imag_1[1]~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[1]~q ),
	.prn(vcc));
defparam \result_imag_1[1] .is_wysiwyg = "true";
defparam \result_imag_1[1] .power_up = "low";

dffeas \result_imag_1[0] (
	.clk(clk),
	.d(\result_imag_1[0]~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[0]~q ),
	.prn(vcc));
defparam \result_imag_1[0] .is_wysiwyg = "true";
defparam \result_imag_1[0] .power_up = "low";

dffeas \result_imag_1[31] (
	.clk(clk),
	.d(\result_imag_1[31]~94_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[31]~q ),
	.prn(vcc));
defparam \result_imag_1[31] .is_wysiwyg = "true";
defparam \result_imag_1[31] .power_up = "low";

dffeas \result_imag_1[17] (
	.clk(clk),
	.d(\result_imag_1[17]~66_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[17]~q ),
	.prn(vcc));
defparam \result_imag_1[17] .is_wysiwyg = "true";
defparam \result_imag_1[17] .power_up = "low";

dffeas \result_imag_1[18] (
	.clk(clk),
	.d(\result_imag_1[18]~68_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[18]~q ),
	.prn(vcc));
defparam \result_imag_1[18] .is_wysiwyg = "true";
defparam \result_imag_1[18] .power_up = "low";

dffeas \result_imag_1[19] (
	.clk(clk),
	.d(\result_imag_1[19]~70_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[19]~q ),
	.prn(vcc));
defparam \result_imag_1[19] .is_wysiwyg = "true";
defparam \result_imag_1[19] .power_up = "low";

dffeas \result_imag_1[20] (
	.clk(clk),
	.d(\result_imag_1[20]~72_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[20]~q ),
	.prn(vcc));
defparam \result_imag_1[20] .is_wysiwyg = "true";
defparam \result_imag_1[20] .power_up = "low";

dffeas \result_imag_1[21] (
	.clk(clk),
	.d(\result_imag_1[21]~74_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[21]~q ),
	.prn(vcc));
defparam \result_imag_1[21] .is_wysiwyg = "true";
defparam \result_imag_1[21] .power_up = "low";

dffeas \result_imag_1[22] (
	.clk(clk),
	.d(\result_imag_1[22]~76_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[22]~q ),
	.prn(vcc));
defparam \result_imag_1[22] .is_wysiwyg = "true";
defparam \result_imag_1[22] .power_up = "low";

dffeas \result_imag_1[23] (
	.clk(clk),
	.d(\result_imag_1[23]~78_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[23]~q ),
	.prn(vcc));
defparam \result_imag_1[23] .is_wysiwyg = "true";
defparam \result_imag_1[23] .power_up = "low";

dffeas \result_imag_1[24] (
	.clk(clk),
	.d(\result_imag_1[24]~80_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[24]~q ),
	.prn(vcc));
defparam \result_imag_1[24] .is_wysiwyg = "true";
defparam \result_imag_1[24] .power_up = "low";

dffeas \result_imag_1[25] (
	.clk(clk),
	.d(\result_imag_1[25]~82_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[25]~q ),
	.prn(vcc));
defparam \result_imag_1[25] .is_wysiwyg = "true";
defparam \result_imag_1[25] .power_up = "low";

dffeas \result_imag_1[26] (
	.clk(clk),
	.d(\result_imag_1[26]~84_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[26]~q ),
	.prn(vcc));
defparam \result_imag_1[26] .is_wysiwyg = "true";
defparam \result_imag_1[26] .power_up = "low";

dffeas \result_imag_1[27] (
	.clk(clk),
	.d(\result_imag_1[27]~86_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[27]~q ),
	.prn(vcc));
defparam \result_imag_1[27] .is_wysiwyg = "true";
defparam \result_imag_1[27] .power_up = "low";

dffeas \result_imag_1[28] (
	.clk(clk),
	.d(\result_imag_1[28]~88_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[28]~q ),
	.prn(vcc));
defparam \result_imag_1[28] .is_wysiwyg = "true";
defparam \result_imag_1[28] .power_up = "low";

dffeas \result_imag_1[29] (
	.clk(clk),
	.d(\result_imag_1[29]~90_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[29]~q ),
	.prn(vcc));
defparam \result_imag_1[29] .is_wysiwyg = "true";
defparam \result_imag_1[29] .power_up = "low";

dffeas \result_imag_1[30] (
	.clk(clk),
	.d(\result_imag_1[30]~92_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_imag_1[30]~q ),
	.prn(vcc));
defparam \result_imag_1[30] .is_wysiwyg = "true";
defparam \result_imag_1[30] .power_up = "low";

dffeas \result_real_1_tmp[16] (
	.clk(clk),
	.d(\result_real_1_tmp[16]~64_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[16]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[16] .is_wysiwyg = "true";
defparam \result_real_1_tmp[16] .power_up = "low";

dffeas \result_real_1_tmp[15] (
	.clk(clk),
	.d(\result_real_1_tmp[15]~62_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[15]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[15] .is_wysiwyg = "true";
defparam \result_real_1_tmp[15] .power_up = "low";

dffeas \result_real_1_tmp[14] (
	.clk(clk),
	.d(\result_real_1_tmp[14]~60_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[14]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[14] .is_wysiwyg = "true";
defparam \result_real_1_tmp[14] .power_up = "low";

dffeas \result_real_1_tmp[13] (
	.clk(clk),
	.d(\result_real_1_tmp[13]~58_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[13]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[13] .is_wysiwyg = "true";
defparam \result_real_1_tmp[13] .power_up = "low";

dffeas \result_real_1_tmp[12] (
	.clk(clk),
	.d(\result_real_1_tmp[12]~56_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[12]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[12] .is_wysiwyg = "true";
defparam \result_real_1_tmp[12] .power_up = "low";

dffeas \result_real_1_tmp[11] (
	.clk(clk),
	.d(\result_real_1_tmp[11]~54_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[11]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[11] .is_wysiwyg = "true";
defparam \result_real_1_tmp[11] .power_up = "low";

dffeas \result_real_1_tmp[10] (
	.clk(clk),
	.d(\result_real_1_tmp[10]~52_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[10]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[10] .is_wysiwyg = "true";
defparam \result_real_1_tmp[10] .power_up = "low";

dffeas \result_real_1_tmp[9] (
	.clk(clk),
	.d(\result_real_1_tmp[9]~50_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[9]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[9] .is_wysiwyg = "true";
defparam \result_real_1_tmp[9] .power_up = "low";

dffeas \result_real_1_tmp[8] (
	.clk(clk),
	.d(\result_real_1_tmp[8]~48_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[8]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[8] .is_wysiwyg = "true";
defparam \result_real_1_tmp[8] .power_up = "low";

dffeas \result_real_1_tmp[7] (
	.clk(clk),
	.d(\result_real_1_tmp[7]~46_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[7]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[7] .is_wysiwyg = "true";
defparam \result_real_1_tmp[7] .power_up = "low";

dffeas \result_real_1_tmp[6] (
	.clk(clk),
	.d(\result_real_1_tmp[6]~44_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[6]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[6] .is_wysiwyg = "true";
defparam \result_real_1_tmp[6] .power_up = "low";

dffeas \result_real_1_tmp[5] (
	.clk(clk),
	.d(\result_real_1_tmp[5]~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[5]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[5] .is_wysiwyg = "true";
defparam \result_real_1_tmp[5] .power_up = "low";

dffeas \result_real_1_tmp[4] (
	.clk(clk),
	.d(\result_real_1_tmp[4]~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[4]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[4] .is_wysiwyg = "true";
defparam \result_real_1_tmp[4] .power_up = "low";

dffeas \result_real_1_tmp[3] (
	.clk(clk),
	.d(\result_real_1_tmp[3]~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[3]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[3] .is_wysiwyg = "true";
defparam \result_real_1_tmp[3] .power_up = "low";

dffeas \result_real_1_tmp[2] (
	.clk(clk),
	.d(\result_real_1_tmp[2]~36_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[2]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[2] .is_wysiwyg = "true";
defparam \result_real_1_tmp[2] .power_up = "low";

dffeas \result_real_1_tmp[1] (
	.clk(clk),
	.d(\result_real_1_tmp[1]~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[1]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[1] .is_wysiwyg = "true";
defparam \result_real_1_tmp[1] .power_up = "low";

dffeas \result_real_1_tmp[0] (
	.clk(clk),
	.d(\result_real_1_tmp[0]~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[0]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[0] .is_wysiwyg = "true";
defparam \result_real_1_tmp[0] .power_up = "low";

dffeas \result_real_1_tmp[31] (
	.clk(clk),
	.d(\result_real_1_tmp[31]~94_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[31]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[31] .is_wysiwyg = "true";
defparam \result_real_1_tmp[31] .power_up = "low";

dffeas \addresult_ac_bd[16] (
	.clk(clk),
	.d(\addresult_ac_bd[16]~64_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[16]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[16] .is_wysiwyg = "true";
defparam \addresult_ac_bd[16] .power_up = "low";

dffeas \addresult_ac_bd[15] (
	.clk(clk),
	.d(\addresult_ac_bd[15]~62_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[15]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[15] .is_wysiwyg = "true";
defparam \addresult_ac_bd[15] .power_up = "low";

dffeas \addresult_ac_bd[14] (
	.clk(clk),
	.d(\addresult_ac_bd[14]~60_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[14]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[14] .is_wysiwyg = "true";
defparam \addresult_ac_bd[14] .power_up = "low";

dffeas \addresult_ac_bd[13] (
	.clk(clk),
	.d(\addresult_ac_bd[13]~58_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[13]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[13] .is_wysiwyg = "true";
defparam \addresult_ac_bd[13] .power_up = "low";

dffeas \addresult_ac_bd[12] (
	.clk(clk),
	.d(\addresult_ac_bd[12]~56_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[12]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[12] .is_wysiwyg = "true";
defparam \addresult_ac_bd[12] .power_up = "low";

dffeas \addresult_ac_bd[11] (
	.clk(clk),
	.d(\addresult_ac_bd[11]~54_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[11]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[11] .is_wysiwyg = "true";
defparam \addresult_ac_bd[11] .power_up = "low";

dffeas \addresult_ac_bd[10] (
	.clk(clk),
	.d(\addresult_ac_bd[10]~52_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[10]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[10] .is_wysiwyg = "true";
defparam \addresult_ac_bd[10] .power_up = "low";

dffeas \addresult_ac_bd[9] (
	.clk(clk),
	.d(\addresult_ac_bd[9]~50_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[9]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[9] .is_wysiwyg = "true";
defparam \addresult_ac_bd[9] .power_up = "low";

dffeas \addresult_ac_bd[8] (
	.clk(clk),
	.d(\addresult_ac_bd[8]~48_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[8]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[8] .is_wysiwyg = "true";
defparam \addresult_ac_bd[8] .power_up = "low";

dffeas \addresult_ac_bd[7] (
	.clk(clk),
	.d(\addresult_ac_bd[7]~46_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[7]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[7] .is_wysiwyg = "true";
defparam \addresult_ac_bd[7] .power_up = "low";

dffeas \addresult_ac_bd[6] (
	.clk(clk),
	.d(\addresult_ac_bd[6]~44_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[6]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[6] .is_wysiwyg = "true";
defparam \addresult_ac_bd[6] .power_up = "low";

dffeas \addresult_ac_bd[5] (
	.clk(clk),
	.d(\addresult_ac_bd[5]~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[5]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[5] .is_wysiwyg = "true";
defparam \addresult_ac_bd[5] .power_up = "low";

dffeas \addresult_ac_bd[4] (
	.clk(clk),
	.d(\addresult_ac_bd[4]~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[4]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[4] .is_wysiwyg = "true";
defparam \addresult_ac_bd[4] .power_up = "low";

dffeas \addresult_ac_bd[3] (
	.clk(clk),
	.d(\addresult_ac_bd[3]~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[3]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[3] .is_wysiwyg = "true";
defparam \addresult_ac_bd[3] .power_up = "low";

dffeas \addresult_ac_bd[2] (
	.clk(clk),
	.d(\addresult_ac_bd[2]~36_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[2]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[2] .is_wysiwyg = "true";
defparam \addresult_ac_bd[2] .power_up = "low";

dffeas \addresult_ac_bd[1] (
	.clk(clk),
	.d(\addresult_ac_bd[1]~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[1]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[1] .is_wysiwyg = "true";
defparam \addresult_ac_bd[1] .power_up = "low";

dffeas \addresult_ac_bd[0] (
	.clk(clk),
	.d(\addresult_ac_bd[0]~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[0]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[0] .is_wysiwyg = "true";
defparam \addresult_ac_bd[0] .power_up = "low";

cycloneive_lcell_comb \result_imag_1[0]~32 (
	.dataa(\addresult_ac_bd[0]~q ),
	.datab(\result_a_b_c_d_se[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\result_imag_1[0]~32_combout ),
	.cout(\result_imag_1[0]~33 ));
defparam \result_imag_1[0]~32 .lut_mask = 16'h66DD;
defparam \result_imag_1[0]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \result_imag_1[1]~34 (
	.dataa(\addresult_ac_bd[1]~q ),
	.datab(\result_a_b_c_d_se[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[0]~33 ),
	.combout(\result_imag_1[1]~34_combout ),
	.cout(\result_imag_1[1]~35 ));
defparam \result_imag_1[1]~34 .lut_mask = 16'h96BF;
defparam \result_imag_1[1]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[2]~36 (
	.dataa(\addresult_ac_bd[2]~q ),
	.datab(\result_a_b_c_d_se[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[1]~35 ),
	.combout(\result_imag_1[2]~36_combout ),
	.cout(\result_imag_1[2]~37 ));
defparam \result_imag_1[2]~36 .lut_mask = 16'h96DF;
defparam \result_imag_1[2]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[3]~38 (
	.dataa(\addresult_ac_bd[3]~q ),
	.datab(\result_a_b_c_d_se[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[2]~37 ),
	.combout(\result_imag_1[3]~38_combout ),
	.cout(\result_imag_1[3]~39 ));
defparam \result_imag_1[3]~38 .lut_mask = 16'h96BF;
defparam \result_imag_1[3]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[4]~40 (
	.dataa(\addresult_ac_bd[4]~q ),
	.datab(\result_a_b_c_d_se[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[3]~39 ),
	.combout(\result_imag_1[4]~40_combout ),
	.cout(\result_imag_1[4]~41 ));
defparam \result_imag_1[4]~40 .lut_mask = 16'h96DF;
defparam \result_imag_1[4]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[5]~42 (
	.dataa(\addresult_ac_bd[5]~q ),
	.datab(\result_a_b_c_d_se[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[4]~41 ),
	.combout(\result_imag_1[5]~42_combout ),
	.cout(\result_imag_1[5]~43 ));
defparam \result_imag_1[5]~42 .lut_mask = 16'h96BF;
defparam \result_imag_1[5]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[6]~44 (
	.dataa(\addresult_ac_bd[6]~q ),
	.datab(\result_a_b_c_d_se[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[5]~43 ),
	.combout(\result_imag_1[6]~44_combout ),
	.cout(\result_imag_1[6]~45 ));
defparam \result_imag_1[6]~44 .lut_mask = 16'h96DF;
defparam \result_imag_1[6]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[7]~46 (
	.dataa(\addresult_ac_bd[7]~q ),
	.datab(\result_a_b_c_d_se[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[6]~45 ),
	.combout(\result_imag_1[7]~46_combout ),
	.cout(\result_imag_1[7]~47 ));
defparam \result_imag_1[7]~46 .lut_mask = 16'h96BF;
defparam \result_imag_1[7]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[8]~48 (
	.dataa(\addresult_ac_bd[8]~q ),
	.datab(\result_a_b_c_d_se[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[7]~47 ),
	.combout(\result_imag_1[8]~48_combout ),
	.cout(\result_imag_1[8]~49 ));
defparam \result_imag_1[8]~48 .lut_mask = 16'h96DF;
defparam \result_imag_1[8]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[9]~50 (
	.dataa(\addresult_ac_bd[9]~q ),
	.datab(\result_a_b_c_d_se[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[8]~49 ),
	.combout(\result_imag_1[9]~50_combout ),
	.cout(\result_imag_1[9]~51 ));
defparam \result_imag_1[9]~50 .lut_mask = 16'h96BF;
defparam \result_imag_1[9]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[10]~52 (
	.dataa(\addresult_ac_bd[10]~q ),
	.datab(\result_a_b_c_d_se[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[9]~51 ),
	.combout(\result_imag_1[10]~52_combout ),
	.cout(\result_imag_1[10]~53 ));
defparam \result_imag_1[10]~52 .lut_mask = 16'h96DF;
defparam \result_imag_1[10]~52 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[11]~54 (
	.dataa(\addresult_ac_bd[11]~q ),
	.datab(\result_a_b_c_d_se[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[10]~53 ),
	.combout(\result_imag_1[11]~54_combout ),
	.cout(\result_imag_1[11]~55 ));
defparam \result_imag_1[11]~54 .lut_mask = 16'h96BF;
defparam \result_imag_1[11]~54 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[12]~56 (
	.dataa(\addresult_ac_bd[12]~q ),
	.datab(\result_a_b_c_d_se[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[11]~55 ),
	.combout(\result_imag_1[12]~56_combout ),
	.cout(\result_imag_1[12]~57 ));
defparam \result_imag_1[12]~56 .lut_mask = 16'h96DF;
defparam \result_imag_1[12]~56 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[13]~58 (
	.dataa(\addresult_ac_bd[13]~q ),
	.datab(\result_a_b_c_d_se[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[12]~57 ),
	.combout(\result_imag_1[13]~58_combout ),
	.cout(\result_imag_1[13]~59 ));
defparam \result_imag_1[13]~58 .lut_mask = 16'h96BF;
defparam \result_imag_1[13]~58 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[14]~60 (
	.dataa(\addresult_ac_bd[14]~q ),
	.datab(\result_a_b_c_d_se[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[13]~59 ),
	.combout(\result_imag_1[14]~60_combout ),
	.cout(\result_imag_1[14]~61 ));
defparam \result_imag_1[14]~60 .lut_mask = 16'h96DF;
defparam \result_imag_1[14]~60 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[15]~62 (
	.dataa(\addresult_ac_bd[15]~q ),
	.datab(\result_a_b_c_d_se[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[14]~61 ),
	.combout(\result_imag_1[15]~62_combout ),
	.cout(\result_imag_1[15]~63 ));
defparam \result_imag_1[15]~62 .lut_mask = 16'h96BF;
defparam \result_imag_1[15]~62 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[16]~64 (
	.dataa(\addresult_ac_bd[16]~q ),
	.datab(\result_a_b_c_d_se[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[15]~63 ),
	.combout(\result_imag_1[16]~64_combout ),
	.cout(\result_imag_1[16]~65 ));
defparam \result_imag_1[16]~64 .lut_mask = 16'h96DF;
defparam \result_imag_1[16]~64 .sum_lutc_input = "cin";

dffeas \addresult_ac_bd[31] (
	.clk(clk),
	.d(\addresult_ac_bd[31]~94_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[31]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[31] .is_wysiwyg = "true";
defparam \addresult_ac_bd[31] .power_up = "low";

dffeas \addresult_ac_bd[30] (
	.clk(clk),
	.d(\addresult_ac_bd[30]~92_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[30]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[30] .is_wysiwyg = "true";
defparam \addresult_ac_bd[30] .power_up = "low";

dffeas \addresult_ac_bd[29] (
	.clk(clk),
	.d(\addresult_ac_bd[29]~90_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[29]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[29] .is_wysiwyg = "true";
defparam \addresult_ac_bd[29] .power_up = "low";

dffeas \addresult_ac_bd[28] (
	.clk(clk),
	.d(\addresult_ac_bd[28]~88_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[28]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[28] .is_wysiwyg = "true";
defparam \addresult_ac_bd[28] .power_up = "low";

dffeas \addresult_ac_bd[27] (
	.clk(clk),
	.d(\addresult_ac_bd[27]~86_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[27]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[27] .is_wysiwyg = "true";
defparam \addresult_ac_bd[27] .power_up = "low";

dffeas \addresult_ac_bd[26] (
	.clk(clk),
	.d(\addresult_ac_bd[26]~84_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[26]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[26] .is_wysiwyg = "true";
defparam \addresult_ac_bd[26] .power_up = "low";

dffeas \addresult_ac_bd[25] (
	.clk(clk),
	.d(\addresult_ac_bd[25]~82_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[25]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[25] .is_wysiwyg = "true";
defparam \addresult_ac_bd[25] .power_up = "low";

dffeas \addresult_ac_bd[24] (
	.clk(clk),
	.d(\addresult_ac_bd[24]~80_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[24]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[24] .is_wysiwyg = "true";
defparam \addresult_ac_bd[24] .power_up = "low";

dffeas \addresult_ac_bd[23] (
	.clk(clk),
	.d(\addresult_ac_bd[23]~78_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[23]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[23] .is_wysiwyg = "true";
defparam \addresult_ac_bd[23] .power_up = "low";

dffeas \addresult_ac_bd[22] (
	.clk(clk),
	.d(\addresult_ac_bd[22]~76_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[22]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[22] .is_wysiwyg = "true";
defparam \addresult_ac_bd[22] .power_up = "low";

dffeas \addresult_ac_bd[21] (
	.clk(clk),
	.d(\addresult_ac_bd[21]~74_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[21]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[21] .is_wysiwyg = "true";
defparam \addresult_ac_bd[21] .power_up = "low";

dffeas \addresult_ac_bd[20] (
	.clk(clk),
	.d(\addresult_ac_bd[20]~72_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[20]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[20] .is_wysiwyg = "true";
defparam \addresult_ac_bd[20] .power_up = "low";

dffeas \addresult_ac_bd[19] (
	.clk(clk),
	.d(\addresult_ac_bd[19]~70_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[19]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[19] .is_wysiwyg = "true";
defparam \addresult_ac_bd[19] .power_up = "low";

dffeas \addresult_ac_bd[18] (
	.clk(clk),
	.d(\addresult_ac_bd[18]~68_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[18]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[18] .is_wysiwyg = "true";
defparam \addresult_ac_bd[18] .power_up = "low";

dffeas \addresult_ac_bd[17] (
	.clk(clk),
	.d(\addresult_ac_bd[17]~66_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_ac_bd[17]~q ),
	.prn(vcc));
defparam \addresult_ac_bd[17] .is_wysiwyg = "true";
defparam \addresult_ac_bd[17] .power_up = "low";

cycloneive_lcell_comb \result_imag_1[17]~66 (
	.dataa(\addresult_ac_bd[17]~q ),
	.datab(\result_a_b_c_d_se[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[16]~65 ),
	.combout(\result_imag_1[17]~66_combout ),
	.cout(\result_imag_1[17]~67 ));
defparam \result_imag_1[17]~66 .lut_mask = 16'h96BF;
defparam \result_imag_1[17]~66 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[18]~68 (
	.dataa(\addresult_ac_bd[18]~q ),
	.datab(\result_a_b_c_d_se[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[17]~67 ),
	.combout(\result_imag_1[18]~68_combout ),
	.cout(\result_imag_1[18]~69 ));
defparam \result_imag_1[18]~68 .lut_mask = 16'h96DF;
defparam \result_imag_1[18]~68 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[19]~70 (
	.dataa(\addresult_ac_bd[19]~q ),
	.datab(\result_a_b_c_d_se[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[18]~69 ),
	.combout(\result_imag_1[19]~70_combout ),
	.cout(\result_imag_1[19]~71 ));
defparam \result_imag_1[19]~70 .lut_mask = 16'h96BF;
defparam \result_imag_1[19]~70 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[20]~72 (
	.dataa(\addresult_ac_bd[20]~q ),
	.datab(\result_a_b_c_d_se[20]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[19]~71 ),
	.combout(\result_imag_1[20]~72_combout ),
	.cout(\result_imag_1[20]~73 ));
defparam \result_imag_1[20]~72 .lut_mask = 16'h96DF;
defparam \result_imag_1[20]~72 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[21]~74 (
	.dataa(\addresult_ac_bd[21]~q ),
	.datab(\result_a_b_c_d_se[21]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[20]~73 ),
	.combout(\result_imag_1[21]~74_combout ),
	.cout(\result_imag_1[21]~75 ));
defparam \result_imag_1[21]~74 .lut_mask = 16'h96BF;
defparam \result_imag_1[21]~74 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[22]~76 (
	.dataa(\addresult_ac_bd[22]~q ),
	.datab(\result_a_b_c_d_se[22]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[21]~75 ),
	.combout(\result_imag_1[22]~76_combout ),
	.cout(\result_imag_1[22]~77 ));
defparam \result_imag_1[22]~76 .lut_mask = 16'h96DF;
defparam \result_imag_1[22]~76 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[23]~78 (
	.dataa(\addresult_ac_bd[23]~q ),
	.datab(\result_a_b_c_d_se[23]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[22]~77 ),
	.combout(\result_imag_1[23]~78_combout ),
	.cout(\result_imag_1[23]~79 ));
defparam \result_imag_1[23]~78 .lut_mask = 16'h96BF;
defparam \result_imag_1[23]~78 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[24]~80 (
	.dataa(\addresult_ac_bd[24]~q ),
	.datab(\result_a_b_c_d_se[24]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[23]~79 ),
	.combout(\result_imag_1[24]~80_combout ),
	.cout(\result_imag_1[24]~81 ));
defparam \result_imag_1[24]~80 .lut_mask = 16'h96DF;
defparam \result_imag_1[24]~80 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[25]~82 (
	.dataa(\addresult_ac_bd[25]~q ),
	.datab(\result_a_b_c_d_se[25]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[24]~81 ),
	.combout(\result_imag_1[25]~82_combout ),
	.cout(\result_imag_1[25]~83 ));
defparam \result_imag_1[25]~82 .lut_mask = 16'h96BF;
defparam \result_imag_1[25]~82 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[26]~84 (
	.dataa(\addresult_ac_bd[26]~q ),
	.datab(\result_a_b_c_d_se[26]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[25]~83 ),
	.combout(\result_imag_1[26]~84_combout ),
	.cout(\result_imag_1[26]~85 ));
defparam \result_imag_1[26]~84 .lut_mask = 16'h96DF;
defparam \result_imag_1[26]~84 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[27]~86 (
	.dataa(\addresult_ac_bd[27]~q ),
	.datab(\result_a_b_c_d_se[27]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[26]~85 ),
	.combout(\result_imag_1[27]~86_combout ),
	.cout(\result_imag_1[27]~87 ));
defparam \result_imag_1[27]~86 .lut_mask = 16'h96BF;
defparam \result_imag_1[27]~86 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[28]~88 (
	.dataa(\addresult_ac_bd[28]~q ),
	.datab(\result_a_b_c_d_se[28]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[27]~87 ),
	.combout(\result_imag_1[28]~88_combout ),
	.cout(\result_imag_1[28]~89 ));
defparam \result_imag_1[28]~88 .lut_mask = 16'h96DF;
defparam \result_imag_1[28]~88 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[29]~90 (
	.dataa(\addresult_ac_bd[29]~q ),
	.datab(\result_a_b_c_d_se[29]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[28]~89 ),
	.combout(\result_imag_1[29]~90_combout ),
	.cout(\result_imag_1[29]~91 ));
defparam \result_imag_1[29]~90 .lut_mask = 16'h96BF;
defparam \result_imag_1[29]~90 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[30]~92 (
	.dataa(\addresult_ac_bd[30]~q ),
	.datab(\result_a_b_c_d_se[30]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_imag_1[29]~91 ),
	.combout(\result_imag_1[30]~92_combout ),
	.cout(\result_imag_1[30]~93 ));
defparam \result_imag_1[30]~92 .lut_mask = 16'h96DF;
defparam \result_imag_1[30]~92 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_imag_1[31]~94 (
	.dataa(\addresult_ac_bd[31]~q ),
	.datab(\result_a_b_c_d_se[31]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\result_imag_1[30]~93 ),
	.combout(\result_imag_1[31]~94_combout ),
	.cout());
defparam \result_imag_1[31]~94 .lut_mask = 16'h9696;
defparam \result_imag_1[31]~94 .sum_lutc_input = "cin";

dffeas \result_real_1_tmp[17] (
	.clk(clk),
	.d(\result_real_1_tmp[17]~66_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[17]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[17] .is_wysiwyg = "true";
defparam \result_real_1_tmp[17] .power_up = "low";

dffeas \result_real_1_tmp[18] (
	.clk(clk),
	.d(\result_real_1_tmp[18]~68_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[18]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[18] .is_wysiwyg = "true";
defparam \result_real_1_tmp[18] .power_up = "low";

dffeas \result_real_1_tmp[19] (
	.clk(clk),
	.d(\result_real_1_tmp[19]~70_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[19]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[19] .is_wysiwyg = "true";
defparam \result_real_1_tmp[19] .power_up = "low";

dffeas \result_real_1_tmp[20] (
	.clk(clk),
	.d(\result_real_1_tmp[20]~72_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[20]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[20] .is_wysiwyg = "true";
defparam \result_real_1_tmp[20] .power_up = "low";

dffeas \result_real_1_tmp[21] (
	.clk(clk),
	.d(\result_real_1_tmp[21]~74_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[21]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[21] .is_wysiwyg = "true";
defparam \result_real_1_tmp[21] .power_up = "low";

dffeas \result_real_1_tmp[22] (
	.clk(clk),
	.d(\result_real_1_tmp[22]~76_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[22]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[22] .is_wysiwyg = "true";
defparam \result_real_1_tmp[22] .power_up = "low";

dffeas \result_real_1_tmp[23] (
	.clk(clk),
	.d(\result_real_1_tmp[23]~78_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[23]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[23] .is_wysiwyg = "true";
defparam \result_real_1_tmp[23] .power_up = "low";

dffeas \result_real_1_tmp[24] (
	.clk(clk),
	.d(\result_real_1_tmp[24]~80_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[24]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[24] .is_wysiwyg = "true";
defparam \result_real_1_tmp[24] .power_up = "low";

dffeas \result_real_1_tmp[25] (
	.clk(clk),
	.d(\result_real_1_tmp[25]~82_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[25]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[25] .is_wysiwyg = "true";
defparam \result_real_1_tmp[25] .power_up = "low";

dffeas \result_real_1_tmp[26] (
	.clk(clk),
	.d(\result_real_1_tmp[26]~84_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[26]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[26] .is_wysiwyg = "true";
defparam \result_real_1_tmp[26] .power_up = "low";

dffeas \result_real_1_tmp[27] (
	.clk(clk),
	.d(\result_real_1_tmp[27]~86_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[27]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[27] .is_wysiwyg = "true";
defparam \result_real_1_tmp[27] .power_up = "low";

dffeas \result_real_1_tmp[28] (
	.clk(clk),
	.d(\result_real_1_tmp[28]~88_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[28]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[28] .is_wysiwyg = "true";
defparam \result_real_1_tmp[28] .power_up = "low";

dffeas \result_real_1_tmp[29] (
	.clk(clk),
	.d(\result_real_1_tmp[29]~90_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[29]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[29] .is_wysiwyg = "true";
defparam \result_real_1_tmp[29] .power_up = "low";

dffeas \result_real_1_tmp[30] (
	.clk(clk),
	.d(\result_real_1_tmp[30]~92_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_real_1_tmp[30]~q ),
	.prn(vcc));
defparam \result_real_1_tmp[30] .is_wysiwyg = "true";
defparam \result_real_1_tmp[30] .power_up = "low";

cycloneive_lcell_comb \result_real_1_tmp[0]~32 (
	.dataa(\result_a_c_se[0]~q ),
	.datab(\result_b_d_se[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\result_real_1_tmp[0]~32_combout ),
	.cout(\result_real_1_tmp[0]~33 ));
defparam \result_real_1_tmp[0]~32 .lut_mask = 16'h66BB;
defparam \result_real_1_tmp[0]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \result_real_1_tmp[1]~34 (
	.dataa(\result_a_c_se[1]~q ),
	.datab(\result_b_d_se[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[0]~33 ),
	.combout(\result_real_1_tmp[1]~34_combout ),
	.cout(\result_real_1_tmp[1]~35 ));
defparam \result_real_1_tmp[1]~34 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[1]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[2]~36 (
	.dataa(\result_a_c_se[2]~q ),
	.datab(\result_b_d_se[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[1]~35 ),
	.combout(\result_real_1_tmp[2]~36_combout ),
	.cout(\result_real_1_tmp[2]~37 ));
defparam \result_real_1_tmp[2]~36 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[2]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[3]~38 (
	.dataa(\result_a_c_se[3]~q ),
	.datab(\result_b_d_se[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[2]~37 ),
	.combout(\result_real_1_tmp[3]~38_combout ),
	.cout(\result_real_1_tmp[3]~39 ));
defparam \result_real_1_tmp[3]~38 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[3]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[4]~40 (
	.dataa(\result_a_c_se[4]~q ),
	.datab(\result_b_d_se[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[3]~39 ),
	.combout(\result_real_1_tmp[4]~40_combout ),
	.cout(\result_real_1_tmp[4]~41 ));
defparam \result_real_1_tmp[4]~40 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[4]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[5]~42 (
	.dataa(\result_a_c_se[5]~q ),
	.datab(\result_b_d_se[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[4]~41 ),
	.combout(\result_real_1_tmp[5]~42_combout ),
	.cout(\result_real_1_tmp[5]~43 ));
defparam \result_real_1_tmp[5]~42 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[5]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[6]~44 (
	.dataa(\result_a_c_se[6]~q ),
	.datab(\result_b_d_se[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[5]~43 ),
	.combout(\result_real_1_tmp[6]~44_combout ),
	.cout(\result_real_1_tmp[6]~45 ));
defparam \result_real_1_tmp[6]~44 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[6]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[7]~46 (
	.dataa(\result_a_c_se[7]~q ),
	.datab(\result_b_d_se[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[6]~45 ),
	.combout(\result_real_1_tmp[7]~46_combout ),
	.cout(\result_real_1_tmp[7]~47 ));
defparam \result_real_1_tmp[7]~46 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[7]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[8]~48 (
	.dataa(\result_a_c_se[8]~q ),
	.datab(\result_b_d_se[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[7]~47 ),
	.combout(\result_real_1_tmp[8]~48_combout ),
	.cout(\result_real_1_tmp[8]~49 ));
defparam \result_real_1_tmp[8]~48 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[8]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[9]~50 (
	.dataa(\result_a_c_se[9]~q ),
	.datab(\result_b_d_se[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[8]~49 ),
	.combout(\result_real_1_tmp[9]~50_combout ),
	.cout(\result_real_1_tmp[9]~51 ));
defparam \result_real_1_tmp[9]~50 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[9]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[10]~52 (
	.dataa(\result_a_c_se[10]~q ),
	.datab(\result_b_d_se[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[9]~51 ),
	.combout(\result_real_1_tmp[10]~52_combout ),
	.cout(\result_real_1_tmp[10]~53 ));
defparam \result_real_1_tmp[10]~52 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[10]~52 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[11]~54 (
	.dataa(\result_a_c_se[11]~q ),
	.datab(\result_b_d_se[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[10]~53 ),
	.combout(\result_real_1_tmp[11]~54_combout ),
	.cout(\result_real_1_tmp[11]~55 ));
defparam \result_real_1_tmp[11]~54 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[11]~54 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[12]~56 (
	.dataa(\result_a_c_se[12]~q ),
	.datab(\result_b_d_se[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[11]~55 ),
	.combout(\result_real_1_tmp[12]~56_combout ),
	.cout(\result_real_1_tmp[12]~57 ));
defparam \result_real_1_tmp[12]~56 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[12]~56 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[13]~58 (
	.dataa(\result_a_c_se[13]~q ),
	.datab(\result_b_d_se[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[12]~57 ),
	.combout(\result_real_1_tmp[13]~58_combout ),
	.cout(\result_real_1_tmp[13]~59 ));
defparam \result_real_1_tmp[13]~58 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[13]~58 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[14]~60 (
	.dataa(\result_a_c_se[14]~q ),
	.datab(\result_b_d_se[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[13]~59 ),
	.combout(\result_real_1_tmp[14]~60_combout ),
	.cout(\result_real_1_tmp[14]~61 ));
defparam \result_real_1_tmp[14]~60 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[14]~60 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[15]~62 (
	.dataa(\result_a_c_se[15]~q ),
	.datab(\result_b_d_se[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[14]~61 ),
	.combout(\result_real_1_tmp[15]~62_combout ),
	.cout(\result_real_1_tmp[15]~63 ));
defparam \result_real_1_tmp[15]~62 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[15]~62 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[16]~64 (
	.dataa(\result_a_c_se[16]~q ),
	.datab(\result_b_d_se[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[15]~63 ),
	.combout(\result_real_1_tmp[16]~64_combout ),
	.cout(\result_real_1_tmp[16]~65 ));
defparam \result_real_1_tmp[16]~64 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[16]~64 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[17]~66 (
	.dataa(\result_a_c_se[17]~q ),
	.datab(\result_b_d_se[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[16]~65 ),
	.combout(\result_real_1_tmp[17]~66_combout ),
	.cout(\result_real_1_tmp[17]~67 ));
defparam \result_real_1_tmp[17]~66 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[17]~66 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[18]~68 (
	.dataa(\result_a_c_se[18]~q ),
	.datab(\result_b_d_se[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[17]~67 ),
	.combout(\result_real_1_tmp[18]~68_combout ),
	.cout(\result_real_1_tmp[18]~69 ));
defparam \result_real_1_tmp[18]~68 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[18]~68 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[19]~70 (
	.dataa(\result_a_c_se[19]~q ),
	.datab(\result_b_d_se[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[18]~69 ),
	.combout(\result_real_1_tmp[19]~70_combout ),
	.cout(\result_real_1_tmp[19]~71 ));
defparam \result_real_1_tmp[19]~70 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[19]~70 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[20]~72 (
	.dataa(\result_a_c_se[20]~q ),
	.datab(\result_b_d_se[20]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[19]~71 ),
	.combout(\result_real_1_tmp[20]~72_combout ),
	.cout(\result_real_1_tmp[20]~73 ));
defparam \result_real_1_tmp[20]~72 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[20]~72 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[21]~74 (
	.dataa(\result_a_c_se[21]~q ),
	.datab(\result_b_d_se[21]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[20]~73 ),
	.combout(\result_real_1_tmp[21]~74_combout ),
	.cout(\result_real_1_tmp[21]~75 ));
defparam \result_real_1_tmp[21]~74 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[21]~74 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[22]~76 (
	.dataa(\result_a_c_se[22]~q ),
	.datab(\result_b_d_se[22]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[21]~75 ),
	.combout(\result_real_1_tmp[22]~76_combout ),
	.cout(\result_real_1_tmp[22]~77 ));
defparam \result_real_1_tmp[22]~76 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[22]~76 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[23]~78 (
	.dataa(\result_a_c_se[23]~q ),
	.datab(\result_b_d_se[23]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[22]~77 ),
	.combout(\result_real_1_tmp[23]~78_combout ),
	.cout(\result_real_1_tmp[23]~79 ));
defparam \result_real_1_tmp[23]~78 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[23]~78 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[24]~80 (
	.dataa(\result_a_c_se[24]~q ),
	.datab(\result_b_d_se[24]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[23]~79 ),
	.combout(\result_real_1_tmp[24]~80_combout ),
	.cout(\result_real_1_tmp[24]~81 ));
defparam \result_real_1_tmp[24]~80 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[24]~80 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[25]~82 (
	.dataa(\result_a_c_se[25]~q ),
	.datab(\result_b_d_se[25]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[24]~81 ),
	.combout(\result_real_1_tmp[25]~82_combout ),
	.cout(\result_real_1_tmp[25]~83 ));
defparam \result_real_1_tmp[25]~82 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[25]~82 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[26]~84 (
	.dataa(\result_a_c_se[26]~q ),
	.datab(\result_b_d_se[26]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[25]~83 ),
	.combout(\result_real_1_tmp[26]~84_combout ),
	.cout(\result_real_1_tmp[26]~85 ));
defparam \result_real_1_tmp[26]~84 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[26]~84 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[27]~86 (
	.dataa(\result_a_c_se[27]~q ),
	.datab(\result_b_d_se[27]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[26]~85 ),
	.combout(\result_real_1_tmp[27]~86_combout ),
	.cout(\result_real_1_tmp[27]~87 ));
defparam \result_real_1_tmp[27]~86 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[27]~86 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[28]~88 (
	.dataa(\result_a_c_se[28]~q ),
	.datab(\result_b_d_se[28]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[27]~87 ),
	.combout(\result_real_1_tmp[28]~88_combout ),
	.cout(\result_real_1_tmp[28]~89 ));
defparam \result_real_1_tmp[28]~88 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[28]~88 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[29]~90 (
	.dataa(\result_a_c_se[29]~q ),
	.datab(\result_b_d_se[29]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[28]~89 ),
	.combout(\result_real_1_tmp[29]~90_combout ),
	.cout(\result_real_1_tmp[29]~91 ));
defparam \result_real_1_tmp[29]~90 .lut_mask = 16'h96DF;
defparam \result_real_1_tmp[29]~90 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[30]~92 (
	.dataa(\result_a_c_se[30]~q ),
	.datab(\result_b_d_se[30]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_real_1_tmp[29]~91 ),
	.combout(\result_real_1_tmp[30]~92_combout ),
	.cout(\result_real_1_tmp[30]~93 ));
defparam \result_real_1_tmp[30]~92 .lut_mask = 16'h96BF;
defparam \result_real_1_tmp[30]~92 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_real_1_tmp[31]~94 (
	.dataa(\result_a_c_se[31]~q ),
	.datab(\result_b_d_se[31]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\result_real_1_tmp[30]~93 ),
	.combout(\result_real_1_tmp[31]~94_combout ),
	.cout());
defparam \result_real_1_tmp[31]~94 .lut_mask = 16'h9696;
defparam \result_real_1_tmp[31]~94 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[0]~32 (
	.dataa(\result_a_c_se[0]~q ),
	.datab(\result_b_d_se[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\addresult_ac_bd[0]~32_combout ),
	.cout(\addresult_ac_bd[0]~33 ));
defparam \addresult_ac_bd[0]~32 .lut_mask = 16'h66EE;
defparam \addresult_ac_bd[0]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addresult_ac_bd[1]~34 (
	.dataa(\result_a_c_se[1]~q ),
	.datab(\result_b_d_se[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[0]~33 ),
	.combout(\addresult_ac_bd[1]~34_combout ),
	.cout(\addresult_ac_bd[1]~35 ));
defparam \addresult_ac_bd[1]~34 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[1]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[2]~36 (
	.dataa(\result_a_c_se[2]~q ),
	.datab(\result_b_d_se[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[1]~35 ),
	.combout(\addresult_ac_bd[2]~36_combout ),
	.cout(\addresult_ac_bd[2]~37 ));
defparam \addresult_ac_bd[2]~36 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[2]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[3]~38 (
	.dataa(\result_a_c_se[3]~q ),
	.datab(\result_b_d_se[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[2]~37 ),
	.combout(\addresult_ac_bd[3]~38_combout ),
	.cout(\addresult_ac_bd[3]~39 ));
defparam \addresult_ac_bd[3]~38 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[3]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[4]~40 (
	.dataa(\result_a_c_se[4]~q ),
	.datab(\result_b_d_se[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[3]~39 ),
	.combout(\addresult_ac_bd[4]~40_combout ),
	.cout(\addresult_ac_bd[4]~41 ));
defparam \addresult_ac_bd[4]~40 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[4]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[5]~42 (
	.dataa(\result_a_c_se[5]~q ),
	.datab(\result_b_d_se[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[4]~41 ),
	.combout(\addresult_ac_bd[5]~42_combout ),
	.cout(\addresult_ac_bd[5]~43 ));
defparam \addresult_ac_bd[5]~42 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[5]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[6]~44 (
	.dataa(\result_a_c_se[6]~q ),
	.datab(\result_b_d_se[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[5]~43 ),
	.combout(\addresult_ac_bd[6]~44_combout ),
	.cout(\addresult_ac_bd[6]~45 ));
defparam \addresult_ac_bd[6]~44 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[6]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[7]~46 (
	.dataa(\result_a_c_se[7]~q ),
	.datab(\result_b_d_se[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[6]~45 ),
	.combout(\addresult_ac_bd[7]~46_combout ),
	.cout(\addresult_ac_bd[7]~47 ));
defparam \addresult_ac_bd[7]~46 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[7]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[8]~48 (
	.dataa(\result_a_c_se[8]~q ),
	.datab(\result_b_d_se[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[7]~47 ),
	.combout(\addresult_ac_bd[8]~48_combout ),
	.cout(\addresult_ac_bd[8]~49 ));
defparam \addresult_ac_bd[8]~48 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[8]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[9]~50 (
	.dataa(\result_a_c_se[9]~q ),
	.datab(\result_b_d_se[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[8]~49 ),
	.combout(\addresult_ac_bd[9]~50_combout ),
	.cout(\addresult_ac_bd[9]~51 ));
defparam \addresult_ac_bd[9]~50 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[9]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[10]~52 (
	.dataa(\result_a_c_se[10]~q ),
	.datab(\result_b_d_se[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[9]~51 ),
	.combout(\addresult_ac_bd[10]~52_combout ),
	.cout(\addresult_ac_bd[10]~53 ));
defparam \addresult_ac_bd[10]~52 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[10]~52 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[11]~54 (
	.dataa(\result_a_c_se[11]~q ),
	.datab(\result_b_d_se[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[10]~53 ),
	.combout(\addresult_ac_bd[11]~54_combout ),
	.cout(\addresult_ac_bd[11]~55 ));
defparam \addresult_ac_bd[11]~54 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[11]~54 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[12]~56 (
	.dataa(\result_a_c_se[12]~q ),
	.datab(\result_b_d_se[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[11]~55 ),
	.combout(\addresult_ac_bd[12]~56_combout ),
	.cout(\addresult_ac_bd[12]~57 ));
defparam \addresult_ac_bd[12]~56 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[12]~56 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[13]~58 (
	.dataa(\result_a_c_se[13]~q ),
	.datab(\result_b_d_se[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[12]~57 ),
	.combout(\addresult_ac_bd[13]~58_combout ),
	.cout(\addresult_ac_bd[13]~59 ));
defparam \addresult_ac_bd[13]~58 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[13]~58 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[14]~60 (
	.dataa(\result_a_c_se[14]~q ),
	.datab(\result_b_d_se[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[13]~59 ),
	.combout(\addresult_ac_bd[14]~60_combout ),
	.cout(\addresult_ac_bd[14]~61 ));
defparam \addresult_ac_bd[14]~60 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[14]~60 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[15]~62 (
	.dataa(\result_a_c_se[15]~q ),
	.datab(\result_b_d_se[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[14]~61 ),
	.combout(\addresult_ac_bd[15]~62_combout ),
	.cout(\addresult_ac_bd[15]~63 ));
defparam \addresult_ac_bd[15]~62 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[15]~62 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[16]~64 (
	.dataa(\result_a_c_se[16]~q ),
	.datab(\result_b_d_se[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[15]~63 ),
	.combout(\addresult_ac_bd[16]~64_combout ),
	.cout(\addresult_ac_bd[16]~65 ));
defparam \addresult_ac_bd[16]~64 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[16]~64 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[17]~66 (
	.dataa(\result_a_c_se[17]~q ),
	.datab(\result_b_d_se[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[16]~65 ),
	.combout(\addresult_ac_bd[17]~66_combout ),
	.cout(\addresult_ac_bd[17]~67 ));
defparam \addresult_ac_bd[17]~66 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[17]~66 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[18]~68 (
	.dataa(\result_a_c_se[18]~q ),
	.datab(\result_b_d_se[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[17]~67 ),
	.combout(\addresult_ac_bd[18]~68_combout ),
	.cout(\addresult_ac_bd[18]~69 ));
defparam \addresult_ac_bd[18]~68 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[18]~68 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[19]~70 (
	.dataa(\result_a_c_se[19]~q ),
	.datab(\result_b_d_se[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[18]~69 ),
	.combout(\addresult_ac_bd[19]~70_combout ),
	.cout(\addresult_ac_bd[19]~71 ));
defparam \addresult_ac_bd[19]~70 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[19]~70 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[20]~72 (
	.dataa(\result_a_c_se[20]~q ),
	.datab(\result_b_d_se[20]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[19]~71 ),
	.combout(\addresult_ac_bd[20]~72_combout ),
	.cout(\addresult_ac_bd[20]~73 ));
defparam \addresult_ac_bd[20]~72 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[20]~72 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[21]~74 (
	.dataa(\result_a_c_se[21]~q ),
	.datab(\result_b_d_se[21]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[20]~73 ),
	.combout(\addresult_ac_bd[21]~74_combout ),
	.cout(\addresult_ac_bd[21]~75 ));
defparam \addresult_ac_bd[21]~74 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[21]~74 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[22]~76 (
	.dataa(\result_a_c_se[22]~q ),
	.datab(\result_b_d_se[22]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[21]~75 ),
	.combout(\addresult_ac_bd[22]~76_combout ),
	.cout(\addresult_ac_bd[22]~77 ));
defparam \addresult_ac_bd[22]~76 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[22]~76 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[23]~78 (
	.dataa(\result_a_c_se[23]~q ),
	.datab(\result_b_d_se[23]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[22]~77 ),
	.combout(\addresult_ac_bd[23]~78_combout ),
	.cout(\addresult_ac_bd[23]~79 ));
defparam \addresult_ac_bd[23]~78 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[23]~78 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[24]~80 (
	.dataa(\result_a_c_se[24]~q ),
	.datab(\result_b_d_se[24]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[23]~79 ),
	.combout(\addresult_ac_bd[24]~80_combout ),
	.cout(\addresult_ac_bd[24]~81 ));
defparam \addresult_ac_bd[24]~80 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[24]~80 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[25]~82 (
	.dataa(\result_a_c_se[25]~q ),
	.datab(\result_b_d_se[25]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[24]~81 ),
	.combout(\addresult_ac_bd[25]~82_combout ),
	.cout(\addresult_ac_bd[25]~83 ));
defparam \addresult_ac_bd[25]~82 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[25]~82 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[26]~84 (
	.dataa(\result_a_c_se[26]~q ),
	.datab(\result_b_d_se[26]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[25]~83 ),
	.combout(\addresult_ac_bd[26]~84_combout ),
	.cout(\addresult_ac_bd[26]~85 ));
defparam \addresult_ac_bd[26]~84 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[26]~84 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[27]~86 (
	.dataa(\result_a_c_se[27]~q ),
	.datab(\result_b_d_se[27]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[26]~85 ),
	.combout(\addresult_ac_bd[27]~86_combout ),
	.cout(\addresult_ac_bd[27]~87 ));
defparam \addresult_ac_bd[27]~86 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[27]~86 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[28]~88 (
	.dataa(\result_a_c_se[28]~q ),
	.datab(\result_b_d_se[28]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[27]~87 ),
	.combout(\addresult_ac_bd[28]~88_combout ),
	.cout(\addresult_ac_bd[28]~89 ));
defparam \addresult_ac_bd[28]~88 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[28]~88 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[29]~90 (
	.dataa(\result_a_c_se[29]~q ),
	.datab(\result_b_d_se[29]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[28]~89 ),
	.combout(\addresult_ac_bd[29]~90_combout ),
	.cout(\addresult_ac_bd[29]~91 ));
defparam \addresult_ac_bd[29]~90 .lut_mask = 16'h967F;
defparam \addresult_ac_bd[29]~90 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[30]~92 (
	.dataa(\result_a_c_se[30]~q ),
	.datab(\result_b_d_se[30]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_ac_bd[29]~91 ),
	.combout(\addresult_ac_bd[30]~92_combout ),
	.cout(\addresult_ac_bd[30]~93 ));
defparam \addresult_ac_bd[30]~92 .lut_mask = 16'h96EF;
defparam \addresult_ac_bd[30]~92 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_ac_bd[31]~94 (
	.dataa(\result_a_c_se[31]~q ),
	.datab(\result_b_d_se[31]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\addresult_ac_bd[30]~93 ),
	.combout(\addresult_ac_bd[31]~94_combout ),
	.cout());
defparam \addresult_ac_bd[31]~94 .lut_mask = 16'h9696;
defparam \addresult_ac_bd[31]~94 .sum_lutc_input = "cin";

dffeas \addresult_a_b[0] (
	.clk(clk),
	.d(\addresult_a_b[0]~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[0]~q ),
	.prn(vcc));
defparam \addresult_a_b[0] .is_wysiwyg = "true";
defparam \addresult_a_b[0] .power_up = "low";

dffeas \addresult_a_b[1] (
	.clk(clk),
	.d(\addresult_a_b[1]~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[1]~q ),
	.prn(vcc));
defparam \addresult_a_b[1] .is_wysiwyg = "true";
defparam \addresult_a_b[1] .power_up = "low";

dffeas \addresult_a_b[2] (
	.clk(clk),
	.d(\addresult_a_b[2]~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[2]~q ),
	.prn(vcc));
defparam \addresult_a_b[2] .is_wysiwyg = "true";
defparam \addresult_a_b[2] .power_up = "low";

dffeas \addresult_a_b[3] (
	.clk(clk),
	.d(\addresult_a_b[3]~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[3]~q ),
	.prn(vcc));
defparam \addresult_a_b[3] .is_wysiwyg = "true";
defparam \addresult_a_b[3] .power_up = "low";

dffeas \addresult_a_b[4] (
	.clk(clk),
	.d(\addresult_a_b[4]~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[4]~q ),
	.prn(vcc));
defparam \addresult_a_b[4] .is_wysiwyg = "true";
defparam \addresult_a_b[4] .power_up = "low";

dffeas \addresult_a_b[5] (
	.clk(clk),
	.d(\addresult_a_b[5]~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[5]~q ),
	.prn(vcc));
defparam \addresult_a_b[5] .is_wysiwyg = "true";
defparam \addresult_a_b[5] .power_up = "low";

dffeas \addresult_a_b[6] (
	.clk(clk),
	.d(\addresult_a_b[6]~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[6]~q ),
	.prn(vcc));
defparam \addresult_a_b[6] .is_wysiwyg = "true";
defparam \addresult_a_b[6] .power_up = "low";

dffeas \addresult_a_b[7] (
	.clk(clk),
	.d(\addresult_a_b[7]~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[7]~q ),
	.prn(vcc));
defparam \addresult_a_b[7] .is_wysiwyg = "true";
defparam \addresult_a_b[7] .power_up = "low";

dffeas \addresult_a_b[8] (
	.clk(clk),
	.d(\addresult_a_b[8]~33_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[8]~q ),
	.prn(vcc));
defparam \addresult_a_b[8] .is_wysiwyg = "true";
defparam \addresult_a_b[8] .power_up = "low";

dffeas \addresult_a_b[9] (
	.clk(clk),
	.d(\addresult_a_b[9]~35_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[9]~q ),
	.prn(vcc));
defparam \addresult_a_b[9] .is_wysiwyg = "true";
defparam \addresult_a_b[9] .power_up = "low";

dffeas \addresult_a_b[10] (
	.clk(clk),
	.d(\addresult_a_b[10]~37_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[10]~q ),
	.prn(vcc));
defparam \addresult_a_b[10] .is_wysiwyg = "true";
defparam \addresult_a_b[10] .power_up = "low";

dffeas \addresult_a_b[11] (
	.clk(clk),
	.d(\addresult_a_b[11]~39_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[11]~q ),
	.prn(vcc));
defparam \addresult_a_b[11] .is_wysiwyg = "true";
defparam \addresult_a_b[11] .power_up = "low";

dffeas \addresult_a_b[12] (
	.clk(clk),
	.d(\addresult_a_b[12]~41_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[12]~q ),
	.prn(vcc));
defparam \addresult_a_b[12] .is_wysiwyg = "true";
defparam \addresult_a_b[12] .power_up = "low";

dffeas \addresult_a_b[13] (
	.clk(clk),
	.d(\addresult_a_b[13]~43_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[13]~q ),
	.prn(vcc));
defparam \addresult_a_b[13] .is_wysiwyg = "true";
defparam \addresult_a_b[13] .power_up = "low";

dffeas \addresult_a_b[14] (
	.clk(clk),
	.d(\addresult_a_b[14]~45_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[14]~q ),
	.prn(vcc));
defparam \addresult_a_b[14] .is_wysiwyg = "true";
defparam \addresult_a_b[14] .power_up = "low";

dffeas \addresult_a_b[15] (
	.clk(clk),
	.d(\addresult_a_b[15]~47_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[15]~q ),
	.prn(vcc));
defparam \addresult_a_b[15] .is_wysiwyg = "true";
defparam \addresult_a_b[15] .power_up = "low";

dffeas \addresult_a_b[16] (
	.clk(clk),
	.d(\addresult_a_b[16]~49_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_a_b[16]~q ),
	.prn(vcc));
defparam \addresult_a_b[16] .is_wysiwyg = "true";
defparam \addresult_a_b[16] .power_up = "low";

dffeas \addresult_c_d[0] (
	.clk(clk),
	.d(\addresult_c_d[0]~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[0]~q ),
	.prn(vcc));
defparam \addresult_c_d[0] .is_wysiwyg = "true";
defparam \addresult_c_d[0] .power_up = "low";

dffeas \addresult_c_d[1] (
	.clk(clk),
	.d(\addresult_c_d[1]~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[1]~q ),
	.prn(vcc));
defparam \addresult_c_d[1] .is_wysiwyg = "true";
defparam \addresult_c_d[1] .power_up = "low";

dffeas \addresult_c_d[2] (
	.clk(clk),
	.d(\addresult_c_d[2]~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[2]~q ),
	.prn(vcc));
defparam \addresult_c_d[2] .is_wysiwyg = "true";
defparam \addresult_c_d[2] .power_up = "low";

dffeas \addresult_c_d[3] (
	.clk(clk),
	.d(\addresult_c_d[3]~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[3]~q ),
	.prn(vcc));
defparam \addresult_c_d[3] .is_wysiwyg = "true";
defparam \addresult_c_d[3] .power_up = "low";

dffeas \addresult_c_d[4] (
	.clk(clk),
	.d(\addresult_c_d[4]~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[4]~q ),
	.prn(vcc));
defparam \addresult_c_d[4] .is_wysiwyg = "true";
defparam \addresult_c_d[4] .power_up = "low";

dffeas \addresult_c_d[5] (
	.clk(clk),
	.d(\addresult_c_d[5]~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[5]~q ),
	.prn(vcc));
defparam \addresult_c_d[5] .is_wysiwyg = "true";
defparam \addresult_c_d[5] .power_up = "low";

dffeas \addresult_c_d[6] (
	.clk(clk),
	.d(\addresult_c_d[6]~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[6]~q ),
	.prn(vcc));
defparam \addresult_c_d[6] .is_wysiwyg = "true";
defparam \addresult_c_d[6] .power_up = "low";

dffeas \addresult_c_d[7] (
	.clk(clk),
	.d(\addresult_c_d[7]~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[7]~q ),
	.prn(vcc));
defparam \addresult_c_d[7] .is_wysiwyg = "true";
defparam \addresult_c_d[7] .power_up = "low";

dffeas \addresult_c_d[8] (
	.clk(clk),
	.d(\addresult_c_d[8]~33_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[8]~q ),
	.prn(vcc));
defparam \addresult_c_d[8] .is_wysiwyg = "true";
defparam \addresult_c_d[8] .power_up = "low";

dffeas \addresult_c_d[9] (
	.clk(clk),
	.d(\addresult_c_d[9]~35_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[9]~q ),
	.prn(vcc));
defparam \addresult_c_d[9] .is_wysiwyg = "true";
defparam \addresult_c_d[9] .power_up = "low";

dffeas \addresult_c_d[10] (
	.clk(clk),
	.d(\addresult_c_d[10]~37_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[10]~q ),
	.prn(vcc));
defparam \addresult_c_d[10] .is_wysiwyg = "true";
defparam \addresult_c_d[10] .power_up = "low";

dffeas \addresult_c_d[11] (
	.clk(clk),
	.d(\addresult_c_d[11]~39_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[11]~q ),
	.prn(vcc));
defparam \addresult_c_d[11] .is_wysiwyg = "true";
defparam \addresult_c_d[11] .power_up = "low";

dffeas \addresult_c_d[12] (
	.clk(clk),
	.d(\addresult_c_d[12]~41_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[12]~q ),
	.prn(vcc));
defparam \addresult_c_d[12] .is_wysiwyg = "true";
defparam \addresult_c_d[12] .power_up = "low";

dffeas \addresult_c_d[13] (
	.clk(clk),
	.d(\addresult_c_d[13]~43_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[13]~q ),
	.prn(vcc));
defparam \addresult_c_d[13] .is_wysiwyg = "true";
defparam \addresult_c_d[13] .power_up = "low";

dffeas \addresult_c_d[14] (
	.clk(clk),
	.d(\addresult_c_d[14]~45_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[14]~q ),
	.prn(vcc));
defparam \addresult_c_d[14] .is_wysiwyg = "true";
defparam \addresult_c_d[14] .power_up = "low";

dffeas \addresult_c_d[15] (
	.clk(clk),
	.d(\addresult_c_d[15]~47_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[15]~q ),
	.prn(vcc));
defparam \addresult_c_d[15] .is_wysiwyg = "true";
defparam \addresult_c_d[15] .power_up = "low";

dffeas \addresult_c_d[16] (
	.clk(clk),
	.d(\addresult_c_d[16]~49_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\addresult_c_d[16]~q ),
	.prn(vcc));
defparam \addresult_c_d[16] .is_wysiwyg = "true";
defparam \addresult_c_d[16] .power_up = "low";

cycloneive_lcell_comb \addresult_a_b[0]~17 (
	.dataa(pipeline_dffe_2),
	.datab(pipeline_dffe_210),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\addresult_a_b[0]~17_combout ),
	.cout(\addresult_a_b[0]~18 ));
defparam \addresult_a_b[0]~17 .lut_mask = 16'h66EE;
defparam \addresult_a_b[0]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addresult_a_b[1]~19 (
	.dataa(pipeline_dffe_3),
	.datab(pipeline_dffe_32),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[0]~18 ),
	.combout(\addresult_a_b[1]~19_combout ),
	.cout(\addresult_a_b[1]~20 ));
defparam \addresult_a_b[1]~19 .lut_mask = 16'h967F;
defparam \addresult_a_b[1]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_a_b[2]~21 (
	.dataa(pipeline_dffe_4),
	.datab(pipeline_dffe_41),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[1]~20 ),
	.combout(\addresult_a_b[2]~21_combout ),
	.cout(\addresult_a_b[2]~22 ));
defparam \addresult_a_b[2]~21 .lut_mask = 16'h96EF;
defparam \addresult_a_b[2]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_a_b[3]~23 (
	.dataa(pipeline_dffe_5),
	.datab(pipeline_dffe_51),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[2]~22 ),
	.combout(\addresult_a_b[3]~23_combout ),
	.cout(\addresult_a_b[3]~24 ));
defparam \addresult_a_b[3]~23 .lut_mask = 16'h967F;
defparam \addresult_a_b[3]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_a_b[4]~25 (
	.dataa(pipeline_dffe_6),
	.datab(pipeline_dffe_61),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[3]~24 ),
	.combout(\addresult_a_b[4]~25_combout ),
	.cout(\addresult_a_b[4]~26 ));
defparam \addresult_a_b[4]~25 .lut_mask = 16'h96EF;
defparam \addresult_a_b[4]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_a_b[5]~27 (
	.dataa(pipeline_dffe_7),
	.datab(pipeline_dffe_71),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[4]~26 ),
	.combout(\addresult_a_b[5]~27_combout ),
	.cout(\addresult_a_b[5]~28 ));
defparam \addresult_a_b[5]~27 .lut_mask = 16'h967F;
defparam \addresult_a_b[5]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_a_b[6]~29 (
	.dataa(pipeline_dffe_8),
	.datab(pipeline_dffe_81),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[5]~28 ),
	.combout(\addresult_a_b[6]~29_combout ),
	.cout(\addresult_a_b[6]~30 ));
defparam \addresult_a_b[6]~29 .lut_mask = 16'h96EF;
defparam \addresult_a_b[6]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_a_b[7]~31 (
	.dataa(pipeline_dffe_9),
	.datab(pipeline_dffe_91),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[6]~30 ),
	.combout(\addresult_a_b[7]~31_combout ),
	.cout(\addresult_a_b[7]~32 ));
defparam \addresult_a_b[7]~31 .lut_mask = 16'h967F;
defparam \addresult_a_b[7]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_a_b[8]~33 (
	.dataa(pipeline_dffe_10),
	.datab(pipeline_dffe_101),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[7]~32 ),
	.combout(\addresult_a_b[8]~33_combout ),
	.cout(\addresult_a_b[8]~34 ));
defparam \addresult_a_b[8]~33 .lut_mask = 16'h96EF;
defparam \addresult_a_b[8]~33 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_a_b[9]~35 (
	.dataa(pipeline_dffe_11),
	.datab(pipeline_dffe_111),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[8]~34 ),
	.combout(\addresult_a_b[9]~35_combout ),
	.cout(\addresult_a_b[9]~36 ));
defparam \addresult_a_b[9]~35 .lut_mask = 16'h967F;
defparam \addresult_a_b[9]~35 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_a_b[10]~37 (
	.dataa(pipeline_dffe_12),
	.datab(pipeline_dffe_121),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[9]~36 ),
	.combout(\addresult_a_b[10]~37_combout ),
	.cout(\addresult_a_b[10]~38 ));
defparam \addresult_a_b[10]~37 .lut_mask = 16'h96EF;
defparam \addresult_a_b[10]~37 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_a_b[11]~39 (
	.dataa(pipeline_dffe_13),
	.datab(pipeline_dffe_131),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[10]~38 ),
	.combout(\addresult_a_b[11]~39_combout ),
	.cout(\addresult_a_b[11]~40 ));
defparam \addresult_a_b[11]~39 .lut_mask = 16'h967F;
defparam \addresult_a_b[11]~39 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_a_b[12]~41 (
	.dataa(pipeline_dffe_14),
	.datab(pipeline_dffe_141),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[11]~40 ),
	.combout(\addresult_a_b[12]~41_combout ),
	.cout(\addresult_a_b[12]~42 ));
defparam \addresult_a_b[12]~41 .lut_mask = 16'h96EF;
defparam \addresult_a_b[12]~41 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_a_b[13]~43 (
	.dataa(pipeline_dffe_15),
	.datab(pipeline_dffe_151),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[12]~42 ),
	.combout(\addresult_a_b[13]~43_combout ),
	.cout(\addresult_a_b[13]~44 ));
defparam \addresult_a_b[13]~43 .lut_mask = 16'h967F;
defparam \addresult_a_b[13]~43 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_a_b[14]~45 (
	.dataa(pipeline_dffe_161),
	.datab(pipeline_dffe_162),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[13]~44 ),
	.combout(\addresult_a_b[14]~45_combout ),
	.cout(\addresult_a_b[14]~46 ));
defparam \addresult_a_b[14]~45 .lut_mask = 16'h96EF;
defparam \addresult_a_b[14]~45 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_a_b[15]~47 (
	.dataa(pipeline_dffe_171),
	.datab(pipeline_dffe_172),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_a_b[14]~46 ),
	.combout(\addresult_a_b[15]~47_combout ),
	.cout(\addresult_a_b[15]~48 ));
defparam \addresult_a_b[15]~47 .lut_mask = 16'h967F;
defparam \addresult_a_b[15]~47 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_a_b[16]~49 (
	.dataa(pipeline_dffe_171),
	.datab(pipeline_dffe_172),
	.datac(gnd),
	.datad(gnd),
	.cin(\addresult_a_b[15]~48 ),
	.combout(\addresult_a_b[16]~49_combout ),
	.cout());
defparam \addresult_a_b[16]~49 .lut_mask = 16'h9696;
defparam \addresult_a_b[16]~49 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_c_d[0]~17 (
	.dataa(twiddle_data_real_0),
	.datab(twiddle_data_imag_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\addresult_c_d[0]~17_combout ),
	.cout(\addresult_c_d[0]~18 ));
defparam \addresult_c_d[0]~17 .lut_mask = 16'h66EE;
defparam \addresult_c_d[0]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addresult_c_d[1]~19 (
	.dataa(twiddle_data_real_1),
	.datab(twiddle_data_imag_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[0]~18 ),
	.combout(\addresult_c_d[1]~19_combout ),
	.cout(\addresult_c_d[1]~20 ));
defparam \addresult_c_d[1]~19 .lut_mask = 16'h967F;
defparam \addresult_c_d[1]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_c_d[2]~21 (
	.dataa(twiddle_data_real_2),
	.datab(twiddle_data_imag_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[1]~20 ),
	.combout(\addresult_c_d[2]~21_combout ),
	.cout(\addresult_c_d[2]~22 ));
defparam \addresult_c_d[2]~21 .lut_mask = 16'h96EF;
defparam \addresult_c_d[2]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_c_d[3]~23 (
	.dataa(twiddle_data_real_3),
	.datab(twiddle_data_imag_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[2]~22 ),
	.combout(\addresult_c_d[3]~23_combout ),
	.cout(\addresult_c_d[3]~24 ));
defparam \addresult_c_d[3]~23 .lut_mask = 16'h967F;
defparam \addresult_c_d[3]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_c_d[4]~25 (
	.dataa(twiddle_data_real_4),
	.datab(twiddle_data_imag_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[3]~24 ),
	.combout(\addresult_c_d[4]~25_combout ),
	.cout(\addresult_c_d[4]~26 ));
defparam \addresult_c_d[4]~25 .lut_mask = 16'h96EF;
defparam \addresult_c_d[4]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_c_d[5]~27 (
	.dataa(twiddle_data_real_5),
	.datab(twiddle_data_imag_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[4]~26 ),
	.combout(\addresult_c_d[5]~27_combout ),
	.cout(\addresult_c_d[5]~28 ));
defparam \addresult_c_d[5]~27 .lut_mask = 16'h967F;
defparam \addresult_c_d[5]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_c_d[6]~29 (
	.dataa(twiddle_data_real_6),
	.datab(twiddle_data_imag_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[5]~28 ),
	.combout(\addresult_c_d[6]~29_combout ),
	.cout(\addresult_c_d[6]~30 ));
defparam \addresult_c_d[6]~29 .lut_mask = 16'h96EF;
defparam \addresult_c_d[6]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_c_d[7]~31 (
	.dataa(twiddle_data_real_7),
	.datab(twiddle_data_imag_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[6]~30 ),
	.combout(\addresult_c_d[7]~31_combout ),
	.cout(\addresult_c_d[7]~32 ));
defparam \addresult_c_d[7]~31 .lut_mask = 16'h967F;
defparam \addresult_c_d[7]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_c_d[8]~33 (
	.dataa(twiddle_data_real_8),
	.datab(twiddle_data_imag_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[7]~32 ),
	.combout(\addresult_c_d[8]~33_combout ),
	.cout(\addresult_c_d[8]~34 ));
defparam \addresult_c_d[8]~33 .lut_mask = 16'h96EF;
defparam \addresult_c_d[8]~33 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_c_d[9]~35 (
	.dataa(twiddle_data_real_9),
	.datab(twiddle_data_imag_9),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[8]~34 ),
	.combout(\addresult_c_d[9]~35_combout ),
	.cout(\addresult_c_d[9]~36 ));
defparam \addresult_c_d[9]~35 .lut_mask = 16'h967F;
defparam \addresult_c_d[9]~35 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_c_d[10]~37 (
	.dataa(twiddle_data_real_10),
	.datab(twiddle_data_imag_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[9]~36 ),
	.combout(\addresult_c_d[10]~37_combout ),
	.cout(\addresult_c_d[10]~38 ));
defparam \addresult_c_d[10]~37 .lut_mask = 16'h96EF;
defparam \addresult_c_d[10]~37 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_c_d[11]~39 (
	.dataa(twiddle_data_real_11),
	.datab(twiddle_data_imag_11),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[10]~38 ),
	.combout(\addresult_c_d[11]~39_combout ),
	.cout(\addresult_c_d[11]~40 ));
defparam \addresult_c_d[11]~39 .lut_mask = 16'h967F;
defparam \addresult_c_d[11]~39 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_c_d[12]~41 (
	.dataa(twiddle_data_real_12),
	.datab(twiddle_data_imag_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[11]~40 ),
	.combout(\addresult_c_d[12]~41_combout ),
	.cout(\addresult_c_d[12]~42 ));
defparam \addresult_c_d[12]~41 .lut_mask = 16'h96EF;
defparam \addresult_c_d[12]~41 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_c_d[13]~43 (
	.dataa(twiddle_data_real_13),
	.datab(twiddle_data_imag_13),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[12]~42 ),
	.combout(\addresult_c_d[13]~43_combout ),
	.cout(\addresult_c_d[13]~44 ));
defparam \addresult_c_d[13]~43 .lut_mask = 16'h967F;
defparam \addresult_c_d[13]~43 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_c_d[14]~45 (
	.dataa(twiddle_data_real_14),
	.datab(twiddle_data_imag_14),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[13]~44 ),
	.combout(\addresult_c_d[14]~45_combout ),
	.cout(\addresult_c_d[14]~46 ));
defparam \addresult_c_d[14]~45 .lut_mask = 16'h96EF;
defparam \addresult_c_d[14]~45 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_c_d[15]~47 (
	.dataa(twiddle_data_imag_15),
	.datab(twiddle_data_real_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\addresult_c_d[14]~46 ),
	.combout(\addresult_c_d[15]~47_combout ),
	.cout(\addresult_c_d[15]~48 ));
defparam \addresult_c_d[15]~47 .lut_mask = 16'h967F;
defparam \addresult_c_d[15]~47 .sum_lutc_input = "cin";

cycloneive_lcell_comb \addresult_c_d[16]~49 (
	.dataa(twiddle_data_imag_15),
	.datab(twiddle_data_real_15),
	.datac(gnd),
	.datad(gnd),
	.cin(\addresult_c_d[15]~48 ),
	.combout(\addresult_c_d[16]~49_combout ),
	.cout());
defparam \addresult_c_d[16]~49 .lut_mask = 16'h9696;
defparam \addresult_c_d[16]~49 .sum_lutc_input = "cin";

dffeas \result_a_b_c_d_se[16] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[16]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[16] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[16] .power_up = "low";

dffeas \result_a_b_c_d_se[15] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[15]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[15] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[15] .power_up = "low";

dffeas \result_a_b_c_d_se[14] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[14]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[14] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[14] .power_up = "low";

dffeas \result_a_b_c_d_se[13] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[13]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[13] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[13] .power_up = "low";

dffeas \result_a_b_c_d_se[12] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[12]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[12] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[12] .power_up = "low";

dffeas \result_a_b_c_d_se[11] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[11]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[11] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[11] .power_up = "low";

dffeas \result_a_b_c_d_se[10] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[10]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[10] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[10] .power_up = "low";

dffeas \result_a_b_c_d_se[9] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[9]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[9] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[9] .power_up = "low";

dffeas \result_a_b_c_d_se[8] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[8]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[8] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[8] .power_up = "low";

dffeas \result_a_b_c_d_se[7] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[7]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[7] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[7] .power_up = "low";

dffeas \result_a_b_c_d_se[6] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[6]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[6] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[6] .power_up = "low";

dffeas \result_a_b_c_d_se[5] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[5]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[5] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[5] .power_up = "low";

dffeas \result_a_b_c_d_se[4] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[4]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[4] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[4] .power_up = "low";

dffeas \result_a_b_c_d_se[3] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[3]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[3] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[3] .power_up = "low";

dffeas \result_a_b_c_d_se[2] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[2]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[2] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[2] .power_up = "low";

dffeas \result_a_b_c_d_se[1] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[1]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[1] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[1] .power_up = "low";

dffeas \result_a_b_c_d_se[0] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[0]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[0] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[0] .power_up = "low";

dffeas \result_a_b_c_d_se[31] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[31]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[31]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[31] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[31] .power_up = "low";

dffeas \result_a_b_c_d_se[30] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[30]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[30]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[30] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[30] .power_up = "low";

dffeas \result_a_b_c_d_se[29] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[29]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[29]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[29] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[29] .power_up = "low";

dffeas \result_a_b_c_d_se[28] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[28]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[28]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[28] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[28] .power_up = "low";

dffeas \result_a_b_c_d_se[27] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[27]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[27]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[27] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[27] .power_up = "low";

dffeas \result_a_b_c_d_se[26] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[26]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[26]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[26] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[26] .power_up = "low";

dffeas \result_a_b_c_d_se[25] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[25]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[25]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[25] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[25] .power_up = "low";

dffeas \result_a_b_c_d_se[24] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[24]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[24]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[24] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[24] .power_up = "low";

dffeas \result_a_b_c_d_se[23] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[23]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[23]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[23] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[23] .power_up = "low";

dffeas \result_a_b_c_d_se[22] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[22]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[22]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[22] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[22] .power_up = "low";

dffeas \result_a_b_c_d_se[21] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[21]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[21]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[21] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[21] .power_up = "low";

dffeas \result_a_b_c_d_se[20] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[20]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[20] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[20] .power_up = "low";

dffeas \result_a_b_c_d_se[19] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[19]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[19] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[19] .power_up = "low";

dffeas \result_a_b_c_d_se[18] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[18]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[18] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[18] .power_up = "low";

dffeas \result_a_b_c_d_se[17] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_b_c_d_se[17]~q ),
	.prn(vcc));
defparam \result_a_b_c_d_se[17] .is_wysiwyg = "true";
defparam \result_a_b_c_d_se[17] .power_up = "low";

dffeas \result_a_c_se[16] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[16]~q ),
	.prn(vcc));
defparam \result_a_c_se[16] .is_wysiwyg = "true";
defparam \result_a_c_se[16] .power_up = "low";

dffeas \result_b_d_se[16] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[16]~q ),
	.prn(vcc));
defparam \result_b_d_se[16] .is_wysiwyg = "true";
defparam \result_b_d_se[16] .power_up = "low";

dffeas \result_a_c_se[15] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[15]~q ),
	.prn(vcc));
defparam \result_a_c_se[15] .is_wysiwyg = "true";
defparam \result_a_c_se[15] .power_up = "low";

dffeas \result_b_d_se[15] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[15]~q ),
	.prn(vcc));
defparam \result_b_d_se[15] .is_wysiwyg = "true";
defparam \result_b_d_se[15] .power_up = "low";

dffeas \result_a_c_se[14] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[14]~q ),
	.prn(vcc));
defparam \result_a_c_se[14] .is_wysiwyg = "true";
defparam \result_a_c_se[14] .power_up = "low";

dffeas \result_b_d_se[14] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[14]~q ),
	.prn(vcc));
defparam \result_b_d_se[14] .is_wysiwyg = "true";
defparam \result_b_d_se[14] .power_up = "low";

dffeas \result_a_c_se[13] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[13]~q ),
	.prn(vcc));
defparam \result_a_c_se[13] .is_wysiwyg = "true";
defparam \result_a_c_se[13] .power_up = "low";

dffeas \result_b_d_se[13] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[13]~q ),
	.prn(vcc));
defparam \result_b_d_se[13] .is_wysiwyg = "true";
defparam \result_b_d_se[13] .power_up = "low";

dffeas \result_a_c_se[12] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[12]~q ),
	.prn(vcc));
defparam \result_a_c_se[12] .is_wysiwyg = "true";
defparam \result_a_c_se[12] .power_up = "low";

dffeas \result_b_d_se[12] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[12]~q ),
	.prn(vcc));
defparam \result_b_d_se[12] .is_wysiwyg = "true";
defparam \result_b_d_se[12] .power_up = "low";

dffeas \result_a_c_se[11] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[11]~q ),
	.prn(vcc));
defparam \result_a_c_se[11] .is_wysiwyg = "true";
defparam \result_a_c_se[11] .power_up = "low";

dffeas \result_b_d_se[11] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[11]~q ),
	.prn(vcc));
defparam \result_b_d_se[11] .is_wysiwyg = "true";
defparam \result_b_d_se[11] .power_up = "low";

dffeas \result_a_c_se[10] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[10]~q ),
	.prn(vcc));
defparam \result_a_c_se[10] .is_wysiwyg = "true";
defparam \result_a_c_se[10] .power_up = "low";

dffeas \result_b_d_se[10] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[10]~q ),
	.prn(vcc));
defparam \result_b_d_se[10] .is_wysiwyg = "true";
defparam \result_b_d_se[10] .power_up = "low";

dffeas \result_a_c_se[9] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[9]~q ),
	.prn(vcc));
defparam \result_a_c_se[9] .is_wysiwyg = "true";
defparam \result_a_c_se[9] .power_up = "low";

dffeas \result_b_d_se[9] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[9]~q ),
	.prn(vcc));
defparam \result_b_d_se[9] .is_wysiwyg = "true";
defparam \result_b_d_se[9] .power_up = "low";

dffeas \result_a_c_se[8] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[8]~q ),
	.prn(vcc));
defparam \result_a_c_se[8] .is_wysiwyg = "true";
defparam \result_a_c_se[8] .power_up = "low";

dffeas \result_b_d_se[8] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[8]~q ),
	.prn(vcc));
defparam \result_b_d_se[8] .is_wysiwyg = "true";
defparam \result_b_d_se[8] .power_up = "low";

dffeas \result_a_c_se[7] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[7]~q ),
	.prn(vcc));
defparam \result_a_c_se[7] .is_wysiwyg = "true";
defparam \result_a_c_se[7] .power_up = "low";

dffeas \result_b_d_se[7] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[7]~q ),
	.prn(vcc));
defparam \result_b_d_se[7] .is_wysiwyg = "true";
defparam \result_b_d_se[7] .power_up = "low";

dffeas \result_a_c_se[6] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[6]~q ),
	.prn(vcc));
defparam \result_a_c_se[6] .is_wysiwyg = "true";
defparam \result_a_c_se[6] .power_up = "low";

dffeas \result_b_d_se[6] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[6]~q ),
	.prn(vcc));
defparam \result_b_d_se[6] .is_wysiwyg = "true";
defparam \result_b_d_se[6] .power_up = "low";

dffeas \result_a_c_se[5] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[5]~q ),
	.prn(vcc));
defparam \result_a_c_se[5] .is_wysiwyg = "true";
defparam \result_a_c_se[5] .power_up = "low";

dffeas \result_b_d_se[5] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[5]~q ),
	.prn(vcc));
defparam \result_b_d_se[5] .is_wysiwyg = "true";
defparam \result_b_d_se[5] .power_up = "low";

dffeas \result_a_c_se[4] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[4]~q ),
	.prn(vcc));
defparam \result_a_c_se[4] .is_wysiwyg = "true";
defparam \result_a_c_se[4] .power_up = "low";

dffeas \result_b_d_se[4] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[4]~q ),
	.prn(vcc));
defparam \result_b_d_se[4] .is_wysiwyg = "true";
defparam \result_b_d_se[4] .power_up = "low";

dffeas \result_a_c_se[3] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[3]~q ),
	.prn(vcc));
defparam \result_a_c_se[3] .is_wysiwyg = "true";
defparam \result_a_c_se[3] .power_up = "low";

dffeas \result_b_d_se[3] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[3]~q ),
	.prn(vcc));
defparam \result_b_d_se[3] .is_wysiwyg = "true";
defparam \result_b_d_se[3] .power_up = "low";

dffeas \result_a_c_se[2] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[2]~q ),
	.prn(vcc));
defparam \result_a_c_se[2] .is_wysiwyg = "true";
defparam \result_a_c_se[2] .power_up = "low";

dffeas \result_b_d_se[2] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[2]~q ),
	.prn(vcc));
defparam \result_b_d_se[2] .is_wysiwyg = "true";
defparam \result_b_d_se[2] .power_up = "low";

dffeas \result_a_c_se[1] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[1]~q ),
	.prn(vcc));
defparam \result_a_c_se[1] .is_wysiwyg = "true";
defparam \result_a_c_se[1] .power_up = "low";

dffeas \result_b_d_se[1] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[1]~q ),
	.prn(vcc));
defparam \result_b_d_se[1] .is_wysiwyg = "true";
defparam \result_b_d_se[1] .power_up = "low";

dffeas \result_a_c_se[0] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[0]~q ),
	.prn(vcc));
defparam \result_a_c_se[0] .is_wysiwyg = "true";
defparam \result_a_c_se[0] .power_up = "low";

dffeas \result_b_d_se[0] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[0]~q ),
	.prn(vcc));
defparam \result_b_d_se[0] .is_wysiwyg = "true";
defparam \result_b_d_se[0] .power_up = "low";

dffeas \result_a_c_se[31] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[31]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[31]~q ),
	.prn(vcc));
defparam \result_a_c_se[31] .is_wysiwyg = "true";
defparam \result_a_c_se[31] .power_up = "low";

dffeas \result_b_d_se[31] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[31]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[31]~q ),
	.prn(vcc));
defparam \result_b_d_se[31] .is_wysiwyg = "true";
defparam \result_b_d_se[31] .power_up = "low";

dffeas \result_a_c_se[30] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[30]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[30]~q ),
	.prn(vcc));
defparam \result_a_c_se[30] .is_wysiwyg = "true";
defparam \result_a_c_se[30] .power_up = "low";

dffeas \result_b_d_se[30] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[30]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[30]~q ),
	.prn(vcc));
defparam \result_b_d_se[30] .is_wysiwyg = "true";
defparam \result_b_d_se[30] .power_up = "low";

dffeas \result_a_c_se[29] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[29]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[29]~q ),
	.prn(vcc));
defparam \result_a_c_se[29] .is_wysiwyg = "true";
defparam \result_a_c_se[29] .power_up = "low";

dffeas \result_b_d_se[29] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[29]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[29]~q ),
	.prn(vcc));
defparam \result_b_d_se[29] .is_wysiwyg = "true";
defparam \result_b_d_se[29] .power_up = "low";

dffeas \result_a_c_se[28] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[28]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[28]~q ),
	.prn(vcc));
defparam \result_a_c_se[28] .is_wysiwyg = "true";
defparam \result_a_c_se[28] .power_up = "low";

dffeas \result_b_d_se[28] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[28]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[28]~q ),
	.prn(vcc));
defparam \result_b_d_se[28] .is_wysiwyg = "true";
defparam \result_b_d_se[28] .power_up = "low";

dffeas \result_a_c_se[27] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[27]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[27]~q ),
	.prn(vcc));
defparam \result_a_c_se[27] .is_wysiwyg = "true";
defparam \result_a_c_se[27] .power_up = "low";

dffeas \result_b_d_se[27] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[27]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[27]~q ),
	.prn(vcc));
defparam \result_b_d_se[27] .is_wysiwyg = "true";
defparam \result_b_d_se[27] .power_up = "low";

dffeas \result_a_c_se[26] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[26]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[26]~q ),
	.prn(vcc));
defparam \result_a_c_se[26] .is_wysiwyg = "true";
defparam \result_a_c_se[26] .power_up = "low";

dffeas \result_b_d_se[26] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[26]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[26]~q ),
	.prn(vcc));
defparam \result_b_d_se[26] .is_wysiwyg = "true";
defparam \result_b_d_se[26] .power_up = "low";

dffeas \result_a_c_se[25] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[25]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[25]~q ),
	.prn(vcc));
defparam \result_a_c_se[25] .is_wysiwyg = "true";
defparam \result_a_c_se[25] .power_up = "low";

dffeas \result_b_d_se[25] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[25]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[25]~q ),
	.prn(vcc));
defparam \result_b_d_se[25] .is_wysiwyg = "true";
defparam \result_b_d_se[25] .power_up = "low";

dffeas \result_a_c_se[24] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[24]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[24]~q ),
	.prn(vcc));
defparam \result_a_c_se[24] .is_wysiwyg = "true";
defparam \result_a_c_se[24] .power_up = "low";

dffeas \result_b_d_se[24] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[24]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[24]~q ),
	.prn(vcc));
defparam \result_b_d_se[24] .is_wysiwyg = "true";
defparam \result_b_d_se[24] .power_up = "low";

dffeas \result_a_c_se[23] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[23]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[23]~q ),
	.prn(vcc));
defparam \result_a_c_se[23] .is_wysiwyg = "true";
defparam \result_a_c_se[23] .power_up = "low";

dffeas \result_b_d_se[23] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[23]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[23]~q ),
	.prn(vcc));
defparam \result_b_d_se[23] .is_wysiwyg = "true";
defparam \result_b_d_se[23] .power_up = "low";

dffeas \result_a_c_se[22] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[22]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[22]~q ),
	.prn(vcc));
defparam \result_a_c_se[22] .is_wysiwyg = "true";
defparam \result_a_c_se[22] .power_up = "low";

dffeas \result_b_d_se[22] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[22]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[22]~q ),
	.prn(vcc));
defparam \result_b_d_se[22] .is_wysiwyg = "true";
defparam \result_b_d_se[22] .power_up = "low";

dffeas \result_a_c_se[21] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[21]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[21]~q ),
	.prn(vcc));
defparam \result_a_c_se[21] .is_wysiwyg = "true";
defparam \result_a_c_se[21] .power_up = "low";

dffeas \result_b_d_se[21] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[21]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[21]~q ),
	.prn(vcc));
defparam \result_b_d_se[21] .is_wysiwyg = "true";
defparam \result_b_d_se[21] .power_up = "low";

dffeas \result_a_c_se[20] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[20]~q ),
	.prn(vcc));
defparam \result_a_c_se[20] .is_wysiwyg = "true";
defparam \result_a_c_se[20] .power_up = "low";

dffeas \result_b_d_se[20] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[20]~q ),
	.prn(vcc));
defparam \result_b_d_se[20] .is_wysiwyg = "true";
defparam \result_b_d_se[20] .power_up = "low";

dffeas \result_a_c_se[19] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[19]~q ),
	.prn(vcc));
defparam \result_a_c_se[19] .is_wysiwyg = "true";
defparam \result_a_c_se[19] .power_up = "low";

dffeas \result_b_d_se[19] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[19]~q ),
	.prn(vcc));
defparam \result_b_d_se[19] .is_wysiwyg = "true";
defparam \result_b_d_se[19] .power_up = "low";

dffeas \result_a_c_se[18] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[18]~q ),
	.prn(vcc));
defparam \result_a_c_se[18] .is_wysiwyg = "true";
defparam \result_a_c_se[18] .power_up = "low";

dffeas \result_b_d_se[18] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[18]~q ),
	.prn(vcc));
defparam \result_b_d_se[18] .is_wysiwyg = "true";
defparam \result_b_d_se[18] .power_up = "low";

dffeas \result_a_c_se[17] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_a_c_se[17]~q ),
	.prn(vcc));
defparam \result_a_c_se[17] .is_wysiwyg = "true";
defparam \result_a_c_se[17] .power_up = "low";

dffeas \result_b_d_se[17] (
	.clk(clk),
	.d(\gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_b_d_se[17]~q ),
	.prn(vcc));
defparam \result_b_d_se[17] .is_wysiwyg = "true";
defparam \result_b_d_se[17] .power_up = "low";

dffeas \real_out[0] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_0),
	.prn(vcc));
defparam \real_out[0] .is_wysiwyg = "true";
defparam \real_out[0] .power_up = "low";

dffeas \real_out[1] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_1),
	.prn(vcc));
defparam \real_out[1] .is_wysiwyg = "true";
defparam \real_out[1] .power_up = "low";

dffeas \real_out[2] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_2),
	.prn(vcc));
defparam \real_out[2] .is_wysiwyg = "true";
defparam \real_out[2] .power_up = "low";

dffeas \real_out[3] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_3),
	.prn(vcc));
defparam \real_out[3] .is_wysiwyg = "true";
defparam \real_out[3] .power_up = "low";

dffeas \real_out[4] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_4),
	.prn(vcc));
defparam \real_out[4] .is_wysiwyg = "true";
defparam \real_out[4] .power_up = "low";

dffeas \real_out[5] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_5),
	.prn(vcc));
defparam \real_out[5] .is_wysiwyg = "true";
defparam \real_out[5] .power_up = "low";

dffeas \real_out[6] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_6),
	.prn(vcc));
defparam \real_out[6] .is_wysiwyg = "true";
defparam \real_out[6] .power_up = "low";

dffeas \real_out[7] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_7),
	.prn(vcc));
defparam \real_out[7] .is_wysiwyg = "true";
defparam \real_out[7] .power_up = "low";

dffeas \real_out[8] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_8),
	.prn(vcc));
defparam \real_out[8] .is_wysiwyg = "true";
defparam \real_out[8] .power_up = "low";

dffeas \real_out[9] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_9),
	.prn(vcc));
defparam \real_out[9] .is_wysiwyg = "true";
defparam \real_out[9] .power_up = "low";

dffeas \real_out[10] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_10),
	.prn(vcc));
defparam \real_out[10] .is_wysiwyg = "true";
defparam \real_out[10] .power_up = "low";

dffeas \real_out[11] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_11),
	.prn(vcc));
defparam \real_out[11] .is_wysiwyg = "true";
defparam \real_out[11] .power_up = "low";

dffeas \real_out[12] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_12),
	.prn(vcc));
defparam \real_out[12] .is_wysiwyg = "true";
defparam \real_out[12] .power_up = "low";

dffeas \real_out[13] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_13),
	.prn(vcc));
defparam \real_out[13] .is_wysiwyg = "true";
defparam \real_out[13] .power_up = "low";

dffeas \real_out[14] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_14),
	.prn(vcc));
defparam \real_out[14] .is_wysiwyg = "true";
defparam \real_out[14] .power_up = "low";

dffeas \real_out[15] (
	.clk(clk),
	.d(\gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(real_out_15),
	.prn(vcc));
defparam \real_out[15] .is_wysiwyg = "true";
defparam \real_out[15] .power_up = "low";

endmodule

module fft256_asj_fft_pround_fft_121 (
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_31,
	result_real_1_tmp_16,
	result_real_1_tmp_15,
	result_real_1_tmp_14,
	result_real_1_tmp_13,
	result_real_1_tmp_12,
	result_real_1_tmp_11,
	result_real_1_tmp_10,
	result_real_1_tmp_9,
	result_real_1_tmp_8,
	result_real_1_tmp_7,
	result_real_1_tmp_6,
	result_real_1_tmp_5,
	result_real_1_tmp_4,
	result_real_1_tmp_3,
	result_real_1_tmp_2,
	result_real_1_tmp_1,
	result_real_1_tmp_0,
	result_real_1_tmp_31,
	result_real_1_tmp_17,
	result_real_1_tmp_18,
	result_real_1_tmp_19,
	result_real_1_tmp_20,
	result_real_1_tmp_21,
	result_real_1_tmp_22,
	result_real_1_tmp_23,
	result_real_1_tmp_24,
	result_real_1_tmp_25,
	result_real_1_tmp_26,
	result_real_1_tmp_27,
	result_real_1_tmp_28,
	result_real_1_tmp_29,
	result_real_1_tmp_30,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_31;
input 	result_real_1_tmp_16;
input 	result_real_1_tmp_15;
input 	result_real_1_tmp_14;
input 	result_real_1_tmp_13;
input 	result_real_1_tmp_12;
input 	result_real_1_tmp_11;
input 	result_real_1_tmp_10;
input 	result_real_1_tmp_9;
input 	result_real_1_tmp_8;
input 	result_real_1_tmp_7;
input 	result_real_1_tmp_6;
input 	result_real_1_tmp_5;
input 	result_real_1_tmp_4;
input 	result_real_1_tmp_3;
input 	result_real_1_tmp_2;
input 	result_real_1_tmp_1;
input 	result_real_1_tmp_0;
input 	result_real_1_tmp_31;
input 	result_real_1_tmp_17;
input 	result_real_1_tmp_18;
input 	result_real_1_tmp_19;
input 	result_real_1_tmp_20;
input 	result_real_1_tmp_21;
input 	result_real_1_tmp_22;
input 	result_real_1_tmp_23;
input 	result_real_1_tmp_24;
input 	result_real_1_tmp_25;
input 	result_real_1_tmp_26;
input 	result_real_1_tmp_27;
input 	result_real_1_tmp_28;
input 	result_real_1_tmp_29;
input 	result_real_1_tmp_30;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_LPM_ADD_SUB_1 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_31(pipeline_dffe_31),
	.result_real_1_tmp_16(result_real_1_tmp_16),
	.result_real_1_tmp_15(result_real_1_tmp_15),
	.result_real_1_tmp_14(result_real_1_tmp_14),
	.result_real_1_tmp_13(result_real_1_tmp_13),
	.result_real_1_tmp_12(result_real_1_tmp_12),
	.result_real_1_tmp_11(result_real_1_tmp_11),
	.result_real_1_tmp_10(result_real_1_tmp_10),
	.result_real_1_tmp_9(result_real_1_tmp_9),
	.result_real_1_tmp_8(result_real_1_tmp_8),
	.result_real_1_tmp_7(result_real_1_tmp_7),
	.result_real_1_tmp_6(result_real_1_tmp_6),
	.result_real_1_tmp_5(result_real_1_tmp_5),
	.result_real_1_tmp_4(result_real_1_tmp_4),
	.result_real_1_tmp_3(result_real_1_tmp_3),
	.result_real_1_tmp_2(result_real_1_tmp_2),
	.result_real_1_tmp_1(result_real_1_tmp_1),
	.result_real_1_tmp_0(result_real_1_tmp_0),
	.result_real_1_tmp_31(result_real_1_tmp_31),
	.result_real_1_tmp_17(result_real_1_tmp_17),
	.result_real_1_tmp_18(result_real_1_tmp_18),
	.result_real_1_tmp_19(result_real_1_tmp_19),
	.result_real_1_tmp_20(result_real_1_tmp_20),
	.result_real_1_tmp_21(result_real_1_tmp_21),
	.result_real_1_tmp_22(result_real_1_tmp_22),
	.result_real_1_tmp_23(result_real_1_tmp_23),
	.result_real_1_tmp_24(result_real_1_tmp_24),
	.result_real_1_tmp_25(result_real_1_tmp_25),
	.result_real_1_tmp_26(result_real_1_tmp_26),
	.result_real_1_tmp_27(result_real_1_tmp_27),
	.result_real_1_tmp_28(result_real_1_tmp_28),
	.result_real_1_tmp_29(result_real_1_tmp_29),
	.result_real_1_tmp_30(result_real_1_tmp_30),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft256_LPM_ADD_SUB_1 (
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_31,
	result_real_1_tmp_16,
	result_real_1_tmp_15,
	result_real_1_tmp_14,
	result_real_1_tmp_13,
	result_real_1_tmp_12,
	result_real_1_tmp_11,
	result_real_1_tmp_10,
	result_real_1_tmp_9,
	result_real_1_tmp_8,
	result_real_1_tmp_7,
	result_real_1_tmp_6,
	result_real_1_tmp_5,
	result_real_1_tmp_4,
	result_real_1_tmp_3,
	result_real_1_tmp_2,
	result_real_1_tmp_1,
	result_real_1_tmp_0,
	result_real_1_tmp_31,
	result_real_1_tmp_17,
	result_real_1_tmp_18,
	result_real_1_tmp_19,
	result_real_1_tmp_20,
	result_real_1_tmp_21,
	result_real_1_tmp_22,
	result_real_1_tmp_23,
	result_real_1_tmp_24,
	result_real_1_tmp_25,
	result_real_1_tmp_26,
	result_real_1_tmp_27,
	result_real_1_tmp_28,
	result_real_1_tmp_29,
	result_real_1_tmp_30,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_31;
input 	result_real_1_tmp_16;
input 	result_real_1_tmp_15;
input 	result_real_1_tmp_14;
input 	result_real_1_tmp_13;
input 	result_real_1_tmp_12;
input 	result_real_1_tmp_11;
input 	result_real_1_tmp_10;
input 	result_real_1_tmp_9;
input 	result_real_1_tmp_8;
input 	result_real_1_tmp_7;
input 	result_real_1_tmp_6;
input 	result_real_1_tmp_5;
input 	result_real_1_tmp_4;
input 	result_real_1_tmp_3;
input 	result_real_1_tmp_2;
input 	result_real_1_tmp_1;
input 	result_real_1_tmp_0;
input 	result_real_1_tmp_31;
input 	result_real_1_tmp_17;
input 	result_real_1_tmp_18;
input 	result_real_1_tmp_19;
input 	result_real_1_tmp_20;
input 	result_real_1_tmp_21;
input 	result_real_1_tmp_22;
input 	result_real_1_tmp_23;
input 	result_real_1_tmp_24;
input 	result_real_1_tmp_25;
input 	result_real_1_tmp_26;
input 	result_real_1_tmp_27;
input 	result_real_1_tmp_28;
input 	result_real_1_tmp_29;
input 	result_real_1_tmp_30;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_add_sub_knj auto_generated(
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_31(pipeline_dffe_31),
	.result_real_1_tmp_16(result_real_1_tmp_16),
	.result_real_1_tmp_15(result_real_1_tmp_15),
	.result_real_1_tmp_14(result_real_1_tmp_14),
	.result_real_1_tmp_13(result_real_1_tmp_13),
	.result_real_1_tmp_12(result_real_1_tmp_12),
	.result_real_1_tmp_11(result_real_1_tmp_11),
	.result_real_1_tmp_10(result_real_1_tmp_10),
	.result_real_1_tmp_9(result_real_1_tmp_9),
	.result_real_1_tmp_8(result_real_1_tmp_8),
	.result_real_1_tmp_7(result_real_1_tmp_7),
	.result_real_1_tmp_6(result_real_1_tmp_6),
	.result_real_1_tmp_5(result_real_1_tmp_5),
	.result_real_1_tmp_4(result_real_1_tmp_4),
	.result_real_1_tmp_3(result_real_1_tmp_3),
	.result_real_1_tmp_2(result_real_1_tmp_2),
	.result_real_1_tmp_1(result_real_1_tmp_1),
	.result_real_1_tmp_0(result_real_1_tmp_0),
	.result_real_1_tmp_31(result_real_1_tmp_31),
	.result_real_1_tmp_17(result_real_1_tmp_17),
	.result_real_1_tmp_18(result_real_1_tmp_18),
	.result_real_1_tmp_19(result_real_1_tmp_19),
	.result_real_1_tmp_20(result_real_1_tmp_20),
	.result_real_1_tmp_21(result_real_1_tmp_21),
	.result_real_1_tmp_22(result_real_1_tmp_22),
	.result_real_1_tmp_23(result_real_1_tmp_23),
	.result_real_1_tmp_24(result_real_1_tmp_24),
	.result_real_1_tmp_25(result_real_1_tmp_25),
	.result_real_1_tmp_26(result_real_1_tmp_26),
	.result_real_1_tmp_27(result_real_1_tmp_27),
	.result_real_1_tmp_28(result_real_1_tmp_28),
	.result_real_1_tmp_29(result_real_1_tmp_29),
	.result_real_1_tmp_30(result_real_1_tmp_30),
	.clken(clken),
	.clock(clock));

endmodule

module fft256_add_sub_knj (
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_31,
	result_real_1_tmp_16,
	result_real_1_tmp_15,
	result_real_1_tmp_14,
	result_real_1_tmp_13,
	result_real_1_tmp_12,
	result_real_1_tmp_11,
	result_real_1_tmp_10,
	result_real_1_tmp_9,
	result_real_1_tmp_8,
	result_real_1_tmp_7,
	result_real_1_tmp_6,
	result_real_1_tmp_5,
	result_real_1_tmp_4,
	result_real_1_tmp_3,
	result_real_1_tmp_2,
	result_real_1_tmp_1,
	result_real_1_tmp_0,
	result_real_1_tmp_31,
	result_real_1_tmp_17,
	result_real_1_tmp_18,
	result_real_1_tmp_19,
	result_real_1_tmp_20,
	result_real_1_tmp_21,
	result_real_1_tmp_22,
	result_real_1_tmp_23,
	result_real_1_tmp_24,
	result_real_1_tmp_25,
	result_real_1_tmp_26,
	result_real_1_tmp_27,
	result_real_1_tmp_28,
	result_real_1_tmp_29,
	result_real_1_tmp_30,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_31;
input 	result_real_1_tmp_16;
input 	result_real_1_tmp_15;
input 	result_real_1_tmp_14;
input 	result_real_1_tmp_13;
input 	result_real_1_tmp_12;
input 	result_real_1_tmp_11;
input 	result_real_1_tmp_10;
input 	result_real_1_tmp_9;
input 	result_real_1_tmp_8;
input 	result_real_1_tmp_7;
input 	result_real_1_tmp_6;
input 	result_real_1_tmp_5;
input 	result_real_1_tmp_4;
input 	result_real_1_tmp_3;
input 	result_real_1_tmp_2;
input 	result_real_1_tmp_1;
input 	result_real_1_tmp_0;
input 	result_real_1_tmp_31;
input 	result_real_1_tmp_17;
input 	result_real_1_tmp_18;
input 	result_real_1_tmp_19;
input 	result_real_1_tmp_20;
input 	result_real_1_tmp_21;
input 	result_real_1_tmp_22;
input 	result_real_1_tmp_23;
input 	result_real_1_tmp_24;
input 	result_real_1_tmp_25;
input 	result_real_1_tmp_26;
input 	result_real_1_tmp_27;
input 	result_real_1_tmp_28;
input 	result_real_1_tmp_29;
input 	result_real_1_tmp_30;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~17_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~19_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~21_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~23_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~25_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~27_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~29_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~31_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~33_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~35_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~37_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~39_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~41_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~43_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~47_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~49_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~51 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~53 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~54_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~55 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~56_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~57 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~58_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~59 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~60_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~61 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~62_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~63 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~64_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~65 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~66_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~67 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~68_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~69 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~70_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~71 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~72_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~73 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~74_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~75 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~76_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~77 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~78_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~79 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~80_combout ;


dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_18),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_19),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_20),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_21),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_22),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~64_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_23),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_24),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~68_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_25),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~70_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_26),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~72_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_27),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~74_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_28),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~76_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_29),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~78_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_30),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~80_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_31),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31] .power_up = "low";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~17 (
	.dataa(result_real_1_tmp_31),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~17_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~17 .lut_mask = 16'h0055;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~19 (
	.dataa(result_real_1_tmp_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~17_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~19_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~19 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~21 (
	.dataa(result_real_1_tmp_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~19_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~21_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~21 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~23 (
	.dataa(result_real_1_tmp_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~21_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~23_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~23 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~25 (
	.dataa(result_real_1_tmp_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~23_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~25_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~25 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~27 (
	.dataa(result_real_1_tmp_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~25_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~27_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~27 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~29 (
	.dataa(result_real_1_tmp_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~27_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~29_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~29 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~31 (
	.dataa(result_real_1_tmp_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~29_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~31_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~31 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~33 (
	.dataa(result_real_1_tmp_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~31_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~33_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~33 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~33 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~35 (
	.dataa(result_real_1_tmp_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~33_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~35_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~35 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~35 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~37 (
	.dataa(result_real_1_tmp_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~35_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~37_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~37 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~37 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~39 (
	.dataa(result_real_1_tmp_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~37_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~39_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~39 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~39 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~41 (
	.dataa(result_real_1_tmp_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~39_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~41_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~41 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~41 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~43 (
	.dataa(result_real_1_tmp_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~41_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~43_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~43 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~43 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 (
	.dataa(result_real_1_tmp_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~43_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~47 (
	.dataa(result_real_1_tmp_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~47_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~47 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~47 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~49 (
	.dataa(result_real_1_tmp_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~47_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~49_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~49 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~49 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50 (
	.dataa(result_real_1_tmp_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~49_cout ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~51 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52 (
	.dataa(result_real_1_tmp_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~51 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~53 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~54 (
	.dataa(result_real_1_tmp_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~53 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~54_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~55 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~54 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~54 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~56 (
	.dataa(result_real_1_tmp_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~55 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~56_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~57 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~56 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~56 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~58 (
	.dataa(result_real_1_tmp_20),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~57 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~58_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~59 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~58 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~58 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~60 (
	.dataa(result_real_1_tmp_21),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~59 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~60_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~61 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~60 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~60 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~62 (
	.dataa(result_real_1_tmp_22),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~61 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~62_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~63 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~62 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~62 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~64 (
	.dataa(result_real_1_tmp_23),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~63 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~64_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~65 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~64 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~64 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~66 (
	.dataa(result_real_1_tmp_24),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~65 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~66_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~67 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~66 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~66 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~68 (
	.dataa(result_real_1_tmp_25),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~67 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~68_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~69 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~68 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~68 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~70 (
	.dataa(result_real_1_tmp_26),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~69 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~70_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~71 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~70 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~70 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~72 (
	.dataa(result_real_1_tmp_27),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~71 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~72_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~73 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~72 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~72 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~74 (
	.dataa(result_real_1_tmp_28),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~73 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~74_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~75 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~74 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~74 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~76 (
	.dataa(result_real_1_tmp_29),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~75 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~76_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~77 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~76 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~76 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~78 (
	.dataa(result_real_1_tmp_30),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~77 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~78_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~79 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~78 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~78 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~80 (
	.dataa(result_real_1_tmp_31),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~79 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~80_combout ),
	.cout());
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~80 .lut_mask = 16'h5A5A;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~80 .sum_lutc_input = "cin";

endmodule

module fft256_asj_fft_pround_fft_121_1 (
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_31,
	result_imag_1_16,
	result_imag_1_15,
	result_imag_1_14,
	result_imag_1_13,
	result_imag_1_12,
	result_imag_1_11,
	result_imag_1_10,
	result_imag_1_9,
	result_imag_1_8,
	result_imag_1_7,
	result_imag_1_6,
	result_imag_1_5,
	result_imag_1_4,
	result_imag_1_3,
	result_imag_1_2,
	result_imag_1_1,
	result_imag_1_0,
	result_imag_1_31,
	result_imag_1_17,
	result_imag_1_18,
	result_imag_1_19,
	result_imag_1_20,
	result_imag_1_21,
	result_imag_1_22,
	result_imag_1_23,
	result_imag_1_24,
	result_imag_1_25,
	result_imag_1_26,
	result_imag_1_27,
	result_imag_1_28,
	result_imag_1_29,
	result_imag_1_30,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_31;
input 	result_imag_1_16;
input 	result_imag_1_15;
input 	result_imag_1_14;
input 	result_imag_1_13;
input 	result_imag_1_12;
input 	result_imag_1_11;
input 	result_imag_1_10;
input 	result_imag_1_9;
input 	result_imag_1_8;
input 	result_imag_1_7;
input 	result_imag_1_6;
input 	result_imag_1_5;
input 	result_imag_1_4;
input 	result_imag_1_3;
input 	result_imag_1_2;
input 	result_imag_1_1;
input 	result_imag_1_0;
input 	result_imag_1_31;
input 	result_imag_1_17;
input 	result_imag_1_18;
input 	result_imag_1_19;
input 	result_imag_1_20;
input 	result_imag_1_21;
input 	result_imag_1_22;
input 	result_imag_1_23;
input 	result_imag_1_24;
input 	result_imag_1_25;
input 	result_imag_1_26;
input 	result_imag_1_27;
input 	result_imag_1_28;
input 	result_imag_1_29;
input 	result_imag_1_30;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_LPM_ADD_SUB_2 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_31(pipeline_dffe_31),
	.result_imag_1_16(result_imag_1_16),
	.result_imag_1_15(result_imag_1_15),
	.result_imag_1_14(result_imag_1_14),
	.result_imag_1_13(result_imag_1_13),
	.result_imag_1_12(result_imag_1_12),
	.result_imag_1_11(result_imag_1_11),
	.result_imag_1_10(result_imag_1_10),
	.result_imag_1_9(result_imag_1_9),
	.result_imag_1_8(result_imag_1_8),
	.result_imag_1_7(result_imag_1_7),
	.result_imag_1_6(result_imag_1_6),
	.result_imag_1_5(result_imag_1_5),
	.result_imag_1_4(result_imag_1_4),
	.result_imag_1_3(result_imag_1_3),
	.result_imag_1_2(result_imag_1_2),
	.result_imag_1_1(result_imag_1_1),
	.result_imag_1_0(result_imag_1_0),
	.result_imag_1_31(result_imag_1_31),
	.result_imag_1_17(result_imag_1_17),
	.result_imag_1_18(result_imag_1_18),
	.result_imag_1_19(result_imag_1_19),
	.result_imag_1_20(result_imag_1_20),
	.result_imag_1_21(result_imag_1_21),
	.result_imag_1_22(result_imag_1_22),
	.result_imag_1_23(result_imag_1_23),
	.result_imag_1_24(result_imag_1_24),
	.result_imag_1_25(result_imag_1_25),
	.result_imag_1_26(result_imag_1_26),
	.result_imag_1_27(result_imag_1_27),
	.result_imag_1_28(result_imag_1_28),
	.result_imag_1_29(result_imag_1_29),
	.result_imag_1_30(result_imag_1_30),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft256_LPM_ADD_SUB_2 (
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_31,
	result_imag_1_16,
	result_imag_1_15,
	result_imag_1_14,
	result_imag_1_13,
	result_imag_1_12,
	result_imag_1_11,
	result_imag_1_10,
	result_imag_1_9,
	result_imag_1_8,
	result_imag_1_7,
	result_imag_1_6,
	result_imag_1_5,
	result_imag_1_4,
	result_imag_1_3,
	result_imag_1_2,
	result_imag_1_1,
	result_imag_1_0,
	result_imag_1_31,
	result_imag_1_17,
	result_imag_1_18,
	result_imag_1_19,
	result_imag_1_20,
	result_imag_1_21,
	result_imag_1_22,
	result_imag_1_23,
	result_imag_1_24,
	result_imag_1_25,
	result_imag_1_26,
	result_imag_1_27,
	result_imag_1_28,
	result_imag_1_29,
	result_imag_1_30,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_31;
input 	result_imag_1_16;
input 	result_imag_1_15;
input 	result_imag_1_14;
input 	result_imag_1_13;
input 	result_imag_1_12;
input 	result_imag_1_11;
input 	result_imag_1_10;
input 	result_imag_1_9;
input 	result_imag_1_8;
input 	result_imag_1_7;
input 	result_imag_1_6;
input 	result_imag_1_5;
input 	result_imag_1_4;
input 	result_imag_1_3;
input 	result_imag_1_2;
input 	result_imag_1_1;
input 	result_imag_1_0;
input 	result_imag_1_31;
input 	result_imag_1_17;
input 	result_imag_1_18;
input 	result_imag_1_19;
input 	result_imag_1_20;
input 	result_imag_1_21;
input 	result_imag_1_22;
input 	result_imag_1_23;
input 	result_imag_1_24;
input 	result_imag_1_25;
input 	result_imag_1_26;
input 	result_imag_1_27;
input 	result_imag_1_28;
input 	result_imag_1_29;
input 	result_imag_1_30;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_add_sub_knj_1 auto_generated(
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_31(pipeline_dffe_31),
	.result_imag_1_16(result_imag_1_16),
	.result_imag_1_15(result_imag_1_15),
	.result_imag_1_14(result_imag_1_14),
	.result_imag_1_13(result_imag_1_13),
	.result_imag_1_12(result_imag_1_12),
	.result_imag_1_11(result_imag_1_11),
	.result_imag_1_10(result_imag_1_10),
	.result_imag_1_9(result_imag_1_9),
	.result_imag_1_8(result_imag_1_8),
	.result_imag_1_7(result_imag_1_7),
	.result_imag_1_6(result_imag_1_6),
	.result_imag_1_5(result_imag_1_5),
	.result_imag_1_4(result_imag_1_4),
	.result_imag_1_3(result_imag_1_3),
	.result_imag_1_2(result_imag_1_2),
	.result_imag_1_1(result_imag_1_1),
	.result_imag_1_0(result_imag_1_0),
	.result_imag_1_31(result_imag_1_31),
	.result_imag_1_17(result_imag_1_17),
	.result_imag_1_18(result_imag_1_18),
	.result_imag_1_19(result_imag_1_19),
	.result_imag_1_20(result_imag_1_20),
	.result_imag_1_21(result_imag_1_21),
	.result_imag_1_22(result_imag_1_22),
	.result_imag_1_23(result_imag_1_23),
	.result_imag_1_24(result_imag_1_24),
	.result_imag_1_25(result_imag_1_25),
	.result_imag_1_26(result_imag_1_26),
	.result_imag_1_27(result_imag_1_27),
	.result_imag_1_28(result_imag_1_28),
	.result_imag_1_29(result_imag_1_29),
	.result_imag_1_30(result_imag_1_30),
	.clken(clken),
	.clock(clock));

endmodule

module fft256_add_sub_knj_1 (
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_31,
	result_imag_1_16,
	result_imag_1_15,
	result_imag_1_14,
	result_imag_1_13,
	result_imag_1_12,
	result_imag_1_11,
	result_imag_1_10,
	result_imag_1_9,
	result_imag_1_8,
	result_imag_1_7,
	result_imag_1_6,
	result_imag_1_5,
	result_imag_1_4,
	result_imag_1_3,
	result_imag_1_2,
	result_imag_1_1,
	result_imag_1_0,
	result_imag_1_31,
	result_imag_1_17,
	result_imag_1_18,
	result_imag_1_19,
	result_imag_1_20,
	result_imag_1_21,
	result_imag_1_22,
	result_imag_1_23,
	result_imag_1_24,
	result_imag_1_25,
	result_imag_1_26,
	result_imag_1_27,
	result_imag_1_28,
	result_imag_1_29,
	result_imag_1_30,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_31;
input 	result_imag_1_16;
input 	result_imag_1_15;
input 	result_imag_1_14;
input 	result_imag_1_13;
input 	result_imag_1_12;
input 	result_imag_1_11;
input 	result_imag_1_10;
input 	result_imag_1_9;
input 	result_imag_1_8;
input 	result_imag_1_7;
input 	result_imag_1_6;
input 	result_imag_1_5;
input 	result_imag_1_4;
input 	result_imag_1_3;
input 	result_imag_1_2;
input 	result_imag_1_1;
input 	result_imag_1_0;
input 	result_imag_1_31;
input 	result_imag_1_17;
input 	result_imag_1_18;
input 	result_imag_1_19;
input 	result_imag_1_20;
input 	result_imag_1_21;
input 	result_imag_1_22;
input 	result_imag_1_23;
input 	result_imag_1_24;
input 	result_imag_1_25;
input 	result_imag_1_26;
input 	result_imag_1_27;
input 	result_imag_1_28;
input 	result_imag_1_29;
input 	result_imag_1_30;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~17_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~19_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~21_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~23_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~25_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~27_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~29_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~31_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~33_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~35_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~37_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~39_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~41_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~43_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~47_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~49_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~51 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~53 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~54_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~55 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~56_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~57 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~58_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~59 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~60_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~61 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~62_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~63 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~64_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~65 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~66_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~67 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~68_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~69 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~70_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~71 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~72_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~73 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~74_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~75 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~76_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~77 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~78_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~79 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~80_combout ;


dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_18),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_19),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_20),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_21),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_22),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~64_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_23),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_24),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~68_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_25),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~70_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_26),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~72_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_27),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~74_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_28),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~76_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_29),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~78_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_30),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~80_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_31),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31] .power_up = "low";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~17 (
	.dataa(result_imag_1_31),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~17_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~17 .lut_mask = 16'h0055;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~19 (
	.dataa(result_imag_1_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~17_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~19_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~19 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~21 (
	.dataa(result_imag_1_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~19_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~21_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~21 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~23 (
	.dataa(result_imag_1_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~21_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~23_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~23 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~25 (
	.dataa(result_imag_1_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~23_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~25_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~25 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~27 (
	.dataa(result_imag_1_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~25_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~27_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~27 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~29 (
	.dataa(result_imag_1_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~27_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~29_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~29 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~31 (
	.dataa(result_imag_1_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~29_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~31_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~31 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~33 (
	.dataa(result_imag_1_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~31_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~33_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~33 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~33 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~35 (
	.dataa(result_imag_1_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~33_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~35_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~35 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~35 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~37 (
	.dataa(result_imag_1_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~35_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~37_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~37 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~37 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~39 (
	.dataa(result_imag_1_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~37_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~39_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~39 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~39 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~41 (
	.dataa(result_imag_1_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~39_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~41_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~41 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~41 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~43 (
	.dataa(result_imag_1_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~41_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~43_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~43 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~43 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 (
	.dataa(result_imag_1_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~43_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~47 (
	.dataa(result_imag_1_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~47_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~47 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~47 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~49 (
	.dataa(result_imag_1_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~47_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~49_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~49 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~49 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50 (
	.dataa(result_imag_1_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~49_cout ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~51 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52 (
	.dataa(result_imag_1_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~51 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~53 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~54 (
	.dataa(result_imag_1_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~53 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~54_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~55 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~54 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~54 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~56 (
	.dataa(result_imag_1_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~55 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~56_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~57 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~56 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~56 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~58 (
	.dataa(result_imag_1_20),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~57 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~58_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~59 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~58 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~58 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~60 (
	.dataa(result_imag_1_21),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[20]~59 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~60_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~61 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~60 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~60 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~62 (
	.dataa(result_imag_1_22),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[21]~61 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~62_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~63 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~62 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~62 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~64 (
	.dataa(result_imag_1_23),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[22]~63 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~64_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~65 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~64 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~64 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~66 (
	.dataa(result_imag_1_24),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[23]~65 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~66_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~67 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~66 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~66 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~68 (
	.dataa(result_imag_1_25),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[24]~67 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~68_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~69 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~68 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~68 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~70 (
	.dataa(result_imag_1_26),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[25]~69 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~70_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~71 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~70 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~70 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~72 (
	.dataa(result_imag_1_27),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[26]~71 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~72_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~73 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~72 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~72 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~74 (
	.dataa(result_imag_1_28),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[27]~73 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~74_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~75 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~74 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~74 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~76 (
	.dataa(result_imag_1_29),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[28]~75 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~76_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~77 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~76 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~76 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~78 (
	.dataa(result_imag_1_30),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[29]~77 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~78_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~79 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~78 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~78 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~80 (
	.dataa(result_imag_1_31),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[30]~79 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~80_combout ),
	.cout());
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~80 .lut_mask = 16'h5A5A;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_unsc:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[31]~80 .sum_lutc_input = "cin";

endmodule

module fft256_LPM_MULT_1 (
	dataa,
	datab,
	clken,
	dffe3a_16,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_31,
	dffe3a_30,
	dffe3a_29,
	dffe3a_28,
	dffe3a_27,
	dffe3a_26,
	dffe3a_25,
	dffe3a_24,
	dffe3a_23,
	dffe3a_22,
	dffe3a_21,
	dffe3a_20,
	dffe3a_19,
	dffe3a_18,
	dffe3a_17,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[16:0] dataa;
input 	[16:0] datab;
input 	clken;
output 	dffe3a_16;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_31;
output 	dffe3a_30;
output 	dffe3a_29;
output 	dffe3a_28;
output 	dffe3a_27;
output 	dffe3a_26;
output 	dffe3a_25;
output 	dffe3a_24;
output 	dffe3a_23;
output 	dffe3a_22;
output 	dffe3a_21;
output 	dffe3a_20;
output 	dffe3a_19;
output 	dffe3a_18;
output 	dffe3a_17;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_mult_9t01 auto_generated(
	.dataa({dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clken(clken),
	.dffe3a_16(dffe3a_16),
	.dffe3a_15(dffe3a_15),
	.dffe3a_14(dffe3a_14),
	.dffe3a_13(dffe3a_13),
	.dffe3a_12(dffe3a_12),
	.dffe3a_11(dffe3a_11),
	.dffe3a_10(dffe3a_10),
	.dffe3a_9(dffe3a_9),
	.dffe3a_8(dffe3a_8),
	.dffe3a_7(dffe3a_7),
	.dffe3a_6(dffe3a_6),
	.dffe3a_5(dffe3a_5),
	.dffe3a_4(dffe3a_4),
	.dffe3a_3(dffe3a_3),
	.dffe3a_2(dffe3a_2),
	.dffe3a_1(dffe3a_1),
	.dffe3a_0(dffe3a_0),
	.dffe3a_31(dffe3a_31),
	.dffe3a_30(dffe3a_30),
	.dffe3a_29(dffe3a_29),
	.dffe3a_28(dffe3a_28),
	.dffe3a_27(dffe3a_27),
	.dffe3a_26(dffe3a_26),
	.dffe3a_25(dffe3a_25),
	.dffe3a_24(dffe3a_24),
	.dffe3a_23(dffe3a_23),
	.dffe3a_22(dffe3a_22),
	.dffe3a_21(dffe3a_21),
	.dffe3a_20(dffe3a_20),
	.dffe3a_19(dffe3a_19),
	.dffe3a_18(dffe3a_18),
	.dffe3a_17(dffe3a_17),
	.clock(clock));

endmodule

module fft256_mult_9t01 (
	dataa,
	datab,
	clken,
	dffe3a_16,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_31,
	dffe3a_30,
	dffe3a_29,
	dffe3a_28,
	dffe3a_27,
	dffe3a_26,
	dffe3a_25,
	dffe3a_24,
	dffe3a_23,
	dffe3a_22,
	dffe3a_21,
	dffe3a_20,
	dffe3a_19,
	dffe3a_18,
	dffe3a_17,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[16:0] dataa;
input 	[16:0] datab;
input 	clken;
output 	dffe3a_16;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_31;
output 	dffe3a_30;
output 	dffe3a_29;
output 	dffe3a_28;
output 	dffe3a_27;
output 	dffe3a_26;
output 	dffe3a_25;
output 	dffe3a_24;
output 	dffe3a_23;
output 	dffe3a_22;
output 	dffe3a_21;
output 	dffe3a_20;
output 	dffe3a_19;
output 	dffe3a_18;
output 	dffe3a_17;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT32 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT33 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~dataout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT1 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT2 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT3 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT4 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT5 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT6 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT7 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT8 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT9 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT10 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT11 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT12 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT13 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT14 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT15 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT16 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT17 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT18 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT19 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT20 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT21 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT22 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT23 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT24 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT25 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT26 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT27 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT28 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT29 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT30 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT31 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT32 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT33 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT16 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT15 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT14 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT13 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT12 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT11 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT10 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT9 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT8 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT7 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT6 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT5 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT4 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT3 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT2 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT1 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~dataout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT31 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT30 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT29 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT28 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT27 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT26 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT25 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT24 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT23 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT22 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT21 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT20 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT19 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT18 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT17 ;

wire [35:0] \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus ;
wire [35:0] \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus ;

assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~dataout  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [0];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT1  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [1];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT2  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [2];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT3  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [3];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT4  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [4];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT5  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [5];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT6  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [6];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT7  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [7];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT8  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [8];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT9  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [9];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT10  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [10];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT11  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [11];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT12  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [12];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT13  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [13];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT14  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [14];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT15  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [15];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT16  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [16];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT17  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [17];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT18  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [18];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT19  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [19];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT20  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [20];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT21  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [21];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT22  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [22];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT23  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [23];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT24  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [24];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT25  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [25];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT26  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [26];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT27  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [27];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT28  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [28];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT29  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [29];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT30  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [30];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT31  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [31];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT32  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [32];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT33  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus [33];

assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~dataout  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [0];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT1  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [1];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT2  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [2];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT3  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [3];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT4  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [4];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT5  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [5];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT6  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [6];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT7  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [7];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT8  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [8];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT9  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [9];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT10  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [10];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT11  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [11];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT12  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [12];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT13  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [13];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT14  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [14];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT15  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [15];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT16  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [16];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT17  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [17];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT18  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [18];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT19  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [19];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT20  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [20];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT21  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [21];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT22  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [22];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT23  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [23];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT24  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [24];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT25  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [25];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT26  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [26];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT27  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [27];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT28  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [28];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT29  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [29];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT30  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [30];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT31  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [31];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT32  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [32];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT33  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus [33];

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[16] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT16 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_16),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[16] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[16] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[15] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT15 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_15),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[15] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[15] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[14] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT14 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_14),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[14] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[14] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[13] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT13 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_13),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[13] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[13] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[12] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT12 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_12),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[12] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[12] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[11] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT11 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_11),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[11] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[11] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[10] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT10 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_10),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[10] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[10] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[9] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT9 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_9),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[9] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[9] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[8] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT8 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_8),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[8] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[8] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[7] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT7 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_7),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[7] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[7] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[6] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT6 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_6),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[6] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[6] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[5] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT5 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_5),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[5] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[5] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[4] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT4 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_4),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[4] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[3] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT3 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_3),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[3] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[2] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT2 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_2),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[2] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[1] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT1 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_1),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[1] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[0] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~dataout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_0),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[0] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[31] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT31 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_31),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[31] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[31] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[30] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT30 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_30),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[30] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[30] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[29] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT29 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_29),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[29] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[29] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[28] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT28 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_28),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[28] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[28] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[27] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT27 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_27),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[27] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[27] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[26] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT26 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_26),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[26] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[26] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[25] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT25 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_25),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[25] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[25] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[24] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT24 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_24),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[24] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[24] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[23] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT23 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_23),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[23] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[23] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[22] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT22 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_22),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[22] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[22] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[21] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT21 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_21),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[21] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[21] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[20] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT20 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_20),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[20] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[20] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[19] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT19 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_19),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[19] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[19] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[18] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT18 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_18),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[18] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[18] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[17] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2~DATAOUT17 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_17),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[17] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|dffe3a[17] .power_up = "low";

cycloneive_mac_mult \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1 (
	.signa(vcc),
	.signb(vcc),
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1_DATAOUT_bus ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1 .dataa_clock = "0";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1 .dataa_width = 17;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1 .datab_clock = "0";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1 .datab_width = 17;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1 .signa_clock = "none";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1 .signb_clock = "none";

cycloneive_mac_out \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2 (
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT33 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT32 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT31 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT30 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT29 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT28 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT27 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT26 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT25 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT24 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT23 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT22 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT21 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT20 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT19 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT18 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT17 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT16 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT15 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT14 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT13 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT12 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT11 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT10 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT9 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT8 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT7 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT6 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT5 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT4 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT3 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT2 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~DATAOUT1 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_mult1~dataout }),
	.dataout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2_DATAOUT_bus ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2 .dataa_width = 34;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_a_b_c_d:m_a_b_c_d|auto_generated|mac_out2 .output_clock = "0";

endmodule

module fft256_LPM_MULT_2 (
	dataa,
	datab,
	clken,
	dffe3a_16,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_31,
	dffe3a_30,
	dffe3a_29,
	dffe3a_28,
	dffe3a_27,
	dffe3a_26,
	dffe3a_25,
	dffe3a_24,
	dffe3a_23,
	dffe3a_22,
	dffe3a_21,
	dffe3a_20,
	dffe3a_19,
	dffe3a_18,
	dffe3a_17,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[16:0] dataa;
input 	[16:0] datab;
input 	clken;
output 	dffe3a_16;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_31;
output 	dffe3a_30;
output 	dffe3a_29;
output 	dffe3a_28;
output 	dffe3a_27;
output 	dffe3a_26;
output 	dffe3a_25;
output 	dffe3a_24;
output 	dffe3a_23;
output 	dffe3a_22;
output 	dffe3a_21;
output 	dffe3a_20;
output 	dffe3a_19;
output 	dffe3a_18;
output 	dffe3a_17;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_mult_5t01 auto_generated(
	.dataa({dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clken(clken),
	.dffe3a_16(dffe3a_16),
	.dffe3a_15(dffe3a_15),
	.dffe3a_14(dffe3a_14),
	.dffe3a_13(dffe3a_13),
	.dffe3a_12(dffe3a_12),
	.dffe3a_11(dffe3a_11),
	.dffe3a_10(dffe3a_10),
	.dffe3a_9(dffe3a_9),
	.dffe3a_8(dffe3a_8),
	.dffe3a_7(dffe3a_7),
	.dffe3a_6(dffe3a_6),
	.dffe3a_5(dffe3a_5),
	.dffe3a_4(dffe3a_4),
	.dffe3a_3(dffe3a_3),
	.dffe3a_2(dffe3a_2),
	.dffe3a_1(dffe3a_1),
	.dffe3a_0(dffe3a_0),
	.dffe3a_31(dffe3a_31),
	.dffe3a_30(dffe3a_30),
	.dffe3a_29(dffe3a_29),
	.dffe3a_28(dffe3a_28),
	.dffe3a_27(dffe3a_27),
	.dffe3a_26(dffe3a_26),
	.dffe3a_25(dffe3a_25),
	.dffe3a_24(dffe3a_24),
	.dffe3a_23(dffe3a_23),
	.dffe3a_22(dffe3a_22),
	.dffe3a_21(dffe3a_21),
	.dffe3a_20(dffe3a_20),
	.dffe3a_19(dffe3a_19),
	.dffe3a_18(dffe3a_18),
	.dffe3a_17(dffe3a_17),
	.clock(clock));

endmodule

module fft256_mult_5t01 (
	dataa,
	datab,
	clken,
	dffe3a_16,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_31,
	dffe3a_30,
	dffe3a_29,
	dffe3a_28,
	dffe3a_27,
	dffe3a_26,
	dffe3a_25,
	dffe3a_24,
	dffe3a_23,
	dffe3a_22,
	dffe3a_21,
	dffe3a_20,
	dffe3a_19,
	dffe3a_18,
	dffe3a_17,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[15:0] dataa;
input 	[15:0] datab;
input 	clken;
output 	dffe3a_16;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_31;
output 	dffe3a_30;
output 	dffe3a_29;
output 	dffe3a_28;
output 	dffe3a_27;
output 	dffe3a_26;
output 	dffe3a_25;
output 	dffe3a_24;
output 	dffe3a_23;
output 	dffe3a_22;
output 	dffe3a_21;
output 	dffe3a_20;
output 	dffe3a_19;
output 	dffe3a_18;
output 	dffe3a_17;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~dataout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT1 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT2 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT3 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT4 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT5 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT6 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT7 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT8 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT9 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT10 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT11 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT12 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT13 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT14 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT15 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT16 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT17 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT18 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT19 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT20 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT21 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT22 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT23 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT24 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT25 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT26 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT27 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT28 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT29 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT30 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT31 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT16 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT15 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT14 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT13 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT12 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT11 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT10 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT9 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT8 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT7 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT6 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT5 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT4 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT3 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT2 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT1 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~dataout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT31 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT30 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT29 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT28 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT27 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT26 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT25 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT24 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT23 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT22 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT21 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT20 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT19 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT18 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT17 ;

wire [35:0] \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus ;
wire [35:0] \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus ;

assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~dataout  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [0];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT1  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [1];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT2  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [2];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT3  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [3];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT4  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [4];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT5  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [5];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT6  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [6];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT7  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [7];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT8  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [8];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT9  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [9];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT10  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [10];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT11  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [11];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT12  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [12];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT13  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [13];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT14  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [14];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT15  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [15];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT16  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [16];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT17  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [17];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT18  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [18];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT19  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [19];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT20  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [20];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT21  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [21];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT22  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [22];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT23  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [23];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT24  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [24];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT25  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [25];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT26  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [26];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT27  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [27];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT28  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [28];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT29  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [29];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT30  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [30];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT31  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus [31];

assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~dataout  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [0];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT1  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [1];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT2  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [2];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT3  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [3];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT4  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [4];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT5  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [5];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT6  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [6];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT7  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [7];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT8  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [8];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT9  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [9];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT10  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [10];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT11  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [11];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT12  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [12];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT13  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [13];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT14  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [14];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT15  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [15];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT16  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [16];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT17  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [17];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT18  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [18];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT19  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [19];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT20  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [20];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT21  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [21];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT22  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [22];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT23  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [23];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT24  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [24];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT25  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [25];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT26  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [26];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT27  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [27];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT28  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [28];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT29  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [29];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT30  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [30];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT31  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus [31];

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[16] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT16 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_16),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[16] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[16] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[15] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT15 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_15),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[15] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[15] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[14] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT14 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_14),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[14] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[14] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[13] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT13 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_13),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[13] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[13] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[12] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT12 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_12),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[12] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[12] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[11] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT11 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_11),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[11] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[11] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[10] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT10 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_10),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[10] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[10] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[9] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT9 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_9),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[9] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[9] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[8] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT8 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_8),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[8] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[8] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[7] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT7 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_7),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[7] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[7] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[6] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT6 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_6),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[6] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[6] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[5] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT5 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_5),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[5] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[5] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[4] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT4 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_4),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[4] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[3] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT3 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_3),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[3] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[2] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT2 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_2),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[2] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[1] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT1 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_1),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[1] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[0] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~dataout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_0),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[0] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[31] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT31 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_31),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[31] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[31] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[30] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT30 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_30),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[30] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[30] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[29] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT29 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_29),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[29] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[29] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[28] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT28 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_28),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[28] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[28] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[27] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT27 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_27),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[27] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[27] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[26] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT26 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_26),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[26] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[26] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[25] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT25 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_25),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[25] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[25] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[24] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT24 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_24),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[24] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[24] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[23] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT23 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_23),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[23] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[23] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[22] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT22 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_22),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[22] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[22] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[21] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT21 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_21),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[21] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[21] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[20] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT20 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_20),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[20] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[20] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[19] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT19 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_19),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[19] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[19] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[18] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT18 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_18),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[18] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[18] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[17] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2~DATAOUT17 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_17),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[17] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|dffe3a[17] .power_up = "low";

cycloneive_mac_mult \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1 (
	.signa(vcc),
	.signb(vcc),
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1_DATAOUT_bus ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1 .dataa_clock = "0";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1 .dataa_width = 16;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1 .datab_clock = "0";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1 .datab_width = 16;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1 .signa_clock = "none";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1 .signb_clock = "none";

cycloneive_mac_out \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2 (
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT31 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT30 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT29 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT28 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT27 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT26 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT25 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT24 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT23 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT22 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT21 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT20 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT19 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT18 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT17 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT16 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT15 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT14 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT13 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT12 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT11 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT10 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT9 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT8 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT7 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT6 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT5 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT4 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT3 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT2 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~DATAOUT1 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_mult1~dataout }),
	.dataout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2_DATAOUT_bus ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2 .dataa_width = 32;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_ac:m_ac|auto_generated|mac_out2 .output_clock = "0";

endmodule

module fft256_LPM_MULT_3 (
	dataa,
	datab,
	clken,
	dffe3a_16,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_31,
	dffe3a_30,
	dffe3a_29,
	dffe3a_28,
	dffe3a_27,
	dffe3a_26,
	dffe3a_25,
	dffe3a_24,
	dffe3a_23,
	dffe3a_22,
	dffe3a_21,
	dffe3a_20,
	dffe3a_19,
	dffe3a_18,
	dffe3a_17,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[16:0] dataa;
input 	[16:0] datab;
input 	clken;
output 	dffe3a_16;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_31;
output 	dffe3a_30;
output 	dffe3a_29;
output 	dffe3a_28;
output 	dffe3a_27;
output 	dffe3a_26;
output 	dffe3a_25;
output 	dffe3a_24;
output 	dffe3a_23;
output 	dffe3a_22;
output 	dffe3a_21;
output 	dffe3a_20;
output 	dffe3a_19;
output 	dffe3a_18;
output 	dffe3a_17;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_mult_5t01_1 auto_generated(
	.dataa({dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clken(clken),
	.dffe3a_16(dffe3a_16),
	.dffe3a_15(dffe3a_15),
	.dffe3a_14(dffe3a_14),
	.dffe3a_13(dffe3a_13),
	.dffe3a_12(dffe3a_12),
	.dffe3a_11(dffe3a_11),
	.dffe3a_10(dffe3a_10),
	.dffe3a_9(dffe3a_9),
	.dffe3a_8(dffe3a_8),
	.dffe3a_7(dffe3a_7),
	.dffe3a_6(dffe3a_6),
	.dffe3a_5(dffe3a_5),
	.dffe3a_4(dffe3a_4),
	.dffe3a_3(dffe3a_3),
	.dffe3a_2(dffe3a_2),
	.dffe3a_1(dffe3a_1),
	.dffe3a_0(dffe3a_0),
	.dffe3a_31(dffe3a_31),
	.dffe3a_30(dffe3a_30),
	.dffe3a_29(dffe3a_29),
	.dffe3a_28(dffe3a_28),
	.dffe3a_27(dffe3a_27),
	.dffe3a_26(dffe3a_26),
	.dffe3a_25(dffe3a_25),
	.dffe3a_24(dffe3a_24),
	.dffe3a_23(dffe3a_23),
	.dffe3a_22(dffe3a_22),
	.dffe3a_21(dffe3a_21),
	.dffe3a_20(dffe3a_20),
	.dffe3a_19(dffe3a_19),
	.dffe3a_18(dffe3a_18),
	.dffe3a_17(dffe3a_17),
	.clock(clock));

endmodule

module fft256_mult_5t01_1 (
	dataa,
	datab,
	clken,
	dffe3a_16,
	dffe3a_15,
	dffe3a_14,
	dffe3a_13,
	dffe3a_12,
	dffe3a_11,
	dffe3a_10,
	dffe3a_9,
	dffe3a_8,
	dffe3a_7,
	dffe3a_6,
	dffe3a_5,
	dffe3a_4,
	dffe3a_3,
	dffe3a_2,
	dffe3a_1,
	dffe3a_0,
	dffe3a_31,
	dffe3a_30,
	dffe3a_29,
	dffe3a_28,
	dffe3a_27,
	dffe3a_26,
	dffe3a_25,
	dffe3a_24,
	dffe3a_23,
	dffe3a_22,
	dffe3a_21,
	dffe3a_20,
	dffe3a_19,
	dffe3a_18,
	dffe3a_17,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[15:0] dataa;
input 	[15:0] datab;
input 	clken;
output 	dffe3a_16;
output 	dffe3a_15;
output 	dffe3a_14;
output 	dffe3a_13;
output 	dffe3a_12;
output 	dffe3a_11;
output 	dffe3a_10;
output 	dffe3a_9;
output 	dffe3a_8;
output 	dffe3a_7;
output 	dffe3a_6;
output 	dffe3a_5;
output 	dffe3a_4;
output 	dffe3a_3;
output 	dffe3a_2;
output 	dffe3a_1;
output 	dffe3a_0;
output 	dffe3a_31;
output 	dffe3a_30;
output 	dffe3a_29;
output 	dffe3a_28;
output 	dffe3a_27;
output 	dffe3a_26;
output 	dffe3a_25;
output 	dffe3a_24;
output 	dffe3a_23;
output 	dffe3a_22;
output 	dffe3a_21;
output 	dffe3a_20;
output 	dffe3a_19;
output 	dffe3a_18;
output 	dffe3a_17;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~dataout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT1 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT2 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT3 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT4 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT5 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT6 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT7 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT8 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT9 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT10 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT11 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT12 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT13 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT14 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT15 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT16 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT17 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT18 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT19 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT20 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT21 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT22 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT23 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT24 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT25 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT26 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT27 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT28 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT29 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT30 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT31 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT16 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT15 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT14 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT13 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT12 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT11 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT10 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT9 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT8 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT7 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT6 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT5 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT4 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT3 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT2 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT1 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~dataout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT31 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT30 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT29 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT28 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT27 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT26 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT25 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT24 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT23 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT22 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT21 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT20 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT19 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT18 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT17 ;

wire [35:0] \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus ;
wire [35:0] \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus ;

assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~dataout  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [0];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT1  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [1];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT2  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [2];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT3  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [3];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT4  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [4];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT5  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [5];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT6  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [6];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT7  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [7];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT8  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [8];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT9  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [9];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT10  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [10];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT11  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [11];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT12  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [12];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT13  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [13];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT14  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [14];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT15  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [15];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT16  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [16];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT17  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [17];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT18  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [18];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT19  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [19];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT20  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [20];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT21  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [21];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT22  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [22];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT23  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [23];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT24  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [24];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT25  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [25];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT26  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [26];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT27  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [27];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT28  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [28];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT29  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [29];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT30  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [30];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT31  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus [31];

assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~dataout  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [0];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT1  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [1];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT2  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [2];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT3  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [3];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT4  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [4];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT5  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [5];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT6  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [6];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT7  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [7];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT8  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [8];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT9  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [9];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT10  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [10];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT11  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [11];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT12  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [12];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT13  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [13];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT14  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [14];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT15  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [15];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT16  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [16];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT17  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [17];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT18  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [18];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT19  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [19];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT20  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [20];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT21  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [21];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT22  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [22];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT23  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [23];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT24  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [24];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT25  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [25];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT26  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [26];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT27  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [27];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT28  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [28];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT29  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [29];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT30  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [30];
assign \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT31  = \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus [31];

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[16] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT16 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_16),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[16] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[16] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[15] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT15 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_15),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[15] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[15] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[14] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT14 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_14),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[14] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[14] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[13] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT13 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_13),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[13] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[13] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[12] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT12 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_12),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[12] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[12] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[11] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT11 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_11),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[11] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[11] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[10] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT10 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_10),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[10] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[10] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[9] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT9 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_9),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[9] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[9] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[8] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT8 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_8),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[8] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[8] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[7] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT7 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_7),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[7] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[7] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[6] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT6 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_6),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[6] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[6] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[5] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT5 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_5),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[5] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[5] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[4] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT4 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_4),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[4] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[3] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT3 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_3),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[3] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[2] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT2 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_2),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[2] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[1] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT1 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_1),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[1] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[0] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~dataout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_0),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[0] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[31] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT31 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_31),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[31] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[31] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[30] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT30 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_30),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[30] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[30] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[29] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT29 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_29),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[29] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[29] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[28] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT28 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_28),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[28] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[28] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[27] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT27 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_27),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[27] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[27] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[26] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT26 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_26),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[26] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[26] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[25] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT25 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_25),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[25] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[25] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[24] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT24 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_24),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[24] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[24] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[23] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT23 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_23),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[23] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[23] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[22] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT22 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_22),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[22] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[22] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[21] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT21 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_21),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[21] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[21] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[20] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT20 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_20),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[20] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[20] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[19] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT19 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_19),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[19] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[19] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[18] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT18 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_18),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[18] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[18] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[17] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2~DATAOUT17 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe3a_17),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[17] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|dffe3a[17] .power_up = "low";

cycloneive_mac_mult \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1 (
	.signa(vcc),
	.signb(vcc),
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1_DATAOUT_bus ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1 .dataa_clock = "0";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1 .dataa_width = 16;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1 .datab_clock = "0";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1 .datab_width = 16;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1 .signa_clock = "none";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1 .signb_clock = "none";

cycloneive_mac_out \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2 (
	.clk(clock),
	.aclr(gnd),
	.ena(clken),
	.dataa({gnd,gnd,gnd,gnd,\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT31 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT30 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT29 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT28 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT27 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT26 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT25 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT24 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT23 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT22 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT21 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT20 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT19 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT18 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT17 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT16 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT15 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT14 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT13 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT12 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT11 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT10 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT9 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT8 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT7 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT6 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT5 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT4 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT3 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT2 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~DATAOUT1 ,
\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_mult1~dataout }),
	.dataout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2_DATAOUT_bus ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2 .dataa_width = 32;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_da0:gen_canonic:cm1|gen_ded_m1:gen_unext_m_bd:m_bd|auto_generated|mac_out2 .output_clock = "0";

endmodule

module fft256_asj_fft_pround_fft_121_2 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_16,
	pipeline_dffe_17,
	butterfly_st_real_2,
	butterfly_st_real_1,
	butterfly_st_real_0,
	butterfly_st_real_17,
	butterfly_st_real_3,
	butterfly_st_real_4,
	butterfly_st_real_5,
	butterfly_st_real_6,
	butterfly_st_real_7,
	butterfly_st_real_8,
	butterfly_st_real_9,
	butterfly_st_real_10,
	butterfly_st_real_11,
	butterfly_st_real_12,
	butterfly_st_real_13,
	butterfly_st_real_14,
	butterfly_st_real_15,
	butterfly_st_real_16,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
input 	butterfly_st_real_2;
input 	butterfly_st_real_1;
input 	butterfly_st_real_0;
input 	butterfly_st_real_17;
input 	butterfly_st_real_3;
input 	butterfly_st_real_4;
input 	butterfly_st_real_5;
input 	butterfly_st_real_6;
input 	butterfly_st_real_7;
input 	butterfly_st_real_8;
input 	butterfly_st_real_9;
input 	butterfly_st_real_10;
input 	butterfly_st_real_11;
input 	butterfly_st_real_12;
input 	butterfly_st_real_13;
input 	butterfly_st_real_14;
input 	butterfly_st_real_15;
input 	butterfly_st_real_16;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_LPM_ADD_SUB_3 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.butterfly_st_real_2(butterfly_st_real_2),
	.butterfly_st_real_1(butterfly_st_real_1),
	.butterfly_st_real_0(butterfly_st_real_0),
	.butterfly_st_real_17(butterfly_st_real_17),
	.butterfly_st_real_3(butterfly_st_real_3),
	.butterfly_st_real_4(butterfly_st_real_4),
	.butterfly_st_real_5(butterfly_st_real_5),
	.butterfly_st_real_6(butterfly_st_real_6),
	.butterfly_st_real_7(butterfly_st_real_7),
	.butterfly_st_real_8(butterfly_st_real_8),
	.butterfly_st_real_9(butterfly_st_real_9),
	.butterfly_st_real_10(butterfly_st_real_10),
	.butterfly_st_real_11(butterfly_st_real_11),
	.butterfly_st_real_12(butterfly_st_real_12),
	.butterfly_st_real_13(butterfly_st_real_13),
	.butterfly_st_real_14(butterfly_st_real_14),
	.butterfly_st_real_15(butterfly_st_real_15),
	.butterfly_st_real_16(butterfly_st_real_16),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft256_LPM_ADD_SUB_3 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_16,
	pipeline_dffe_17,
	butterfly_st_real_2,
	butterfly_st_real_1,
	butterfly_st_real_0,
	butterfly_st_real_17,
	butterfly_st_real_3,
	butterfly_st_real_4,
	butterfly_st_real_5,
	butterfly_st_real_6,
	butterfly_st_real_7,
	butterfly_st_real_8,
	butterfly_st_real_9,
	butterfly_st_real_10,
	butterfly_st_real_11,
	butterfly_st_real_12,
	butterfly_st_real_13,
	butterfly_st_real_14,
	butterfly_st_real_15,
	butterfly_st_real_16,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
input 	butterfly_st_real_2;
input 	butterfly_st_real_1;
input 	butterfly_st_real_0;
input 	butterfly_st_real_17;
input 	butterfly_st_real_3;
input 	butterfly_st_real_4;
input 	butterfly_st_real_5;
input 	butterfly_st_real_6;
input 	butterfly_st_real_7;
input 	butterfly_st_real_8;
input 	butterfly_st_real_9;
input 	butterfly_st_real_10;
input 	butterfly_st_real_11;
input 	butterfly_st_real_12;
input 	butterfly_st_real_13;
input 	butterfly_st_real_14;
input 	butterfly_st_real_15;
input 	butterfly_st_real_16;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_add_sub_onj auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.butterfly_st_real_2(butterfly_st_real_2),
	.butterfly_st_real_1(butterfly_st_real_1),
	.butterfly_st_real_0(butterfly_st_real_0),
	.butterfly_st_real_17(butterfly_st_real_17),
	.butterfly_st_real_3(butterfly_st_real_3),
	.butterfly_st_real_4(butterfly_st_real_4),
	.butterfly_st_real_5(butterfly_st_real_5),
	.butterfly_st_real_6(butterfly_st_real_6),
	.butterfly_st_real_7(butterfly_st_real_7),
	.butterfly_st_real_8(butterfly_st_real_8),
	.butterfly_st_real_9(butterfly_st_real_9),
	.butterfly_st_real_10(butterfly_st_real_10),
	.butterfly_st_real_11(butterfly_st_real_11),
	.butterfly_st_real_12(butterfly_st_real_12),
	.butterfly_st_real_13(butterfly_st_real_13),
	.butterfly_st_real_14(butterfly_st_real_14),
	.butterfly_st_real_15(butterfly_st_real_15),
	.butterfly_st_real_16(butterfly_st_real_16),
	.clken(clken),
	.clock(clock));

endmodule

module fft256_add_sub_onj (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_16,
	pipeline_dffe_17,
	butterfly_st_real_2,
	butterfly_st_real_1,
	butterfly_st_real_0,
	butterfly_st_real_17,
	butterfly_st_real_3,
	butterfly_st_real_4,
	butterfly_st_real_5,
	butterfly_st_real_6,
	butterfly_st_real_7,
	butterfly_st_real_8,
	butterfly_st_real_9,
	butterfly_st_real_10,
	butterfly_st_real_11,
	butterfly_st_real_12,
	butterfly_st_real_13,
	butterfly_st_real_14,
	butterfly_st_real_15,
	butterfly_st_real_16,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
input 	butterfly_st_real_2;
input 	butterfly_st_real_1;
input 	butterfly_st_real_0;
input 	butterfly_st_real_17;
input 	butterfly_st_real_3;
input 	butterfly_st_real_4;
input 	butterfly_st_real_5;
input 	butterfly_st_real_6;
input 	butterfly_st_real_7;
input 	butterfly_st_real_8;
input 	butterfly_st_real_9;
input 	butterfly_st_real_10;
input 	butterfly_st_real_11;
input 	butterfly_st_real_12;
input 	butterfly_st_real_13;
input 	butterfly_st_real_14;
input 	butterfly_st_real_15;
input 	butterfly_st_real_16;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~19_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~21_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~22_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~23 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~24_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~25 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~26_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~27 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~28_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~29 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~30_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~31 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~32_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~33 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~34_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~35 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~36_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~37 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~38_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~39 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~40_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~41 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~42_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~43 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~44_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~45 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~46_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~47 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~48_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~49 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~51 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52_combout ;


dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .power_up = "low";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 (
	.dataa(butterfly_st_real_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 .lut_mask = 16'h0055;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~19 (
	.dataa(butterfly_st_real_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~19_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~19 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~21 (
	.dataa(butterfly_st_real_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~19_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~21_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~21 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~22 (
	.dataa(butterfly_st_real_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~21_cout ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~22_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~23 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~22 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~24 (
	.dataa(butterfly_st_real_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~23 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~24_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~25 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~24 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~26 (
	.dataa(butterfly_st_real_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~25 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~26_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~27 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~26 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~28 (
	.dataa(butterfly_st_real_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~27 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~28_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~29 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~28 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~30 (
	.dataa(butterfly_st_real_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~29 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~30_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~31 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~30 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~32 (
	.dataa(butterfly_st_real_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~31 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~32_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~33 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~32 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~34 (
	.dataa(butterfly_st_real_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~33 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~34_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~35 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~34 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~36 (
	.dataa(butterfly_st_real_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~35 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~36_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~37 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~36 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~38 (
	.dataa(butterfly_st_real_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~37 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~38_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~39 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~38 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~40 (
	.dataa(butterfly_st_real_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~39 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~40_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~41 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~40 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~42 (
	.dataa(butterfly_st_real_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~41 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~42_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~43 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~42 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~44 (
	.dataa(butterfly_st_real_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~43 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~44_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~45 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~44 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~46 (
	.dataa(butterfly_st_real_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~45 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~46_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~47 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~46 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~48 (
	.dataa(butterfly_st_real_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~47 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~48_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~49 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~48 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50 (
	.dataa(butterfly_st_real_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~49 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~51 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52 (
	.dataa(butterfly_st_real_17),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~51 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52_combout ),
	.cout());
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52 .lut_mask = 16'h5A5A;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52 .sum_lutc_input = "cin";

endmodule

module fft256_asj_fft_pround_fft_121_3 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_16,
	pipeline_dffe_17,
	butterfly_st_imag_2,
	butterfly_st_imag_1,
	butterfly_st_imag_0,
	butterfly_st_imag_17,
	butterfly_st_imag_3,
	butterfly_st_imag_4,
	butterfly_st_imag_5,
	butterfly_st_imag_6,
	butterfly_st_imag_7,
	butterfly_st_imag_8,
	butterfly_st_imag_9,
	butterfly_st_imag_10,
	butterfly_st_imag_11,
	butterfly_st_imag_12,
	butterfly_st_imag_13,
	butterfly_st_imag_14,
	butterfly_st_imag_15,
	butterfly_st_imag_16,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
input 	butterfly_st_imag_2;
input 	butterfly_st_imag_1;
input 	butterfly_st_imag_0;
input 	butterfly_st_imag_17;
input 	butterfly_st_imag_3;
input 	butterfly_st_imag_4;
input 	butterfly_st_imag_5;
input 	butterfly_st_imag_6;
input 	butterfly_st_imag_7;
input 	butterfly_st_imag_8;
input 	butterfly_st_imag_9;
input 	butterfly_st_imag_10;
input 	butterfly_st_imag_11;
input 	butterfly_st_imag_12;
input 	butterfly_st_imag_13;
input 	butterfly_st_imag_14;
input 	butterfly_st_imag_15;
input 	butterfly_st_imag_16;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_LPM_ADD_SUB_4 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.butterfly_st_imag_2(butterfly_st_imag_2),
	.butterfly_st_imag_1(butterfly_st_imag_1),
	.butterfly_st_imag_0(butterfly_st_imag_0),
	.butterfly_st_imag_17(butterfly_st_imag_17),
	.butterfly_st_imag_3(butterfly_st_imag_3),
	.butterfly_st_imag_4(butterfly_st_imag_4),
	.butterfly_st_imag_5(butterfly_st_imag_5),
	.butterfly_st_imag_6(butterfly_st_imag_6),
	.butterfly_st_imag_7(butterfly_st_imag_7),
	.butterfly_st_imag_8(butterfly_st_imag_8),
	.butterfly_st_imag_9(butterfly_st_imag_9),
	.butterfly_st_imag_10(butterfly_st_imag_10),
	.butterfly_st_imag_11(butterfly_st_imag_11),
	.butterfly_st_imag_12(butterfly_st_imag_12),
	.butterfly_st_imag_13(butterfly_st_imag_13),
	.butterfly_st_imag_14(butterfly_st_imag_14),
	.butterfly_st_imag_15(butterfly_st_imag_15),
	.butterfly_st_imag_16(butterfly_st_imag_16),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fft256_LPM_ADD_SUB_4 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_16,
	pipeline_dffe_17,
	butterfly_st_imag_2,
	butterfly_st_imag_1,
	butterfly_st_imag_0,
	butterfly_st_imag_17,
	butterfly_st_imag_3,
	butterfly_st_imag_4,
	butterfly_st_imag_5,
	butterfly_st_imag_6,
	butterfly_st_imag_7,
	butterfly_st_imag_8,
	butterfly_st_imag_9,
	butterfly_st_imag_10,
	butterfly_st_imag_11,
	butterfly_st_imag_12,
	butterfly_st_imag_13,
	butterfly_st_imag_14,
	butterfly_st_imag_15,
	butterfly_st_imag_16,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
input 	butterfly_st_imag_2;
input 	butterfly_st_imag_1;
input 	butterfly_st_imag_0;
input 	butterfly_st_imag_17;
input 	butterfly_st_imag_3;
input 	butterfly_st_imag_4;
input 	butterfly_st_imag_5;
input 	butterfly_st_imag_6;
input 	butterfly_st_imag_7;
input 	butterfly_st_imag_8;
input 	butterfly_st_imag_9;
input 	butterfly_st_imag_10;
input 	butterfly_st_imag_11;
input 	butterfly_st_imag_12;
input 	butterfly_st_imag_13;
input 	butterfly_st_imag_14;
input 	butterfly_st_imag_15;
input 	butterfly_st_imag_16;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_add_sub_onj_1 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.butterfly_st_imag_2(butterfly_st_imag_2),
	.butterfly_st_imag_1(butterfly_st_imag_1),
	.butterfly_st_imag_0(butterfly_st_imag_0),
	.butterfly_st_imag_17(butterfly_st_imag_17),
	.butterfly_st_imag_3(butterfly_st_imag_3),
	.butterfly_st_imag_4(butterfly_st_imag_4),
	.butterfly_st_imag_5(butterfly_st_imag_5),
	.butterfly_st_imag_6(butterfly_st_imag_6),
	.butterfly_st_imag_7(butterfly_st_imag_7),
	.butterfly_st_imag_8(butterfly_st_imag_8),
	.butterfly_st_imag_9(butterfly_st_imag_9),
	.butterfly_st_imag_10(butterfly_st_imag_10),
	.butterfly_st_imag_11(butterfly_st_imag_11),
	.butterfly_st_imag_12(butterfly_st_imag_12),
	.butterfly_st_imag_13(butterfly_st_imag_13),
	.butterfly_st_imag_14(butterfly_st_imag_14),
	.butterfly_st_imag_15(butterfly_st_imag_15),
	.butterfly_st_imag_16(butterfly_st_imag_16),
	.clken(clken),
	.clock(clock));

endmodule

module fft256_add_sub_onj_1 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_16,
	pipeline_dffe_17,
	butterfly_st_imag_2,
	butterfly_st_imag_1,
	butterfly_st_imag_0,
	butterfly_st_imag_17,
	butterfly_st_imag_3,
	butterfly_st_imag_4,
	butterfly_st_imag_5,
	butterfly_st_imag_6,
	butterfly_st_imag_7,
	butterfly_st_imag_8,
	butterfly_st_imag_9,
	butterfly_st_imag_10,
	butterfly_st_imag_11,
	butterfly_st_imag_12,
	butterfly_st_imag_13,
	butterfly_st_imag_14,
	butterfly_st_imag_15,
	butterfly_st_imag_16,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
input 	butterfly_st_imag_2;
input 	butterfly_st_imag_1;
input 	butterfly_st_imag_0;
input 	butterfly_st_imag_17;
input 	butterfly_st_imag_3;
input 	butterfly_st_imag_4;
input 	butterfly_st_imag_5;
input 	butterfly_st_imag_6;
input 	butterfly_st_imag_7;
input 	butterfly_st_imag_8;
input 	butterfly_st_imag_9;
input 	butterfly_st_imag_10;
input 	butterfly_st_imag_11;
input 	butterfly_st_imag_12;
input 	butterfly_st_imag_13;
input 	butterfly_st_imag_14;
input 	butterfly_st_imag_15;
input 	butterfly_st_imag_16;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~19_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~21_cout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~22_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~23 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~24_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~25 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~26_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~27 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~28_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~29 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~30_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~31 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~32_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~33 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~34_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~35 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~36_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~37 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~38_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~39 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~40_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~41 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~42_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~43 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~44_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~45 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~46_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~47 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~48_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~49 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50_combout ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~51 ;
wire \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52_combout ;


dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .power_up = "low";

dffeas \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] (
	.clk(clock),
	.d(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .is_wysiwyg = "true";
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .power_up = "low";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 (
	.dataa(butterfly_st_imag_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 .lut_mask = 16'h0055;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~19 (
	.dataa(butterfly_st_imag_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~19_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~19 .lut_mask = 16'h005F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~21 (
	.dataa(butterfly_st_imag_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~19_cout ),
	.combout(),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~21_cout ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~21 .lut_mask = 16'h00AF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~22 (
	.dataa(butterfly_st_imag_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~21_cout ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~22_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~23 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~22 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~24 (
	.dataa(butterfly_st_imag_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~23 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~24_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~25 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~24 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~26 (
	.dataa(butterfly_st_imag_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~25 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~26_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~27 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~26 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~28 (
	.dataa(butterfly_st_imag_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~27 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~28_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~29 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~28 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~30 (
	.dataa(butterfly_st_imag_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~29 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~30_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~31 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~30 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~32 (
	.dataa(butterfly_st_imag_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~31 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~32_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~33 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~32 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~34 (
	.dataa(butterfly_st_imag_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~33 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~34_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~35 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~34 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~36 (
	.dataa(butterfly_st_imag_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~35 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~36_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~37 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~36 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~38 (
	.dataa(butterfly_st_imag_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~37 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~38_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~39 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~38 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~40 (
	.dataa(butterfly_st_imag_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~39 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~40_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~41 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~40 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~42 (
	.dataa(butterfly_st_imag_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~41 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~42_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~43 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~42 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~44 (
	.dataa(butterfly_st_imag_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~43 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~44_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~45 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~44 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~46 (
	.dataa(butterfly_st_imag_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~45 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~46_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~47 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~46 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~48 (
	.dataa(butterfly_st_imag_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~47 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~48_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~49 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~48 .lut_mask = 16'h5AAF;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50 (
	.dataa(butterfly_st_imag_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~49 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50_combout ),
	.cout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~51 ));
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50 .lut_mask = 16'h5A5F;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52 (
	.dataa(butterfly_st_imag_17),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~51 ),
	.combout(\asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52_combout ),
	.cout());
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52 .lut_mask = 16'h5A5A;
defparam \asj_fft_si_sose_so_b_fft_121_inst|gen_se:bfpdft|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~52 .sum_lutc_input = "cin";

endmodule

module fft256_asj_fft_in_write_sgl_fft_121 (
	disable_wr1,
	rdy_for_next_block1,
	core_imag_in_0,
	core_real_in_0,
	core_imag_in_1,
	core_real_in_1,
	core_imag_in_2,
	core_real_in_2,
	core_imag_in_3,
	core_real_in_3,
	core_imag_in_4,
	core_real_in_4,
	core_imag_in_5,
	core_real_in_5,
	core_imag_in_6,
	core_real_in_6,
	core_imag_in_7,
	core_real_in_7,
	core_imag_in_8,
	core_real_in_8,
	core_imag_in_9,
	core_real_in_9,
	core_imag_in_10,
	core_real_in_10,
	core_imag_in_11,
	core_real_in_11,
	core_imag_in_12,
	core_real_in_12,
	core_imag_in_13,
	core_real_in_13,
	core_imag_in_14,
	core_real_in_14,
	core_imag_in_15,
	core_real_in_15,
	data_rdy_int1,
	send_sop_s,
	global_clock_enable,
	blk_done,
	tdl_arr_0,
	data_in_i_0,
	wr_address_i_int_0,
	wr_address_i_int_1,
	wr_address_i_int_2,
	wr_address_i_int_3,
	wr_address_i_int_4,
	wr_address_i_int_5,
	wr_address_i_int_6,
	wr_address_i_int_7,
	data_in_r_0,
	data_in_i_1,
	data_in_r_1,
	data_in_i_2,
	data_in_r_2,
	data_in_i_3,
	data_in_r_3,
	data_in_i_4,
	data_in_r_4,
	data_in_i_5,
	data_in_r_5,
	data_in_i_6,
	data_in_r_6,
	data_in_i_7,
	data_in_r_7,
	data_in_i_8,
	data_in_r_8,
	data_in_i_9,
	data_in_r_9,
	data_in_i_10,
	data_in_r_10,
	data_in_i_11,
	data_in_r_11,
	data_in_i_12,
	data_in_r_12,
	data_in_i_13,
	data_in_r_13,
	data_in_i_14,
	data_in_r_14,
	data_in_i_15,
	data_in_r_15,
	counter_i,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	disable_wr1;
output 	rdy_for_next_block1;
input 	core_imag_in_0;
input 	core_real_in_0;
input 	core_imag_in_1;
input 	core_real_in_1;
input 	core_imag_in_2;
input 	core_real_in_2;
input 	core_imag_in_3;
input 	core_real_in_3;
input 	core_imag_in_4;
input 	core_real_in_4;
input 	core_imag_in_5;
input 	core_real_in_5;
input 	core_imag_in_6;
input 	core_real_in_6;
input 	core_imag_in_7;
input 	core_real_in_7;
input 	core_imag_in_8;
input 	core_real_in_8;
input 	core_imag_in_9;
input 	core_real_in_9;
input 	core_imag_in_10;
input 	core_real_in_10;
input 	core_imag_in_11;
input 	core_real_in_11;
input 	core_imag_in_12;
input 	core_real_in_12;
input 	core_imag_in_13;
input 	core_real_in_13;
input 	core_imag_in_14;
input 	core_real_in_14;
input 	core_imag_in_15;
input 	core_real_in_15;
output 	data_rdy_int1;
input 	send_sop_s;
input 	global_clock_enable;
input 	blk_done;
output 	tdl_arr_0;
output 	data_in_i_0;
output 	wr_address_i_int_0;
output 	wr_address_i_int_1;
output 	wr_address_i_int_2;
output 	wr_address_i_int_3;
output 	wr_address_i_int_4;
output 	wr_address_i_int_5;
output 	wr_address_i_int_6;
output 	wr_address_i_int_7;
output 	data_in_r_0;
output 	data_in_i_1;
output 	data_in_r_1;
output 	data_in_i_2;
output 	data_in_r_2;
output 	data_in_i_3;
output 	data_in_r_3;
output 	data_in_i_4;
output 	data_in_r_4;
output 	data_in_i_5;
output 	data_in_r_5;
output 	data_in_i_6;
output 	data_in_r_6;
output 	data_in_i_7;
output 	data_in_r_7;
output 	data_in_i_8;
output 	data_in_r_8;
output 	data_in_i_9;
output 	data_in_r_9;
output 	data_in_i_10;
output 	data_in_r_10;
output 	data_in_i_11;
output 	data_in_r_11;
output 	data_in_i_12;
output 	data_in_r_12;
output 	data_in_i_13;
output 	data_in_r_13;
output 	data_in_i_14;
output 	data_in_r_14;
output 	data_in_i_15;
output 	data_in_r_15;
output 	counter_i;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal0~0_combout ;
wire \so_count[0]~9 ;
wire \so_count[1]~12 ;
wire \so_count[2]~14 ;
wire \so_count[3]~16 ;
wire \so_count[4]~18 ;
wire \so_count[5]~19_combout ;
wire \burst_count_en~0_combout ;
wire \burst_count_en~q ;
wire \so_count[0]~10_combout ;
wire \so_count[5]~q ;
wire \so_count[5]~20 ;
wire \so_count[6]~21_combout ;
wire \so_count[6]~q ;
wire \so_count[6]~22 ;
wire \so_count[7]~23_combout ;
wire \so_count[7]~q ;
wire \Equal0~1_combout ;
wire \so_count[2]~13_combout ;
wire \so_count[2]~q ;
wire \Equal1~0_combout ;
wire \Equal0~2_combout ;
wire \data_rdy_int~0_combout ;
wire \data_in_i~0_combout ;
wire \so_count[0]~8_combout ;
wire \so_count[0]~q ;
wire \wr_address_i_early~0_combout ;
wire \wr_address_i_early[0]~q ;
wire \wr_address_i_int~0_combout ;
wire \so_count[1]~11_combout ;
wire \so_count[1]~q ;
wire \wr_address_i_early~1_combout ;
wire \wr_address_i_early[1]~q ;
wire \wr_address_i_int~1_combout ;
wire \wr_address_i_early~2_combout ;
wire \wr_address_i_early[2]~q ;
wire \wr_address_i_int~2_combout ;
wire \so_count[3]~15_combout ;
wire \so_count[3]~q ;
wire \wr_address_i_early~3_combout ;
wire \wr_address_i_early[3]~q ;
wire \wr_address_i_int~3_combout ;
wire \so_count[4]~17_combout ;
wire \so_count[4]~q ;
wire \wr_address_i_early~4_combout ;
wire \wr_address_i_early[4]~q ;
wire \wr_address_i_int~4_combout ;
wire \wr_address_i_early~5_combout ;
wire \wr_address_i_early[5]~q ;
wire \wr_address_i_int~5_combout ;
wire \wr_address_i_early~6_combout ;
wire \wr_address_i_early[6]~q ;
wire \wr_address_i_int~6_combout ;
wire \wr_address_i_early~7_combout ;
wire \wr_address_i_early[7]~q ;
wire \wr_address_i_int~7_combout ;
wire \data_in_r~0_combout ;
wire \data_in_i~1_combout ;
wire \data_in_r~1_combout ;
wire \data_in_i~2_combout ;
wire \data_in_r~2_combout ;
wire \data_in_i~3_combout ;
wire \data_in_r~3_combout ;
wire \data_in_i~4_combout ;
wire \data_in_r~4_combout ;
wire \data_in_i~5_combout ;
wire \data_in_r~5_combout ;
wire \data_in_i~6_combout ;
wire \data_in_r~6_combout ;
wire \data_in_i~7_combout ;
wire \data_in_r~7_combout ;
wire \data_in_i~8_combout ;
wire \data_in_r~8_combout ;
wire \data_in_i~9_combout ;
wire \data_in_r~9_combout ;
wire \data_in_i~10_combout ;
wire \data_in_r~10_combout ;
wire \data_in_i~11_combout ;
wire \data_in_r~11_combout ;
wire \data_in_i~12_combout ;
wire \data_in_r~12_combout ;
wire \data_in_i~13_combout ;
wire \data_in_r~13_combout ;
wire \data_in_i~14_combout ;
wire \data_in_r~14_combout ;
wire \data_in_i~15_combout ;
wire \data_in_r~15_combout ;


fft256_asj_fft_tdl_bit_rst_fft_121_1 \gen_soe:delay_swd (
	.global_clock_enable(global_clock_enable),
	.tdl_arr_0(tdl_arr_0),
	.clk(clk),
	.reset_n(reset_n));

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\so_count[0]~q ),
	.datab(\so_count[1]~q ),
	.datac(\so_count[3]~q ),
	.datad(\so_count[4]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hFFFE;
defparam \Equal0~0 .sum_lutc_input = "datac";

dffeas disable_wr(
	.clk(clk),
	.d(\Equal1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(disable_wr1),
	.prn(vcc));
defparam disable_wr.is_wysiwyg = "true";
defparam disable_wr.power_up = "low";

dffeas rdy_for_next_block(
	.clk(clk),
	.d(\Equal0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdy_for_next_block1),
	.prn(vcc));
defparam rdy_for_next_block.is_wysiwyg = "true";
defparam rdy_for_next_block.power_up = "low";

dffeas data_rdy_int(
	.clk(clk),
	.d(\data_rdy_int~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_rdy_int1),
	.prn(vcc));
defparam data_rdy_int.is_wysiwyg = "true";
defparam data_rdy_int.power_up = "low";

dffeas \data_in_i[0] (
	.clk(clk),
	.d(\data_in_i~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_0),
	.prn(vcc));
defparam \data_in_i[0] .is_wysiwyg = "true";
defparam \data_in_i[0] .power_up = "low";

dffeas \wr_address_i_int[0] (
	.clk(clk),
	.d(\wr_address_i_int~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_0),
	.prn(vcc));
defparam \wr_address_i_int[0] .is_wysiwyg = "true";
defparam \wr_address_i_int[0] .power_up = "low";

dffeas \wr_address_i_int[1] (
	.clk(clk),
	.d(\wr_address_i_int~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_1),
	.prn(vcc));
defparam \wr_address_i_int[1] .is_wysiwyg = "true";
defparam \wr_address_i_int[1] .power_up = "low";

dffeas \wr_address_i_int[2] (
	.clk(clk),
	.d(\wr_address_i_int~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_2),
	.prn(vcc));
defparam \wr_address_i_int[2] .is_wysiwyg = "true";
defparam \wr_address_i_int[2] .power_up = "low";

dffeas \wr_address_i_int[3] (
	.clk(clk),
	.d(\wr_address_i_int~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_3),
	.prn(vcc));
defparam \wr_address_i_int[3] .is_wysiwyg = "true";
defparam \wr_address_i_int[3] .power_up = "low";

dffeas \wr_address_i_int[4] (
	.clk(clk),
	.d(\wr_address_i_int~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_4),
	.prn(vcc));
defparam \wr_address_i_int[4] .is_wysiwyg = "true";
defparam \wr_address_i_int[4] .power_up = "low";

dffeas \wr_address_i_int[5] (
	.clk(clk),
	.d(\wr_address_i_int~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_5),
	.prn(vcc));
defparam \wr_address_i_int[5] .is_wysiwyg = "true";
defparam \wr_address_i_int[5] .power_up = "low";

dffeas \wr_address_i_int[6] (
	.clk(clk),
	.d(\wr_address_i_int~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_6),
	.prn(vcc));
defparam \wr_address_i_int[6] .is_wysiwyg = "true";
defparam \wr_address_i_int[6] .power_up = "low";

dffeas \wr_address_i_int[7] (
	.clk(clk),
	.d(\wr_address_i_int~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_7),
	.prn(vcc));
defparam \wr_address_i_int[7] .is_wysiwyg = "true";
defparam \wr_address_i_int[7] .power_up = "low";

dffeas \data_in_r[0] (
	.clk(clk),
	.d(\data_in_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_0),
	.prn(vcc));
defparam \data_in_r[0] .is_wysiwyg = "true";
defparam \data_in_r[0] .power_up = "low";

dffeas \data_in_i[1] (
	.clk(clk),
	.d(\data_in_i~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_1),
	.prn(vcc));
defparam \data_in_i[1] .is_wysiwyg = "true";
defparam \data_in_i[1] .power_up = "low";

dffeas \data_in_r[1] (
	.clk(clk),
	.d(\data_in_r~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_1),
	.prn(vcc));
defparam \data_in_r[1] .is_wysiwyg = "true";
defparam \data_in_r[1] .power_up = "low";

dffeas \data_in_i[2] (
	.clk(clk),
	.d(\data_in_i~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_2),
	.prn(vcc));
defparam \data_in_i[2] .is_wysiwyg = "true";
defparam \data_in_i[2] .power_up = "low";

dffeas \data_in_r[2] (
	.clk(clk),
	.d(\data_in_r~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_2),
	.prn(vcc));
defparam \data_in_r[2] .is_wysiwyg = "true";
defparam \data_in_r[2] .power_up = "low";

dffeas \data_in_i[3] (
	.clk(clk),
	.d(\data_in_i~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_3),
	.prn(vcc));
defparam \data_in_i[3] .is_wysiwyg = "true";
defparam \data_in_i[3] .power_up = "low";

dffeas \data_in_r[3] (
	.clk(clk),
	.d(\data_in_r~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_3),
	.prn(vcc));
defparam \data_in_r[3] .is_wysiwyg = "true";
defparam \data_in_r[3] .power_up = "low";

dffeas \data_in_i[4] (
	.clk(clk),
	.d(\data_in_i~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_4),
	.prn(vcc));
defparam \data_in_i[4] .is_wysiwyg = "true";
defparam \data_in_i[4] .power_up = "low";

dffeas \data_in_r[4] (
	.clk(clk),
	.d(\data_in_r~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_4),
	.prn(vcc));
defparam \data_in_r[4] .is_wysiwyg = "true";
defparam \data_in_r[4] .power_up = "low";

dffeas \data_in_i[5] (
	.clk(clk),
	.d(\data_in_i~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_5),
	.prn(vcc));
defparam \data_in_i[5] .is_wysiwyg = "true";
defparam \data_in_i[5] .power_up = "low";

dffeas \data_in_r[5] (
	.clk(clk),
	.d(\data_in_r~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_5),
	.prn(vcc));
defparam \data_in_r[5] .is_wysiwyg = "true";
defparam \data_in_r[5] .power_up = "low";

dffeas \data_in_i[6] (
	.clk(clk),
	.d(\data_in_i~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_6),
	.prn(vcc));
defparam \data_in_i[6] .is_wysiwyg = "true";
defparam \data_in_i[6] .power_up = "low";

dffeas \data_in_r[6] (
	.clk(clk),
	.d(\data_in_r~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_6),
	.prn(vcc));
defparam \data_in_r[6] .is_wysiwyg = "true";
defparam \data_in_r[6] .power_up = "low";

dffeas \data_in_i[7] (
	.clk(clk),
	.d(\data_in_i~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_7),
	.prn(vcc));
defparam \data_in_i[7] .is_wysiwyg = "true";
defparam \data_in_i[7] .power_up = "low";

dffeas \data_in_r[7] (
	.clk(clk),
	.d(\data_in_r~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_7),
	.prn(vcc));
defparam \data_in_r[7] .is_wysiwyg = "true";
defparam \data_in_r[7] .power_up = "low";

dffeas \data_in_i[8] (
	.clk(clk),
	.d(\data_in_i~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_8),
	.prn(vcc));
defparam \data_in_i[8] .is_wysiwyg = "true";
defparam \data_in_i[8] .power_up = "low";

dffeas \data_in_r[8] (
	.clk(clk),
	.d(\data_in_r~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_8),
	.prn(vcc));
defparam \data_in_r[8] .is_wysiwyg = "true";
defparam \data_in_r[8] .power_up = "low";

dffeas \data_in_i[9] (
	.clk(clk),
	.d(\data_in_i~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_9),
	.prn(vcc));
defparam \data_in_i[9] .is_wysiwyg = "true";
defparam \data_in_i[9] .power_up = "low";

dffeas \data_in_r[9] (
	.clk(clk),
	.d(\data_in_r~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_9),
	.prn(vcc));
defparam \data_in_r[9] .is_wysiwyg = "true";
defparam \data_in_r[9] .power_up = "low";

dffeas \data_in_i[10] (
	.clk(clk),
	.d(\data_in_i~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_10),
	.prn(vcc));
defparam \data_in_i[10] .is_wysiwyg = "true";
defparam \data_in_i[10] .power_up = "low";

dffeas \data_in_r[10] (
	.clk(clk),
	.d(\data_in_r~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_10),
	.prn(vcc));
defparam \data_in_r[10] .is_wysiwyg = "true";
defparam \data_in_r[10] .power_up = "low";

dffeas \data_in_i[11] (
	.clk(clk),
	.d(\data_in_i~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_11),
	.prn(vcc));
defparam \data_in_i[11] .is_wysiwyg = "true";
defparam \data_in_i[11] .power_up = "low";

dffeas \data_in_r[11] (
	.clk(clk),
	.d(\data_in_r~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_11),
	.prn(vcc));
defparam \data_in_r[11] .is_wysiwyg = "true";
defparam \data_in_r[11] .power_up = "low";

dffeas \data_in_i[12] (
	.clk(clk),
	.d(\data_in_i~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_12),
	.prn(vcc));
defparam \data_in_i[12] .is_wysiwyg = "true";
defparam \data_in_i[12] .power_up = "low";

dffeas \data_in_r[12] (
	.clk(clk),
	.d(\data_in_r~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_12),
	.prn(vcc));
defparam \data_in_r[12] .is_wysiwyg = "true";
defparam \data_in_r[12] .power_up = "low";

dffeas \data_in_i[13] (
	.clk(clk),
	.d(\data_in_i~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_13),
	.prn(vcc));
defparam \data_in_i[13] .is_wysiwyg = "true";
defparam \data_in_i[13] .power_up = "low";

dffeas \data_in_r[13] (
	.clk(clk),
	.d(\data_in_r~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_13),
	.prn(vcc));
defparam \data_in_r[13] .is_wysiwyg = "true";
defparam \data_in_r[13] .power_up = "low";

dffeas \data_in_i[14] (
	.clk(clk),
	.d(\data_in_i~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_14),
	.prn(vcc));
defparam \data_in_i[14] .is_wysiwyg = "true";
defparam \data_in_i[14] .power_up = "low";

dffeas \data_in_r[14] (
	.clk(clk),
	.d(\data_in_r~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_14),
	.prn(vcc));
defparam \data_in_r[14] .is_wysiwyg = "true";
defparam \data_in_r[14] .power_up = "low";

dffeas \data_in_i[15] (
	.clk(clk),
	.d(\data_in_i~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_15),
	.prn(vcc));
defparam \data_in_i[15] .is_wysiwyg = "true";
defparam \data_in_i[15] .power_up = "low";

dffeas \data_in_r[15] (
	.clk(clk),
	.d(\data_in_r~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_15),
	.prn(vcc));
defparam \data_in_r[15] .is_wysiwyg = "true";
defparam \data_in_r[15] .power_up = "low";

cycloneive_lcell_comb \counter_i~0 (
	.dataa(send_sop_s),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(counter_i),
	.cout());
defparam \counter_i~0 .lut_mask = 16'hAAFF;
defparam \counter_i~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \so_count[0]~8 (
	.dataa(\so_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\so_count[0]~8_combout ),
	.cout(\so_count[0]~9 ));
defparam \so_count[0]~8 .lut_mask = 16'h55AA;
defparam \so_count[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \so_count[1]~11 (
	.dataa(\so_count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\so_count[0]~9 ),
	.combout(\so_count[1]~11_combout ),
	.cout(\so_count[1]~12 ));
defparam \so_count[1]~11 .lut_mask = 16'h5A5F;
defparam \so_count[1]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \so_count[2]~13 (
	.dataa(\so_count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\so_count[1]~12 ),
	.combout(\so_count[2]~13_combout ),
	.cout(\so_count[2]~14 ));
defparam \so_count[2]~13 .lut_mask = 16'h5AAF;
defparam \so_count[2]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \so_count[3]~15 (
	.dataa(\so_count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\so_count[2]~14 ),
	.combout(\so_count[3]~15_combout ),
	.cout(\so_count[3]~16 ));
defparam \so_count[3]~15 .lut_mask = 16'h5A5F;
defparam \so_count[3]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \so_count[4]~17 (
	.dataa(\so_count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\so_count[3]~16 ),
	.combout(\so_count[4]~17_combout ),
	.cout(\so_count[4]~18 ));
defparam \so_count[4]~17 .lut_mask = 16'h5AAF;
defparam \so_count[4]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \so_count[5]~19 (
	.dataa(\so_count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\so_count[4]~18 ),
	.combout(\so_count[5]~19_combout ),
	.cout(\so_count[5]~20 ));
defparam \so_count[5]~19 .lut_mask = 16'h5A5F;
defparam \so_count[5]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \burst_count_en~0 (
	.dataa(send_sop_s),
	.datab(\burst_count_en~q ),
	.datac(gnd),
	.datad(rdy_for_next_block1),
	.cin(gnd),
	.combout(\burst_count_en~0_combout ),
	.cout());
defparam \burst_count_en~0 .lut_mask = 16'hEEFF;
defparam \burst_count_en~0 .sum_lutc_input = "datac";

dffeas burst_count_en(
	.clk(clk),
	.d(\burst_count_en~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\burst_count_en~q ),
	.prn(vcc));
defparam burst_count_en.is_wysiwyg = "true";
defparam burst_count_en.power_up = "low";

cycloneive_lcell_comb \so_count[0]~10 (
	.dataa(global_clock_enable),
	.datab(tdl_arr_0),
	.datac(\burst_count_en~q ),
	.datad(counter_i),
	.cin(gnd),
	.combout(\so_count[0]~10_combout ),
	.cout());
defparam \so_count[0]~10 .lut_mask = 16'hFFFE;
defparam \so_count[0]~10 .sum_lutc_input = "datac";

dffeas \so_count[5] (
	.clk(clk),
	.d(\so_count[5]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(counter_i),
	.sload(gnd),
	.ena(\so_count[0]~10_combout ),
	.q(\so_count[5]~q ),
	.prn(vcc));
defparam \so_count[5] .is_wysiwyg = "true";
defparam \so_count[5] .power_up = "low";

cycloneive_lcell_comb \so_count[6]~21 (
	.dataa(\so_count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\so_count[5]~20 ),
	.combout(\so_count[6]~21_combout ),
	.cout(\so_count[6]~22 ));
defparam \so_count[6]~21 .lut_mask = 16'h5AAF;
defparam \so_count[6]~21 .sum_lutc_input = "cin";

dffeas \so_count[6] (
	.clk(clk),
	.d(\so_count[6]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(counter_i),
	.sload(gnd),
	.ena(\so_count[0]~10_combout ),
	.q(\so_count[6]~q ),
	.prn(vcc));
defparam \so_count[6] .is_wysiwyg = "true";
defparam \so_count[6] .power_up = "low";

cycloneive_lcell_comb \so_count[7]~23 (
	.dataa(\so_count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\so_count[6]~22 ),
	.combout(\so_count[7]~23_combout ),
	.cout());
defparam \so_count[7]~23 .lut_mask = 16'h5A5A;
defparam \so_count[7]~23 .sum_lutc_input = "cin";

dffeas \so_count[7] (
	.clk(clk),
	.d(\so_count[7]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(counter_i),
	.sload(gnd),
	.ena(\so_count[0]~10_combout ),
	.q(\so_count[7]~q ),
	.prn(vcc));
defparam \so_count[7] .is_wysiwyg = "true";
defparam \so_count[7] .power_up = "low";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\Equal0~0_combout ),
	.datab(\so_count[5]~q ),
	.datac(\so_count[6]~q ),
	.datad(\so_count[7]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hFFFE;
defparam \Equal0~1 .sum_lutc_input = "datac";

dffeas \so_count[2] (
	.clk(clk),
	.d(\so_count[2]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(counter_i),
	.sload(gnd),
	.ena(\so_count[0]~10_combout ),
	.q(\so_count[2]~q ),
	.prn(vcc));
defparam \so_count[2] .is_wysiwyg = "true";
defparam \so_count[2] .power_up = "low";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(\Equal0~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\so_count[2]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hAAFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\so_count[2]~q ),
	.datab(\Equal0~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hEEEE;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_rdy_int~0 (
	.dataa(rdy_for_next_block1),
	.datab(data_rdy_int1),
	.datac(gnd),
	.datad(blk_done),
	.cin(gnd),
	.combout(\data_rdy_int~0_combout ),
	.cout());
defparam \data_rdy_int~0 .lut_mask = 16'hEEFF;
defparam \data_rdy_int~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~0 (
	.dataa(reset_n),
	.datab(core_imag_in_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~0_combout ),
	.cout());
defparam \data_in_i~0 .lut_mask = 16'hEEEE;
defparam \data_in_i~0 .sum_lutc_input = "datac";

dffeas \so_count[0] (
	.clk(clk),
	.d(\so_count[0]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(counter_i),
	.sload(gnd),
	.ena(\so_count[0]~10_combout ),
	.q(\so_count[0]~q ),
	.prn(vcc));
defparam \so_count[0] .is_wysiwyg = "true";
defparam \so_count[0] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_early~0 (
	.dataa(reset_n),
	.datab(\so_count[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_early~0_combout ),
	.cout());
defparam \wr_address_i_early~0 .lut_mask = 16'hEEEE;
defparam \wr_address_i_early~0 .sum_lutc_input = "datac";

dffeas \wr_address_i_early[0] (
	.clk(clk),
	.d(\wr_address_i_early~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_address_i_early[0]~q ),
	.prn(vcc));
defparam \wr_address_i_early[0] .is_wysiwyg = "true";
defparam \wr_address_i_early[0] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_int~0 (
	.dataa(reset_n),
	.datab(\wr_address_i_early[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~0_combout ),
	.cout());
defparam \wr_address_i_int~0 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~0 .sum_lutc_input = "datac";

dffeas \so_count[1] (
	.clk(clk),
	.d(\so_count[1]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(counter_i),
	.sload(gnd),
	.ena(\so_count[0]~10_combout ),
	.q(\so_count[1]~q ),
	.prn(vcc));
defparam \so_count[1] .is_wysiwyg = "true";
defparam \so_count[1] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_early~1 (
	.dataa(reset_n),
	.datab(\so_count[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_early~1_combout ),
	.cout());
defparam \wr_address_i_early~1 .lut_mask = 16'hEEEE;
defparam \wr_address_i_early~1 .sum_lutc_input = "datac";

dffeas \wr_address_i_early[1] (
	.clk(clk),
	.d(\wr_address_i_early~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_address_i_early[1]~q ),
	.prn(vcc));
defparam \wr_address_i_early[1] .is_wysiwyg = "true";
defparam \wr_address_i_early[1] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_int~1 (
	.dataa(reset_n),
	.datab(\wr_address_i_early[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~1_combout ),
	.cout());
defparam \wr_address_i_int~1 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_address_i_early~2 (
	.dataa(reset_n),
	.datab(\so_count[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_early~2_combout ),
	.cout());
defparam \wr_address_i_early~2 .lut_mask = 16'hEEEE;
defparam \wr_address_i_early~2 .sum_lutc_input = "datac";

dffeas \wr_address_i_early[2] (
	.clk(clk),
	.d(\wr_address_i_early~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_address_i_early[2]~q ),
	.prn(vcc));
defparam \wr_address_i_early[2] .is_wysiwyg = "true";
defparam \wr_address_i_early[2] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_int~2 (
	.dataa(reset_n),
	.datab(\wr_address_i_early[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~2_combout ),
	.cout());
defparam \wr_address_i_int~2 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~2 .sum_lutc_input = "datac";

dffeas \so_count[3] (
	.clk(clk),
	.d(\so_count[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(counter_i),
	.sload(gnd),
	.ena(\so_count[0]~10_combout ),
	.q(\so_count[3]~q ),
	.prn(vcc));
defparam \so_count[3] .is_wysiwyg = "true";
defparam \so_count[3] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_early~3 (
	.dataa(reset_n),
	.datab(\so_count[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_early~3_combout ),
	.cout());
defparam \wr_address_i_early~3 .lut_mask = 16'hEEEE;
defparam \wr_address_i_early~3 .sum_lutc_input = "datac";

dffeas \wr_address_i_early[3] (
	.clk(clk),
	.d(\wr_address_i_early~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_address_i_early[3]~q ),
	.prn(vcc));
defparam \wr_address_i_early[3] .is_wysiwyg = "true";
defparam \wr_address_i_early[3] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_int~3 (
	.dataa(reset_n),
	.datab(\wr_address_i_early[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~3_combout ),
	.cout());
defparam \wr_address_i_int~3 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~3 .sum_lutc_input = "datac";

dffeas \so_count[4] (
	.clk(clk),
	.d(\so_count[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(counter_i),
	.sload(gnd),
	.ena(\so_count[0]~10_combout ),
	.q(\so_count[4]~q ),
	.prn(vcc));
defparam \so_count[4] .is_wysiwyg = "true";
defparam \so_count[4] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_early~4 (
	.dataa(reset_n),
	.datab(\so_count[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_early~4_combout ),
	.cout());
defparam \wr_address_i_early~4 .lut_mask = 16'hEEEE;
defparam \wr_address_i_early~4 .sum_lutc_input = "datac";

dffeas \wr_address_i_early[4] (
	.clk(clk),
	.d(\wr_address_i_early~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_address_i_early[4]~q ),
	.prn(vcc));
defparam \wr_address_i_early[4] .is_wysiwyg = "true";
defparam \wr_address_i_early[4] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_int~4 (
	.dataa(reset_n),
	.datab(\wr_address_i_early[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~4_combout ),
	.cout());
defparam \wr_address_i_int~4 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_address_i_early~5 (
	.dataa(reset_n),
	.datab(\so_count[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_early~5_combout ),
	.cout());
defparam \wr_address_i_early~5 .lut_mask = 16'hEEEE;
defparam \wr_address_i_early~5 .sum_lutc_input = "datac";

dffeas \wr_address_i_early[5] (
	.clk(clk),
	.d(\wr_address_i_early~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_address_i_early[5]~q ),
	.prn(vcc));
defparam \wr_address_i_early[5] .is_wysiwyg = "true";
defparam \wr_address_i_early[5] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_int~5 (
	.dataa(reset_n),
	.datab(\wr_address_i_early[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~5_combout ),
	.cout());
defparam \wr_address_i_int~5 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_address_i_early~6 (
	.dataa(reset_n),
	.datab(\so_count[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_early~6_combout ),
	.cout());
defparam \wr_address_i_early~6 .lut_mask = 16'hEEEE;
defparam \wr_address_i_early~6 .sum_lutc_input = "datac";

dffeas \wr_address_i_early[6] (
	.clk(clk),
	.d(\wr_address_i_early~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_address_i_early[6]~q ),
	.prn(vcc));
defparam \wr_address_i_early[6] .is_wysiwyg = "true";
defparam \wr_address_i_early[6] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_int~6 (
	.dataa(reset_n),
	.datab(\wr_address_i_early[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~6_combout ),
	.cout());
defparam \wr_address_i_int~6 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_address_i_early~7 (
	.dataa(reset_n),
	.datab(\so_count[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_early~7_combout ),
	.cout());
defparam \wr_address_i_early~7 .lut_mask = 16'hEEEE;
defparam \wr_address_i_early~7 .sum_lutc_input = "datac";

dffeas \wr_address_i_early[7] (
	.clk(clk),
	.d(\wr_address_i_early~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_address_i_early[7]~q ),
	.prn(vcc));
defparam \wr_address_i_early[7] .is_wysiwyg = "true";
defparam \wr_address_i_early[7] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_int~7 (
	.dataa(reset_n),
	.datab(\wr_address_i_early[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~7_combout ),
	.cout());
defparam \wr_address_i_int~7 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~0 (
	.dataa(reset_n),
	.datab(core_real_in_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~0_combout ),
	.cout());
defparam \data_in_r~0 .lut_mask = 16'hEEEE;
defparam \data_in_r~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~1 (
	.dataa(reset_n),
	.datab(core_imag_in_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~1_combout ),
	.cout());
defparam \data_in_i~1 .lut_mask = 16'hEEEE;
defparam \data_in_i~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~1 (
	.dataa(reset_n),
	.datab(core_real_in_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~1_combout ),
	.cout());
defparam \data_in_r~1 .lut_mask = 16'hEEEE;
defparam \data_in_r~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~2 (
	.dataa(reset_n),
	.datab(core_imag_in_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~2_combout ),
	.cout());
defparam \data_in_i~2 .lut_mask = 16'hEEEE;
defparam \data_in_i~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~2 (
	.dataa(reset_n),
	.datab(core_real_in_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~2_combout ),
	.cout());
defparam \data_in_r~2 .lut_mask = 16'hEEEE;
defparam \data_in_r~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~3 (
	.dataa(reset_n),
	.datab(core_imag_in_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~3_combout ),
	.cout());
defparam \data_in_i~3 .lut_mask = 16'hEEEE;
defparam \data_in_i~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~3 (
	.dataa(reset_n),
	.datab(core_real_in_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~3_combout ),
	.cout());
defparam \data_in_r~3 .lut_mask = 16'hEEEE;
defparam \data_in_r~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~4 (
	.dataa(reset_n),
	.datab(core_imag_in_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~4_combout ),
	.cout());
defparam \data_in_i~4 .lut_mask = 16'hEEEE;
defparam \data_in_i~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~4 (
	.dataa(reset_n),
	.datab(core_real_in_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~4_combout ),
	.cout());
defparam \data_in_r~4 .lut_mask = 16'hEEEE;
defparam \data_in_r~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~5 (
	.dataa(reset_n),
	.datab(core_imag_in_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~5_combout ),
	.cout());
defparam \data_in_i~5 .lut_mask = 16'hEEEE;
defparam \data_in_i~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~5 (
	.dataa(reset_n),
	.datab(core_real_in_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~5_combout ),
	.cout());
defparam \data_in_r~5 .lut_mask = 16'hEEEE;
defparam \data_in_r~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~6 (
	.dataa(reset_n),
	.datab(core_imag_in_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~6_combout ),
	.cout());
defparam \data_in_i~6 .lut_mask = 16'hEEEE;
defparam \data_in_i~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~6 (
	.dataa(reset_n),
	.datab(core_real_in_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~6_combout ),
	.cout());
defparam \data_in_r~6 .lut_mask = 16'hEEEE;
defparam \data_in_r~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~7 (
	.dataa(reset_n),
	.datab(core_imag_in_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~7_combout ),
	.cout());
defparam \data_in_i~7 .lut_mask = 16'hEEEE;
defparam \data_in_i~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~7 (
	.dataa(reset_n),
	.datab(core_real_in_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~7_combout ),
	.cout());
defparam \data_in_r~7 .lut_mask = 16'hEEEE;
defparam \data_in_r~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~8 (
	.dataa(reset_n),
	.datab(core_imag_in_8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~8_combout ),
	.cout());
defparam \data_in_i~8 .lut_mask = 16'hEEEE;
defparam \data_in_i~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~8 (
	.dataa(reset_n),
	.datab(core_real_in_8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~8_combout ),
	.cout());
defparam \data_in_r~8 .lut_mask = 16'hEEEE;
defparam \data_in_r~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~9 (
	.dataa(reset_n),
	.datab(core_imag_in_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~9_combout ),
	.cout());
defparam \data_in_i~9 .lut_mask = 16'hEEEE;
defparam \data_in_i~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~9 (
	.dataa(reset_n),
	.datab(core_real_in_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~9_combout ),
	.cout());
defparam \data_in_r~9 .lut_mask = 16'hEEEE;
defparam \data_in_r~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~10 (
	.dataa(reset_n),
	.datab(core_imag_in_10),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~10_combout ),
	.cout());
defparam \data_in_i~10 .lut_mask = 16'hEEEE;
defparam \data_in_i~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~10 (
	.dataa(reset_n),
	.datab(core_real_in_10),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~10_combout ),
	.cout());
defparam \data_in_r~10 .lut_mask = 16'hEEEE;
defparam \data_in_r~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~11 (
	.dataa(reset_n),
	.datab(core_imag_in_11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~11_combout ),
	.cout());
defparam \data_in_i~11 .lut_mask = 16'hEEEE;
defparam \data_in_i~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~11 (
	.dataa(reset_n),
	.datab(core_real_in_11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~11_combout ),
	.cout());
defparam \data_in_r~11 .lut_mask = 16'hEEEE;
defparam \data_in_r~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~12 (
	.dataa(reset_n),
	.datab(core_imag_in_12),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~12_combout ),
	.cout());
defparam \data_in_i~12 .lut_mask = 16'hEEEE;
defparam \data_in_i~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~12 (
	.dataa(reset_n),
	.datab(core_real_in_12),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~12_combout ),
	.cout());
defparam \data_in_r~12 .lut_mask = 16'hEEEE;
defparam \data_in_r~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~13 (
	.dataa(reset_n),
	.datab(core_imag_in_13),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~13_combout ),
	.cout());
defparam \data_in_i~13 .lut_mask = 16'hEEEE;
defparam \data_in_i~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~13 (
	.dataa(reset_n),
	.datab(core_real_in_13),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~13_combout ),
	.cout());
defparam \data_in_r~13 .lut_mask = 16'hEEEE;
defparam \data_in_r~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~14 (
	.dataa(reset_n),
	.datab(core_imag_in_14),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~14_combout ),
	.cout());
defparam \data_in_i~14 .lut_mask = 16'hEEEE;
defparam \data_in_i~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~14 (
	.dataa(reset_n),
	.datab(core_real_in_14),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~14_combout ),
	.cout());
defparam \data_in_r~14 .lut_mask = 16'hEEEE;
defparam \data_in_r~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~15 (
	.dataa(reset_n),
	.datab(core_imag_in_15),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~15_combout ),
	.cout());
defparam \data_in_i~15 .lut_mask = 16'hEEEE;
defparam \data_in_i~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~15 (
	.dataa(reset_n),
	.datab(core_real_in_15),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~15_combout ),
	.cout());
defparam \data_in_r~15 .lut_mask = 16'hEEEE;
defparam \data_in_r~15 .sum_lutc_input = "datac";

endmodule

module fft256_asj_fft_tdl_bit_rst_fft_121_1 (
	global_clock_enable,
	tdl_arr_0,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_0;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \tdl_arr[0] (
	.clk(clk),
	.d(reset_n),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_0),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

endmodule

module fft256_asj_fft_m_k_counter_fft_121 (
	rdy_for_next_block,
	send_sop_s,
	global_clock_enable,
	blk_done1,
	counter_i,
	p_2,
	p_0,
	p_1,
	rd_addr_a_0,
	k_count_2,
	k_count_0,
	k_count_6,
	k_count_3,
	k_count_1,
	k_count_7,
	k_count_4,
	k_count_5,
	data_rdy_vec_4,
	next_pass_i1,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	rdy_for_next_block;
input 	send_sop_s;
input 	global_clock_enable;
output 	blk_done1;
input 	counter_i;
output 	p_2;
output 	p_0;
output 	p_1;
input 	rd_addr_a_0;
output 	k_count_2;
output 	k_count_0;
output 	k_count_6;
output 	k_count_3;
output 	k_count_1;
output 	k_count_7;
output 	k_count_4;
output 	k_count_5;
input 	data_rdy_vec_4;
output 	next_pass_i1;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \del_npi_cnt[0]~q ;
wire \del_npi_cnt[1]~q ;
wire \del_npi_cnt[2]~q ;
wire \del_npi_cnt[4]~q ;
wire \del_npi_cnt[3]~q ;
wire \del_npi_cnt[0]~7 ;
wire \del_npi_cnt[0]~6_combout ;
wire \del_npi_cnt[1]~9 ;
wire \del_npi_cnt[1]~8_combout ;
wire \del_npi_cnt[2]~11 ;
wire \del_npi_cnt[2]~10_combout ;
wire \del_npi_cnt[3]~13 ;
wire \del_npi_cnt[3]~12_combout ;
wire \del_npi_cnt[4]~14_combout ;
wire \Add1~0_combout ;
wire \next_pass_id~q ;
wire \k_state.HOLD~q ;
wire \k_state.IDLE~q ;
wire \k_state~10_combout ;
wire \next_pass_id~0_combout ;
wire \next_pass_id~1_combout ;
wire \k_state.HOLD~2_combout ;
wire \k_state.IDLE~2_combout ;
wire \k_state.HOLD~3_combout ;
wire \k_state.IDLE~3_combout ;
wire \p[0]~1_combout ;
wire \p~2_combout ;
wire \p[0]~0_combout ;
wire \p[0]~3_combout ;
wire \p[3]~q ;
wire \k[0]~11 ;
wire \k[1]~13 ;
wire \k[2]~15 ;
wire \k[3]~17 ;
wire \k[4]~19 ;
wire \k[5]~20_combout ;
wire \k[1]~12_combout ;
wire \k[1]~q ;
wire \k[2]~14_combout ;
wire \k[2]~q ;
wire \k[3]~16_combout ;
wire \k[3]~q ;
wire \Equal2~0_combout ;
wire \k_state~11_combout ;
wire \k_state~12_combout ;
wire \k_state.RUN_CNT~q ;
wire \k[0]~26_combout ;
wire \k[5]~q ;
wire \k[5]~21 ;
wire \k[6]~22_combout ;
wire \k[6]~q ;
wire \k[6]~23 ;
wire \k[7]~24_combout ;
wire \k[7]~q ;
wire \Equal2~1_combout ;
wire \k_state~9_combout ;
wire \k_state.NEXT_PASS_UPD~q ;
wire \blk_done~0_combout ;
wire \blk_done~1_combout ;
wire \p~4_combout ;
wire \p~5_combout ;
wire \p~6_combout ;
wire \k[0]~10_combout ;
wire \k[0]~q ;
wire \k[4]~18_combout ;
wire \k[4]~q ;


dffeas \del_npi_cnt[0] (
	.clk(clk),
	.d(\del_npi_cnt[0]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_state.HOLD~q ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_npi_cnt[0]~q ),
	.prn(vcc));
defparam \del_npi_cnt[0] .is_wysiwyg = "true";
defparam \del_npi_cnt[0] .power_up = "low";

dffeas \del_npi_cnt[1] (
	.clk(clk),
	.d(\del_npi_cnt[1]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_state.HOLD~q ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_npi_cnt[1]~q ),
	.prn(vcc));
defparam \del_npi_cnt[1] .is_wysiwyg = "true";
defparam \del_npi_cnt[1] .power_up = "low";

dffeas \del_npi_cnt[2] (
	.clk(clk),
	.d(\del_npi_cnt[2]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_state.HOLD~q ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_npi_cnt[2]~q ),
	.prn(vcc));
defparam \del_npi_cnt[2] .is_wysiwyg = "true";
defparam \del_npi_cnt[2] .power_up = "low";

dffeas \del_npi_cnt[4] (
	.clk(clk),
	.d(\del_npi_cnt[4]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_state.HOLD~q ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_npi_cnt[4]~q ),
	.prn(vcc));
defparam \del_npi_cnt[4] .is_wysiwyg = "true";
defparam \del_npi_cnt[4] .power_up = "low";

dffeas \del_npi_cnt[3] (
	.clk(clk),
	.d(\del_npi_cnt[3]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_state.HOLD~q ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_npi_cnt[3]~q ),
	.prn(vcc));
defparam \del_npi_cnt[3] .is_wysiwyg = "true";
defparam \del_npi_cnt[3] .power_up = "low";

cycloneive_lcell_comb \del_npi_cnt[0]~6 (
	.dataa(\del_npi_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\del_npi_cnt[0]~6_combout ),
	.cout(\del_npi_cnt[0]~7 ));
defparam \del_npi_cnt[0]~6 .lut_mask = 16'h55AA;
defparam \del_npi_cnt[0]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \del_npi_cnt[1]~8 (
	.dataa(\del_npi_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_npi_cnt[0]~7 ),
	.combout(\del_npi_cnt[1]~8_combout ),
	.cout(\del_npi_cnt[1]~9 ));
defparam \del_npi_cnt[1]~8 .lut_mask = 16'h5A5F;
defparam \del_npi_cnt[1]~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \del_npi_cnt[2]~10 (
	.dataa(\del_npi_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_npi_cnt[1]~9 ),
	.combout(\del_npi_cnt[2]~10_combout ),
	.cout(\del_npi_cnt[2]~11 ));
defparam \del_npi_cnt[2]~10 .lut_mask = 16'h5AAF;
defparam \del_npi_cnt[2]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \del_npi_cnt[3]~12 (
	.dataa(\del_npi_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_npi_cnt[2]~11 ),
	.combout(\del_npi_cnt[3]~12_combout ),
	.cout(\del_npi_cnt[3]~13 ));
defparam \del_npi_cnt[3]~12 .lut_mask = 16'h5A5F;
defparam \del_npi_cnt[3]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \del_npi_cnt[4]~14 (
	.dataa(\del_npi_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\del_npi_cnt[3]~13 ),
	.combout(\del_npi_cnt[4]~14_combout ),
	.cout());
defparam \del_npi_cnt[4]~14 .lut_mask = 16'h5A5A;
defparam \del_npi_cnt[4]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~0 (
	.dataa(\p[3]~q ),
	.datab(p_2),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h6996;
defparam \Add1~0 .sum_lutc_input = "datac";

dffeas next_pass_id(
	.clk(clk),
	.d(\next_pass_id~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\next_pass_id~q ),
	.prn(vcc));
defparam next_pass_id.is_wysiwyg = "true";
defparam next_pass_id.power_up = "low";

dffeas \k_state.HOLD (
	.clk(clk),
	.d(\k_state.HOLD~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\k_state.HOLD~q ),
	.prn(vcc));
defparam \k_state.HOLD .is_wysiwyg = "true";
defparam \k_state.HOLD .power_up = "low";

dffeas \k_state.IDLE (
	.clk(clk),
	.d(\k_state.IDLE~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\k_state.IDLE~q ),
	.prn(vcc));
defparam \k_state.IDLE .is_wysiwyg = "true";
defparam \k_state.IDLE .power_up = "low";

cycloneive_lcell_comb \k_state~10 (
	.dataa(\next_pass_id~q ),
	.datab(\k_state.HOLD~q ),
	.datac(data_rdy_vec_4),
	.datad(\k_state.IDLE~q ),
	.cin(gnd),
	.combout(\k_state~10_combout ),
	.cout());
defparam \k_state~10 .lut_mask = 16'hFEFF;
defparam \k_state~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_pass_id~0 (
	.dataa(\k_state.HOLD~q ),
	.datab(\del_npi_cnt[0]~q ),
	.datac(\del_npi_cnt[1]~q ),
	.datad(\del_npi_cnt[2]~q ),
	.cin(gnd),
	.combout(\next_pass_id~0_combout ),
	.cout());
defparam \next_pass_id~0 .lut_mask = 16'hEFFF;
defparam \next_pass_id~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_pass_id~1 (
	.dataa(\next_pass_id~0_combout ),
	.datab(\del_npi_cnt[4]~q ),
	.datac(gnd),
	.datad(\del_npi_cnt[3]~q ),
	.cin(gnd),
	.combout(\next_pass_id~1_combout ),
	.cout());
defparam \next_pass_id~1 .lut_mask = 16'hEEFF;
defparam \next_pass_id~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \k_state.HOLD~2 (
	.dataa(\k_state.HOLD~q ),
	.datab(data_rdy_vec_4),
	.datac(next_pass_i1),
	.datad(\next_pass_id~q ),
	.cin(gnd),
	.combout(\k_state.HOLD~2_combout ),
	.cout());
defparam \k_state.HOLD~2 .lut_mask = 16'hEFFF;
defparam \k_state.HOLD~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \k_state.IDLE~2 (
	.dataa(next_pass_i1),
	.datab(\k_state.HOLD~q ),
	.datac(\next_pass_id~q ),
	.datad(\k_state.IDLE~q ),
	.cin(gnd),
	.combout(\k_state.IDLE~2_combout ),
	.cout());
defparam \k_state.IDLE~2 .lut_mask = 16'hEFFF;
defparam \k_state.IDLE~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \k_state.HOLD~3 (
	.dataa(send_sop_s),
	.datab(reset_n),
	.datac(\k_state.NEXT_PASS_UPD~q ),
	.datad(\k_state.HOLD~2_combout ),
	.cin(gnd),
	.combout(\k_state.HOLD~3_combout ),
	.cout());
defparam \k_state.HOLD~3 .lut_mask = 16'hFFFD;
defparam \k_state.HOLD~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \k_state.IDLE~3 (
	.dataa(send_sop_s),
	.datab(reset_n),
	.datac(\k_state.IDLE~2_combout ),
	.datad(data_rdy_vec_4),
	.cin(gnd),
	.combout(\k_state.IDLE~3_combout ),
	.cout());
defparam \k_state.IDLE~3 .lut_mask = 16'hFFDF;
defparam \k_state.IDLE~3 .sum_lutc_input = "datac";

dffeas blk_done(
	.clk(clk),
	.d(\blk_done~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(blk_done1),
	.prn(vcc));
defparam blk_done.is_wysiwyg = "true";
defparam blk_done.power_up = "low";

dffeas \p[2] (
	.clk(clk),
	.d(\p~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p[0]~3_combout ),
	.q(p_2),
	.prn(vcc));
defparam \p[2] .is_wysiwyg = "true";
defparam \p[2] .power_up = "low";

dffeas \p[0] (
	.clk(clk),
	.d(\p~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p[0]~3_combout ),
	.q(p_0),
	.prn(vcc));
defparam \p[0] .is_wysiwyg = "true";
defparam \p[0] .power_up = "low";

dffeas \p[1] (
	.clk(clk),
	.d(\p~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p[0]~3_combout ),
	.q(p_1),
	.prn(vcc));
defparam \p[1] .is_wysiwyg = "true";
defparam \p[1] .power_up = "low";

dffeas \k_count[2] (
	.clk(clk),
	.d(\k[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_2),
	.prn(vcc));
defparam \k_count[2] .is_wysiwyg = "true";
defparam \k_count[2] .power_up = "low";

dffeas \k_count[0] (
	.clk(clk),
	.d(\k[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_0),
	.prn(vcc));
defparam \k_count[0] .is_wysiwyg = "true";
defparam \k_count[0] .power_up = "low";

dffeas \k_count[6] (
	.clk(clk),
	.d(\k[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_6),
	.prn(vcc));
defparam \k_count[6] .is_wysiwyg = "true";
defparam \k_count[6] .power_up = "low";

dffeas \k_count[3] (
	.clk(clk),
	.d(\k[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_3),
	.prn(vcc));
defparam \k_count[3] .is_wysiwyg = "true";
defparam \k_count[3] .power_up = "low";

dffeas \k_count[1] (
	.clk(clk),
	.d(\k[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_1),
	.prn(vcc));
defparam \k_count[1] .is_wysiwyg = "true";
defparam \k_count[1] .power_up = "low";

dffeas \k_count[7] (
	.clk(clk),
	.d(\k[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_7),
	.prn(vcc));
defparam \k_count[7] .is_wysiwyg = "true";
defparam \k_count[7] .power_up = "low";

dffeas \k_count[4] (
	.clk(clk),
	.d(\k[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_4),
	.prn(vcc));
defparam \k_count[4] .is_wysiwyg = "true";
defparam \k_count[4] .power_up = "low";

dffeas \k_count[5] (
	.clk(clk),
	.d(\k[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_5),
	.prn(vcc));
defparam \k_count[5] .is_wysiwyg = "true";
defparam \k_count[5] .power_up = "low";

dffeas next_pass_i(
	.clk(clk),
	.d(\blk_done~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(next_pass_i1),
	.prn(vcc));
defparam next_pass_i.is_wysiwyg = "true";
defparam next_pass_i.power_up = "low";

cycloneive_lcell_comb \p[0]~1 (
	.dataa(\p[0]~0_combout ),
	.datab(\p[3]~q ),
	.datac(p_2),
	.datad(rd_addr_a_0),
	.cin(gnd),
	.combout(\p[0]~1_combout ),
	.cout());
defparam \p[0]~1 .lut_mask = 16'hDFFF;
defparam \p[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p~2 (
	.dataa(\Add1~0_combout ),
	.datab(\p[0]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p~2_combout ),
	.cout());
defparam \p~2 .lut_mask = 16'hEEEE;
defparam \p~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p[0]~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(rdy_for_next_block),
	.cin(gnd),
	.combout(\p[0]~0_combout ),
	.cout());
defparam \p[0]~0 .lut_mask = 16'hFF55;
defparam \p[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p[0]~3 (
	.dataa(global_clock_enable),
	.datab(\p[0]~0_combout ),
	.datac(data_rdy_vec_4),
	.datad(next_pass_i1),
	.cin(gnd),
	.combout(\p[0]~3_combout ),
	.cout());
defparam \p[0]~3 .lut_mask = 16'hFFFE;
defparam \p[0]~3 .sum_lutc_input = "datac";

dffeas \p[3] (
	.clk(clk),
	.d(\p~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p[0]~3_combout ),
	.q(\p[3]~q ),
	.prn(vcc));
defparam \p[3] .is_wysiwyg = "true";
defparam \p[3] .power_up = "low";

cycloneive_lcell_comb \k[0]~10 (
	.dataa(\k[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\k[0]~10_combout ),
	.cout(\k[0]~11 ));
defparam \k[0]~10 .lut_mask = 16'h55AA;
defparam \k[0]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \k[1]~12 (
	.dataa(\k[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k[0]~11 ),
	.combout(\k[1]~12_combout ),
	.cout(\k[1]~13 ));
defparam \k[1]~12 .lut_mask = 16'h5A5F;
defparam \k[1]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \k[2]~14 (
	.dataa(\k[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k[1]~13 ),
	.combout(\k[2]~14_combout ),
	.cout(\k[2]~15 ));
defparam \k[2]~14 .lut_mask = 16'h5AAF;
defparam \k[2]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \k[3]~16 (
	.dataa(\k[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k[2]~15 ),
	.combout(\k[3]~16_combout ),
	.cout(\k[3]~17 ));
defparam \k[3]~16 .lut_mask = 16'h5A5F;
defparam \k[3]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \k[4]~18 (
	.dataa(\k[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k[3]~17 ),
	.combout(\k[4]~18_combout ),
	.cout(\k[4]~19 ));
defparam \k[4]~18 .lut_mask = 16'h5AAF;
defparam \k[4]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \k[5]~20 (
	.dataa(\k[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k[4]~19 ),
	.combout(\k[5]~20_combout ),
	.cout(\k[5]~21 ));
defparam \k[5]~20 .lut_mask = 16'h5A5F;
defparam \k[5]~20 .sum_lutc_input = "cin";

dffeas \k[1] (
	.clk(clk),
	.d(\k[1]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\p[0]~0_combout ),
	.sload(gnd),
	.ena(\k[0]~26_combout ),
	.q(\k[1]~q ),
	.prn(vcc));
defparam \k[1] .is_wysiwyg = "true";
defparam \k[1] .power_up = "low";

dffeas \k[2] (
	.clk(clk),
	.d(\k[2]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\p[0]~0_combout ),
	.sload(gnd),
	.ena(\k[0]~26_combout ),
	.q(\k[2]~q ),
	.prn(vcc));
defparam \k[2] .is_wysiwyg = "true";
defparam \k[2] .power_up = "low";

dffeas \k[3] (
	.clk(clk),
	.d(\k[3]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\p[0]~0_combout ),
	.sload(gnd),
	.ena(\k[0]~26_combout ),
	.q(\k[3]~q ),
	.prn(vcc));
defparam \k[3] .is_wysiwyg = "true";
defparam \k[3] .power_up = "low";

cycloneive_lcell_comb \Equal2~0 (
	.dataa(\k[0]~q ),
	.datab(\k[1]~q ),
	.datac(\k[2]~q ),
	.datad(\k[3]~q ),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hFFFE;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \k_state~11 (
	.dataa(\k_state~10_combout ),
	.datab(\k_state.RUN_CNT~q ),
	.datac(\Equal2~0_combout ),
	.datad(\Equal2~1_combout ),
	.cin(gnd),
	.combout(\k_state~11_combout ),
	.cout());
defparam \k_state~11 .lut_mask = 16'hEFFF;
defparam \k_state~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \k_state~12 (
	.dataa(send_sop_s),
	.datab(reset_n),
	.datac(\k_state~11_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\k_state~12_combout ),
	.cout());
defparam \k_state~12 .lut_mask = 16'hFDFD;
defparam \k_state~12 .sum_lutc_input = "datac";

dffeas \k_state.RUN_CNT (
	.clk(clk),
	.d(\k_state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\k_state.RUN_CNT~q ),
	.prn(vcc));
defparam \k_state.RUN_CNT .is_wysiwyg = "true";
defparam \k_state.RUN_CNT .power_up = "low";

cycloneive_lcell_comb \k[0]~26 (
	.dataa(reset_n),
	.datab(rdy_for_next_block),
	.datac(\k_state.RUN_CNT~q ),
	.datad(global_clock_enable),
	.cin(gnd),
	.combout(\k[0]~26_combout ),
	.cout());
defparam \k[0]~26 .lut_mask = 16'hFFFD;
defparam \k[0]~26 .sum_lutc_input = "datac";

dffeas \k[5] (
	.clk(clk),
	.d(\k[5]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\p[0]~0_combout ),
	.sload(gnd),
	.ena(\k[0]~26_combout ),
	.q(\k[5]~q ),
	.prn(vcc));
defparam \k[5] .is_wysiwyg = "true";
defparam \k[5] .power_up = "low";

cycloneive_lcell_comb \k[6]~22 (
	.dataa(\k[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k[5]~21 ),
	.combout(\k[6]~22_combout ),
	.cout(\k[6]~23 ));
defparam \k[6]~22 .lut_mask = 16'h5AAF;
defparam \k[6]~22 .sum_lutc_input = "cin";

dffeas \k[6] (
	.clk(clk),
	.d(\k[6]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\p[0]~0_combout ),
	.sload(gnd),
	.ena(\k[0]~26_combout ),
	.q(\k[6]~q ),
	.prn(vcc));
defparam \k[6] .is_wysiwyg = "true";
defparam \k[6] .power_up = "low";

cycloneive_lcell_comb \k[7]~24 (
	.dataa(\k[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\k[6]~23 ),
	.combout(\k[7]~24_combout ),
	.cout());
defparam \k[7]~24 .lut_mask = 16'h5A5A;
defparam \k[7]~24 .sum_lutc_input = "cin";

dffeas \k[7] (
	.clk(clk),
	.d(\k[7]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\p[0]~0_combout ),
	.sload(gnd),
	.ena(\k[0]~26_combout ),
	.q(\k[7]~q ),
	.prn(vcc));
defparam \k[7] .is_wysiwyg = "true";
defparam \k[7] .power_up = "low";

cycloneive_lcell_comb \Equal2~1 (
	.dataa(\k[4]~q ),
	.datab(\k[5]~q ),
	.datac(\k[6]~q ),
	.datad(\k[7]~q ),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
defparam \Equal2~1 .lut_mask = 16'hFFFE;
defparam \Equal2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \k_state~9 (
	.dataa(\Equal2~0_combout ),
	.datab(\Equal2~1_combout ),
	.datac(\k_state.RUN_CNT~q ),
	.datad(counter_i),
	.cin(gnd),
	.combout(\k_state~9_combout ),
	.cout());
defparam \k_state~9 .lut_mask = 16'hFEFF;
defparam \k_state~9 .sum_lutc_input = "datac";

dffeas \k_state.NEXT_PASS_UPD (
	.clk(clk),
	.d(\k_state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\k_state.NEXT_PASS_UPD~q ),
	.prn(vcc));
defparam \k_state.NEXT_PASS_UPD .is_wysiwyg = "true";
defparam \k_state.NEXT_PASS_UPD .power_up = "low";

cycloneive_lcell_comb \blk_done~0 (
	.dataa(reset_n),
	.datab(\k_state.NEXT_PASS_UPD~q ),
	.datac(gnd),
	.datad(send_sop_s),
	.cin(gnd),
	.combout(\blk_done~0_combout ),
	.cout());
defparam \blk_done~0 .lut_mask = 16'hEEFF;
defparam \blk_done~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_done~1 (
	.dataa(\p[3]~q ),
	.datab(\blk_done~0_combout ),
	.datac(p_2),
	.datad(rd_addr_a_0),
	.cin(gnd),
	.combout(\blk_done~1_combout ),
	.cout());
defparam \blk_done~1 .lut_mask = 16'hFFFD;
defparam \blk_done~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p~4 (
	.dataa(\p[0]~1_combout ),
	.datab(p_2),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\p~4_combout ),
	.cout());
defparam \p~4 .lut_mask = 16'hEBBE;
defparam \p~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p~5 (
	.dataa(reset_n),
	.datab(rdy_for_next_block),
	.datac(\p[0]~1_combout ),
	.datad(p_0),
	.cin(gnd),
	.combout(\p~5_combout ),
	.cout());
defparam \p~5 .lut_mask = 16'hFEFF;
defparam \p~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p~6 (
	.dataa(\p[0]~1_combout ),
	.datab(gnd),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\p~6_combout ),
	.cout());
defparam \p~6 .lut_mask = 16'hAFFA;
defparam \p~6 .sum_lutc_input = "datac";

dffeas \k[0] (
	.clk(clk),
	.d(\k[0]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\p[0]~0_combout ),
	.sload(gnd),
	.ena(\k[0]~26_combout ),
	.q(\k[0]~q ),
	.prn(vcc));
defparam \k[0] .is_wysiwyg = "true";
defparam \k[0] .power_up = "low";

dffeas \k[4] (
	.clk(clk),
	.d(\k[4]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\p[0]~0_combout ),
	.sload(gnd),
	.ena(\k[0]~26_combout ),
	.q(\k[4]~q ),
	.prn(vcc));
defparam \k[4] .is_wysiwyg = "true";
defparam \k[4] .power_up = "low";

endmodule

module fft256_asj_fft_tdl_bit_fft_121_3 (
	data_in,
	global_clock_enable,
	tdl_arr_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	data_in;
input 	global_clock_enable;
output 	tdl_arr_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \tdl_arr[0] (
	.clk(clk),
	.d(data_in),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_0),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

endmodule

module fft256_asj_fft_tdl_bit_rst_fft_121_2 (
	global_clock_enable,
	tdl_arr_9,
	next_pass,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_9;
input 	next_pass;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0]~q ;
wire \tdl_arr~8_combout ;
wire \tdl_arr[1]~q ;
wire \tdl_arr~7_combout ;
wire \tdl_arr[2]~q ;
wire \tdl_arr~6_combout ;
wire \tdl_arr[3]~q ;
wire \tdl_arr~5_combout ;
wire \tdl_arr[4]~q ;
wire \tdl_arr~4_combout ;
wire \tdl_arr[5]~q ;
wire \tdl_arr~3_combout ;
wire \tdl_arr[6]~q ;
wire \tdl_arr~2_combout ;
wire \tdl_arr[7]~q ;
wire \tdl_arr~1_combout ;
wire \tdl_arr[8]~q ;
wire \tdl_arr~0_combout ;


dffeas \tdl_arr[9] (
	.clk(clk),
	.d(\tdl_arr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_9),
	.prn(vcc));
defparam \tdl_arr[9] .is_wysiwyg = "true";
defparam \tdl_arr[9] .power_up = "low";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(next_pass),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~8 (
	.dataa(reset_n),
	.datab(\tdl_arr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~8_combout ),
	.cout());
defparam \tdl_arr~8 .lut_mask = 16'hEEEE;
defparam \tdl_arr~8 .sum_lutc_input = "datac";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~7 (
	.dataa(reset_n),
	.datab(\tdl_arr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~7_combout ),
	.cout());
defparam \tdl_arr~7 .lut_mask = 16'hEEEE;
defparam \tdl_arr~7 .sum_lutc_input = "datac";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~6 (
	.dataa(reset_n),
	.datab(\tdl_arr[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~6_combout ),
	.cout());
defparam \tdl_arr~6 .lut_mask = 16'hEEEE;
defparam \tdl_arr~6 .sum_lutc_input = "datac";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~5 (
	.dataa(reset_n),
	.datab(\tdl_arr[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~5_combout ),
	.cout());
defparam \tdl_arr~5 .lut_mask = 16'hEEEE;
defparam \tdl_arr~5 .sum_lutc_input = "datac";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~4 (
	.dataa(reset_n),
	.datab(\tdl_arr[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~4_combout ),
	.cout());
defparam \tdl_arr~4 .lut_mask = 16'hEEEE;
defparam \tdl_arr~4 .sum_lutc_input = "datac";

dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5]~q ),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~3 (
	.dataa(reset_n),
	.datab(\tdl_arr[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~3_combout ),
	.cout());
defparam \tdl_arr~3 .lut_mask = 16'hEEEE;
defparam \tdl_arr~3 .sum_lutc_input = "datac";

dffeas \tdl_arr[6] (
	.clk(clk),
	.d(\tdl_arr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[6]~q ),
	.prn(vcc));
defparam \tdl_arr[6] .is_wysiwyg = "true";
defparam \tdl_arr[6] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~2 (
	.dataa(reset_n),
	.datab(\tdl_arr[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~2_combout ),
	.cout());
defparam \tdl_arr~2 .lut_mask = 16'hEEEE;
defparam \tdl_arr~2 .sum_lutc_input = "datac";

dffeas \tdl_arr[7] (
	.clk(clk),
	.d(\tdl_arr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[7]~q ),
	.prn(vcc));
defparam \tdl_arr[7] .is_wysiwyg = "true";
defparam \tdl_arr[7] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~1 (
	.dataa(reset_n),
	.datab(\tdl_arr[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~1_combout ),
	.cout());
defparam \tdl_arr~1 .lut_mask = 16'hEEEE;
defparam \tdl_arr~1 .sum_lutc_input = "datac";

dffeas \tdl_arr[8] (
	.clk(clk),
	.d(\tdl_arr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[8]~q ),
	.prn(vcc));
defparam \tdl_arr[8] .is_wysiwyg = "true";
defparam \tdl_arr[8] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~0 (
	.dataa(reset_n),
	.datab(\tdl_arr[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~0_combout ),
	.cout());
defparam \tdl_arr~0 .lut_mask = 16'hEEEE;
defparam \tdl_arr~0 .sum_lutc_input = "datac";

endmodule

module fft256_asj_fft_twadsogen_q_fft_121 (
	twad_tempo_0,
	twad_tempe_1,
	twad_tempe_2,
	twad_tempe_3,
	twad_tempe_4,
	twad_tempe_5,
	twad_tempo_1,
	twad_tempo_2,
	twad_tempo_3,
	twad_tempo_4,
	twad_tempo_5,
	k_count_tw_0,
	k_count_tw_2,
	k_count_tw_1,
	k_count_tw_3,
	k_count_tw_5,
	k_count_tw_4,
	k_count_tw_7,
	k_count_tw_6,
	global_clock_enable,
	quad_reg_2,
	quad_reg_0,
	quad_reg_1,
	p_tdl_0_10,
	p_tdl_1_10,
	p_tdl_2_10,
	data_addr_held_by1,
	data_addr_held_by2,
	clk)/* synthesis synthesis_greybox=1 */;
output 	twad_tempo_0;
output 	twad_tempe_1;
output 	twad_tempe_2;
output 	twad_tempe_3;
output 	twad_tempe_4;
output 	twad_tempe_5;
output 	twad_tempo_1;
output 	twad_tempo_2;
output 	twad_tempo_3;
output 	twad_tempo_4;
output 	twad_tempo_5;
input 	k_count_tw_0;
input 	k_count_tw_2;
input 	k_count_tw_1;
input 	k_count_tw_3;
input 	k_count_tw_5;
input 	k_count_tw_4;
input 	k_count_tw_7;
input 	k_count_tw_6;
input 	global_clock_enable;
output 	quad_reg_2;
output 	quad_reg_0;
output 	quad_reg_1;
input 	p_tdl_0_10;
input 	p_tdl_1_10;
input 	p_tdl_2_10;
output 	data_addr_held_by1;
output 	data_addr_held_by2;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add2~1 ;
wire \Add2~0_combout ;
wire \Add2~3 ;
wire \Add2~2_combout ;
wire \Add2~5 ;
wire \Add2~4_combout ;
wire \Add2~7 ;
wire \Add2~6_combout ;
wire \Add1~4_combout ;
wire \Add2~8_combout ;
wire \data_addr_held_by1[1]~q ;
wire \Mux1~0_combout ;
wire \data_addr_held_by1[3]~q ;
wire \data_addr_held_by1[2]~q ;
wire \Mux1~1_combout ;
wire \data_addr_held_by2[5]~q ;
wire \data_addr_held_by1[5]~q ;
wire \data_addr_held_by1[4]~q ;
wire \Mux5~0_combout ;
wire \Mux4~0_combout ;
wire \Mux3~0_combout ;
wire \Mux2~0_combout ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \data_addr_held_by1~1_combout ;
wire \data_addr_held_by1~2_combout ;
wire \data_addr_held_by1~3_combout ;
wire \data_addr_held_by2~4_combout ;
wire \data_addr_held_by1~4_combout ;
wire \data_addr_held_by1~5_combout ;
wire \data_addr_held_by1[0]~q ;
wire \Mux7~0_combout ;
wire \perm_addr[0]~q ;
wire \Mux7~1_combout ;
wire \data_addr_held_by2~5_combout ;
wire \data_addr_held_by2[4]~q ;
wire \data_addr_held_by2~2_combout ;
wire \data_addr_held_by2[3]~q ;
wire \data_addr_held_by2~3_combout ;
wire \data_addr_held_by2[2]~q ;
wire \data_addr_held_by2[1]~q ;
wire \data_addr_held_by2~1_combout ;
wire \data_addr_held_by2[0]~q ;
wire \Add1~1 ;
wire \Add1~3 ;
wire \Add1~5 ;
wire \Add1~7 ;
wire \Add1~9 ;
wire \Add1~10_combout ;
wire \Mux1~2_combout ;
wire \perm_addr[6]~q ;
wire \Add0~2_combout ;
wire \twad_tempo[0]~6_combout ;
wire \Add1~0_combout ;
wire \Mux6~2_combout ;
wire \perm_addr[1]~q ;
wire \twad_tempe[1]~5_combout ;
wire \Add1~2_combout ;
wire \Mux5~1_combout ;
wire \perm_addr[2]~q ;
wire \twad_tempe[1]~6 ;
wire \twad_tempe[2]~7_combout ;
wire \Mux4~1_combout ;
wire \perm_addr[3]~q ;
wire \twad_tempe[2]~8 ;
wire \twad_tempe[3]~9_combout ;
wire \Add1~6_combout ;
wire \Mux3~1_combout ;
wire \perm_addr[4]~q ;
wire \twad_tempe[3]~10 ;
wire \twad_tempe[4]~11_combout ;
wire \Add1~8_combout ;
wire \Mux2~1_combout ;
wire \perm_addr[5]~q ;
wire \twad_tempe[4]~12 ;
wire \twad_tempe[5]~13_combout ;
wire \twad_tempo[0]~7 ;
wire \twad_tempo[1]~8_combout ;
wire \twad_tempo[1]~9 ;
wire \twad_tempo[2]~10_combout ;
wire \twad_tempo[2]~11 ;
wire \twad_tempo[3]~12_combout ;
wire \twad_tempo[3]~13 ;
wire \twad_tempo[4]~14_combout ;
wire \twad_tempo[4]~15 ;
wire \twad_tempo[5]~16_combout ;
wire \Add1~11 ;
wire \Add1~12_combout ;
wire \Mux0~2_combout ;
wire \perm_addr[7]~q ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;


cycloneive_lcell_comb \Add2~0 (
	.dataa(\data_addr_held_by1[1]~q ),
	.datab(\data_addr_held_by2[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout(\Add2~1 ));
defparam \Add2~0 .lut_mask = 16'h66EE;
defparam \Add2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add2~2 (
	.dataa(\data_addr_held_by1[2]~q ),
	.datab(\data_addr_held_by2[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~1 ),
	.combout(\Add2~2_combout ),
	.cout(\Add2~3 ));
defparam \Add2~2 .lut_mask = 16'h967F;
defparam \Add2~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~4 (
	.dataa(\data_addr_held_by1[3]~q ),
	.datab(\data_addr_held_by2[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~3 ),
	.combout(\Add2~4_combout ),
	.cout(\Add2~5 ));
defparam \Add2~4 .lut_mask = 16'h96EF;
defparam \Add2~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~6 (
	.dataa(\data_addr_held_by2[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~5 ),
	.combout(\Add2~6_combout ),
	.cout(\Add2~7 ));
defparam \Add2~6 .lut_mask = 16'h5A5F;
defparam \Add2~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~4 (
	.dataa(\data_addr_held_by1[3]~q ),
	.datab(\data_addr_held_by2[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
defparam \Add1~4 .lut_mask = 16'h96EF;
defparam \Add1~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add2~7 ),
	.combout(\Add2~8_combout ),
	.cout());
defparam \Add2~8 .lut_mask = 16'h0F0F;
defparam \Add2~8 .sum_lutc_input = "cin";

dffeas \data_addr_held_by1[1] (
	.clk(clk),
	.d(\data_addr_held_by1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\data_addr_held_by1[1]~q ),
	.prn(vcc));
defparam \data_addr_held_by1[1] .is_wysiwyg = "true";
defparam \data_addr_held_by1[1] .power_up = "low";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(p_tdl_0_10),
	.datab(\data_addr_held_by2[1]~q ),
	.datac(\data_addr_held_by1[1]~q ),
	.datad(\data_addr_held_by2[0]~q ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hEBBE;
defparam \Mux1~0 .sum_lutc_input = "datac";

dffeas \data_addr_held_by1[3] (
	.clk(clk),
	.d(\data_addr_held_by1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\data_addr_held_by1[3]~q ),
	.prn(vcc));
defparam \data_addr_held_by1[3] .is_wysiwyg = "true";
defparam \data_addr_held_by1[3] .power_up = "low";

dffeas \data_addr_held_by1[2] (
	.clk(clk),
	.d(\data_addr_held_by1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\data_addr_held_by1[2]~q ),
	.prn(vcc));
defparam \data_addr_held_by1[2] .is_wysiwyg = "true";
defparam \data_addr_held_by1[2] .power_up = "low";

cycloneive_lcell_comb \Mux1~1 (
	.dataa(p_tdl_1_10),
	.datab(\Mux1~0_combout ),
	.datac(\Add2~6_combout ),
	.datad(p_tdl_0_10),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hFEFF;
defparam \Mux1~1 .sum_lutc_input = "datac";

dffeas \data_addr_held_by2[5] (
	.clk(clk),
	.d(\data_addr_held_by2~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\data_addr_held_by2[5]~q ),
	.prn(vcc));
defparam \data_addr_held_by2[5] .is_wysiwyg = "true";
defparam \data_addr_held_by2[5] .power_up = "low";

dffeas \data_addr_held_by1[5] (
	.clk(clk),
	.d(\data_addr_held_by1~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\data_addr_held_by1[5]~q ),
	.prn(vcc));
defparam \data_addr_held_by1[5] .is_wysiwyg = "true";
defparam \data_addr_held_by1[5] .power_up = "low";

dffeas \data_addr_held_by1[4] (
	.clk(clk),
	.d(\data_addr_held_by1~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\data_addr_held_by1[4]~q ),
	.prn(vcc));
defparam \data_addr_held_by1[4] .is_wysiwyg = "true";
defparam \data_addr_held_by1[4] .power_up = "low";

cycloneive_lcell_comb \Mux5~0 (
	.dataa(p_tdl_1_10),
	.datab(\data_addr_held_by1[0]~q ),
	.datac(gnd),
	.datad(p_tdl_0_10),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'hEEFF;
defparam \Mux5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~0 (
	.dataa(\Add2~0_combout ),
	.datab(\Add1~4_combout ),
	.datac(p_tdl_0_10),
	.datad(p_tdl_1_10),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'hEFFE;
defparam \Mux4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~0 (
	.dataa(p_tdl_1_10),
	.datab(\data_addr_held_by1[0]~q ),
	.datac(\Add2~2_combout ),
	.datad(p_tdl_0_10),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hFAFC;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~0 (
	.dataa(p_tdl_1_10),
	.datab(\Add1~0_combout ),
	.datac(\Add2~4_combout ),
	.datad(p_tdl_0_10),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFAFC;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(p_tdl_0_10),
	.datab(\data_addr_held_by2[1]~q ),
	.datac(\data_addr_held_by1[1]~q ),
	.datad(\data_addr_held_by2[0]~q ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hFFFE;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~1 (
	.dataa(p_tdl_1_10),
	.datab(\Mux0~0_combout ),
	.datac(\Add2~8_combout ),
	.datad(p_tdl_0_10),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hFEFF;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_addr_held_by1~1 (
	.dataa(k_count_tw_0),
	.datab(k_count_tw_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_addr_held_by1~1_combout ),
	.cout());
defparam \data_addr_held_by1~1 .lut_mask = 16'hEEEE;
defparam \data_addr_held_by1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_addr_held_by1~2 (
	.dataa(k_count_tw_0),
	.datab(k_count_tw_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_addr_held_by1~2_combout ),
	.cout());
defparam \data_addr_held_by1~2 .lut_mask = 16'hEEEE;
defparam \data_addr_held_by1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_addr_held_by1~3 (
	.dataa(k_count_tw_0),
	.datab(k_count_tw_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_addr_held_by1~3_combout ),
	.cout());
defparam \data_addr_held_by1~3 .lut_mask = 16'hEEEE;
defparam \data_addr_held_by1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_addr_held_by2~4 (
	.dataa(k_count_tw_1),
	.datab(k_count_tw_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_addr_held_by2~4_combout ),
	.cout());
defparam \data_addr_held_by2~4 .lut_mask = 16'hEEEE;
defparam \data_addr_held_by2~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_addr_held_by1~4 (
	.dataa(k_count_tw_0),
	.datab(k_count_tw_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_addr_held_by1~4_combout ),
	.cout());
defparam \data_addr_held_by1~4 .lut_mask = 16'hEEEE;
defparam \data_addr_held_by1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_addr_held_by1~5 (
	.dataa(k_count_tw_0),
	.datab(k_count_tw_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_addr_held_by1~5_combout ),
	.cout());
defparam \data_addr_held_by1~5 .lut_mask = 16'hEEEE;
defparam \data_addr_held_by1~5 .sum_lutc_input = "datac";

dffeas \twad_tempo[0] (
	.clk(clk),
	.d(\twad_tempo[0]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(twad_tempo_0),
	.prn(vcc));
defparam \twad_tempo[0] .is_wysiwyg = "true";
defparam \twad_tempo[0] .power_up = "low";

dffeas \twad_tempe[1] (
	.clk(clk),
	.d(\twad_tempe[1]~5_combout ),
	.asdata(\perm_addr[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\perm_addr[6]~q ),
	.ena(global_clock_enable),
	.q(twad_tempe_1),
	.prn(vcc));
defparam \twad_tempe[1] .is_wysiwyg = "true";
defparam \twad_tempe[1] .power_up = "low";

dffeas \twad_tempe[2] (
	.clk(clk),
	.d(\twad_tempe[2]~7_combout ),
	.asdata(\perm_addr[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\perm_addr[6]~q ),
	.ena(global_clock_enable),
	.q(twad_tempe_2),
	.prn(vcc));
defparam \twad_tempe[2] .is_wysiwyg = "true";
defparam \twad_tempe[2] .power_up = "low";

dffeas \twad_tempe[3] (
	.clk(clk),
	.d(\twad_tempe[3]~9_combout ),
	.asdata(\perm_addr[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\perm_addr[6]~q ),
	.ena(global_clock_enable),
	.q(twad_tempe_3),
	.prn(vcc));
defparam \twad_tempe[3] .is_wysiwyg = "true";
defparam \twad_tempe[3] .power_up = "low";

dffeas \twad_tempe[4] (
	.clk(clk),
	.d(\twad_tempe[4]~11_combout ),
	.asdata(\perm_addr[4]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\perm_addr[6]~q ),
	.ena(global_clock_enable),
	.q(twad_tempe_4),
	.prn(vcc));
defparam \twad_tempe[4] .is_wysiwyg = "true";
defparam \twad_tempe[4] .power_up = "low";

dffeas \twad_tempe[5] (
	.clk(clk),
	.d(\twad_tempe[5]~13_combout ),
	.asdata(\perm_addr[5]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\perm_addr[6]~q ),
	.ena(global_clock_enable),
	.q(twad_tempe_5),
	.prn(vcc));
defparam \twad_tempe[5] .is_wysiwyg = "true";
defparam \twad_tempe[5] .power_up = "low";

dffeas \twad_tempo[1] (
	.clk(clk),
	.d(\twad_tempo[1]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(twad_tempo_1),
	.prn(vcc));
defparam \twad_tempo[1] .is_wysiwyg = "true";
defparam \twad_tempo[1] .power_up = "low";

dffeas \twad_tempo[2] (
	.clk(clk),
	.d(\twad_tempo[2]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(twad_tempo_2),
	.prn(vcc));
defparam \twad_tempo[2] .is_wysiwyg = "true";
defparam \twad_tempo[2] .power_up = "low";

dffeas \twad_tempo[3] (
	.clk(clk),
	.d(\twad_tempo[3]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(twad_tempo_3),
	.prn(vcc));
defparam \twad_tempo[3] .is_wysiwyg = "true";
defparam \twad_tempo[3] .power_up = "low";

dffeas \twad_tempo[4] (
	.clk(clk),
	.d(\twad_tempo[4]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(twad_tempo_4),
	.prn(vcc));
defparam \twad_tempo[4] .is_wysiwyg = "true";
defparam \twad_tempo[4] .power_up = "low";

dffeas \twad_tempo[5] (
	.clk(clk),
	.d(\twad_tempo[5]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(twad_tempo_5),
	.prn(vcc));
defparam \twad_tempo[5] .is_wysiwyg = "true";
defparam \twad_tempo[5] .power_up = "low";

dffeas \quad_reg[2] (
	.clk(clk),
	.d(\perm_addr[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(quad_reg_2),
	.prn(vcc));
defparam \quad_reg[2] .is_wysiwyg = "true";
defparam \quad_reg[2] .power_up = "low";

dffeas \quad_reg[0] (
	.clk(clk),
	.d(\Equal0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(quad_reg_0),
	.prn(vcc));
defparam \quad_reg[0] .is_wysiwyg = "true";
defparam \quad_reg[0] .power_up = "low";

dffeas \quad_reg[1] (
	.clk(clk),
	.d(\perm_addr[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(quad_reg_1),
	.prn(vcc));
defparam \quad_reg[1] .is_wysiwyg = "true";
defparam \quad_reg[1] .power_up = "low";

cycloneive_lcell_comb \data_addr_held_by1~0 (
	.dataa(k_count_tw_0),
	.datab(k_count_tw_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(data_addr_held_by1),
	.cout());
defparam \data_addr_held_by1~0 .lut_mask = 16'hEEEE;
defparam \data_addr_held_by1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_addr_held_by2~0 (
	.dataa(k_count_tw_1),
	.datab(k_count_tw_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(data_addr_held_by2),
	.cout());
defparam \data_addr_held_by2~0 .lut_mask = 16'hEEEE;
defparam \data_addr_held_by2~0 .sum_lutc_input = "datac";

dffeas \data_addr_held_by1[0] (
	.clk(clk),
	.d(data_addr_held_by1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\data_addr_held_by1[0]~q ),
	.prn(vcc));
defparam \data_addr_held_by1[0] .is_wysiwyg = "true";
defparam \data_addr_held_by1[0] .power_up = "low";

cycloneive_lcell_comb \Mux7~0 (
	.dataa(p_tdl_0_10),
	.datab(\data_addr_held_by1[0]~q ),
	.datac(p_tdl_2_10),
	.datad(p_tdl_1_10),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'hEFFF;
defparam \Mux7~0 .sum_lutc_input = "datac";

dffeas \perm_addr[0] (
	.clk(clk),
	.d(\Mux7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\perm_addr[0]~q ),
	.prn(vcc));
defparam \perm_addr[0] .is_wysiwyg = "true";
defparam \perm_addr[0] .power_up = "low";

cycloneive_lcell_comb \Mux7~1 (
	.dataa(p_tdl_0_10),
	.datab(gnd),
	.datac(gnd),
	.datad(p_tdl_1_10),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
defparam \Mux7~1 .lut_mask = 16'hAAFF;
defparam \Mux7~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_addr_held_by2~5 (
	.dataa(k_count_tw_1),
	.datab(k_count_tw_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_addr_held_by2~5_combout ),
	.cout());
defparam \data_addr_held_by2~5 .lut_mask = 16'hEEEE;
defparam \data_addr_held_by2~5 .sum_lutc_input = "datac";

dffeas \data_addr_held_by2[4] (
	.clk(clk),
	.d(\data_addr_held_by2~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\data_addr_held_by2[4]~q ),
	.prn(vcc));
defparam \data_addr_held_by2[4] .is_wysiwyg = "true";
defparam \data_addr_held_by2[4] .power_up = "low";

cycloneive_lcell_comb \data_addr_held_by2~2 (
	.dataa(k_count_tw_1),
	.datab(k_count_tw_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_addr_held_by2~2_combout ),
	.cout());
defparam \data_addr_held_by2~2 .lut_mask = 16'hEEEE;
defparam \data_addr_held_by2~2 .sum_lutc_input = "datac";

dffeas \data_addr_held_by2[3] (
	.clk(clk),
	.d(\data_addr_held_by2~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\data_addr_held_by2[3]~q ),
	.prn(vcc));
defparam \data_addr_held_by2[3] .is_wysiwyg = "true";
defparam \data_addr_held_by2[3] .power_up = "low";

cycloneive_lcell_comb \data_addr_held_by2~3 (
	.dataa(k_count_tw_1),
	.datab(k_count_tw_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_addr_held_by2~3_combout ),
	.cout());
defparam \data_addr_held_by2~3 .lut_mask = 16'hEEEE;
defparam \data_addr_held_by2~3 .sum_lutc_input = "datac";

dffeas \data_addr_held_by2[2] (
	.clk(clk),
	.d(\data_addr_held_by2~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\data_addr_held_by2[2]~q ),
	.prn(vcc));
defparam \data_addr_held_by2[2] .is_wysiwyg = "true";
defparam \data_addr_held_by2[2] .power_up = "low";

dffeas \data_addr_held_by2[1] (
	.clk(clk),
	.d(data_addr_held_by2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\data_addr_held_by2[1]~q ),
	.prn(vcc));
defparam \data_addr_held_by2[1] .is_wysiwyg = "true";
defparam \data_addr_held_by2[1] .power_up = "low";

cycloneive_lcell_comb \data_addr_held_by2~1 (
	.dataa(k_count_tw_2),
	.datab(k_count_tw_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_addr_held_by2~1_combout ),
	.cout());
defparam \data_addr_held_by2~1 .lut_mask = 16'hEEEE;
defparam \data_addr_held_by2~1 .sum_lutc_input = "datac";

dffeas \data_addr_held_by2[0] (
	.clk(clk),
	.d(\data_addr_held_by2~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\data_addr_held_by2[0]~q ),
	.prn(vcc));
defparam \data_addr_held_by2[0] .is_wysiwyg = "true";
defparam \data_addr_held_by2[0] .power_up = "low";

cycloneive_lcell_comb \Add1~0 (
	.dataa(\data_addr_held_by1[1]~q ),
	.datab(\data_addr_held_by2[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
defparam \Add1~0 .lut_mask = 16'h66EE;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~2 (
	.dataa(\data_addr_held_by1[2]~q ),
	.datab(\data_addr_held_by2[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
defparam \Add1~2 .lut_mask = 16'h967F;
defparam \Add1~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~6 (
	.dataa(\data_addr_held_by1[4]~q ),
	.datab(\data_addr_held_by2[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
defparam \Add1~6 .lut_mask = 16'h967F;
defparam \Add1~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~8 (
	.dataa(\data_addr_held_by1[5]~q ),
	.datab(\data_addr_held_by2[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
defparam \Add1~8 .lut_mask = 16'h96EF;
defparam \Add1~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~10 (
	.dataa(\data_addr_held_by2[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout(\Add1~11 ));
defparam \Add1~10 .lut_mask = 16'h5A5F;
defparam \Add1~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mux1~2 (
	.dataa(\Mux1~1_combout ),
	.datab(\Mux7~1_combout ),
	.datac(\Add1~10_combout ),
	.datad(p_tdl_2_10),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
defparam \Mux1~2 .lut_mask = 16'hFEFF;
defparam \Mux1~2 .sum_lutc_input = "datac";

dffeas \perm_addr[6] (
	.clk(clk),
	.d(\Mux1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\perm_addr[6]~q ),
	.prn(vcc));
defparam \perm_addr[6] .is_wysiwyg = "true";
defparam \perm_addr[6] .power_up = "low";

cycloneive_lcell_comb \Add0~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\perm_addr[0]~q ),
	.datad(\perm_addr[6]~q ),
	.cin(gnd),
	.combout(\Add0~2_combout ),
	.cout());
defparam \Add0~2 .lut_mask = 16'h0FF0;
defparam \Add0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twad_tempo[0]~6 (
	.dataa(\Add0~2_combout ),
	.datab(\perm_addr[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\twad_tempo[0]~6_combout ),
	.cout(\twad_tempo[0]~7 ));
defparam \twad_tempo[0]~6 .lut_mask = 16'h6677;
defparam \twad_tempo[0]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~2 (
	.dataa(p_tdl_0_10),
	.datab(p_tdl_1_10),
	.datac(\Add1~0_combout ),
	.datad(p_tdl_2_10),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
defparam \Mux6~2 .lut_mask = 16'hFBFF;
defparam \Mux6~2 .sum_lutc_input = "datac";

dffeas \perm_addr[1] (
	.clk(clk),
	.d(\Mux6~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\perm_addr[1]~q ),
	.prn(vcc));
defparam \perm_addr[1] .is_wysiwyg = "true";
defparam \perm_addr[1] .power_up = "low";

cycloneive_lcell_comb \twad_tempe[1]~5 (
	.dataa(\perm_addr[1]~q ),
	.datab(\perm_addr[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\twad_tempe[1]~5_combout ),
	.cout(\twad_tempe[1]~6 ));
defparam \twad_tempe[1]~5 .lut_mask = 16'h6677;
defparam \twad_tempe[1]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~1 (
	.dataa(\Mux5~0_combout ),
	.datab(\Mux7~1_combout ),
	.datac(\Add1~2_combout ),
	.datad(p_tdl_2_10),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
defparam \Mux5~1 .lut_mask = 16'hFEFF;
defparam \Mux5~1 .sum_lutc_input = "datac";

dffeas \perm_addr[2] (
	.clk(clk),
	.d(\Mux5~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\perm_addr[2]~q ),
	.prn(vcc));
defparam \perm_addr[2] .is_wysiwyg = "true";
defparam \perm_addr[2] .power_up = "low";

cycloneive_lcell_comb \twad_tempe[2]~7 (
	.dataa(\perm_addr[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\twad_tempe[1]~6 ),
	.combout(\twad_tempe[2]~7_combout ),
	.cout(\twad_tempe[2]~8 ));
defparam \twad_tempe[2]~7 .lut_mask = 16'h5AAF;
defparam \twad_tempe[2]~7 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mux4~1 (
	.dataa(\Mux4~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(p_tdl_2_10),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
defparam \Mux4~1 .lut_mask = 16'hAAFF;
defparam \Mux4~1 .sum_lutc_input = "datac";

dffeas \perm_addr[3] (
	.clk(clk),
	.d(\Mux4~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\perm_addr[3]~q ),
	.prn(vcc));
defparam \perm_addr[3] .is_wysiwyg = "true";
defparam \perm_addr[3] .power_up = "low";

cycloneive_lcell_comb \twad_tempe[3]~9 (
	.dataa(\perm_addr[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\twad_tempe[2]~8 ),
	.combout(\twad_tempe[3]~9_combout ),
	.cout(\twad_tempe[3]~10 ));
defparam \twad_tempe[3]~9 .lut_mask = 16'h5A5F;
defparam \twad_tempe[3]~9 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mux3~1 (
	.dataa(\Mux3~0_combout ),
	.datab(\Mux7~1_combout ),
	.datac(\Add1~6_combout ),
	.datad(p_tdl_2_10),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
defparam \Mux3~1 .lut_mask = 16'hFEFF;
defparam \Mux3~1 .sum_lutc_input = "datac";

dffeas \perm_addr[4] (
	.clk(clk),
	.d(\Mux3~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\perm_addr[4]~q ),
	.prn(vcc));
defparam \perm_addr[4] .is_wysiwyg = "true";
defparam \perm_addr[4] .power_up = "low";

cycloneive_lcell_comb \twad_tempe[4]~11 (
	.dataa(\perm_addr[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\twad_tempe[3]~10 ),
	.combout(\twad_tempe[4]~11_combout ),
	.cout(\twad_tempe[4]~12 ));
defparam \twad_tempe[4]~11 .lut_mask = 16'h5AAF;
defparam \twad_tempe[4]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mux2~1 (
	.dataa(\Mux2~0_combout ),
	.datab(\Mux7~1_combout ),
	.datac(\Add1~8_combout ),
	.datad(p_tdl_2_10),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
defparam \Mux2~1 .lut_mask = 16'hFEFF;
defparam \Mux2~1 .sum_lutc_input = "datac";

dffeas \perm_addr[5] (
	.clk(clk),
	.d(\Mux2~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\perm_addr[5]~q ),
	.prn(vcc));
defparam \perm_addr[5] .is_wysiwyg = "true";
defparam \perm_addr[5] .power_up = "low";

cycloneive_lcell_comb \twad_tempe[5]~13 (
	.dataa(\perm_addr[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\twad_tempe[4]~12 ),
	.combout(\twad_tempe[5]~13_combout ),
	.cout());
defparam \twad_tempe[5]~13 .lut_mask = 16'h5A5A;
defparam \twad_tempe[5]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twad_tempo[1]~8 (
	.dataa(\perm_addr[1]~q ),
	.datab(\perm_addr[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\twad_tempo[0]~7 ),
	.combout(\twad_tempo[1]~8_combout ),
	.cout(\twad_tempo[1]~9 ));
defparam \twad_tempo[1]~8 .lut_mask = 16'h966F;
defparam \twad_tempo[1]~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twad_tempo[2]~10 (
	.dataa(\perm_addr[2]~q ),
	.datab(\perm_addr[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\twad_tempo[1]~9 ),
	.combout(\twad_tempo[2]~10_combout ),
	.cout(\twad_tempo[2]~11 ));
defparam \twad_tempo[2]~10 .lut_mask = 16'h966F;
defparam \twad_tempo[2]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twad_tempo[3]~12 (
	.dataa(\perm_addr[3]~q ),
	.datab(\perm_addr[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\twad_tempo[2]~11 ),
	.combout(\twad_tempo[3]~12_combout ),
	.cout(\twad_tempo[3]~13 ));
defparam \twad_tempo[3]~12 .lut_mask = 16'h966F;
defparam \twad_tempo[3]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twad_tempo[4]~14 (
	.dataa(\perm_addr[4]~q ),
	.datab(\perm_addr[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\twad_tempo[3]~13 ),
	.combout(\twad_tempo[4]~14_combout ),
	.cout(\twad_tempo[4]~15 ));
defparam \twad_tempo[4]~14 .lut_mask = 16'h966F;
defparam \twad_tempo[4]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twad_tempo[5]~16 (
	.dataa(\perm_addr[5]~q ),
	.datab(\perm_addr[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\twad_tempo[4]~15 ),
	.combout(\twad_tempo[5]~16_combout ),
	.cout());
defparam \twad_tempo[5]~16 .lut_mask = 16'h9696;
defparam \twad_tempo[5]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~11 ),
	.combout(\Add1~12_combout ),
	.cout());
defparam \Add1~12 .lut_mask = 16'h0F0F;
defparam \Add1~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mux0~2 (
	.dataa(\Mux0~1_combout ),
	.datab(\Mux7~1_combout ),
	.datac(\Add1~12_combout ),
	.datad(p_tdl_2_10),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
defparam \Mux0~2 .lut_mask = 16'hFEFF;
defparam \Mux0~2 .sum_lutc_input = "datac";

dffeas \perm_addr[7] (
	.clk(clk),
	.d(\Mux0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\perm_addr[7]~q ),
	.prn(vcc));
defparam \perm_addr[7] .is_wysiwyg = "true";
defparam \perm_addr[7] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\perm_addr[0]~q ),
	.datab(\perm_addr[1]~q ),
	.datac(\perm_addr[2]~q ),
	.datad(\perm_addr[3]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h7FFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\Equal0~0_combout ),
	.datab(gnd),
	.datac(\perm_addr[4]~q ),
	.datad(\perm_addr[5]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hAFFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

endmodule

module fft256_asj_fft_unbburst_sose_ctrl_fft_121 (
	q_b_0,
	q_b_16,
	q_b_1,
	q_b_17,
	q_b_2,
	q_b_18,
	q_b_3,
	q_b_19,
	q_b_4,
	q_b_20,
	q_b_5,
	q_b_21,
	q_b_6,
	q_b_22,
	q_b_7,
	q_b_23,
	q_b_8,
	q_b_24,
	q_b_9,
	q_b_25,
	q_b_10,
	q_b_26,
	q_b_11,
	q_b_27,
	q_b_12,
	q_b_28,
	q_b_13,
	q_b_29,
	q_b_14,
	q_b_30,
	q_b_15,
	q_b_31,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_31,
	global_clock_enable,
	a_ram_data_in_bus_0,
	wraddress_a_bus_0,
	wraddress_a_bus_1,
	wraddress_a_bus_2,
	wraddress_a_bus_3,
	wraddress_a_bus_4,
	wraddress_a_bus_5,
	wraddress_a_bus_6,
	wraddress_a_bus_7,
	rdaddress_a_bus_0,
	rdaddress_a_bus_1,
	rdaddress_a_bus_2,
	rdaddress_a_bus_3,
	rdaddress_a_bus_4,
	rdaddress_a_bus_5,
	rdaddress_a_bus_6,
	rdaddress_a_bus_7,
	a_ram_data_in_bus_16,
	a_ram_data_in_bus_1,
	a_ram_data_in_bus_17,
	a_ram_data_in_bus_2,
	a_ram_data_in_bus_18,
	a_ram_data_in_bus_3,
	a_ram_data_in_bus_19,
	a_ram_data_in_bus_4,
	a_ram_data_in_bus_20,
	a_ram_data_in_bus_5,
	a_ram_data_in_bus_21,
	a_ram_data_in_bus_6,
	a_ram_data_in_bus_22,
	a_ram_data_in_bus_7,
	a_ram_data_in_bus_23,
	a_ram_data_in_bus_8,
	a_ram_data_in_bus_24,
	a_ram_data_in_bus_9,
	a_ram_data_in_bus_25,
	a_ram_data_in_bus_10,
	a_ram_data_in_bus_26,
	a_ram_data_in_bus_11,
	a_ram_data_in_bus_27,
	a_ram_data_in_bus_12,
	a_ram_data_in_bus_28,
	a_ram_data_in_bus_13,
	a_ram_data_in_bus_29,
	a_ram_data_in_bus_14,
	a_ram_data_in_bus_30,
	a_ram_data_in_bus_15,
	a_ram_data_in_bus_31,
	data_rdy_vec_21,
	real_out_0,
	data_in_i_0,
	sel_ram_in,
	wraddress_a_bus_ctrl_i_0,
	wr_address_i_int_0,
	wraddress_a_bus_ctrl_i_1,
	wr_address_i_int_1,
	wraddress_a_bus_ctrl_i_2,
	wr_address_i_int_2,
	wraddress_a_bus_ctrl_i_3,
	wr_address_i_int_3,
	wraddress_a_bus_ctrl_i_4,
	wr_address_i_int_4,
	wraddress_a_bus_ctrl_i_5,
	wr_address_i_int_5,
	wraddress_a_bus_ctrl_i_6,
	wr_address_i_int_6,
	wraddress_a_bus_ctrl_i_7,
	wr_address_i_int_7,
	rd_addr_a_0,
	rd_addr_a_1,
	rd_addr_a_2,
	rd_addr_a_3,
	rd_addr_a_4,
	rd_addr_a_5,
	rd_addr_a_6,
	rd_addr_a_7,
	data_in_r_0,
	real_out_1,
	data_in_i_1,
	data_in_r_1,
	real_out_2,
	data_in_i_2,
	data_in_r_2,
	real_out_3,
	data_in_i_3,
	data_in_r_3,
	real_out_4,
	data_in_i_4,
	data_in_r_4,
	real_out_5,
	data_in_i_5,
	data_in_r_5,
	real_out_6,
	data_in_i_6,
	data_in_r_6,
	real_out_7,
	data_in_i_7,
	data_in_r_7,
	real_out_8,
	data_in_i_8,
	data_in_r_8,
	real_out_9,
	data_in_i_9,
	data_in_r_9,
	real_out_10,
	data_in_i_10,
	data_in_r_10,
	real_out_11,
	data_in_i_11,
	data_in_r_11,
	real_out_12,
	data_in_i_12,
	data_in_r_12,
	real_out_13,
	data_in_i_13,
	data_in_r_13,
	real_out_14,
	data_in_i_14,
	data_in_r_14,
	real_out_15,
	data_in_i_15,
	data_in_r_15,
	ram_data_out_0,
	ram_data_out_2,
	ram_data_out_1,
	ram_data_out_14,
	ram_data_out_12,
	ram_data_out_13,
	ram_data_out_15,
	ram_data_out_11,
	ram_data_out_10,
	ram_data_out_9,
	ram_data_out_8,
	ram_data_out_7,
	ram_data_out_6,
	ram_data_out_5,
	ram_data_out_4,
	ram_data_out_3,
	ram_data_out_16,
	ram_data_out_18,
	ram_data_out_17,
	ram_data_out_28,
	ram_data_out_29,
	ram_data_out_30,
	ram_data_out_31,
	ram_data_out_27,
	ram_data_out_26,
	ram_data_out_25,
	ram_data_out_24,
	ram_data_out_23,
	ram_data_out_22,
	ram_data_out_21,
	ram_data_out_20,
	ram_data_out_19,
	clk)/* synthesis synthesis_greybox=1 */;
input 	q_b_0;
input 	q_b_16;
input 	q_b_1;
input 	q_b_17;
input 	q_b_2;
input 	q_b_18;
input 	q_b_3;
input 	q_b_19;
input 	q_b_4;
input 	q_b_20;
input 	q_b_5;
input 	q_b_21;
input 	q_b_6;
input 	q_b_22;
input 	q_b_7;
input 	q_b_23;
input 	q_b_8;
input 	q_b_24;
input 	q_b_9;
input 	q_b_25;
input 	q_b_10;
input 	q_b_26;
input 	q_b_11;
input 	q_b_27;
input 	q_b_12;
input 	q_b_28;
input 	q_b_13;
input 	q_b_29;
input 	q_b_14;
input 	q_b_30;
input 	q_b_15;
input 	q_b_31;
input 	pipeline_dffe_16;
input 	pipeline_dffe_17;
input 	pipeline_dffe_18;
input 	pipeline_dffe_19;
input 	pipeline_dffe_20;
input 	pipeline_dffe_21;
input 	pipeline_dffe_22;
input 	pipeline_dffe_23;
input 	pipeline_dffe_24;
input 	pipeline_dffe_25;
input 	pipeline_dffe_26;
input 	pipeline_dffe_27;
input 	pipeline_dffe_28;
input 	pipeline_dffe_29;
input 	pipeline_dffe_30;
input 	pipeline_dffe_31;
input 	global_clock_enable;
output 	a_ram_data_in_bus_0;
output 	wraddress_a_bus_0;
output 	wraddress_a_bus_1;
output 	wraddress_a_bus_2;
output 	wraddress_a_bus_3;
output 	wraddress_a_bus_4;
output 	wraddress_a_bus_5;
output 	wraddress_a_bus_6;
output 	wraddress_a_bus_7;
output 	rdaddress_a_bus_0;
output 	rdaddress_a_bus_1;
output 	rdaddress_a_bus_2;
output 	rdaddress_a_bus_3;
output 	rdaddress_a_bus_4;
output 	rdaddress_a_bus_5;
output 	rdaddress_a_bus_6;
output 	rdaddress_a_bus_7;
output 	a_ram_data_in_bus_16;
output 	a_ram_data_in_bus_1;
output 	a_ram_data_in_bus_17;
output 	a_ram_data_in_bus_2;
output 	a_ram_data_in_bus_18;
output 	a_ram_data_in_bus_3;
output 	a_ram_data_in_bus_19;
output 	a_ram_data_in_bus_4;
output 	a_ram_data_in_bus_20;
output 	a_ram_data_in_bus_5;
output 	a_ram_data_in_bus_21;
output 	a_ram_data_in_bus_6;
output 	a_ram_data_in_bus_22;
output 	a_ram_data_in_bus_7;
output 	a_ram_data_in_bus_23;
output 	a_ram_data_in_bus_8;
output 	a_ram_data_in_bus_24;
output 	a_ram_data_in_bus_9;
output 	a_ram_data_in_bus_25;
output 	a_ram_data_in_bus_10;
output 	a_ram_data_in_bus_26;
output 	a_ram_data_in_bus_11;
output 	a_ram_data_in_bus_27;
output 	a_ram_data_in_bus_12;
output 	a_ram_data_in_bus_28;
output 	a_ram_data_in_bus_13;
output 	a_ram_data_in_bus_29;
output 	a_ram_data_in_bus_14;
output 	a_ram_data_in_bus_30;
output 	a_ram_data_in_bus_15;
output 	a_ram_data_in_bus_31;
input 	data_rdy_vec_21;
input 	real_out_0;
input 	data_in_i_0;
input 	sel_ram_in;
input 	wraddress_a_bus_ctrl_i_0;
input 	wr_address_i_int_0;
input 	wraddress_a_bus_ctrl_i_1;
input 	wr_address_i_int_1;
input 	wraddress_a_bus_ctrl_i_2;
input 	wr_address_i_int_2;
input 	wraddress_a_bus_ctrl_i_3;
input 	wr_address_i_int_3;
input 	wraddress_a_bus_ctrl_i_4;
input 	wr_address_i_int_4;
input 	wraddress_a_bus_ctrl_i_5;
input 	wr_address_i_int_5;
input 	wraddress_a_bus_ctrl_i_6;
input 	wr_address_i_int_6;
input 	wraddress_a_bus_ctrl_i_7;
input 	wr_address_i_int_7;
input 	rd_addr_a_0;
input 	rd_addr_a_1;
input 	rd_addr_a_2;
input 	rd_addr_a_3;
input 	rd_addr_a_4;
input 	rd_addr_a_5;
input 	rd_addr_a_6;
input 	rd_addr_a_7;
input 	data_in_r_0;
input 	real_out_1;
input 	data_in_i_1;
input 	data_in_r_1;
input 	real_out_2;
input 	data_in_i_2;
input 	data_in_r_2;
input 	real_out_3;
input 	data_in_i_3;
input 	data_in_r_3;
input 	real_out_4;
input 	data_in_i_4;
input 	data_in_r_4;
input 	real_out_5;
input 	data_in_i_5;
input 	data_in_r_5;
input 	real_out_6;
input 	data_in_i_6;
input 	data_in_r_6;
input 	real_out_7;
input 	data_in_i_7;
input 	data_in_r_7;
input 	real_out_8;
input 	data_in_i_8;
input 	data_in_r_8;
input 	real_out_9;
input 	data_in_i_9;
input 	data_in_r_9;
input 	real_out_10;
input 	data_in_i_10;
input 	data_in_r_10;
input 	real_out_11;
input 	data_in_i_11;
input 	data_in_r_11;
input 	real_out_12;
input 	data_in_i_12;
input 	data_in_r_12;
input 	real_out_13;
input 	data_in_i_13;
input 	data_in_r_13;
input 	real_out_14;
input 	data_in_i_14;
input 	data_in_r_14;
input 	real_out_15;
input 	data_in_i_15;
input 	data_in_r_15;
output 	ram_data_out_0;
output 	ram_data_out_2;
output 	ram_data_out_1;
output 	ram_data_out_14;
output 	ram_data_out_12;
output 	ram_data_out_13;
output 	ram_data_out_15;
output 	ram_data_out_11;
output 	ram_data_out_10;
output 	ram_data_out_9;
output 	ram_data_out_8;
output 	ram_data_out_7;
output 	ram_data_out_6;
output 	ram_data_out_5;
output 	ram_data_out_4;
output 	ram_data_out_3;
output 	ram_data_out_16;
output 	ram_data_out_18;
output 	ram_data_out_17;
output 	ram_data_out_28;
output 	ram_data_out_29;
output 	ram_data_out_30;
output 	ram_data_out_31;
output 	ram_data_out_27;
output 	ram_data_out_26;
output 	ram_data_out_25;
output 	ram_data_out_24;
output 	ram_data_out_23;
output 	ram_data_out_22;
output 	ram_data_out_21;
output 	ram_data_out_20;
output 	ram_data_out_19;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a_ram_data_in_bus~0_combout ;
wire \wraddress_a_bus~0_combout ;
wire \wraddress_a_bus~1_combout ;
wire \wraddress_a_bus~2_combout ;
wire \wraddress_a_bus~3_combout ;
wire \wraddress_a_bus~4_combout ;
wire \wraddress_a_bus~5_combout ;
wire \wraddress_a_bus~6_combout ;
wire \wraddress_a_bus~7_combout ;
wire \a_ram_data_in_bus~1_combout ;
wire \a_ram_data_in_bus~2_combout ;
wire \a_ram_data_in_bus~3_combout ;
wire \a_ram_data_in_bus~4_combout ;
wire \a_ram_data_in_bus~5_combout ;
wire \a_ram_data_in_bus~6_combout ;
wire \a_ram_data_in_bus~7_combout ;
wire \a_ram_data_in_bus~8_combout ;
wire \a_ram_data_in_bus~9_combout ;
wire \a_ram_data_in_bus~10_combout ;
wire \a_ram_data_in_bus~11_combout ;
wire \a_ram_data_in_bus~12_combout ;
wire \a_ram_data_in_bus~13_combout ;
wire \a_ram_data_in_bus~14_combout ;
wire \a_ram_data_in_bus~15_combout ;
wire \a_ram_data_in_bus~16_combout ;
wire \a_ram_data_in_bus~17_combout ;
wire \a_ram_data_in_bus~18_combout ;
wire \a_ram_data_in_bus~19_combout ;
wire \a_ram_data_in_bus~20_combout ;
wire \a_ram_data_in_bus~21_combout ;
wire \a_ram_data_in_bus~22_combout ;
wire \a_ram_data_in_bus~23_combout ;
wire \a_ram_data_in_bus~24_combout ;
wire \a_ram_data_in_bus~25_combout ;
wire \a_ram_data_in_bus~26_combout ;
wire \a_ram_data_in_bus~27_combout ;
wire \a_ram_data_in_bus~28_combout ;
wire \a_ram_data_in_bus~29_combout ;
wire \a_ram_data_in_bus~30_combout ;
wire \a_ram_data_in_bus~31_combout ;


dffeas \a_ram_data_in_bus[0] (
	.clk(clk),
	.d(\a_ram_data_in_bus~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_0),
	.prn(vcc));
defparam \a_ram_data_in_bus[0] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[0] .power_up = "low";

dffeas \wraddress_a_bus[0] (
	.clk(clk),
	.d(\wraddress_a_bus~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_0),
	.prn(vcc));
defparam \wraddress_a_bus[0] .is_wysiwyg = "true";
defparam \wraddress_a_bus[0] .power_up = "low";

dffeas \wraddress_a_bus[1] (
	.clk(clk),
	.d(\wraddress_a_bus~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_1),
	.prn(vcc));
defparam \wraddress_a_bus[1] .is_wysiwyg = "true";
defparam \wraddress_a_bus[1] .power_up = "low";

dffeas \wraddress_a_bus[2] (
	.clk(clk),
	.d(\wraddress_a_bus~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_2),
	.prn(vcc));
defparam \wraddress_a_bus[2] .is_wysiwyg = "true";
defparam \wraddress_a_bus[2] .power_up = "low";

dffeas \wraddress_a_bus[3] (
	.clk(clk),
	.d(\wraddress_a_bus~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_3),
	.prn(vcc));
defparam \wraddress_a_bus[3] .is_wysiwyg = "true";
defparam \wraddress_a_bus[3] .power_up = "low";

dffeas \wraddress_a_bus[4] (
	.clk(clk),
	.d(\wraddress_a_bus~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_4),
	.prn(vcc));
defparam \wraddress_a_bus[4] .is_wysiwyg = "true";
defparam \wraddress_a_bus[4] .power_up = "low";

dffeas \wraddress_a_bus[5] (
	.clk(clk),
	.d(\wraddress_a_bus~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_5),
	.prn(vcc));
defparam \wraddress_a_bus[5] .is_wysiwyg = "true";
defparam \wraddress_a_bus[5] .power_up = "low";

dffeas \wraddress_a_bus[6] (
	.clk(clk),
	.d(\wraddress_a_bus~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_6),
	.prn(vcc));
defparam \wraddress_a_bus[6] .is_wysiwyg = "true";
defparam \wraddress_a_bus[6] .power_up = "low";

dffeas \wraddress_a_bus[7] (
	.clk(clk),
	.d(\wraddress_a_bus~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_7),
	.prn(vcc));
defparam \wraddress_a_bus[7] .is_wysiwyg = "true";
defparam \wraddress_a_bus[7] .power_up = "low";

dffeas \rdaddress_a_bus[0] (
	.clk(clk),
	.d(rd_addr_a_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_0),
	.prn(vcc));
defparam \rdaddress_a_bus[0] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[0] .power_up = "low";

dffeas \rdaddress_a_bus[1] (
	.clk(clk),
	.d(rd_addr_a_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_1),
	.prn(vcc));
defparam \rdaddress_a_bus[1] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[1] .power_up = "low";

dffeas \rdaddress_a_bus[2] (
	.clk(clk),
	.d(rd_addr_a_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_2),
	.prn(vcc));
defparam \rdaddress_a_bus[2] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[2] .power_up = "low";

dffeas \rdaddress_a_bus[3] (
	.clk(clk),
	.d(rd_addr_a_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_3),
	.prn(vcc));
defparam \rdaddress_a_bus[3] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[3] .power_up = "low";

dffeas \rdaddress_a_bus[4] (
	.clk(clk),
	.d(rd_addr_a_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_4),
	.prn(vcc));
defparam \rdaddress_a_bus[4] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[4] .power_up = "low";

dffeas \rdaddress_a_bus[5] (
	.clk(clk),
	.d(rd_addr_a_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_5),
	.prn(vcc));
defparam \rdaddress_a_bus[5] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[5] .power_up = "low";

dffeas \rdaddress_a_bus[6] (
	.clk(clk),
	.d(rd_addr_a_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_6),
	.prn(vcc));
defparam \rdaddress_a_bus[6] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[6] .power_up = "low";

dffeas \rdaddress_a_bus[7] (
	.clk(clk),
	.d(rd_addr_a_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_7),
	.prn(vcc));
defparam \rdaddress_a_bus[7] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[7] .power_up = "low";

dffeas \a_ram_data_in_bus[16] (
	.clk(clk),
	.d(\a_ram_data_in_bus~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_16),
	.prn(vcc));
defparam \a_ram_data_in_bus[16] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[16] .power_up = "low";

dffeas \a_ram_data_in_bus[1] (
	.clk(clk),
	.d(\a_ram_data_in_bus~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_1),
	.prn(vcc));
defparam \a_ram_data_in_bus[1] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[1] .power_up = "low";

dffeas \a_ram_data_in_bus[17] (
	.clk(clk),
	.d(\a_ram_data_in_bus~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_17),
	.prn(vcc));
defparam \a_ram_data_in_bus[17] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[17] .power_up = "low";

dffeas \a_ram_data_in_bus[2] (
	.clk(clk),
	.d(\a_ram_data_in_bus~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_2),
	.prn(vcc));
defparam \a_ram_data_in_bus[2] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[2] .power_up = "low";

dffeas \a_ram_data_in_bus[18] (
	.clk(clk),
	.d(\a_ram_data_in_bus~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_18),
	.prn(vcc));
defparam \a_ram_data_in_bus[18] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[18] .power_up = "low";

dffeas \a_ram_data_in_bus[3] (
	.clk(clk),
	.d(\a_ram_data_in_bus~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_3),
	.prn(vcc));
defparam \a_ram_data_in_bus[3] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[3] .power_up = "low";

dffeas \a_ram_data_in_bus[19] (
	.clk(clk),
	.d(\a_ram_data_in_bus~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_19),
	.prn(vcc));
defparam \a_ram_data_in_bus[19] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[19] .power_up = "low";

dffeas \a_ram_data_in_bus[4] (
	.clk(clk),
	.d(\a_ram_data_in_bus~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_4),
	.prn(vcc));
defparam \a_ram_data_in_bus[4] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[4] .power_up = "low";

dffeas \a_ram_data_in_bus[20] (
	.clk(clk),
	.d(\a_ram_data_in_bus~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_20),
	.prn(vcc));
defparam \a_ram_data_in_bus[20] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[20] .power_up = "low";

dffeas \a_ram_data_in_bus[5] (
	.clk(clk),
	.d(\a_ram_data_in_bus~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_5),
	.prn(vcc));
defparam \a_ram_data_in_bus[5] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[5] .power_up = "low";

dffeas \a_ram_data_in_bus[21] (
	.clk(clk),
	.d(\a_ram_data_in_bus~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_21),
	.prn(vcc));
defparam \a_ram_data_in_bus[21] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[21] .power_up = "low";

dffeas \a_ram_data_in_bus[6] (
	.clk(clk),
	.d(\a_ram_data_in_bus~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_6),
	.prn(vcc));
defparam \a_ram_data_in_bus[6] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[6] .power_up = "low";

dffeas \a_ram_data_in_bus[22] (
	.clk(clk),
	.d(\a_ram_data_in_bus~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_22),
	.prn(vcc));
defparam \a_ram_data_in_bus[22] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[22] .power_up = "low";

dffeas \a_ram_data_in_bus[7] (
	.clk(clk),
	.d(\a_ram_data_in_bus~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_7),
	.prn(vcc));
defparam \a_ram_data_in_bus[7] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[7] .power_up = "low";

dffeas \a_ram_data_in_bus[23] (
	.clk(clk),
	.d(\a_ram_data_in_bus~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_23),
	.prn(vcc));
defparam \a_ram_data_in_bus[23] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[23] .power_up = "low";

dffeas \a_ram_data_in_bus[8] (
	.clk(clk),
	.d(\a_ram_data_in_bus~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_8),
	.prn(vcc));
defparam \a_ram_data_in_bus[8] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[8] .power_up = "low";

dffeas \a_ram_data_in_bus[24] (
	.clk(clk),
	.d(\a_ram_data_in_bus~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_24),
	.prn(vcc));
defparam \a_ram_data_in_bus[24] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[24] .power_up = "low";

dffeas \a_ram_data_in_bus[9] (
	.clk(clk),
	.d(\a_ram_data_in_bus~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_9),
	.prn(vcc));
defparam \a_ram_data_in_bus[9] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[9] .power_up = "low";

dffeas \a_ram_data_in_bus[25] (
	.clk(clk),
	.d(\a_ram_data_in_bus~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_25),
	.prn(vcc));
defparam \a_ram_data_in_bus[25] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[25] .power_up = "low";

dffeas \a_ram_data_in_bus[10] (
	.clk(clk),
	.d(\a_ram_data_in_bus~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_10),
	.prn(vcc));
defparam \a_ram_data_in_bus[10] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[10] .power_up = "low";

dffeas \a_ram_data_in_bus[26] (
	.clk(clk),
	.d(\a_ram_data_in_bus~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_26),
	.prn(vcc));
defparam \a_ram_data_in_bus[26] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[26] .power_up = "low";

dffeas \a_ram_data_in_bus[11] (
	.clk(clk),
	.d(\a_ram_data_in_bus~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_11),
	.prn(vcc));
defparam \a_ram_data_in_bus[11] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[11] .power_up = "low";

dffeas \a_ram_data_in_bus[27] (
	.clk(clk),
	.d(\a_ram_data_in_bus~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_27),
	.prn(vcc));
defparam \a_ram_data_in_bus[27] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[27] .power_up = "low";

dffeas \a_ram_data_in_bus[12] (
	.clk(clk),
	.d(\a_ram_data_in_bus~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_12),
	.prn(vcc));
defparam \a_ram_data_in_bus[12] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[12] .power_up = "low";

dffeas \a_ram_data_in_bus[28] (
	.clk(clk),
	.d(\a_ram_data_in_bus~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_28),
	.prn(vcc));
defparam \a_ram_data_in_bus[28] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[28] .power_up = "low";

dffeas \a_ram_data_in_bus[13] (
	.clk(clk),
	.d(\a_ram_data_in_bus~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_13),
	.prn(vcc));
defparam \a_ram_data_in_bus[13] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[13] .power_up = "low";

dffeas \a_ram_data_in_bus[29] (
	.clk(clk),
	.d(\a_ram_data_in_bus~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_29),
	.prn(vcc));
defparam \a_ram_data_in_bus[29] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[29] .power_up = "low";

dffeas \a_ram_data_in_bus[14] (
	.clk(clk),
	.d(\a_ram_data_in_bus~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_14),
	.prn(vcc));
defparam \a_ram_data_in_bus[14] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[14] .power_up = "low";

dffeas \a_ram_data_in_bus[30] (
	.clk(clk),
	.d(\a_ram_data_in_bus~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_30),
	.prn(vcc));
defparam \a_ram_data_in_bus[30] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[30] .power_up = "low";

dffeas \a_ram_data_in_bus[15] (
	.clk(clk),
	.d(\a_ram_data_in_bus~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_15),
	.prn(vcc));
defparam \a_ram_data_in_bus[15] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[15] .power_up = "low";

dffeas \a_ram_data_in_bus[31] (
	.clk(clk),
	.d(\a_ram_data_in_bus~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_31),
	.prn(vcc));
defparam \a_ram_data_in_bus[31] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[31] .power_up = "low";

dffeas \ram_data_out[0] (
	.clk(clk),
	.d(q_b_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_0),
	.prn(vcc));
defparam \ram_data_out[0] .is_wysiwyg = "true";
defparam \ram_data_out[0] .power_up = "low";

dffeas \ram_data_out[2] (
	.clk(clk),
	.d(q_b_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_2),
	.prn(vcc));
defparam \ram_data_out[2] .is_wysiwyg = "true";
defparam \ram_data_out[2] .power_up = "low";

dffeas \ram_data_out[1] (
	.clk(clk),
	.d(q_b_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_1),
	.prn(vcc));
defparam \ram_data_out[1] .is_wysiwyg = "true";
defparam \ram_data_out[1] .power_up = "low";

dffeas \ram_data_out[14] (
	.clk(clk),
	.d(q_b_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_14),
	.prn(vcc));
defparam \ram_data_out[14] .is_wysiwyg = "true";
defparam \ram_data_out[14] .power_up = "low";

dffeas \ram_data_out[12] (
	.clk(clk),
	.d(q_b_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_12),
	.prn(vcc));
defparam \ram_data_out[12] .is_wysiwyg = "true";
defparam \ram_data_out[12] .power_up = "low";

dffeas \ram_data_out[13] (
	.clk(clk),
	.d(q_b_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_13),
	.prn(vcc));
defparam \ram_data_out[13] .is_wysiwyg = "true";
defparam \ram_data_out[13] .power_up = "low";

dffeas \ram_data_out[15] (
	.clk(clk),
	.d(q_b_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_15),
	.prn(vcc));
defparam \ram_data_out[15] .is_wysiwyg = "true";
defparam \ram_data_out[15] .power_up = "low";

dffeas \ram_data_out[11] (
	.clk(clk),
	.d(q_b_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_11),
	.prn(vcc));
defparam \ram_data_out[11] .is_wysiwyg = "true";
defparam \ram_data_out[11] .power_up = "low";

dffeas \ram_data_out[10] (
	.clk(clk),
	.d(q_b_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_10),
	.prn(vcc));
defparam \ram_data_out[10] .is_wysiwyg = "true";
defparam \ram_data_out[10] .power_up = "low";

dffeas \ram_data_out[9] (
	.clk(clk),
	.d(q_b_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_9),
	.prn(vcc));
defparam \ram_data_out[9] .is_wysiwyg = "true";
defparam \ram_data_out[9] .power_up = "low";

dffeas \ram_data_out[8] (
	.clk(clk),
	.d(q_b_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_8),
	.prn(vcc));
defparam \ram_data_out[8] .is_wysiwyg = "true";
defparam \ram_data_out[8] .power_up = "low";

dffeas \ram_data_out[7] (
	.clk(clk),
	.d(q_b_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_7),
	.prn(vcc));
defparam \ram_data_out[7] .is_wysiwyg = "true";
defparam \ram_data_out[7] .power_up = "low";

dffeas \ram_data_out[6] (
	.clk(clk),
	.d(q_b_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_6),
	.prn(vcc));
defparam \ram_data_out[6] .is_wysiwyg = "true";
defparam \ram_data_out[6] .power_up = "low";

dffeas \ram_data_out[5] (
	.clk(clk),
	.d(q_b_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_5),
	.prn(vcc));
defparam \ram_data_out[5] .is_wysiwyg = "true";
defparam \ram_data_out[5] .power_up = "low";

dffeas \ram_data_out[4] (
	.clk(clk),
	.d(q_b_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_4),
	.prn(vcc));
defparam \ram_data_out[4] .is_wysiwyg = "true";
defparam \ram_data_out[4] .power_up = "low";

dffeas \ram_data_out[3] (
	.clk(clk),
	.d(q_b_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_3),
	.prn(vcc));
defparam \ram_data_out[3] .is_wysiwyg = "true";
defparam \ram_data_out[3] .power_up = "low";

dffeas \ram_data_out[16] (
	.clk(clk),
	.d(q_b_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_16),
	.prn(vcc));
defparam \ram_data_out[16] .is_wysiwyg = "true";
defparam \ram_data_out[16] .power_up = "low";

dffeas \ram_data_out[18] (
	.clk(clk),
	.d(q_b_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_18),
	.prn(vcc));
defparam \ram_data_out[18] .is_wysiwyg = "true";
defparam \ram_data_out[18] .power_up = "low";

dffeas \ram_data_out[17] (
	.clk(clk),
	.d(q_b_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_17),
	.prn(vcc));
defparam \ram_data_out[17] .is_wysiwyg = "true";
defparam \ram_data_out[17] .power_up = "low";

dffeas \ram_data_out[28] (
	.clk(clk),
	.d(q_b_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_28),
	.prn(vcc));
defparam \ram_data_out[28] .is_wysiwyg = "true";
defparam \ram_data_out[28] .power_up = "low";

dffeas \ram_data_out[29] (
	.clk(clk),
	.d(q_b_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_29),
	.prn(vcc));
defparam \ram_data_out[29] .is_wysiwyg = "true";
defparam \ram_data_out[29] .power_up = "low";

dffeas \ram_data_out[30] (
	.clk(clk),
	.d(q_b_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_30),
	.prn(vcc));
defparam \ram_data_out[30] .is_wysiwyg = "true";
defparam \ram_data_out[30] .power_up = "low";

dffeas \ram_data_out[31] (
	.clk(clk),
	.d(q_b_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_31),
	.prn(vcc));
defparam \ram_data_out[31] .is_wysiwyg = "true";
defparam \ram_data_out[31] .power_up = "low";

dffeas \ram_data_out[27] (
	.clk(clk),
	.d(q_b_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_27),
	.prn(vcc));
defparam \ram_data_out[27] .is_wysiwyg = "true";
defparam \ram_data_out[27] .power_up = "low";

dffeas \ram_data_out[26] (
	.clk(clk),
	.d(q_b_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_26),
	.prn(vcc));
defparam \ram_data_out[26] .is_wysiwyg = "true";
defparam \ram_data_out[26] .power_up = "low";

dffeas \ram_data_out[25] (
	.clk(clk),
	.d(q_b_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_25),
	.prn(vcc));
defparam \ram_data_out[25] .is_wysiwyg = "true";
defparam \ram_data_out[25] .power_up = "low";

dffeas \ram_data_out[24] (
	.clk(clk),
	.d(q_b_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_24),
	.prn(vcc));
defparam \ram_data_out[24] .is_wysiwyg = "true";
defparam \ram_data_out[24] .power_up = "low";

dffeas \ram_data_out[23] (
	.clk(clk),
	.d(q_b_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_23),
	.prn(vcc));
defparam \ram_data_out[23] .is_wysiwyg = "true";
defparam \ram_data_out[23] .power_up = "low";

dffeas \ram_data_out[22] (
	.clk(clk),
	.d(q_b_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_22),
	.prn(vcc));
defparam \ram_data_out[22] .is_wysiwyg = "true";
defparam \ram_data_out[22] .power_up = "low";

dffeas \ram_data_out[21] (
	.clk(clk),
	.d(q_b_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_21),
	.prn(vcc));
defparam \ram_data_out[21] .is_wysiwyg = "true";
defparam \ram_data_out[21] .power_up = "low";

dffeas \ram_data_out[20] (
	.clk(clk),
	.d(q_b_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_20),
	.prn(vcc));
defparam \ram_data_out[20] .is_wysiwyg = "true";
defparam \ram_data_out[20] .power_up = "low";

dffeas \ram_data_out[19] (
	.clk(clk),
	.d(q_b_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out_19),
	.prn(vcc));
defparam \ram_data_out[19] .is_wysiwyg = "true";
defparam \ram_data_out[19] .power_up = "low";

cycloneive_lcell_comb \a_ram_data_in_bus~0 (
	.dataa(real_out_0),
	.datab(data_in_i_0),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~0_combout ),
	.cout());
defparam \a_ram_data_in_bus~0 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~0 (
	.dataa(wraddress_a_bus_ctrl_i_0),
	.datab(wr_address_i_int_0),
	.datac(gnd),
	.datad(data_rdy_vec_21),
	.cin(gnd),
	.combout(\wraddress_a_bus~0_combout ),
	.cout());
defparam \wraddress_a_bus~0 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~1 (
	.dataa(wraddress_a_bus_ctrl_i_1),
	.datab(wr_address_i_int_1),
	.datac(gnd),
	.datad(data_rdy_vec_21),
	.cin(gnd),
	.combout(\wraddress_a_bus~1_combout ),
	.cout());
defparam \wraddress_a_bus~1 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~2 (
	.dataa(wraddress_a_bus_ctrl_i_2),
	.datab(wr_address_i_int_2),
	.datac(gnd),
	.datad(data_rdy_vec_21),
	.cin(gnd),
	.combout(\wraddress_a_bus~2_combout ),
	.cout());
defparam \wraddress_a_bus~2 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~3 (
	.dataa(wraddress_a_bus_ctrl_i_3),
	.datab(wr_address_i_int_3),
	.datac(gnd),
	.datad(data_rdy_vec_21),
	.cin(gnd),
	.combout(\wraddress_a_bus~3_combout ),
	.cout());
defparam \wraddress_a_bus~3 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~4 (
	.dataa(wraddress_a_bus_ctrl_i_4),
	.datab(wr_address_i_int_4),
	.datac(gnd),
	.datad(data_rdy_vec_21),
	.cin(gnd),
	.combout(\wraddress_a_bus~4_combout ),
	.cout());
defparam \wraddress_a_bus~4 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~5 (
	.dataa(wraddress_a_bus_ctrl_i_5),
	.datab(wr_address_i_int_5),
	.datac(gnd),
	.datad(data_rdy_vec_21),
	.cin(gnd),
	.combout(\wraddress_a_bus~5_combout ),
	.cout());
defparam \wraddress_a_bus~5 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~6 (
	.dataa(wraddress_a_bus_ctrl_i_6),
	.datab(wr_address_i_int_6),
	.datac(gnd),
	.datad(data_rdy_vec_21),
	.cin(gnd),
	.combout(\wraddress_a_bus~6_combout ),
	.cout());
defparam \wraddress_a_bus~6 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~7 (
	.dataa(wraddress_a_bus_ctrl_i_7),
	.datab(wr_address_i_int_7),
	.datac(gnd),
	.datad(data_rdy_vec_21),
	.cin(gnd),
	.combout(\wraddress_a_bus~7_combout ),
	.cout());
defparam \wraddress_a_bus~7 .lut_mask = 16'hAACC;
defparam \wraddress_a_bus~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~1 (
	.dataa(pipeline_dffe_16),
	.datab(data_in_r_0),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~1_combout ),
	.cout());
defparam \a_ram_data_in_bus~1 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~2 (
	.dataa(real_out_1),
	.datab(data_in_i_1),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~2_combout ),
	.cout());
defparam \a_ram_data_in_bus~2 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~3 (
	.dataa(pipeline_dffe_17),
	.datab(data_in_r_1),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~3_combout ),
	.cout());
defparam \a_ram_data_in_bus~3 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~4 (
	.dataa(real_out_2),
	.datab(data_in_i_2),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~4_combout ),
	.cout());
defparam \a_ram_data_in_bus~4 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~5 (
	.dataa(pipeline_dffe_18),
	.datab(data_in_r_2),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~5_combout ),
	.cout());
defparam \a_ram_data_in_bus~5 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~6 (
	.dataa(real_out_3),
	.datab(data_in_i_3),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~6_combout ),
	.cout());
defparam \a_ram_data_in_bus~6 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~7 (
	.dataa(pipeline_dffe_19),
	.datab(data_in_r_3),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~7_combout ),
	.cout());
defparam \a_ram_data_in_bus~7 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~8 (
	.dataa(real_out_4),
	.datab(data_in_i_4),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~8_combout ),
	.cout());
defparam \a_ram_data_in_bus~8 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~9 (
	.dataa(pipeline_dffe_20),
	.datab(data_in_r_4),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~9_combout ),
	.cout());
defparam \a_ram_data_in_bus~9 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~10 (
	.dataa(real_out_5),
	.datab(data_in_i_5),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~10_combout ),
	.cout());
defparam \a_ram_data_in_bus~10 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~11 (
	.dataa(pipeline_dffe_21),
	.datab(data_in_r_5),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~11_combout ),
	.cout());
defparam \a_ram_data_in_bus~11 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~12 (
	.dataa(real_out_6),
	.datab(data_in_i_6),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~12_combout ),
	.cout());
defparam \a_ram_data_in_bus~12 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~13 (
	.dataa(pipeline_dffe_22),
	.datab(data_in_r_6),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~13_combout ),
	.cout());
defparam \a_ram_data_in_bus~13 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~14 (
	.dataa(real_out_7),
	.datab(data_in_i_7),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~14_combout ),
	.cout());
defparam \a_ram_data_in_bus~14 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~15 (
	.dataa(pipeline_dffe_23),
	.datab(data_in_r_7),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~15_combout ),
	.cout());
defparam \a_ram_data_in_bus~15 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~16 (
	.dataa(real_out_8),
	.datab(data_in_i_8),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~16_combout ),
	.cout());
defparam \a_ram_data_in_bus~16 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~17 (
	.dataa(pipeline_dffe_24),
	.datab(data_in_r_8),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~17_combout ),
	.cout());
defparam \a_ram_data_in_bus~17 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~18 (
	.dataa(real_out_9),
	.datab(data_in_i_9),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~18_combout ),
	.cout());
defparam \a_ram_data_in_bus~18 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~19 (
	.dataa(pipeline_dffe_25),
	.datab(data_in_r_9),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~19_combout ),
	.cout());
defparam \a_ram_data_in_bus~19 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~20 (
	.dataa(real_out_10),
	.datab(data_in_i_10),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~20_combout ),
	.cout());
defparam \a_ram_data_in_bus~20 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~21 (
	.dataa(pipeline_dffe_26),
	.datab(data_in_r_10),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~21_combout ),
	.cout());
defparam \a_ram_data_in_bus~21 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~22 (
	.dataa(real_out_11),
	.datab(data_in_i_11),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~22_combout ),
	.cout());
defparam \a_ram_data_in_bus~22 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~23 (
	.dataa(pipeline_dffe_27),
	.datab(data_in_r_11),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~23_combout ),
	.cout());
defparam \a_ram_data_in_bus~23 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~24 (
	.dataa(real_out_12),
	.datab(data_in_i_12),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~24_combout ),
	.cout());
defparam \a_ram_data_in_bus~24 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~25 (
	.dataa(pipeline_dffe_28),
	.datab(data_in_r_12),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~25_combout ),
	.cout());
defparam \a_ram_data_in_bus~25 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~26 (
	.dataa(real_out_13),
	.datab(data_in_i_13),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~26_combout ),
	.cout());
defparam \a_ram_data_in_bus~26 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~27 (
	.dataa(pipeline_dffe_29),
	.datab(data_in_r_13),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~27_combout ),
	.cout());
defparam \a_ram_data_in_bus~27 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~28 (
	.dataa(real_out_14),
	.datab(data_in_i_14),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~28_combout ),
	.cout());
defparam \a_ram_data_in_bus~28 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~29 (
	.dataa(pipeline_dffe_30),
	.datab(data_in_r_14),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~29_combout ),
	.cout());
defparam \a_ram_data_in_bus~29 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~30 (
	.dataa(real_out_15),
	.datab(data_in_i_15),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~30_combout ),
	.cout());
defparam \a_ram_data_in_bus~30 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~31 (
	.dataa(pipeline_dffe_31),
	.datab(data_in_r_15),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~31_combout ),
	.cout());
defparam \a_ram_data_in_bus~31 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~31 .sum_lutc_input = "datac";

endmodule

module fft256_auk_dspip_avalon_streaming_controller_fft_121 (
	master_sink_ena,
	source_packet_error_0,
	source_packet_error_1,
	source_stall_reg1,
	sink_stall_reg1,
	sink_ready_ctrl,
	sink_start,
	empty_dff,
	sink_stall,
	packet_error_s_0,
	packet_error_s_1,
	stall_reg1,
	Mux0,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	master_sink_ena;
output 	source_packet_error_0;
output 	source_packet_error_1;
output 	source_stall_reg1;
output 	sink_stall_reg1;
output 	sink_ready_ctrl;
input 	sink_start;
input 	empty_dff;
input 	sink_stall;
input 	packet_error_s_0;
input 	packet_error_s_1;
output 	stall_reg1;
input 	Mux0;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \source_stall_reg~0_combout ;
wire \sink_stall_reg~0_combout ;
wire \stall_int~combout ;


dffeas \source_packet_error[0] (
	.clk(clk),
	.d(packet_error_s_0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(source_packet_error_0),
	.prn(vcc));
defparam \source_packet_error[0] .is_wysiwyg = "true";
defparam \source_packet_error[0] .power_up = "low";

dffeas \source_packet_error[1] (
	.clk(clk),
	.d(packet_error_s_1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(source_packet_error_1),
	.prn(vcc));
defparam \source_packet_error[1] .is_wysiwyg = "true";
defparam \source_packet_error[1] .power_up = "low";

dffeas source_stall_reg(
	.clk(clk),
	.d(\source_stall_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(source_stall_reg1),
	.prn(vcc));
defparam source_stall_reg.is_wysiwyg = "true";
defparam source_stall_reg.power_up = "low";

dffeas sink_stall_reg(
	.clk(clk),
	.d(\sink_stall_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sink_stall_reg1),
	.prn(vcc));
defparam sink_stall_reg.is_wysiwyg = "true";
defparam sink_stall_reg.power_up = "low";

cycloneive_lcell_comb \sink_ready_ctrl~0 (
	.dataa(master_sink_ena),
	.datab(source_stall_reg1),
	.datac(gnd),
	.datad(sink_stall_reg1),
	.cin(gnd),
	.combout(sink_ready_ctrl),
	.cout());
defparam \sink_ready_ctrl~0 .lut_mask = 16'hEEFF;
defparam \sink_ready_ctrl~0 .sum_lutc_input = "datac";

dffeas stall_reg(
	.clk(clk),
	.d(\stall_int~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stall_reg1),
	.prn(vcc));
defparam stall_reg.is_wysiwyg = "true";
defparam stall_reg.power_up = "low";

cycloneive_lcell_comb \source_stall_reg~0 (
	.dataa(Mux0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\source_stall_reg~0_combout ),
	.cout());
defparam \source_stall_reg~0 .lut_mask = 16'h5555;
defparam \source_stall_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_stall_reg~0 (
	.dataa(sink_stall),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sink_stall_reg~0_combout ),
	.cout());
defparam \sink_stall_reg~0 .lut_mask = 16'h5555;
defparam \sink_stall_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb stall_int(
	.dataa(sink_start),
	.datab(empty_dff),
	.datac(Mux0),
	.datad(gnd),
	.cin(gnd),
	.combout(\stall_int~combout ),
	.cout());
defparam stall_int.lut_mask = 16'hEFEF;
defparam stall_int.sum_lutc_input = "datac";

endmodule

module fft256_auk_dspip_avalon_streaming_sink_fft_121 (
	master_sink_ena,
	q_b_16,
	q_b_0,
	q_b_17,
	q_b_1,
	q_b_18,
	q_b_2,
	q_b_19,
	q_b_3,
	q_b_20,
	q_b_4,
	q_b_21,
	q_b_5,
	q_b_22,
	q_b_6,
	q_b_23,
	q_b_7,
	q_b_24,
	q_b_8,
	q_b_25,
	q_b_9,
	q_b_26,
	q_b_10,
	q_b_27,
	q_b_11,
	q_b_28,
	q_b_12,
	q_b_29,
	q_b_13,
	q_b_30,
	q_b_14,
	q_b_31,
	q_b_15,
	at_sink_ready_s1,
	source_stall_reg,
	sink_stall_reg,
	sink_ready_ctrl,
	sink_start1,
	empty_dff,
	sink_stall1,
	packet_error_s_0,
	packet_error_s_1,
	send_sop_s1,
	send_eop_s1,
	clk,
	reset_n,
	sink_valid,
	sink_sop,
	sink_eop,
	sink_error_0,
	sink_error_1,
	at_sink_data)/* synthesis synthesis_greybox=1 */;
input 	master_sink_ena;
output 	q_b_16;
output 	q_b_0;
output 	q_b_17;
output 	q_b_1;
output 	q_b_18;
output 	q_b_2;
output 	q_b_19;
output 	q_b_3;
output 	q_b_20;
output 	q_b_4;
output 	q_b_21;
output 	q_b_5;
output 	q_b_22;
output 	q_b_6;
output 	q_b_23;
output 	q_b_7;
output 	q_b_24;
output 	q_b_8;
output 	q_b_25;
output 	q_b_9;
output 	q_b_26;
output 	q_b_10;
output 	q_b_27;
output 	q_b_11;
output 	q_b_28;
output 	q_b_12;
output 	q_b_29;
output 	q_b_13;
output 	q_b_30;
output 	q_b_14;
output 	q_b_31;
output 	q_b_15;
output 	at_sink_ready_s1;
input 	source_stall_reg;
input 	sink_stall_reg;
input 	sink_ready_ctrl;
output 	sink_start1;
output 	empty_dff;
output 	sink_stall1;
output 	packet_error_s_0;
output 	packet_error_s_1;
output 	send_sop_s1;
output 	send_eop_s1;
input 	clk;
input 	reset_n;
input 	sink_valid;
input 	sink_sop;
input 	sink_eop;
input 	sink_error_0;
input 	sink_error_1;
input 	[31:0] at_sink_data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \out_cnt[0]~q ;
wire \out_cnt[4]~q ;
wire \count[1]~q ;
wire \count[2]~q ;
wire \count[3]~q ;
wire \count[0]~q ;
wire \count[4]~q ;
wire \out_cnt[0]~8_combout ;
wire \out_cnt[4]~16_combout ;
wire \count[0]~8_combout ;
wire \count[1]~10_combout ;
wire \count[2]~14_combout ;
wire \count[3]~16_combout ;
wire \count[4]~18_combout ;
wire \normal_fifo:fifo_eab_on:in_fifo|auto_generated|dffe_af~q ;
wire \normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \Selector3~1_combout ;
wire \Selector3~2_combout ;
wire \max_reached~0_combout ;
wire \LessThan0~0_combout ;
wire \at_sink_data_int[16]~q ;
wire \at_sink_data_int[0]~q ;
wire \at_sink_data_int[17]~q ;
wire \at_sink_data_int[1]~q ;
wire \at_sink_data_int[18]~q ;
wire \at_sink_data_int[2]~q ;
wire \at_sink_data_int[19]~q ;
wire \at_sink_data_int[3]~q ;
wire \at_sink_data_int[20]~q ;
wire \at_sink_data_int[4]~q ;
wire \at_sink_data_int[21]~q ;
wire \at_sink_data_int[5]~q ;
wire \at_sink_data_int[22]~q ;
wire \at_sink_data_int[6]~q ;
wire \at_sink_data_int[23]~q ;
wire \at_sink_data_int[7]~q ;
wire \at_sink_data_int[24]~q ;
wire \at_sink_data_int[8]~q ;
wire \at_sink_data_int[25]~q ;
wire \at_sink_data_int[9]~q ;
wire \at_sink_data_int[26]~q ;
wire \at_sink_data_int[10]~q ;
wire \at_sink_data_int[27]~q ;
wire \at_sink_data_int[11]~q ;
wire \at_sink_data_int[28]~q ;
wire \at_sink_data_int[12]~q ;
wire \at_sink_data_int[29]~q ;
wire \at_sink_data_int[13]~q ;
wire \at_sink_data_int[30]~q ;
wire \at_sink_data_int[14]~q ;
wire \at_sink_data_int[31]~q ;
wire \at_sink_data_int[15]~q ;
wire \data_take~combout ;
wire \fifo_wrreq~0_wirecell_combout ;
wire \at_sink_ready_s~0_combout ;
wire \sink_start~0_combout ;
wire \count[0]~9 ;
wire \count[1]~11 ;
wire \count[2]~15 ;
wire \count[3]~17 ;
wire \count[4]~19 ;
wire \count[5]~20_combout ;
wire \sink_comb_update_2~2_combout ;
wire \Selector4~0_combout ;
wire \sink_state.end1~q ;
wire \sink_state.st_err~q ;
wire \Selector5~0_combout ;
wire \Selector3~3_combout ;
wire \Selector2~2_combout ;
wire \Selector1~2_combout ;
wire \Selector1~3_combout ;
wire \sink_state.stall~q ;
wire \Selector4~1_combout ;
wire \Selector3~4_combout ;
wire \Selector2~5_combout ;
wire \Selector3~5_combout ;
wire \count[0]~12_combout ;
wire \sink_comb_update_2~0_combout ;
wire \Selector0~0_combout ;
wire \Selector0~1_combout ;
wire \sink_state.start~q ;
wire \Selector2~3_combout ;
wire \sink_comb_update_2~1_combout ;
wire \Selector2~4_combout ;
wire \data_take~2_combout ;
wire \count[0]~13_combout ;
wire \count[5]~q ;
wire \count[5]~21 ;
wire \count[6]~22_combout ;
wire \count[6]~q ;
wire \count[6]~23 ;
wire \count[7]~24_combout ;
wire \count[7]~q ;
wire \max_reached~1_combout ;
wire \max_reached~2_combout ;
wire \max_reached~3_combout ;
wire \max_reached~q ;
wire \sink_comb_update_2~3_combout ;
wire \Selector6~0_combout ;
wire \Selector6~1_combout ;
wire \Selector3~0_combout ;
wire \Selector6~2_combout ;
wire \Selector6~3_combout ;
wire \Selector6~4_combout ;
wire \Selector2~6_combout ;
wire \sink_state.run1~q ;
wire \fifo_wrreq~0_combout ;
wire \Selector5~1_combout ;
wire \Selector5~2_combout ;
wire \sink_comb_update_2~4_combout ;
wire \Selector5~3_combout ;
wire \out_cnt[0]~9 ;
wire \out_cnt[1]~10_combout ;
wire \out_cnt[1]~11 ;
wire \out_cnt[2]~13 ;
wire \out_cnt[3]~15 ;
wire \out_cnt[4]~17 ;
wire \out_cnt[5]~18_combout ;
wire \sink_stall_s~q ;
wire \Selector8~0_combout ;
wire \sink_out_state.normal~q ;
wire \Selector7~0_combout ;
wire \out_cnt[5]~q ;
wire \out_cnt[5]~19 ;
wire \out_cnt[6]~20_combout ;
wire \out_cnt[6]~q ;
wire \out_cnt[6]~21 ;
wire \out_cnt[7]~22_combout ;
wire \out_cnt[7]~q ;
wire \LessThan0~1_combout ;
wire \LessThan0~2_combout ;
wire \out_cnt[1]~q ;
wire \out_cnt[2]~12_combout ;
wire \out_cnt[2]~q ;
wire \out_cnt[3]~14_combout ;
wire \out_cnt[3]~q ;
wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \Equal1~2_combout ;
wire \Selector10~0_combout ;
wire \Selector10~1_combout ;
wire \sink_out_state.empty_and_ready~q ;
wire \send_sop_eop_p~0_combout ;


fft256_scfifo_1 \normal_fifo:fifo_eab_on:in_fifo (
	.q({q_unconnected_wire_33,q_unconnected_wire_32,q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.dffe_af(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dffe_af~q ),
	.empty_dff(empty_dff),
	.rdreq(\Selector7~0_combout ),
	.sink_staterun1(\sink_state.run1~q ),
	.sink_stateend1(\sink_state.end1~q ),
	.wrreq(\fifo_wrreq~0_combout ),
	.counter_reg_bit_0(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.data({gnd,gnd,\at_sink_data_int[31]~q ,\at_sink_data_int[30]~q ,\at_sink_data_int[29]~q ,\at_sink_data_int[28]~q ,\at_sink_data_int[27]~q ,\at_sink_data_int[26]~q ,\at_sink_data_int[25]~q ,\at_sink_data_int[24]~q ,\at_sink_data_int[23]~q ,\at_sink_data_int[22]~q ,
\at_sink_data_int[21]~q ,\at_sink_data_int[20]~q ,\at_sink_data_int[19]~q ,\at_sink_data_int[18]~q ,\at_sink_data_int[17]~q ,\at_sink_data_int[16]~q ,\at_sink_data_int[15]~q ,\at_sink_data_int[14]~q ,\at_sink_data_int[13]~q ,\at_sink_data_int[12]~q ,
\at_sink_data_int[11]~q ,\at_sink_data_int[10]~q ,\at_sink_data_int[9]~q ,\at_sink_data_int[8]~q ,\at_sink_data_int[7]~q ,\at_sink_data_int[6]~q ,\at_sink_data_int[5]~q ,\at_sink_data_int[4]~q ,\at_sink_data_int[3]~q ,\at_sink_data_int[2]~q ,\at_sink_data_int[1]~q ,
\at_sink_data_int[0]~q }),
	.fifo_wrreq(\fifo_wrreq~0_wirecell_combout ),
	.clock(clk),
	.reset_n(reset_n));

dffeas \out_cnt[0] (
	.clk(clk),
	.d(\out_cnt[0]~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[0]~q ),
	.prn(vcc));
defparam \out_cnt[0] .is_wysiwyg = "true";
defparam \out_cnt[0] .power_up = "low";

dffeas \out_cnt[4] (
	.clk(clk),
	.d(\out_cnt[4]~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[4]~q ),
	.prn(vcc));
defparam \out_cnt[4] .is_wysiwyg = "true";
defparam \out_cnt[4] .power_up = "low";

dffeas \count[1] (
	.clk(clk),
	.d(\count[1]~10_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[0]~12_combout ),
	.sload(gnd),
	.ena(\count[0]~13_combout ),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

dffeas \count[2] (
	.clk(clk),
	.d(\count[2]~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[0]~12_combout ),
	.sload(gnd),
	.ena(\count[0]~13_combout ),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

dffeas \count[3] (
	.clk(clk),
	.d(\count[3]~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[0]~12_combout ),
	.sload(gnd),
	.ena(\count[0]~13_combout ),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

dffeas \count[0] (
	.clk(clk),
	.d(\count[0]~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[0]~12_combout ),
	.sload(gnd),
	.ena(\count[0]~13_combout ),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

dffeas \count[4] (
	.clk(clk),
	.d(\count[4]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[0]~12_combout ),
	.sload(gnd),
	.ena(\count[0]~13_combout ),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

cycloneive_lcell_comb \out_cnt[0]~8 (
	.dataa(\out_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\out_cnt[0]~8_combout ),
	.cout(\out_cnt[0]~9 ));
defparam \out_cnt[0]~8 .lut_mask = 16'h55AA;
defparam \out_cnt[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_cnt[4]~16 (
	.dataa(\out_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[3]~15 ),
	.combout(\out_cnt[4]~16_combout ),
	.cout(\out_cnt[4]~17 ));
defparam \out_cnt[4]~16 .lut_mask = 16'h5AAF;
defparam \out_cnt[4]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \count[0]~8 (
	.dataa(\count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\count[0]~8_combout ),
	.cout(\count[0]~9 ));
defparam \count[0]~8 .lut_mask = 16'h55AA;
defparam \count[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[1]~10 (
	.dataa(\count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[0]~9 ),
	.combout(\count[1]~10_combout ),
	.cout(\count[1]~11 ));
defparam \count[1]~10 .lut_mask = 16'h5A5F;
defparam \count[1]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \count[2]~14 (
	.dataa(\count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[1]~11 ),
	.combout(\count[2]~14_combout ),
	.cout(\count[2]~15 ));
defparam \count[2]~14 .lut_mask = 16'h5AAF;
defparam \count[2]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \count[3]~16 (
	.dataa(\count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[2]~15 ),
	.combout(\count[3]~16_combout ),
	.cout(\count[3]~17 ));
defparam \count[3]~16 .lut_mask = 16'h5A5F;
defparam \count[3]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \count[4]~18 (
	.dataa(\count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[3]~17 ),
	.combout(\count[4]~18_combout ),
	.cout(\count[4]~19 ));
defparam \count[4]~18 .lut_mask = 16'h5AAF;
defparam \count[4]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Selector3~1 (
	.dataa(sink_valid),
	.datab(at_sink_ready_s1),
	.datac(\max_reached~q ),
	.datad(sink_eop),
	.cin(gnd),
	.combout(\Selector3~1_combout ),
	.cout());
defparam \Selector3~1 .lut_mask = 16'h6996;
defparam \Selector3~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~2 (
	.dataa(\sink_state.stall~q ),
	.datab(\sink_state.run1~q ),
	.datac(\Selector3~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector3~2_combout ),
	.cout());
defparam \Selector3~2 .lut_mask = 16'hFEFE;
defparam \Selector3~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \max_reached~0 (
	.dataa(\count[1]~q ),
	.datab(\count[2]~q ),
	.datac(\count[3]~q ),
	.datad(\count[0]~q ),
	.cin(gnd),
	.combout(\max_reached~0_combout ),
	.cout());
defparam \max_reached~0 .lut_mask = 16'hFEFF;
defparam \max_reached~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \LessThan0~0 (
	.dataa(\out_cnt[0]~q ),
	.datab(\out_cnt[1]~q ),
	.datac(\out_cnt[2]~q ),
	.datad(\out_cnt[3]~q ),
	.cin(gnd),
	.combout(\LessThan0~0_combout ),
	.cout());
defparam \LessThan0~0 .lut_mask = 16'h7FFF;
defparam \LessThan0~0 .sum_lutc_input = "datac";

dffeas \at_sink_data_int[16] (
	.clk(clk),
	.d(at_sink_data[16]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[16]~q ),
	.prn(vcc));
defparam \at_sink_data_int[16] .is_wysiwyg = "true";
defparam \at_sink_data_int[16] .power_up = "low";

dffeas \at_sink_data_int[0] (
	.clk(clk),
	.d(at_sink_data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[0]~q ),
	.prn(vcc));
defparam \at_sink_data_int[0] .is_wysiwyg = "true";
defparam \at_sink_data_int[0] .power_up = "low";

dffeas \at_sink_data_int[17] (
	.clk(clk),
	.d(at_sink_data[17]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[17]~q ),
	.prn(vcc));
defparam \at_sink_data_int[17] .is_wysiwyg = "true";
defparam \at_sink_data_int[17] .power_up = "low";

dffeas \at_sink_data_int[1] (
	.clk(clk),
	.d(at_sink_data[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[1]~q ),
	.prn(vcc));
defparam \at_sink_data_int[1] .is_wysiwyg = "true";
defparam \at_sink_data_int[1] .power_up = "low";

dffeas \at_sink_data_int[18] (
	.clk(clk),
	.d(at_sink_data[18]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[18]~q ),
	.prn(vcc));
defparam \at_sink_data_int[18] .is_wysiwyg = "true";
defparam \at_sink_data_int[18] .power_up = "low";

dffeas \at_sink_data_int[2] (
	.clk(clk),
	.d(at_sink_data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[2]~q ),
	.prn(vcc));
defparam \at_sink_data_int[2] .is_wysiwyg = "true";
defparam \at_sink_data_int[2] .power_up = "low";

dffeas \at_sink_data_int[19] (
	.clk(clk),
	.d(at_sink_data[19]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[19]~q ),
	.prn(vcc));
defparam \at_sink_data_int[19] .is_wysiwyg = "true";
defparam \at_sink_data_int[19] .power_up = "low";

dffeas \at_sink_data_int[3] (
	.clk(clk),
	.d(at_sink_data[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[3]~q ),
	.prn(vcc));
defparam \at_sink_data_int[3] .is_wysiwyg = "true";
defparam \at_sink_data_int[3] .power_up = "low";

dffeas \at_sink_data_int[20] (
	.clk(clk),
	.d(at_sink_data[20]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[20]~q ),
	.prn(vcc));
defparam \at_sink_data_int[20] .is_wysiwyg = "true";
defparam \at_sink_data_int[20] .power_up = "low";

dffeas \at_sink_data_int[4] (
	.clk(clk),
	.d(at_sink_data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[4]~q ),
	.prn(vcc));
defparam \at_sink_data_int[4] .is_wysiwyg = "true";
defparam \at_sink_data_int[4] .power_up = "low";

dffeas \at_sink_data_int[21] (
	.clk(clk),
	.d(at_sink_data[21]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[21]~q ),
	.prn(vcc));
defparam \at_sink_data_int[21] .is_wysiwyg = "true";
defparam \at_sink_data_int[21] .power_up = "low";

dffeas \at_sink_data_int[5] (
	.clk(clk),
	.d(at_sink_data[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[5]~q ),
	.prn(vcc));
defparam \at_sink_data_int[5] .is_wysiwyg = "true";
defparam \at_sink_data_int[5] .power_up = "low";

dffeas \at_sink_data_int[22] (
	.clk(clk),
	.d(at_sink_data[22]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[22]~q ),
	.prn(vcc));
defparam \at_sink_data_int[22] .is_wysiwyg = "true";
defparam \at_sink_data_int[22] .power_up = "low";

dffeas \at_sink_data_int[6] (
	.clk(clk),
	.d(at_sink_data[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[6]~q ),
	.prn(vcc));
defparam \at_sink_data_int[6] .is_wysiwyg = "true";
defparam \at_sink_data_int[6] .power_up = "low";

dffeas \at_sink_data_int[23] (
	.clk(clk),
	.d(at_sink_data[23]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[23]~q ),
	.prn(vcc));
defparam \at_sink_data_int[23] .is_wysiwyg = "true";
defparam \at_sink_data_int[23] .power_up = "low";

dffeas \at_sink_data_int[7] (
	.clk(clk),
	.d(at_sink_data[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[7]~q ),
	.prn(vcc));
defparam \at_sink_data_int[7] .is_wysiwyg = "true";
defparam \at_sink_data_int[7] .power_up = "low";

dffeas \at_sink_data_int[24] (
	.clk(clk),
	.d(at_sink_data[24]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[24]~q ),
	.prn(vcc));
defparam \at_sink_data_int[24] .is_wysiwyg = "true";
defparam \at_sink_data_int[24] .power_up = "low";

dffeas \at_sink_data_int[8] (
	.clk(clk),
	.d(at_sink_data[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[8]~q ),
	.prn(vcc));
defparam \at_sink_data_int[8] .is_wysiwyg = "true";
defparam \at_sink_data_int[8] .power_up = "low";

dffeas \at_sink_data_int[25] (
	.clk(clk),
	.d(at_sink_data[25]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[25]~q ),
	.prn(vcc));
defparam \at_sink_data_int[25] .is_wysiwyg = "true";
defparam \at_sink_data_int[25] .power_up = "low";

dffeas \at_sink_data_int[9] (
	.clk(clk),
	.d(at_sink_data[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[9]~q ),
	.prn(vcc));
defparam \at_sink_data_int[9] .is_wysiwyg = "true";
defparam \at_sink_data_int[9] .power_up = "low";

dffeas \at_sink_data_int[26] (
	.clk(clk),
	.d(at_sink_data[26]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[26]~q ),
	.prn(vcc));
defparam \at_sink_data_int[26] .is_wysiwyg = "true";
defparam \at_sink_data_int[26] .power_up = "low";

dffeas \at_sink_data_int[10] (
	.clk(clk),
	.d(at_sink_data[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[10]~q ),
	.prn(vcc));
defparam \at_sink_data_int[10] .is_wysiwyg = "true";
defparam \at_sink_data_int[10] .power_up = "low";

dffeas \at_sink_data_int[27] (
	.clk(clk),
	.d(at_sink_data[27]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[27]~q ),
	.prn(vcc));
defparam \at_sink_data_int[27] .is_wysiwyg = "true";
defparam \at_sink_data_int[27] .power_up = "low";

dffeas \at_sink_data_int[11] (
	.clk(clk),
	.d(at_sink_data[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[11]~q ),
	.prn(vcc));
defparam \at_sink_data_int[11] .is_wysiwyg = "true";
defparam \at_sink_data_int[11] .power_up = "low";

dffeas \at_sink_data_int[28] (
	.clk(clk),
	.d(at_sink_data[28]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[28]~q ),
	.prn(vcc));
defparam \at_sink_data_int[28] .is_wysiwyg = "true";
defparam \at_sink_data_int[28] .power_up = "low";

dffeas \at_sink_data_int[12] (
	.clk(clk),
	.d(at_sink_data[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[12]~q ),
	.prn(vcc));
defparam \at_sink_data_int[12] .is_wysiwyg = "true";
defparam \at_sink_data_int[12] .power_up = "low";

dffeas \at_sink_data_int[29] (
	.clk(clk),
	.d(at_sink_data[29]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[29]~q ),
	.prn(vcc));
defparam \at_sink_data_int[29] .is_wysiwyg = "true";
defparam \at_sink_data_int[29] .power_up = "low";

dffeas \at_sink_data_int[13] (
	.clk(clk),
	.d(at_sink_data[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[13]~q ),
	.prn(vcc));
defparam \at_sink_data_int[13] .is_wysiwyg = "true";
defparam \at_sink_data_int[13] .power_up = "low";

dffeas \at_sink_data_int[30] (
	.clk(clk),
	.d(at_sink_data[30]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[30]~q ),
	.prn(vcc));
defparam \at_sink_data_int[30] .is_wysiwyg = "true";
defparam \at_sink_data_int[30] .power_up = "low";

dffeas \at_sink_data_int[14] (
	.clk(clk),
	.d(at_sink_data[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[14]~q ),
	.prn(vcc));
defparam \at_sink_data_int[14] .is_wysiwyg = "true";
defparam \at_sink_data_int[14] .power_up = "low";

dffeas \at_sink_data_int[31] (
	.clk(clk),
	.d(at_sink_data[31]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[31]~q ),
	.prn(vcc));
defparam \at_sink_data_int[31] .is_wysiwyg = "true";
defparam \at_sink_data_int[31] .power_up = "low";

dffeas \at_sink_data_int[15] (
	.clk(clk),
	.d(at_sink_data[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[15]~q ),
	.prn(vcc));
defparam \at_sink_data_int[15] .is_wysiwyg = "true";
defparam \at_sink_data_int[15] .power_up = "low";

cycloneive_lcell_comb data_take(
	.dataa(\Selector4~0_combout ),
	.datab(\Selector2~4_combout ),
	.datac(\Selector2~5_combout ),
	.datad(\fifo_wrreq~0_combout ),
	.cin(gnd),
	.combout(\data_take~combout ),
	.cout());
defparam data_take.lut_mask = 16'hFFFE;
defparam data_take.sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_wrreq~0_wirecell (
	.dataa(\fifo_wrreq~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_wrreq~0_wirecell_combout ),
	.cout());
defparam \fifo_wrreq~0_wirecell .lut_mask = 16'h5555;
defparam \fifo_wrreq~0_wirecell .sum_lutc_input = "datac";

dffeas at_sink_ready_s(
	.clk(clk),
	.d(\at_sink_ready_s~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_sink_ready_s1),
	.prn(vcc));
defparam at_sink_ready_s.is_wysiwyg = "true";
defparam at_sink_ready_s.power_up = "low";

dffeas sink_start(
	.clk(clk),
	.d(\sink_start~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sink_start1),
	.prn(vcc));
defparam sink_start.is_wysiwyg = "true";
defparam sink_start.power_up = "low";

cycloneive_lcell_comb sink_stall(
	.dataa(gnd),
	.datab(gnd),
	.datac(sink_start1),
	.datad(empty_dff),
	.cin(gnd),
	.combout(sink_stall1),
	.cout());
defparam sink_stall.lut_mask = 16'h0FFF;
defparam sink_stall.sum_lutc_input = "datac";

dffeas \packet_error_s[0] (
	.clk(clk),
	.d(\Selector6~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(packet_error_s_0),
	.prn(vcc));
defparam \packet_error_s[0] .is_wysiwyg = "true";
defparam \packet_error_s[0] .power_up = "low";

dffeas \packet_error_s[1] (
	.clk(clk),
	.d(\Selector5~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(packet_error_s_1),
	.prn(vcc));
defparam \packet_error_s[1] .is_wysiwyg = "true";
defparam \packet_error_s[1] .power_up = "low";

dffeas send_sop_s(
	.clk(clk),
	.d(\Equal1~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\send_sop_eop_p~0_combout ),
	.q(send_sop_s1),
	.prn(vcc));
defparam send_sop_s.is_wysiwyg = "true";
defparam send_sop_s.power_up = "low";

dffeas send_eop_s(
	.clk(clk),
	.d(\LessThan0~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\send_sop_eop_p~0_combout ),
	.q(send_eop_s1),
	.prn(vcc));
defparam send_eop_s.is_wysiwyg = "true";
defparam send_eop_s.power_up = "low";

cycloneive_lcell_comb \at_sink_ready_s~0 (
	.dataa(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dffe_af~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\at_sink_ready_s~0_combout ),
	.cout());
defparam \at_sink_ready_s~0 .lut_mask = 16'h5555;
defparam \at_sink_ready_s~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_start~0 (
	.dataa(sink_start1),
	.datab(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sink_start~0_combout ),
	.cout());
defparam \sink_start~0 .lut_mask = 16'hEEEE;
defparam \sink_start~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[5]~20 (
	.dataa(\count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[4]~19 ),
	.combout(\count[5]~20_combout ),
	.cout(\count[5]~21 ));
defparam \count[5]~20 .lut_mask = 16'h5A5F;
defparam \count[5]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \sink_comb_update_2~2 (
	.dataa(at_sink_ready_s1),
	.datab(sink_valid),
	.datac(sink_eop),
	.datad(\max_reached~q ),
	.cin(gnd),
	.combout(\sink_comb_update_2~2_combout ),
	.cout());
defparam \sink_comb_update_2~2 .lut_mask = 16'hFFFE;
defparam \sink_comb_update_2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector4~0 (
	.dataa(\Selector2~2_combout ),
	.datab(\sink_comb_update_2~2_combout ),
	.datac(sink_error_0),
	.datad(sink_error_1),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hEFFF;
defparam \Selector4~0 .sum_lutc_input = "datac";

dffeas \sink_state.end1 (
	.clk(clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.end1~q ),
	.prn(vcc));
defparam \sink_state.end1 .is_wysiwyg = "true";
defparam \sink_state.end1 .power_up = "low";

dffeas \sink_state.st_err (
	.clk(clk),
	.d(\Selector3~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.st_err~q ),
	.prn(vcc));
defparam \sink_state.st_err .is_wysiwyg = "true";
defparam \sink_state.st_err .power_up = "low";

cycloneive_lcell_comb \Selector5~0 (
	.dataa(\sink_state.start~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sink_state.st_err~q ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hAAFF;
defparam \Selector5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~3 (
	.dataa(\Selector3~0_combout ),
	.datab(\sink_state.end1~q ),
	.datac(at_sink_ready_s1),
	.datad(\Selector5~0_combout ),
	.cin(gnd),
	.combout(\Selector3~3_combout ),
	.cout());
defparam \Selector3~3 .lut_mask = 16'hFEFF;
defparam \Selector3~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~2 (
	.dataa(\sink_state.run1~q ),
	.datab(\sink_state.stall~q ),
	.datac(sink_valid),
	.datad(sink_sop),
	.cin(gnd),
	.combout(\Selector2~2_combout ),
	.cout());
defparam \Selector2~2 .lut_mask = 16'hEFFF;
defparam \Selector2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~2 (
	.dataa(\max_reached~q ),
	.datab(sink_eop),
	.datac(at_sink_ready_s1),
	.datad(sink_valid),
	.cin(gnd),
	.combout(\Selector1~2_combout ),
	.cout());
defparam \Selector1~2 .lut_mask = 16'hDFD5;
defparam \Selector1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~3 (
	.dataa(sink_error_0),
	.datab(sink_error_1),
	.datac(\Selector2~2_combout ),
	.datad(\Selector1~2_combout ),
	.cin(gnd),
	.combout(\Selector1~3_combout ),
	.cout());
defparam \Selector1~3 .lut_mask = 16'hF7FF;
defparam \Selector1~3 .sum_lutc_input = "datac";

dffeas \sink_state.stall (
	.clk(clk),
	.d(\Selector1~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.stall~q ),
	.prn(vcc));
defparam \sink_state.stall .is_wysiwyg = "true";
defparam \sink_state.stall .power_up = "low";

cycloneive_lcell_comb \Selector4~1 (
	.dataa(\sink_state.run1~q ),
	.datab(\sink_state.stall~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector4~1_combout ),
	.cout());
defparam \Selector4~1 .lut_mask = 16'hEEEE;
defparam \Selector4~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~4 (
	.dataa(sink_valid),
	.datab(\Selector4~1_combout ),
	.datac(sink_sop),
	.datad(\sink_comb_update_2~3_combout ),
	.cin(gnd),
	.combout(\Selector3~4_combout ),
	.cout());
defparam \Selector3~4 .lut_mask = 16'hFFFE;
defparam \Selector3~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(sink_error_0),
	.datad(sink_error_1),
	.cin(gnd),
	.combout(\Selector2~5_combout ),
	.cout());
defparam \Selector2~5 .lut_mask = 16'h0FFF;
defparam \Selector2~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~5 (
	.dataa(\Selector3~2_combout ),
	.datab(\Selector3~3_combout ),
	.datac(\Selector3~4_combout ),
	.datad(\Selector2~5_combout ),
	.cin(gnd),
	.combout(\Selector3~5_combout ),
	.cout());
defparam \Selector3~5 .lut_mask = 16'hFEFF;
defparam \Selector3~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[0]~12 (
	.dataa(\max_reached~q ),
	.datab(\Selector3~5_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count[0]~12_combout ),
	.cout());
defparam \count[0]~12 .lut_mask = 16'hEEEE;
defparam \count[0]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_comb_update_2~0 (
	.dataa(at_sink_ready_s1),
	.datab(sink_valid),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sink_comb_update_2~0_combout ),
	.cout());
defparam \sink_comb_update_2~0 .lut_mask = 16'hEEEE;
defparam \sink_comb_update_2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector0~0 (
	.dataa(\sink_state.end1~q ),
	.datab(sink_sop),
	.datac(at_sink_ready_s1),
	.datad(sink_valid),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hEFFF;
defparam \Selector0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector0~1 (
	.dataa(\Selector2~5_combout ),
	.datab(\Selector0~0_combout ),
	.datac(\sink_comb_update_2~0_combout ),
	.datad(\Selector5~0_combout ),
	.cin(gnd),
	.combout(\Selector0~1_combout ),
	.cout());
defparam \Selector0~1 .lut_mask = 16'hFFF7;
defparam \Selector0~1 .sum_lutc_input = "datac";

dffeas \sink_state.start (
	.clk(clk),
	.d(\Selector0~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.start~q ),
	.prn(vcc));
defparam \sink_state.start .is_wysiwyg = "true";
defparam \sink_state.start .power_up = "low";

cycloneive_lcell_comb \Selector2~3 (
	.dataa(sink_sop),
	.datab(\sink_state.end1~q ),
	.datac(\sink_state.st_err~q ),
	.datad(\sink_state.start~q ),
	.cin(gnd),
	.combout(\Selector2~3_combout ),
	.cout());
defparam \Selector2~3 .lut_mask = 16'hFEFF;
defparam \Selector2~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_comb_update_2~1 (
	.dataa(at_sink_ready_s1),
	.datab(sink_valid),
	.datac(sink_eop),
	.datad(\max_reached~q ),
	.cin(gnd),
	.combout(\sink_comb_update_2~1_combout ),
	.cout());
defparam \sink_comb_update_2~1 .lut_mask = 16'hEFFF;
defparam \sink_comb_update_2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~4 (
	.dataa(\Selector2~2_combout ),
	.datab(\sink_comb_update_2~0_combout ),
	.datac(\Selector2~3_combout ),
	.datad(\sink_comb_update_2~1_combout ),
	.cin(gnd),
	.combout(\Selector2~4_combout ),
	.cout());
defparam \Selector2~4 .lut_mask = 16'hFFFE;
defparam \Selector2~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_take~2 (
	.dataa(\Selector2~2_combout ),
	.datab(\sink_comb_update_2~2_combout ),
	.datac(\Selector2~4_combout ),
	.datad(\Selector2~5_combout ),
	.cin(gnd),
	.combout(\data_take~2_combout ),
	.cout());
defparam \data_take~2 .lut_mask = 16'h7FFF;
defparam \data_take~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[0]~13 (
	.dataa(\Selector3~5_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\data_take~2_combout ),
	.cin(gnd),
	.combout(\count[0]~13_combout ),
	.cout());
defparam \count[0]~13 .lut_mask = 16'hAAFF;
defparam \count[0]~13 .sum_lutc_input = "datac";

dffeas \count[5] (
	.clk(clk),
	.d(\count[5]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[0]~12_combout ),
	.sload(gnd),
	.ena(\count[0]~13_combout ),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

cycloneive_lcell_comb \count[6]~22 (
	.dataa(\count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[5]~21 ),
	.combout(\count[6]~22_combout ),
	.cout(\count[6]~23 ));
defparam \count[6]~22 .lut_mask = 16'h5AAF;
defparam \count[6]~22 .sum_lutc_input = "cin";

dffeas \count[6] (
	.clk(clk),
	.d(\count[6]~22_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[0]~12_combout ),
	.sload(gnd),
	.ena(\count[0]~13_combout ),
	.q(\count[6]~q ),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

cycloneive_lcell_comb \count[7]~24 (
	.dataa(\count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\count[6]~23 ),
	.combout(\count[7]~24_combout ),
	.cout());
defparam \count[7]~24 .lut_mask = 16'h5A5A;
defparam \count[7]~24 .sum_lutc_input = "cin";

dffeas \count[7] (
	.clk(clk),
	.d(\count[7]~24_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[0]~12_combout ),
	.sload(gnd),
	.ena(\count[0]~13_combout ),
	.q(\count[7]~q ),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

cycloneive_lcell_comb \max_reached~1 (
	.dataa(\count[4]~q ),
	.datab(\count[5]~q ),
	.datac(\count[6]~q ),
	.datad(\count[7]~q ),
	.cin(gnd),
	.combout(\max_reached~1_combout ),
	.cout());
defparam \max_reached~1 .lut_mask = 16'hFFFE;
defparam \max_reached~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \max_reached~2 (
	.dataa(\max_reached~0_combout ),
	.datab(\max_reached~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\max_reached~2_combout ),
	.cout());
defparam \max_reached~2 .lut_mask = 16'hEEEE;
defparam \max_reached~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \max_reached~3 (
	.dataa(\max_reached~q ),
	.datab(\max_reached~2_combout ),
	.datac(\data_take~2_combout ),
	.datad(\Selector3~5_combout ),
	.cin(gnd),
	.combout(\max_reached~3_combout ),
	.cout());
defparam \max_reached~3 .lut_mask = 16'hEFFE;
defparam \max_reached~3 .sum_lutc_input = "datac";

dffeas max_reached(
	.clk(clk),
	.d(\max_reached~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\max_reached~q ),
	.prn(vcc));
defparam max_reached.is_wysiwyg = "true";
defparam max_reached.power_up = "low";

cycloneive_lcell_comb \sink_comb_update_2~3 (
	.dataa(sink_eop),
	.datab(gnd),
	.datac(gnd),
	.datad(\max_reached~q ),
	.cin(gnd),
	.combout(\sink_comb_update_2~3_combout ),
	.cout());
defparam \sink_comb_update_2~3 .lut_mask = 16'hAAFF;
defparam \sink_comb_update_2~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector6~0 (
	.dataa(sink_valid),
	.datab(\sink_comb_update_2~3_combout ),
	.datac(sink_sop),
	.datad(at_sink_ready_s1),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
defparam \Selector6~0 .lut_mask = 16'hFEFF;
defparam \Selector6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector6~1 (
	.dataa(\Selector4~1_combout ),
	.datab(sink_error_0),
	.datac(\Selector6~0_combout ),
	.datad(sink_error_1),
	.cin(gnd),
	.combout(\Selector6~1_combout ),
	.cout());
defparam \Selector6~1 .lut_mask = 16'hFEFF;
defparam \Selector6~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~0 (
	.dataa(sink_valid),
	.datab(gnd),
	.datac(gnd),
	.datad(sink_sop),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'hAAFF;
defparam \Selector3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector6~2 (
	.dataa(\sink_state.end1~q ),
	.datab(sink_error_0),
	.datac(\Selector3~0_combout ),
	.datad(sink_error_1),
	.cin(gnd),
	.combout(\Selector6~2_combout ),
	.cout());
defparam \Selector6~2 .lut_mask = 16'hFEFF;
defparam \Selector6~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector6~3 (
	.dataa(sink_error_0),
	.datab(\sink_comb_update_2~0_combout ),
	.datac(sink_sop),
	.datad(sink_error_1),
	.cin(gnd),
	.combout(\Selector6~3_combout ),
	.cout());
defparam \Selector6~3 .lut_mask = 16'hEFFF;
defparam \Selector6~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector6~4 (
	.dataa(\Selector6~1_combout ),
	.datab(\Selector6~2_combout ),
	.datac(\Selector6~3_combout ),
	.datad(\Selector5~0_combout ),
	.cin(gnd),
	.combout(\Selector6~4_combout ),
	.cout());
defparam \Selector6~4 .lut_mask = 16'hFEFF;
defparam \Selector6~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~6 (
	.dataa(sink_error_0),
	.datab(sink_error_1),
	.datac(\Selector2~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector2~6_combout ),
	.cout());
defparam \Selector2~6 .lut_mask = 16'hF7F7;
defparam \Selector2~6 .sum_lutc_input = "datac";

dffeas \sink_state.run1 (
	.clk(clk),
	.d(\Selector2~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.run1~q ),
	.prn(vcc));
defparam \sink_state.run1 .is_wysiwyg = "true";
defparam \sink_state.run1 .power_up = "low";

cycloneive_lcell_comb \fifo_wrreq~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sink_state.run1~q ),
	.datad(\sink_state.end1~q ),
	.cin(gnd),
	.combout(\fifo_wrreq~0_combout ),
	.cout());
defparam \fifo_wrreq~0 .lut_mask = 16'hFFF0;
defparam \fifo_wrreq~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector5~1 (
	.dataa(sink_error_1),
	.datab(\sink_state.stall~q ),
	.datac(\fifo_wrreq~0_combout ),
	.datad(\Selector5~0_combout ),
	.cin(gnd),
	.combout(\Selector5~1_combout ),
	.cout());
defparam \Selector5~1 .lut_mask = 16'hFEFF;
defparam \Selector5~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector5~2 (
	.dataa(\Selector3~2_combout ),
	.datab(sink_valid),
	.datac(\Selector4~1_combout ),
	.datad(\sink_comb_update_2~3_combout ),
	.cin(gnd),
	.combout(\Selector5~2_combout ),
	.cout());
defparam \Selector5~2 .lut_mask = 16'hFFFE;
defparam \Selector5~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_comb_update_2~4 (
	.dataa(sink_valid),
	.datab(sink_sop),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sink_comb_update_2~4_combout ),
	.cout());
defparam \sink_comb_update_2~4 .lut_mask = 16'hEEEE;
defparam \sink_comb_update_2~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector5~3 (
	.dataa(\Selector5~1_combout ),
	.datab(\Selector5~2_combout ),
	.datac(\sink_comb_update_2~4_combout ),
	.datad(sink_error_0),
	.cin(gnd),
	.combout(\Selector5~3_combout ),
	.cout());
defparam \Selector5~3 .lut_mask = 16'hEFFF;
defparam \Selector5~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_cnt[1]~10 (
	.dataa(\out_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[0]~9 ),
	.combout(\out_cnt[1]~10_combout ),
	.cout(\out_cnt[1]~11 ));
defparam \out_cnt[1]~10 .lut_mask = 16'h5A5F;
defparam \out_cnt[1]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \out_cnt[2]~12 (
	.dataa(\out_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[1]~11 ),
	.combout(\out_cnt[2]~12_combout ),
	.cout(\out_cnt[2]~13 ));
defparam \out_cnt[2]~12 .lut_mask = 16'h5AAF;
defparam \out_cnt[2]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \out_cnt[3]~14 (
	.dataa(\out_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[2]~13 ),
	.combout(\out_cnt[3]~14_combout ),
	.cout(\out_cnt[3]~15 ));
defparam \out_cnt[3]~14 .lut_mask = 16'h5A5F;
defparam \out_cnt[3]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \out_cnt[5]~18 (
	.dataa(\out_cnt[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[4]~17 ),
	.combout(\out_cnt[5]~18_combout ),
	.cout(\out_cnt[5]~19 ));
defparam \out_cnt[5]~18 .lut_mask = 16'h5A5F;
defparam \out_cnt[5]~18 .sum_lutc_input = "cin";

dffeas sink_stall_s(
	.clk(clk),
	.d(sink_stall1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_stall_s~q ),
	.prn(vcc));
defparam sink_stall_s.is_wysiwyg = "true";
defparam sink_stall_s.power_up = "low";

cycloneive_lcell_comb \Selector8~0 (
	.dataa(sink_ready_ctrl),
	.datab(\sink_stall_s~q ),
	.datac(\sink_out_state.normal~q ),
	.datad(sink_stall1),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
defparam \Selector8~0 .lut_mask = 16'hFFF7;
defparam \Selector8~0 .sum_lutc_input = "datac";

dffeas \sink_out_state.normal (
	.clk(clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_out_state.normal~q ),
	.prn(vcc));
defparam \sink_out_state.normal .is_wysiwyg = "true";
defparam \sink_out_state.normal .power_up = "low";

cycloneive_lcell_comb \Selector7~0 (
	.dataa(\sink_out_state.empty_and_ready~q ),
	.datab(sink_ready_ctrl),
	.datac(\sink_out_state.normal~q ),
	.datad(sink_stall1),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
defparam \Selector7~0 .lut_mask = 16'hEFFF;
defparam \Selector7~0 .sum_lutc_input = "datac";

dffeas \out_cnt[5] (
	.clk(clk),
	.d(\out_cnt[5]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[5]~q ),
	.prn(vcc));
defparam \out_cnt[5] .is_wysiwyg = "true";
defparam \out_cnt[5] .power_up = "low";

cycloneive_lcell_comb \out_cnt[6]~20 (
	.dataa(\out_cnt[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[5]~19 ),
	.combout(\out_cnt[6]~20_combout ),
	.cout(\out_cnt[6]~21 ));
defparam \out_cnt[6]~20 .lut_mask = 16'h5AAF;
defparam \out_cnt[6]~20 .sum_lutc_input = "cin";

dffeas \out_cnt[6] (
	.clk(clk),
	.d(\out_cnt[6]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[6]~q ),
	.prn(vcc));
defparam \out_cnt[6] .is_wysiwyg = "true";
defparam \out_cnt[6] .power_up = "low";

cycloneive_lcell_comb \out_cnt[7]~22 (
	.dataa(\out_cnt[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\out_cnt[6]~21 ),
	.combout(\out_cnt[7]~22_combout ),
	.cout());
defparam \out_cnt[7]~22 .lut_mask = 16'h5A5A;
defparam \out_cnt[7]~22 .sum_lutc_input = "cin";

dffeas \out_cnt[7] (
	.clk(clk),
	.d(\out_cnt[7]~22_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[7]~q ),
	.prn(vcc));
defparam \out_cnt[7] .is_wysiwyg = "true";
defparam \out_cnt[7] .power_up = "low";

cycloneive_lcell_comb \LessThan0~1 (
	.dataa(\out_cnt[4]~q ),
	.datab(\out_cnt[5]~q ),
	.datac(\out_cnt[6]~q ),
	.datad(\out_cnt[7]~q ),
	.cin(gnd),
	.combout(\LessThan0~1_combout ),
	.cout());
defparam \LessThan0~1 .lut_mask = 16'h7FFF;
defparam \LessThan0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \LessThan0~2 (
	.dataa(\LessThan0~0_combout ),
	.datab(\LessThan0~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\LessThan0~2_combout ),
	.cout());
defparam \LessThan0~2 .lut_mask = 16'h7777;
defparam \LessThan0~2 .sum_lutc_input = "datac";

dffeas \out_cnt[1] (
	.clk(clk),
	.d(\out_cnt[1]~10_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[1]~q ),
	.prn(vcc));
defparam \out_cnt[1] .is_wysiwyg = "true";
defparam \out_cnt[1] .power_up = "low";

dffeas \out_cnt[2] (
	.clk(clk),
	.d(\out_cnt[2]~12_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[2]~q ),
	.prn(vcc));
defparam \out_cnt[2] .is_wysiwyg = "true";
defparam \out_cnt[2] .power_up = "low";

dffeas \out_cnt[3] (
	.clk(clk),
	.d(\out_cnt[3]~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[3]~q ),
	.prn(vcc));
defparam \out_cnt[3] .is_wysiwyg = "true";
defparam \out_cnt[3] .power_up = "low";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(\out_cnt[0]~q ),
	.datab(\out_cnt[1]~q ),
	.datac(\out_cnt[2]~q ),
	.datad(\out_cnt[3]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'h7FFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~1 (
	.dataa(\out_cnt[4]~q ),
	.datab(\out_cnt[5]~q ),
	.datac(\out_cnt[6]~q ),
	.datad(\out_cnt[7]~q ),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'h7FFF;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~2 (
	.dataa(\Equal1~0_combout ),
	.datab(\Equal1~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal1~2_combout ),
	.cout());
defparam \Equal1~2 .lut_mask = 16'hEEEE;
defparam \Equal1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector10~0 (
	.dataa(sink_stall_reg),
	.datab(source_stall_reg),
	.datac(\sink_stall_s~q ),
	.datad(master_sink_ena),
	.cin(gnd),
	.combout(\Selector10~0_combout ),
	.cout());
defparam \Selector10~0 .lut_mask = 16'h6996;
defparam \Selector10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector10~1 (
	.dataa(sink_stall1),
	.datab(\sink_out_state.empty_and_ready~q ),
	.datac(\Selector10~0_combout ),
	.datad(\sink_out_state.normal~q ),
	.cin(gnd),
	.combout(\Selector10~1_combout ),
	.cout());
defparam \Selector10~1 .lut_mask = 16'hFEFF;
defparam \Selector10~1 .sum_lutc_input = "datac";

dffeas \sink_out_state.empty_and_ready (
	.clk(clk),
	.d(\Selector10~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_out_state.empty_and_ready~q ),
	.prn(vcc));
defparam \sink_out_state.empty_and_ready .is_wysiwyg = "true";
defparam \sink_out_state.empty_and_ready .power_up = "low";

cycloneive_lcell_comb \send_sop_eop_p~0 (
	.dataa(sink_ready_ctrl),
	.datab(\sink_out_state.empty_and_ready~q ),
	.datac(\sink_out_state.normal~q ),
	.datad(sink_stall1),
	.cin(gnd),
	.combout(\send_sop_eop_p~0_combout ),
	.cout());
defparam \send_sop_eop_p~0 .lut_mask = 16'hEFFF;
defparam \send_sop_eop_p~0 .sum_lutc_input = "datac";

endmodule

module fft256_scfifo_1 (
	q,
	dffe_af,
	empty_dff,
	rdreq,
	sink_staterun1,
	sink_stateend1,
	wrreq,
	counter_reg_bit_0,
	data,
	fifo_wrreq,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[33:0] q;
output 	dffe_af;
output 	empty_dff;
input 	rdreq;
input 	sink_staterun1;
input 	sink_stateend1;
input 	wrreq;
output 	counter_reg_bit_0;
input 	[33:0] data;
input 	fifo_wrreq;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fft256_scfifo_udh1 auto_generated(
	.q({q_unconnected_wire_33,q_unconnected_wire_32,q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.dffe_af1(dffe_af),
	.empty_dff(empty_dff),
	.rdreq(rdreq),
	.sink_staterun1(sink_staterun1),
	.sink_stateend1(sink_stateend1),
	.wrreq(wrreq),
	.counter_reg_bit_0(counter_reg_bit_0),
	.data({gnd,gnd,data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.fifo_wrreq(fifo_wrreq),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module fft256_scfifo_udh1 (
	q,
	dffe_af1,
	empty_dff,
	rdreq,
	sink_staterun1,
	sink_stateend1,
	wrreq,
	counter_reg_bit_0,
	data,
	fifo_wrreq,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[33:0] q;
output 	dffe_af1;
output 	empty_dff;
input 	rdreq;
input 	sink_staterun1;
input 	sink_stateend1;
input 	wrreq;
output 	counter_reg_bit_0;
input 	[33:0] data;
input 	fifo_wrreq;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \dffe_af~0_combout ;
wire \dffe_af~1_combout ;


fft256_a_dpfifo_no81 dpfifo(
	.q({q_unconnected_wire_33,q_unconnected_wire_32,q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.empty_dff1(empty_dff),
	.rreq(rdreq),
	.sink_staterun1(sink_staterun1),
	.sink_stateend1(sink_stateend1),
	.wreq(wrreq),
	.counter_reg_bit_1(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.data({gnd,gnd,data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.wreq1(fifo_wrreq),
	.clock(clock),
	.reset_n(reset_n));

dffeas dffe_af(
	.clk(clock),
	.d(\dffe_af~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe_af1),
	.prn(vcc));
defparam dffe_af.is_wysiwyg = "true";
defparam dffe_af.power_up = "low";

cycloneive_lcell_comb \dffe_af~0 (
	.dataa(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datab(counter_reg_bit_0),
	.datac(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datad(dffe_af1),
	.cin(gnd),
	.combout(\dffe_af~0_combout ),
	.cout());
defparam \dffe_af~0 .lut_mask = 16'hF7FD;
defparam \dffe_af~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \dffe_af~1 (
	.dataa(rdreq),
	.datab(wrreq),
	.datac(dffe_af1),
	.datad(\dffe_af~0_combout ),
	.cin(gnd),
	.combout(\dffe_af~1_combout ),
	.cout());
defparam \dffe_af~1 .lut_mask = 16'hDDF5;
defparam \dffe_af~1 .sum_lutc_input = "datac";

endmodule

module fft256_a_dpfifo_no81 (
	q,
	empty_dff1,
	rreq,
	sink_staterun1,
	sink_stateend1,
	wreq,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_2,
	data,
	wreq1,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[33:0] q;
output 	empty_dff1;
input 	rreq;
input 	sink_staterun1;
input 	sink_stateend1;
input 	wreq;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
input 	[33:0] data;
input 	wreq1;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \usedw_is_1_dff~q ;
wire \usedw_will_be_1~1_combout ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \_~6_combout ;
wire \_~7_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \usedw_is_0_dff~q ;
wire \_~2_combout ;
wire \_~3_combout ;
wire \_~4_combout ;
wire \usedw_will_be_1~0_combout ;
wire \_~5_combout ;


fft256_cntr_unb wr_ptr(
	.fifo_wrreq(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.clock(clock),
	.reset_n(reset_n));

fft256_cntr_ao7 usedw_counter(
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	._(\_~7_combout ),
	.updown(wreq1),
	.clock(clock),
	.reset_n(reset_n));

fft256_cntr_tnb rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	._(\_~6_combout ),
	.clock(clock),
	.reset_n(reset_n));

fft256_altsyncram_ssf1 FIFOram(
	.q_b({q_b_unconnected_wire_33,q_b_unconnected_wire_32,q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.clocken1(rreq),
	.wren_a(wreq),
	.data_a({gnd,gnd,data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock0(clock),
	.clock1(clock));

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_will_be_1~0_combout ),
	.datab(rreq),
	.datac(wreq),
	.datad(\_~3_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFFEF;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\ram_read_address[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rreq),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(rreq),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\ram_read_address[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(rreq),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\ram_read_address[2]~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(rreq),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~6 (
	.dataa(rreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\_~6_combout ),
	.cout());
defparam \_~6 .lut_mask = 16'hAAFF;
defparam \_~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~7 (
	.dataa(sink_staterun1),
	.datab(sink_stateend1),
	.datac(rreq),
	.datad(gnd),
	.cin(gnd),
	.combout(\_~7_combout ),
	.cout());
defparam \_~7 .lut_mask = 16'h9696;
defparam \_~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(\rd_ptr_lsb~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'h5555;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\_~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_dff1),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

cycloneive_lcell_comb \_~2 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(rreq),
	.datac(wreq),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFF7D;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~3 (
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(counter_reg_bit_0),
	.datad(counter_reg_bit_2),
	.cin(gnd),
	.combout(\_~3_combout ),
	.cout());
defparam \_~3 .lut_mask = 16'hAFFF;
defparam \_~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~4 (
	.dataa(rreq),
	.datab(\_~3_combout ),
	.datac(sink_staterun1),
	.datad(sink_stateend1),
	.cin(gnd),
	.combout(\_~4_combout ),
	.cout());
defparam \_~4 .lut_mask = 16'hEFFF;
defparam \_~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\usedw_is_0_dff~q ),
	.datac(rreq),
	.datad(wreq),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFB;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~5 (
	.dataa(\_~2_combout ),
	.datab(\_~4_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(wreq),
	.cin(gnd),
	.combout(\_~5_combout ),
	.cout());
defparam \_~5 .lut_mask = 16'hBFFF;
defparam \_~5 .sum_lutc_input = "datac";

endmodule

module fft256_altsyncram_ssf1 (
	q_b,
	clocken1,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[33:0] q_b;
input 	clocken1;
input 	wren_a;
input 	[33:0] data_a;
input 	[2:0] address_a;
input 	[2:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 3;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 7;
defparam ram_block1a16.port_a_logical_ram_depth = 8;
defparam ram_block1a16.port_a_logical_ram_width = 34;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 3;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 7;
defparam ram_block1a16.port_b_logical_ram_depth = 8;
defparam ram_block1a16.port_b_logical_ram_width = 34;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 3;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 7;
defparam ram_block1a0.port_a_logical_ram_depth = 8;
defparam ram_block1a0.port_a_logical_ram_width = 34;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 3;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 7;
defparam ram_block1a0.port_b_logical_ram_depth = 8;
defparam ram_block1a0.port_b_logical_ram_width = 34;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 3;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 7;
defparam ram_block1a17.port_a_logical_ram_depth = 8;
defparam ram_block1a17.port_a_logical_ram_width = 34;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 3;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 7;
defparam ram_block1a17.port_b_logical_ram_depth = 8;
defparam ram_block1a17.port_b_logical_ram_width = 34;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 3;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 7;
defparam ram_block1a1.port_a_logical_ram_depth = 8;
defparam ram_block1a1.port_a_logical_ram_width = 34;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 3;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 7;
defparam ram_block1a1.port_b_logical_ram_depth = 8;
defparam ram_block1a1.port_b_logical_ram_width = 34;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 3;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 7;
defparam ram_block1a18.port_a_logical_ram_depth = 8;
defparam ram_block1a18.port_a_logical_ram_width = 34;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 3;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 7;
defparam ram_block1a18.port_b_logical_ram_depth = 8;
defparam ram_block1a18.port_b_logical_ram_width = 34;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 3;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 7;
defparam ram_block1a2.port_a_logical_ram_depth = 8;
defparam ram_block1a2.port_a_logical_ram_width = 34;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 3;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 7;
defparam ram_block1a2.port_b_logical_ram_depth = 8;
defparam ram_block1a2.port_b_logical_ram_width = 34;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 3;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 7;
defparam ram_block1a19.port_a_logical_ram_depth = 8;
defparam ram_block1a19.port_a_logical_ram_width = 34;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 3;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 7;
defparam ram_block1a19.port_b_logical_ram_depth = 8;
defparam ram_block1a19.port_b_logical_ram_width = 34;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 3;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 7;
defparam ram_block1a3.port_a_logical_ram_depth = 8;
defparam ram_block1a3.port_a_logical_ram_width = 34;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 3;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 7;
defparam ram_block1a3.port_b_logical_ram_depth = 8;
defparam ram_block1a3.port_b_logical_ram_width = 34;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 3;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 7;
defparam ram_block1a20.port_a_logical_ram_depth = 8;
defparam ram_block1a20.port_a_logical_ram_width = 34;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 3;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 7;
defparam ram_block1a20.port_b_logical_ram_depth = 8;
defparam ram_block1a20.port_b_logical_ram_width = 34;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 3;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 7;
defparam ram_block1a4.port_a_logical_ram_depth = 8;
defparam ram_block1a4.port_a_logical_ram_width = 34;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 3;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 7;
defparam ram_block1a4.port_b_logical_ram_depth = 8;
defparam ram_block1a4.port_b_logical_ram_width = 34;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 3;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 7;
defparam ram_block1a21.port_a_logical_ram_depth = 8;
defparam ram_block1a21.port_a_logical_ram_width = 34;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 3;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 7;
defparam ram_block1a21.port_b_logical_ram_depth = 8;
defparam ram_block1a21.port_b_logical_ram_width = 34;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 3;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 7;
defparam ram_block1a5.port_a_logical_ram_depth = 8;
defparam ram_block1a5.port_a_logical_ram_width = 34;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 3;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 7;
defparam ram_block1a5.port_b_logical_ram_depth = 8;
defparam ram_block1a5.port_b_logical_ram_width = 34;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.clk1_output_clock_enable = "ena1";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 3;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 7;
defparam ram_block1a22.port_a_logical_ram_depth = 8;
defparam ram_block1a22.port_a_logical_ram_width = 34;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 3;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "clock1";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 7;
defparam ram_block1a22.port_b_logical_ram_depth = 8;
defparam ram_block1a22.port_b_logical_ram_width = 34;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 3;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 7;
defparam ram_block1a6.port_a_logical_ram_depth = 8;
defparam ram_block1a6.port_a_logical_ram_width = 34;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 3;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 7;
defparam ram_block1a6.port_b_logical_ram_depth = 8;
defparam ram_block1a6.port_b_logical_ram_width = 34;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.clk1_output_clock_enable = "ena1";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 3;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 7;
defparam ram_block1a23.port_a_logical_ram_depth = 8;
defparam ram_block1a23.port_a_logical_ram_width = 34;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 3;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "clock1";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 7;
defparam ram_block1a23.port_b_logical_ram_depth = 8;
defparam ram_block1a23.port_b_logical_ram_width = 34;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 3;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 7;
defparam ram_block1a7.port_a_logical_ram_depth = 8;
defparam ram_block1a7.port_a_logical_ram_width = 34;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 3;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 7;
defparam ram_block1a7.port_b_logical_ram_depth = 8;
defparam ram_block1a7.port_b_logical_ram_width = 34;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.clk1_output_clock_enable = "ena1";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 3;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 7;
defparam ram_block1a24.port_a_logical_ram_depth = 8;
defparam ram_block1a24.port_a_logical_ram_width = 34;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 3;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "clock1";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 7;
defparam ram_block1a24.port_b_logical_ram_depth = 8;
defparam ram_block1a24.port_b_logical_ram_width = 34;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 3;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 7;
defparam ram_block1a8.port_a_logical_ram_depth = 8;
defparam ram_block1a8.port_a_logical_ram_width = 34;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 3;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 7;
defparam ram_block1a8.port_b_logical_ram_depth = 8;
defparam ram_block1a8.port_b_logical_ram_width = 34;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.clk1_output_clock_enable = "ena1";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 3;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 7;
defparam ram_block1a25.port_a_logical_ram_depth = 8;
defparam ram_block1a25.port_a_logical_ram_width = 34;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 3;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "clock1";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 7;
defparam ram_block1a25.port_b_logical_ram_depth = 8;
defparam ram_block1a25.port_b_logical_ram_width = 34;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 3;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 7;
defparam ram_block1a9.port_a_logical_ram_depth = 8;
defparam ram_block1a9.port_a_logical_ram_width = 34;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 3;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 7;
defparam ram_block1a9.port_b_logical_ram_depth = 8;
defparam ram_block1a9.port_b_logical_ram_width = 34;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.clk1_output_clock_enable = "ena1";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 3;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 7;
defparam ram_block1a26.port_a_logical_ram_depth = 8;
defparam ram_block1a26.port_a_logical_ram_width = 34;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 3;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "clock1";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 7;
defparam ram_block1a26.port_b_logical_ram_depth = 8;
defparam ram_block1a26.port_b_logical_ram_width = 34;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 3;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 7;
defparam ram_block1a10.port_a_logical_ram_depth = 8;
defparam ram_block1a10.port_a_logical_ram_width = 34;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 3;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 7;
defparam ram_block1a10.port_b_logical_ram_depth = 8;
defparam ram_block1a10.port_b_logical_ram_width = 34;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.clk1_output_clock_enable = "ena1";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 3;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 7;
defparam ram_block1a27.port_a_logical_ram_depth = 8;
defparam ram_block1a27.port_a_logical_ram_width = 34;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 3;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "clock1";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 7;
defparam ram_block1a27.port_b_logical_ram_depth = 8;
defparam ram_block1a27.port_b_logical_ram_width = 34;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 3;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 7;
defparam ram_block1a11.port_a_logical_ram_depth = 8;
defparam ram_block1a11.port_a_logical_ram_width = 34;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 3;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 7;
defparam ram_block1a11.port_b_logical_ram_depth = 8;
defparam ram_block1a11.port_b_logical_ram_width = 34;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.clk1_output_clock_enable = "ena1";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 3;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 7;
defparam ram_block1a28.port_a_logical_ram_depth = 8;
defparam ram_block1a28.port_a_logical_ram_width = 34;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 3;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "clock1";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 7;
defparam ram_block1a28.port_b_logical_ram_depth = 8;
defparam ram_block1a28.port_b_logical_ram_width = 34;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 3;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 7;
defparam ram_block1a12.port_a_logical_ram_depth = 8;
defparam ram_block1a12.port_a_logical_ram_width = 34;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 3;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 7;
defparam ram_block1a12.port_b_logical_ram_depth = 8;
defparam ram_block1a12.port_b_logical_ram_width = 34;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.clk1_output_clock_enable = "ena1";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 3;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 7;
defparam ram_block1a29.port_a_logical_ram_depth = 8;
defparam ram_block1a29.port_a_logical_ram_width = 34;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 3;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "clock1";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 7;
defparam ram_block1a29.port_b_logical_ram_depth = 8;
defparam ram_block1a29.port_b_logical_ram_width = 34;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 3;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 7;
defparam ram_block1a13.port_a_logical_ram_depth = 8;
defparam ram_block1a13.port_a_logical_ram_width = 34;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 3;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 7;
defparam ram_block1a13.port_b_logical_ram_depth = 8;
defparam ram_block1a13.port_b_logical_ram_width = 34;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.clk1_output_clock_enable = "ena1";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 3;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 7;
defparam ram_block1a30.port_a_logical_ram_depth = 8;
defparam ram_block1a30.port_a_logical_ram_width = 34;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 3;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "clock1";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 7;
defparam ram_block1a30.port_b_logical_ram_depth = 8;
defparam ram_block1a30.port_b_logical_ram_width = 34;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 3;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 7;
defparam ram_block1a14.port_a_logical_ram_depth = 8;
defparam ram_block1a14.port_a_logical_ram_width = 34;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 3;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 7;
defparam ram_block1a14.port_b_logical_ram_depth = 8;
defparam ram_block1a14.port_b_logical_ram_width = 34;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.clk1_output_clock_enable = "ena1";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 3;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 7;
defparam ram_block1a31.port_a_logical_ram_depth = 8;
defparam ram_block1a31.port_a_logical_ram_width = 34;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 3;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "clock1";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 7;
defparam ram_block1a31.port_b_logical_ram_depth = 8;
defparam ram_block1a31.port_b_logical_ram_width = 34;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "asj_fft_si_sose_so_b_fft_121:asj_fft_si_sose_so_b_fft_121_inst|auk_dspip_avalon_streaming_sink_fft_121:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_udh1:auto_generated|a_dpfifo_no81:dpfifo|altsyncram_ssf1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 3;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 7;
defparam ram_block1a15.port_a_logical_ram_depth = 8;
defparam ram_block1a15.port_a_logical_ram_width = 34;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 3;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 7;
defparam ram_block1a15.port_b_logical_ram_depth = 8;
defparam ram_block1a15.port_b_logical_ram_width = 34;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

endmodule

module fft256_cntr_ao7 (
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_2,
	_,
	updown,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
input 	_;
input 	updown;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

endmodule

module fft256_cntr_tnb (
	counter_reg_bit_0,
	counter_reg_bit_1,
	_,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
input 	_;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout());
defparam counter_comb_bita1.lut_mask = 16'h5A5A;
defparam counter_comb_bita1.sum_lutc_input = "cin";

endmodule

module fft256_cntr_unb (
	fifo_wrreq,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	fifo_wrreq;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wrreq),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wrreq),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wrreq),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

endmodule

module fft256_auk_dspip_avalon_streaming_source_fft_121 (
	data_count,
	at_source_error_0,
	at_source_error_1,
	at_source_sop_s1,
	at_source_eop_s1,
	at_source_valid_s1,
	at_source_data_0,
	at_source_data_1,
	at_source_data_2,
	at_source_data_3,
	at_source_data_4,
	at_source_data_5,
	at_source_data_22,
	at_source_data_23,
	at_source_data_24,
	at_source_data_25,
	at_source_data_26,
	at_source_data_27,
	at_source_data_28,
	at_source_data_29,
	at_source_data_30,
	at_source_data_31,
	at_source_data_32,
	at_source_data_33,
	at_source_data_34,
	at_source_data_35,
	at_source_data_36,
	at_source_data_37,
	at_source_data_6,
	at_source_data_7,
	at_source_data_8,
	at_source_data_9,
	at_source_data_10,
	at_source_data_11,
	at_source_data_12,
	at_source_data_13,
	at_source_data_14,
	at_source_data_15,
	at_source_data_16,
	at_source_data_17,
	at_source_data_18,
	at_source_data_19,
	at_source_data_20,
	at_source_data_21,
	source_packet_error_0,
	source_packet_error_1,
	source_stall_reg,
	master_source_ena,
	source_valid_ctrl_sop,
	source_valid_ctrl_sop1,
	stall_reg,
	source_stall_int_d1,
	data,
	Mux0,
	clk,
	reset_n,
	source_ready)/* synthesis synthesis_greybox=1 */;
input 	[7:0] data_count;
output 	at_source_error_0;
output 	at_source_error_1;
output 	at_source_sop_s1;
output 	at_source_eop_s1;
output 	at_source_valid_s1;
output 	at_source_data_0;
output 	at_source_data_1;
output 	at_source_data_2;
output 	at_source_data_3;
output 	at_source_data_4;
output 	at_source_data_5;
output 	at_source_data_22;
output 	at_source_data_23;
output 	at_source_data_24;
output 	at_source_data_25;
output 	at_source_data_26;
output 	at_source_data_27;
output 	at_source_data_28;
output 	at_source_data_29;
output 	at_source_data_30;
output 	at_source_data_31;
output 	at_source_data_32;
output 	at_source_data_33;
output 	at_source_data_34;
output 	at_source_data_35;
output 	at_source_data_36;
output 	at_source_data_37;
output 	at_source_data_6;
output 	at_source_data_7;
output 	at_source_data_8;
output 	at_source_data_9;
output 	at_source_data_10;
output 	at_source_data_11;
output 	at_source_data_12;
output 	at_source_data_13;
output 	at_source_data_14;
output 	at_source_data_15;
output 	at_source_data_16;
output 	at_source_data_17;
output 	at_source_data_18;
output 	at_source_data_19;
output 	at_source_data_20;
output 	at_source_data_21;
input 	source_packet_error_0;
input 	source_packet_error_1;
input 	source_stall_reg;
input 	master_source_ena;
input 	source_valid_ctrl_sop;
input 	source_valid_ctrl_sop1;
input 	stall_reg;
output 	source_stall_int_d1;
input 	[37:0] data;
output 	Mux0;
input 	clk;
input 	reset_n;
input 	source_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Selector1~1_combout ;
wire \data_count_int[4]~q ;
wire \source_comb_update_2~0_combout ;
wire \data_count_int1[4]~q ;
wire \source_comb_update_2~1_combout ;
wire \source_comb_update_2~2_combout ;
wire \data_count_int[7]~q ;
wire \data_count_int1[7]~q ;
wire \Selector1~3_combout ;
wire \Mux2~1_combout ;
wire \Mux2~2_combout ;
wire \valid_ctrl_inter~0_combout ;
wire \source_state.st_err~q ;
wire \first_data~0_combout ;
wire \first_data~q ;
wire \data_select~0_combout ;
wire \Mux2~3_combout ;
wire \Mux2~0_combout ;
wire \Mux2~4_combout ;
wire \was_stalled~0_combout ;
wire \was_stalled~1_combout ;
wire \was_stalled~q ;
wire \valid_ctrl_inter~1_combout ;
wire \valid_ctrl_int~q ;
wire \Mux1~0_combout ;
wire \valid_ctrl_inter1~0_combout ;
wire \valid_ctrl_int1~q ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \data_count_int1[1]~q ;
wire \data_count_int[3]~q ;
wire \data_count_int[1]~q ;
wire \data_count_int[2]~q ;
wire \source_comb_update_2~3_combout ;
wire \data_count_int1[3]~q ;
wire \data_count_int1[2]~q ;
wire \source_comb_update_2~4_combout ;
wire \source_comb_update_2~5_combout ;
wire \source_comb_update_2~6_combout ;
wire \data_count_int1[6]~q ;
wire \data_count_int[5]~q ;
wire \data_count_int[0]~q ;
wire \data_count_int[6]~q ;
wire \count_finished~0_combout ;
wire \data_count_int1[5]~q ;
wire \data_count_int1[0]~q ;
wire \count_finished~1_combout ;
wire \count_finished~2_combout ;
wire \count_finished~3_combout ;
wire \count_finished~4_combout ;
wire \count_finished~5_combout ;
wire \Selector1~0_combout ;
wire \source_comb_update_2~7_combout ;
wire \Selector2~4_combout ;
wire \Selector1~5_combout ;
wire \Selector2~3_combout ;
wire \source_state.run1~q ;
wire \Selector3~0_combout ;
wire \Selector3~1_combout ;
wire \Selector3~2_combout ;
wire \source_state.end1~q ;
wire \packet_error0~combout ;
wire \Selector0~1_combout ;
wire \source_state.start~q ;
wire \Selector0~0_combout ;
wire \Selector1~2_combout ;
wire \valid_ctrl_int_selected~0_combout ;
wire \Selector2~2_combout ;
wire \Selector1~4_combout ;
wire \Selector5~0_combout ;
wire \source_state.sop~q ;
wire \Selector5~1_combout ;
wire \at_source_valid_int~0_combout ;
wire \at_source_valid_int~1_combout ;
wire \at_source_valid_int~2_combout ;
wire \data_int1[0]~q ;
wire \data_int[0]~q ;
wire \data_int_selected[0]~0_combout ;
wire \data_int1[1]~q ;
wire \data_int[1]~q ;
wire \data_int_selected[1]~1_combout ;
wire \data_int1[2]~q ;
wire \data_int[2]~q ;
wire \data_int_selected[2]~2_combout ;
wire \data_int1[3]~q ;
wire \data_int[3]~q ;
wire \data_int_selected[3]~3_combout ;
wire \data_int1[4]~q ;
wire \data_int[4]~q ;
wire \data_int_selected[4]~4_combout ;
wire \data_int1[5]~q ;
wire \data_int[5]~q ;
wire \data_int_selected[5]~5_combout ;
wire \data_int1[22]~q ;
wire \data_int[22]~q ;
wire \data_int_selected[22]~6_combout ;
wire \data_int1[23]~q ;
wire \data_int[23]~q ;
wire \data_int_selected[23]~7_combout ;
wire \data_int1[24]~q ;
wire \data_int[24]~q ;
wire \data_int_selected[24]~8_combout ;
wire \data_int1[25]~q ;
wire \data_int[25]~q ;
wire \data_int_selected[25]~9_combout ;
wire \data_int1[26]~q ;
wire \data_int[26]~q ;
wire \data_int_selected[26]~10_combout ;
wire \data_int1[27]~q ;
wire \data_int[27]~q ;
wire \data_int_selected[27]~11_combout ;
wire \data_int1[28]~q ;
wire \data_int[28]~q ;
wire \data_int_selected[28]~12_combout ;
wire \data_int1[29]~q ;
wire \data_int[29]~q ;
wire \data_int_selected[29]~13_combout ;
wire \data_int1[30]~q ;
wire \data_int[30]~q ;
wire \data_int_selected[30]~14_combout ;
wire \data_int1[31]~q ;
wire \data_int[31]~q ;
wire \data_int_selected[31]~15_combout ;
wire \data_int1[32]~q ;
wire \data_int[32]~q ;
wire \data_int_selected[32]~16_combout ;
wire \data_int1[33]~q ;
wire \data_int[33]~q ;
wire \data_int_selected[33]~17_combout ;
wire \data_int1[34]~q ;
wire \data_int[34]~q ;
wire \data_int_selected[34]~18_combout ;
wire \data_int1[35]~q ;
wire \data_int[35]~q ;
wire \data_int_selected[35]~19_combout ;
wire \data_int1[36]~q ;
wire \data_int[36]~q ;
wire \data_int_selected[36]~20_combout ;
wire \data_int1[37]~q ;
wire \data_int[37]~q ;
wire \data_int_selected[37]~21_combout ;
wire \data_int1[6]~q ;
wire \data_int[6]~q ;
wire \data_int_selected[6]~22_combout ;
wire \data_int1[7]~q ;
wire \data_int[7]~q ;
wire \data_int_selected[7]~23_combout ;
wire \data_int1[8]~q ;
wire \data_int[8]~q ;
wire \data_int_selected[8]~24_combout ;
wire \data_int1[9]~q ;
wire \data_int[9]~q ;
wire \data_int_selected[9]~25_combout ;
wire \data_int1[10]~q ;
wire \data_int[10]~q ;
wire \data_int_selected[10]~26_combout ;
wire \data_int1[11]~q ;
wire \data_int[11]~q ;
wire \data_int_selected[11]~27_combout ;
wire \data_int1[12]~q ;
wire \data_int[12]~q ;
wire \data_int_selected[12]~28_combout ;
wire \data_int1[13]~q ;
wire \data_int[13]~q ;
wire \data_int_selected[13]~29_combout ;
wire \data_int1[14]~q ;
wire \data_int[14]~q ;
wire \data_int_selected[14]~30_combout ;
wire \data_int1[15]~q ;
wire \data_int[15]~q ;
wire \data_int_selected[15]~31_combout ;
wire \data_int1[16]~q ;
wire \data_int[16]~q ;
wire \data_int_selected[16]~32_combout ;
wire \data_int1[17]~q ;
wire \data_int[17]~q ;
wire \data_int_selected[17]~33_combout ;
wire \data_int1[18]~q ;
wire \data_int[18]~q ;
wire \data_int_selected[18]~34_combout ;
wire \data_int1[19]~q ;
wire \data_int[19]~q ;
wire \data_int_selected[19]~35_combout ;
wire \data_int1[20]~q ;
wire \data_int[20]~q ;
wire \data_int_selected[20]~36_combout ;
wire \data_int1[21]~q ;
wire \data_int[21]~q ;
wire \data_int_selected[21]~37_combout ;
wire \Mux0~0_combout ;


cycloneive_lcell_comb \Selector1~1 (
	.dataa(\source_state.sop~q ),
	.datab(\Selector1~0_combout ),
	.datac(source_packet_error_0),
	.datad(source_packet_error_1),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
defparam \Selector1~1 .lut_mask = 16'hEFFF;
defparam \Selector1~1 .sum_lutc_input = "datac";

dffeas \data_count_int[4] (
	.clk(clk),
	.d(data_count[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_count_int[4]~q ),
	.prn(vcc));
defparam \data_count_int[4] .is_wysiwyg = "true";
defparam \data_count_int[4] .power_up = "low";

cycloneive_lcell_comb \source_comb_update_2~0 (
	.dataa(\data_count_int[4]~q ),
	.datab(\data_count_int[0]~q ),
	.datac(\data_count_int[6]~q ),
	.datad(\data_count_int[5]~q ),
	.cin(gnd),
	.combout(\source_comb_update_2~0_combout ),
	.cout());
defparam \source_comb_update_2~0 .lut_mask = 16'h7FFF;
defparam \source_comb_update_2~0 .sum_lutc_input = "datac";

dffeas \data_count_int1[4] (
	.clk(clk),
	.d(data_count[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[4]~q ),
	.prn(vcc));
defparam \data_count_int1[4] .is_wysiwyg = "true";
defparam \data_count_int1[4] .power_up = "low";

cycloneive_lcell_comb \source_comb_update_2~1 (
	.dataa(\data_count_int1[4]~q ),
	.datab(\data_count_int1[0]~q ),
	.datac(\data_count_int1[5]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\source_comb_update_2~1_combout ),
	.cout());
defparam \source_comb_update_2~1 .lut_mask = 16'h7F7F;
defparam \source_comb_update_2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \source_comb_update_2~2 (
	.dataa(\data_select~0_combout ),
	.datab(\data_count_int1[6]~q ),
	.datac(\source_comb_update_2~0_combout ),
	.datad(\source_comb_update_2~1_combout ),
	.cin(gnd),
	.combout(\source_comb_update_2~2_combout ),
	.cout());
defparam \source_comb_update_2~2 .lut_mask = 16'hF7B3;
defparam \source_comb_update_2~2 .sum_lutc_input = "datac";

dffeas \data_count_int[7] (
	.clk(clk),
	.d(data_count[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_count_int[7]~q ),
	.prn(vcc));
defparam \data_count_int[7] .is_wysiwyg = "true";
defparam \data_count_int[7] .power_up = "low";

dffeas \data_count_int1[7] (
	.clk(clk),
	.d(data_count[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[7]~q ),
	.prn(vcc));
defparam \data_count_int1[7] .is_wysiwyg = "true";
defparam \data_count_int1[7] .power_up = "low";

cycloneive_lcell_comb \Selector1~3 (
	.dataa(\source_state.sop~q ),
	.datab(gnd),
	.datac(source_packet_error_0),
	.datad(source_packet_error_1),
	.cin(gnd),
	.combout(\Selector1~3_combout ),
	.cout());
defparam \Selector1~3 .lut_mask = 16'hAFFF;
defparam \Selector1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~1 (
	.dataa(master_source_ena),
	.datab(gnd),
	.datac(gnd),
	.datad(\was_stalled~q ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
defparam \Mux2~1 .lut_mask = 16'hAAFF;
defparam \Mux2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~2 (
	.dataa(master_source_ena),
	.datab(source_valid_ctrl_sop),
	.datac(source_stall_reg),
	.datad(\was_stalled~q ),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
defparam \Mux2~2 .lut_mask = 16'hEFFF;
defparam \Mux2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \valid_ctrl_inter~0 (
	.dataa(\valid_ctrl_int~q ),
	.datab(\data_select~0_combout ),
	.datac(\Mux1~0_combout ),
	.datad(\packet_error0~combout ),
	.cin(gnd),
	.combout(\valid_ctrl_inter~0_combout ),
	.cout());
defparam \valid_ctrl_inter~0 .lut_mask = 16'hEFFF;
defparam \valid_ctrl_inter~0 .sum_lutc_input = "datac";

dffeas \source_state.st_err (
	.clk(clk),
	.d(\packet_error0~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\source_state.st_err~q ),
	.prn(vcc));
defparam \source_state.st_err .is_wysiwyg = "true";
defparam \source_state.st_err .power_up = "low";

dffeas \at_source_error[0] (
	.clk(clk),
	.d(source_packet_error_0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_error_0),
	.prn(vcc));
defparam \at_source_error[0] .is_wysiwyg = "true";
defparam \at_source_error[0] .power_up = "low";

dffeas \at_source_error[1] (
	.clk(clk),
	.d(source_packet_error_1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_error_1),
	.prn(vcc));
defparam \at_source_error[1] .is_wysiwyg = "true";
defparam \at_source_error[1] .power_up = "low";

dffeas at_source_sop_s(
	.clk(clk),
	.d(\Selector1~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_sop_s1),
	.prn(vcc));
defparam at_source_sop_s.is_wysiwyg = "true";
defparam at_source_sop_s.power_up = "low";

dffeas at_source_eop_s(
	.clk(clk),
	.d(\Selector5~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_eop_s1),
	.prn(vcc));
defparam at_source_eop_s.is_wysiwyg = "true";
defparam at_source_eop_s.power_up = "low";

dffeas at_source_valid_s(
	.clk(clk),
	.d(\at_source_valid_int~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_valid_s1),
	.prn(vcc));
defparam at_source_valid_s.is_wysiwyg = "true";
defparam at_source_valid_s.power_up = "low";

dffeas \at_source_data[0] (
	.clk(clk),
	.d(\data_int_selected[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_0),
	.prn(vcc));
defparam \at_source_data[0] .is_wysiwyg = "true";
defparam \at_source_data[0] .power_up = "low";

dffeas \at_source_data[1] (
	.clk(clk),
	.d(\data_int_selected[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_1),
	.prn(vcc));
defparam \at_source_data[1] .is_wysiwyg = "true";
defparam \at_source_data[1] .power_up = "low";

dffeas \at_source_data[2] (
	.clk(clk),
	.d(\data_int_selected[2]~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_2),
	.prn(vcc));
defparam \at_source_data[2] .is_wysiwyg = "true";
defparam \at_source_data[2] .power_up = "low";

dffeas \at_source_data[3] (
	.clk(clk),
	.d(\data_int_selected[3]~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_3),
	.prn(vcc));
defparam \at_source_data[3] .is_wysiwyg = "true";
defparam \at_source_data[3] .power_up = "low";

dffeas \at_source_data[4] (
	.clk(clk),
	.d(\data_int_selected[4]~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_4),
	.prn(vcc));
defparam \at_source_data[4] .is_wysiwyg = "true";
defparam \at_source_data[4] .power_up = "low";

dffeas \at_source_data[5] (
	.clk(clk),
	.d(\data_int_selected[5]~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_5),
	.prn(vcc));
defparam \at_source_data[5] .is_wysiwyg = "true";
defparam \at_source_data[5] .power_up = "low";

dffeas \at_source_data[22] (
	.clk(clk),
	.d(\data_int_selected[22]~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_22),
	.prn(vcc));
defparam \at_source_data[22] .is_wysiwyg = "true";
defparam \at_source_data[22] .power_up = "low";

dffeas \at_source_data[23] (
	.clk(clk),
	.d(\data_int_selected[23]~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_23),
	.prn(vcc));
defparam \at_source_data[23] .is_wysiwyg = "true";
defparam \at_source_data[23] .power_up = "low";

dffeas \at_source_data[24] (
	.clk(clk),
	.d(\data_int_selected[24]~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_24),
	.prn(vcc));
defparam \at_source_data[24] .is_wysiwyg = "true";
defparam \at_source_data[24] .power_up = "low";

dffeas \at_source_data[25] (
	.clk(clk),
	.d(\data_int_selected[25]~9_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_25),
	.prn(vcc));
defparam \at_source_data[25] .is_wysiwyg = "true";
defparam \at_source_data[25] .power_up = "low";

dffeas \at_source_data[26] (
	.clk(clk),
	.d(\data_int_selected[26]~10_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_26),
	.prn(vcc));
defparam \at_source_data[26] .is_wysiwyg = "true";
defparam \at_source_data[26] .power_up = "low";

dffeas \at_source_data[27] (
	.clk(clk),
	.d(\data_int_selected[27]~11_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_27),
	.prn(vcc));
defparam \at_source_data[27] .is_wysiwyg = "true";
defparam \at_source_data[27] .power_up = "low";

dffeas \at_source_data[28] (
	.clk(clk),
	.d(\data_int_selected[28]~12_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_28),
	.prn(vcc));
defparam \at_source_data[28] .is_wysiwyg = "true";
defparam \at_source_data[28] .power_up = "low";

dffeas \at_source_data[29] (
	.clk(clk),
	.d(\data_int_selected[29]~13_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_29),
	.prn(vcc));
defparam \at_source_data[29] .is_wysiwyg = "true";
defparam \at_source_data[29] .power_up = "low";

dffeas \at_source_data[30] (
	.clk(clk),
	.d(\data_int_selected[30]~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_30),
	.prn(vcc));
defparam \at_source_data[30] .is_wysiwyg = "true";
defparam \at_source_data[30] .power_up = "low";

dffeas \at_source_data[31] (
	.clk(clk),
	.d(\data_int_selected[31]~15_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_31),
	.prn(vcc));
defparam \at_source_data[31] .is_wysiwyg = "true";
defparam \at_source_data[31] .power_up = "low";

dffeas \at_source_data[32] (
	.clk(clk),
	.d(\data_int_selected[32]~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_32),
	.prn(vcc));
defparam \at_source_data[32] .is_wysiwyg = "true";
defparam \at_source_data[32] .power_up = "low";

dffeas \at_source_data[33] (
	.clk(clk),
	.d(\data_int_selected[33]~17_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_33),
	.prn(vcc));
defparam \at_source_data[33] .is_wysiwyg = "true";
defparam \at_source_data[33] .power_up = "low";

dffeas \at_source_data[34] (
	.clk(clk),
	.d(\data_int_selected[34]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_34),
	.prn(vcc));
defparam \at_source_data[34] .is_wysiwyg = "true";
defparam \at_source_data[34] .power_up = "low";

dffeas \at_source_data[35] (
	.clk(clk),
	.d(\data_int_selected[35]~19_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_35),
	.prn(vcc));
defparam \at_source_data[35] .is_wysiwyg = "true";
defparam \at_source_data[35] .power_up = "low";

dffeas \at_source_data[36] (
	.clk(clk),
	.d(\data_int_selected[36]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_36),
	.prn(vcc));
defparam \at_source_data[36] .is_wysiwyg = "true";
defparam \at_source_data[36] .power_up = "low";

dffeas \at_source_data[37] (
	.clk(clk),
	.d(\data_int_selected[37]~21_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_37),
	.prn(vcc));
defparam \at_source_data[37] .is_wysiwyg = "true";
defparam \at_source_data[37] .power_up = "low";

dffeas \at_source_data[6] (
	.clk(clk),
	.d(\data_int_selected[6]~22_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_6),
	.prn(vcc));
defparam \at_source_data[6] .is_wysiwyg = "true";
defparam \at_source_data[6] .power_up = "low";

dffeas \at_source_data[7] (
	.clk(clk),
	.d(\data_int_selected[7]~23_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_7),
	.prn(vcc));
defparam \at_source_data[7] .is_wysiwyg = "true";
defparam \at_source_data[7] .power_up = "low";

dffeas \at_source_data[8] (
	.clk(clk),
	.d(\data_int_selected[8]~24_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_8),
	.prn(vcc));
defparam \at_source_data[8] .is_wysiwyg = "true";
defparam \at_source_data[8] .power_up = "low";

dffeas \at_source_data[9] (
	.clk(clk),
	.d(\data_int_selected[9]~25_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_9),
	.prn(vcc));
defparam \at_source_data[9] .is_wysiwyg = "true";
defparam \at_source_data[9] .power_up = "low";

dffeas \at_source_data[10] (
	.clk(clk),
	.d(\data_int_selected[10]~26_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_10),
	.prn(vcc));
defparam \at_source_data[10] .is_wysiwyg = "true";
defparam \at_source_data[10] .power_up = "low";

dffeas \at_source_data[11] (
	.clk(clk),
	.d(\data_int_selected[11]~27_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_11),
	.prn(vcc));
defparam \at_source_data[11] .is_wysiwyg = "true";
defparam \at_source_data[11] .power_up = "low";

dffeas \at_source_data[12] (
	.clk(clk),
	.d(\data_int_selected[12]~28_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_12),
	.prn(vcc));
defparam \at_source_data[12] .is_wysiwyg = "true";
defparam \at_source_data[12] .power_up = "low";

dffeas \at_source_data[13] (
	.clk(clk),
	.d(\data_int_selected[13]~29_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_13),
	.prn(vcc));
defparam \at_source_data[13] .is_wysiwyg = "true";
defparam \at_source_data[13] .power_up = "low";

dffeas \at_source_data[14] (
	.clk(clk),
	.d(\data_int_selected[14]~30_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_14),
	.prn(vcc));
defparam \at_source_data[14] .is_wysiwyg = "true";
defparam \at_source_data[14] .power_up = "low";

dffeas \at_source_data[15] (
	.clk(clk),
	.d(\data_int_selected[15]~31_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_15),
	.prn(vcc));
defparam \at_source_data[15] .is_wysiwyg = "true";
defparam \at_source_data[15] .power_up = "low";

dffeas \at_source_data[16] (
	.clk(clk),
	.d(\data_int_selected[16]~32_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_16),
	.prn(vcc));
defparam \at_source_data[16] .is_wysiwyg = "true";
defparam \at_source_data[16] .power_up = "low";

dffeas \at_source_data[17] (
	.clk(clk),
	.d(\data_int_selected[17]~33_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_17),
	.prn(vcc));
defparam \at_source_data[17] .is_wysiwyg = "true";
defparam \at_source_data[17] .power_up = "low";

dffeas \at_source_data[18] (
	.clk(clk),
	.d(\data_int_selected[18]~34_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_18),
	.prn(vcc));
defparam \at_source_data[18] .is_wysiwyg = "true";
defparam \at_source_data[18] .power_up = "low";

dffeas \at_source_data[19] (
	.clk(clk),
	.d(\data_int_selected[19]~35_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_19),
	.prn(vcc));
defparam \at_source_data[19] .is_wysiwyg = "true";
defparam \at_source_data[19] .power_up = "low";

dffeas \at_source_data[20] (
	.clk(clk),
	.d(\data_int_selected[20]~36_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_20),
	.prn(vcc));
defparam \at_source_data[20] .is_wysiwyg = "true";
defparam \at_source_data[20] .power_up = "low";

dffeas \at_source_data[21] (
	.clk(clk),
	.d(\data_int_selected[21]~37_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_21),
	.prn(vcc));
defparam \at_source_data[21] .is_wysiwyg = "true";
defparam \at_source_data[21] .power_up = "low";

dffeas source_stall_int_d(
	.clk(clk),
	.d(Mux0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(source_stall_int_d1),
	.prn(vcc));
defparam source_stall_int_d.is_wysiwyg = "true";
defparam source_stall_int_d.power_up = "low";

cycloneive_lcell_comb \Mux0~1 (
	.dataa(\valid_ctrl_int~q ),
	.datab(\Mux3~0_combout ),
	.datac(\valid_ctrl_int1~q ),
	.datad(\Mux0~0_combout ),
	.cin(gnd),
	.combout(Mux0),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hFFFE;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \first_data~0 (
	.dataa(\valid_ctrl_int1~q ),
	.datab(\first_data~q ),
	.datac(at_source_valid_s1),
	.datad(source_ready),
	.cin(gnd),
	.combout(\first_data~0_combout ),
	.cout());
defparam \first_data~0 .lut_mask = 16'hEBBE;
defparam \first_data~0 .sum_lutc_input = "datac";

dffeas first_data(
	.clk(clk),
	.d(\first_data~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\first_data~q ),
	.prn(vcc));
defparam first_data.is_wysiwyg = "true";
defparam first_data.power_up = "low";

cycloneive_lcell_comb \data_select~0 (
	.dataa(at_source_valid_s1),
	.datab(\first_data~q ),
	.datac(\valid_ctrl_int1~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_select~0_combout ),
	.cout());
defparam \data_select~0 .lut_mask = 16'hFEFE;
defparam \data_select~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~3 (
	.dataa(source_ready),
	.datab(at_source_valid_s1),
	.datac(\first_data~q ),
	.datad(\valid_ctrl_int1~q ),
	.cin(gnd),
	.combout(\Mux2~3_combout ),
	.cout());
defparam \Mux2~3 .lut_mask = 16'hFEFF;
defparam \Mux2~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~0 (
	.dataa(at_source_valid_s1),
	.datab(\valid_ctrl_int~q ),
	.datac(\valid_ctrl_int1~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFEFE;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~4 (
	.dataa(\Mux2~2_combout ),
	.datab(\Mux2~3_combout ),
	.datac(gnd),
	.datad(\Mux2~0_combout ),
	.cin(gnd),
	.combout(\Mux2~4_combout ),
	.cout());
defparam \Mux2~4 .lut_mask = 16'hEEFF;
defparam \Mux2~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \was_stalled~0 (
	.dataa(source_valid_ctrl_sop1),
	.datab(stall_reg),
	.datac(gnd),
	.datad(source_stall_int_d1),
	.cin(gnd),
	.combout(\was_stalled~0_combout ),
	.cout());
defparam \was_stalled~0 .lut_mask = 16'hEEFF;
defparam \was_stalled~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \was_stalled~1 (
	.dataa(\was_stalled~q ),
	.datab(\Mux2~4_combout ),
	.datac(\Mux3~1_combout ),
	.datad(\was_stalled~0_combout ),
	.cin(gnd),
	.combout(\was_stalled~1_combout ),
	.cout());
defparam \was_stalled~1 .lut_mask = 16'hFEFF;
defparam \was_stalled~1 .sum_lutc_input = "datac";

dffeas was_stalled(
	.clk(clk),
	.d(\was_stalled~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\was_stalled~q ),
	.prn(vcc));
defparam was_stalled.is_wysiwyg = "true";
defparam was_stalled.power_up = "low";

cycloneive_lcell_comb \valid_ctrl_inter~1 (
	.dataa(\valid_ctrl_inter~0_combout ),
	.datab(\Mux2~4_combout ),
	.datac(\was_stalled~q ),
	.datad(\was_stalled~0_combout ),
	.cin(gnd),
	.combout(\valid_ctrl_inter~1_combout ),
	.cout());
defparam \valid_ctrl_inter~1 .lut_mask = 16'h8BFF;
defparam \valid_ctrl_inter~1 .sum_lutc_input = "datac";

dffeas valid_ctrl_int(
	.clk(clk),
	.d(\valid_ctrl_inter~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\valid_ctrl_int~q ),
	.prn(vcc));
defparam valid_ctrl_int.is_wysiwyg = "true";
defparam valid_ctrl_int.power_up = "low";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(source_ready),
	.datab(\valid_ctrl_int~q ),
	.datac(\valid_ctrl_int1~q ),
	.datad(at_source_valid_s1),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hFAFC;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \valid_ctrl_inter1~0 (
	.dataa(\Mux3~1_combout ),
	.datab(\valid_ctrl_int1~q ),
	.datac(\data_select~0_combout ),
	.datad(\Mux1~0_combout ),
	.cin(gnd),
	.combout(\valid_ctrl_inter1~0_combout ),
	.cout());
defparam \valid_ctrl_inter1~0 .lut_mask = 16'hEFFF;
defparam \valid_ctrl_inter1~0 .sum_lutc_input = "datac";

dffeas valid_ctrl_int1(
	.clk(clk),
	.d(\valid_ctrl_inter1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\valid_ctrl_int1~q ),
	.prn(vcc));
defparam valid_ctrl_int1.is_wysiwyg = "true";
defparam valid_ctrl_int1.power_up = "low";

cycloneive_lcell_comb \Mux3~0 (
	.dataa(\Mux2~1_combout ),
	.datab(source_valid_ctrl_sop),
	.datac(source_stall_reg),
	.datad(\valid_ctrl_int1~q ),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hEFFF;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~1 (
	.dataa(\Mux2~0_combout ),
	.datab(\Mux3~0_combout ),
	.datac(gnd),
	.datad(source_ready),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
defparam \Mux3~1 .lut_mask = 16'hEEFF;
defparam \Mux3~1 .sum_lutc_input = "datac";

dffeas \data_count_int1[1] (
	.clk(clk),
	.d(data_count[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[1]~q ),
	.prn(vcc));
defparam \data_count_int1[1] .is_wysiwyg = "true";
defparam \data_count_int1[1] .power_up = "low";

dffeas \data_count_int[3] (
	.clk(clk),
	.d(data_count[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_count_int[3]~q ),
	.prn(vcc));
defparam \data_count_int[3] .is_wysiwyg = "true";
defparam \data_count_int[3] .power_up = "low";

dffeas \data_count_int[1] (
	.clk(clk),
	.d(data_count[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_count_int[1]~q ),
	.prn(vcc));
defparam \data_count_int[1] .is_wysiwyg = "true";
defparam \data_count_int[1] .power_up = "low";

dffeas \data_count_int[2] (
	.clk(clk),
	.d(data_count[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_count_int[2]~q ),
	.prn(vcc));
defparam \data_count_int[2] .is_wysiwyg = "true";
defparam \data_count_int[2] .power_up = "low";

cycloneive_lcell_comb \source_comb_update_2~3 (
	.dataa(\data_count_int[7]~q ),
	.datab(\data_count_int[3]~q ),
	.datac(\data_count_int[1]~q ),
	.datad(\data_count_int[2]~q ),
	.cin(gnd),
	.combout(\source_comb_update_2~3_combout ),
	.cout());
defparam \source_comb_update_2~3 .lut_mask = 16'h7FFF;
defparam \source_comb_update_2~3 .sum_lutc_input = "datac";

dffeas \data_count_int1[3] (
	.clk(clk),
	.d(data_count[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[3]~q ),
	.prn(vcc));
defparam \data_count_int1[3] .is_wysiwyg = "true";
defparam \data_count_int1[3] .power_up = "low";

dffeas \data_count_int1[2] (
	.clk(clk),
	.d(data_count[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[2]~q ),
	.prn(vcc));
defparam \data_count_int1[2] .is_wysiwyg = "true";
defparam \data_count_int1[2] .power_up = "low";

cycloneive_lcell_comb \source_comb_update_2~4 (
	.dataa(\data_count_int1[7]~q ),
	.datab(\data_count_int1[3]~q ),
	.datac(\data_count_int1[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\source_comb_update_2~4_combout ),
	.cout());
defparam \source_comb_update_2~4 .lut_mask = 16'h7F7F;
defparam \source_comb_update_2~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \source_comb_update_2~5 (
	.dataa(\data_select~0_combout ),
	.datab(\data_count_int1[1]~q ),
	.datac(\source_comb_update_2~3_combout ),
	.datad(\source_comb_update_2~4_combout ),
	.cin(gnd),
	.combout(\source_comb_update_2~5_combout ),
	.cout());
defparam \source_comb_update_2~5 .lut_mask = 16'hF7B3;
defparam \source_comb_update_2~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \source_comb_update_2~6 (
	.dataa(\source_comb_update_2~2_combout ),
	.datab(\source_comb_update_2~5_combout ),
	.datac(\valid_ctrl_int~q ),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\source_comb_update_2~6_combout ),
	.cout());
defparam \source_comb_update_2~6 .lut_mask = 16'hFFFE;
defparam \source_comb_update_2~6 .sum_lutc_input = "datac";

dffeas \data_count_int1[6] (
	.clk(clk),
	.d(data_count[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[6]~q ),
	.prn(vcc));
defparam \data_count_int1[6] .is_wysiwyg = "true";
defparam \data_count_int1[6] .power_up = "low";

dffeas \data_count_int[5] (
	.clk(clk),
	.d(data_count[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_count_int[5]~q ),
	.prn(vcc));
defparam \data_count_int[5] .is_wysiwyg = "true";
defparam \data_count_int[5] .power_up = "low";

dffeas \data_count_int[0] (
	.clk(clk),
	.d(data_count[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_count_int[0]~q ),
	.prn(vcc));
defparam \data_count_int[0] .is_wysiwyg = "true";
defparam \data_count_int[0] .power_up = "low";

dffeas \data_count_int[6] (
	.clk(clk),
	.d(data_count[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_count_int[6]~q ),
	.prn(vcc));
defparam \data_count_int[6] .is_wysiwyg = "true";
defparam \data_count_int[6] .power_up = "low";

cycloneive_lcell_comb \count_finished~0 (
	.dataa(\data_count_int[4]~q ),
	.datab(\data_count_int[5]~q ),
	.datac(\data_count_int[0]~q ),
	.datad(\data_count_int[6]~q ),
	.cin(gnd),
	.combout(\count_finished~0_combout ),
	.cout());
defparam \count_finished~0 .lut_mask = 16'h7FFF;
defparam \count_finished~0 .sum_lutc_input = "datac";

dffeas \data_count_int1[5] (
	.clk(clk),
	.d(data_count[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[5]~q ),
	.prn(vcc));
defparam \data_count_int1[5] .is_wysiwyg = "true";
defparam \data_count_int1[5] .power_up = "low";

dffeas \data_count_int1[0] (
	.clk(clk),
	.d(data_count[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[0]~q ),
	.prn(vcc));
defparam \data_count_int1[0] .is_wysiwyg = "true";
defparam \data_count_int1[0] .power_up = "low";

cycloneive_lcell_comb \count_finished~1 (
	.dataa(\data_count_int1[4]~q ),
	.datab(\data_count_int1[5]~q ),
	.datac(\data_count_int1[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_finished~1_combout ),
	.cout());
defparam \count_finished~1 .lut_mask = 16'h7F7F;
defparam \count_finished~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count_finished~2 (
	.dataa(\data_select~0_combout ),
	.datab(\data_count_int1[6]~q ),
	.datac(\count_finished~0_combout ),
	.datad(\count_finished~1_combout ),
	.cin(gnd),
	.combout(\count_finished~2_combout ),
	.cout());
defparam \count_finished~2 .lut_mask = 16'hF7B3;
defparam \count_finished~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count_finished~3 (
	.dataa(\data_count_int[7]~q ),
	.datab(\data_count_int[1]~q ),
	.datac(\data_count_int[3]~q ),
	.datad(\data_count_int[2]~q ),
	.cin(gnd),
	.combout(\count_finished~3_combout ),
	.cout());
defparam \count_finished~3 .lut_mask = 16'h7FFF;
defparam \count_finished~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count_finished~4 (
	.dataa(\data_count_int1[7]~q ),
	.datab(\data_count_int1[3]~q ),
	.datac(\data_count_int1[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\count_finished~4_combout ),
	.cout());
defparam \count_finished~4 .lut_mask = 16'h7F7F;
defparam \count_finished~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count_finished~5 (
	.dataa(\data_select~0_combout ),
	.datab(\data_count_int1[1]~q ),
	.datac(\count_finished~3_combout ),
	.datad(\count_finished~4_combout ),
	.cin(gnd),
	.combout(\count_finished~5_combout ),
	.cout());
defparam \count_finished~5 .lut_mask = 16'hF7B3;
defparam \count_finished~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~0 (
	.dataa(at_source_valid_s1),
	.datab(gnd),
	.datac(gnd),
	.datad(source_ready),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hAAFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \source_comb_update_2~7 (
	.dataa(\valid_ctrl_int_selected~0_combout ),
	.datab(\count_finished~2_combout ),
	.datac(\count_finished~5_combout ),
	.datad(\Selector1~0_combout ),
	.cin(gnd),
	.combout(\source_comb_update_2~7_combout ),
	.cout());
defparam \source_comb_update_2~7 .lut_mask = 16'hBFFF;
defparam \source_comb_update_2~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~4 (
	.dataa(source_packet_error_0),
	.datab(source_packet_error_1),
	.datac(\source_comb_update_2~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector2~4_combout ),
	.cout());
defparam \Selector2~4 .lut_mask = 16'h7F7F;
defparam \Selector2~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~5 (
	.dataa(at_source_valid_s1),
	.datab(source_ready),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector1~5_combout ),
	.cout());
defparam \Selector1~5 .lut_mask = 16'hEEEE;
defparam \Selector1~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~3 (
	.dataa(\Selector2~2_combout ),
	.datab(\source_state.run1~q ),
	.datac(\Selector2~4_combout ),
	.datad(\Selector1~5_combout ),
	.cin(gnd),
	.combout(\Selector2~3_combout ),
	.cout());
defparam \Selector2~3 .lut_mask = 16'hFFFE;
defparam \Selector2~3 .sum_lutc_input = "datac";

dffeas \source_state.run1 (
	.clk(clk),
	.d(\Selector2~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\source_state.run1~q ),
	.prn(vcc));
defparam \source_state.run1 .is_wysiwyg = "true";
defparam \source_state.run1 .power_up = "low";

cycloneive_lcell_comb \Selector3~0 (
	.dataa(\source_state.sop~q ),
	.datab(\source_state.run1~q ),
	.datac(source_packet_error_0),
	.datad(source_packet_error_1),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'hEFFF;
defparam \Selector3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~1 (
	.dataa(at_source_valid_s1),
	.datab(source_ready),
	.datac(source_packet_error_0),
	.datad(source_packet_error_1),
	.cin(gnd),
	.combout(\Selector3~1_combout ),
	.cout());
defparam \Selector3~1 .lut_mask = 16'h7FFF;
defparam \Selector3~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~2 (
	.dataa(\source_state.end1~q ),
	.datab(\source_comb_update_2~7_combout ),
	.datac(\Selector3~0_combout ),
	.datad(\Selector3~1_combout ),
	.cin(gnd),
	.combout(\Selector3~2_combout ),
	.cout());
defparam \Selector3~2 .lut_mask = 16'hFFFE;
defparam \Selector3~2 .sum_lutc_input = "datac";

dffeas \source_state.end1 (
	.clk(clk),
	.d(\Selector3~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\source_state.end1~q ),
	.prn(vcc));
defparam \source_state.end1 .is_wysiwyg = "true";
defparam \source_state.end1 .power_up = "low";

cycloneive_lcell_comb packet_error0(
	.dataa(source_packet_error_0),
	.datab(source_packet_error_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_error0~combout ),
	.cout());
defparam packet_error0.lut_mask = 16'hEEEE;
defparam packet_error0.sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector0~1 (
	.dataa(\source_state.st_err~q ),
	.datab(\Selector0~0_combout ),
	.datac(\source_comb_update_2~6_combout ),
	.datad(\packet_error0~combout ),
	.cin(gnd),
	.combout(\Selector0~1_combout ),
	.cout());
defparam \Selector0~1 .lut_mask = 16'hFFF7;
defparam \Selector0~1 .sum_lutc_input = "datac";

dffeas \source_state.start (
	.clk(clk),
	.d(\Selector0~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\source_state.start~q ),
	.prn(vcc));
defparam \source_state.start .is_wysiwyg = "true";
defparam \source_state.start .power_up = "low";

cycloneive_lcell_comb \Selector0~0 (
	.dataa(at_source_valid_s1),
	.datab(source_ready),
	.datac(\source_state.end1~q ),
	.datad(\source_state.start~q ),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hFEFF;
defparam \Selector0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~2 (
	.dataa(\Selector1~1_combout ),
	.datab(\source_comb_update_2~6_combout ),
	.datac(\Selector0~0_combout ),
	.datad(\packet_error0~combout ),
	.cin(gnd),
	.combout(\Selector1~2_combout ),
	.cout());
defparam \Selector1~2 .lut_mask = 16'hFEFF;
defparam \Selector1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \valid_ctrl_int_selected~0 (
	.dataa(\valid_ctrl_int~q ),
	.datab(at_source_valid_s1),
	.datac(\first_data~q ),
	.datad(\valid_ctrl_int1~q ),
	.cin(gnd),
	.combout(\valid_ctrl_int_selected~0_combout ),
	.cout());
defparam \valid_ctrl_int_selected~0 .lut_mask = 16'hFFFE;
defparam \valid_ctrl_int_selected~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~2 (
	.dataa(\Selector1~3_combout ),
	.datab(\count_finished~2_combout ),
	.datac(\count_finished~5_combout ),
	.datad(\valid_ctrl_int_selected~0_combout ),
	.cin(gnd),
	.combout(\Selector2~2_combout ),
	.cout());
defparam \Selector2~2 .lut_mask = 16'hFEFF;
defparam \Selector2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~4 (
	.dataa(\Selector1~2_combout ),
	.datab(\Selector2~2_combout ),
	.datac(gnd),
	.datad(at_source_valid_s1),
	.cin(gnd),
	.combout(\Selector1~4_combout ),
	.cout());
defparam \Selector1~4 .lut_mask = 16'hEEFF;
defparam \Selector1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector5~0 (
	.dataa(\packet_error0~combout ),
	.datab(\source_state.end1~q ),
	.datac(\source_state.start~q ),
	.datad(\Selector1~5_combout ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hEFFF;
defparam \Selector5~0 .sum_lutc_input = "datac";

dffeas \source_state.sop (
	.clk(clk),
	.d(\Selector1~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\source_state.sop~q ),
	.prn(vcc));
defparam \source_state.sop .is_wysiwyg = "true";
defparam \source_state.sop .power_up = "low";

cycloneive_lcell_comb \Selector5~1 (
	.dataa(\Selector5~0_combout ),
	.datab(\source_state.sop~q ),
	.datac(\source_state.run1~q ),
	.datad(\Selector2~4_combout ),
	.cin(gnd),
	.combout(\Selector5~1_combout ),
	.cout());
defparam \Selector5~1 .lut_mask = 16'hFEFF;
defparam \Selector5~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \at_source_valid_int~0 (
	.dataa(at_source_valid_s1),
	.datab(source_packet_error_0),
	.datac(source_packet_error_1),
	.datad(source_ready),
	.cin(gnd),
	.combout(\at_source_valid_int~0_combout ),
	.cout());
defparam \at_source_valid_int~0 .lut_mask = 16'hBFFF;
defparam \at_source_valid_int~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \at_source_valid_int~1 (
	.dataa(at_source_valid_s1),
	.datab(\Selector1~4_combout ),
	.datac(\Selector2~3_combout ),
	.datad(\Selector3~2_combout ),
	.cin(gnd),
	.combout(\at_source_valid_int~1_combout ),
	.cout());
defparam \at_source_valid_int~1 .lut_mask = 16'hFFFE;
defparam \at_source_valid_int~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \at_source_valid_int~2 (
	.dataa(\at_source_valid_int~0_combout ),
	.datab(\valid_ctrl_int_selected~0_combout ),
	.datac(\at_source_valid_int~1_combout ),
	.datad(\packet_error0~combout ),
	.cin(gnd),
	.combout(\at_source_valid_int~2_combout ),
	.cout());
defparam \at_source_valid_int~2 .lut_mask = 16'hFEFF;
defparam \at_source_valid_int~2 .sum_lutc_input = "datac";

dffeas \data_int1[0] (
	.clk(clk),
	.d(data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[0]~q ),
	.prn(vcc));
defparam \data_int1[0] .is_wysiwyg = "true";
defparam \data_int1[0] .power_up = "low";

dffeas \data_int[0] (
	.clk(clk),
	.d(data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[0]~q ),
	.prn(vcc));
defparam \data_int[0] .is_wysiwyg = "true";
defparam \data_int[0] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[0]~0 (
	.dataa(\data_int1[0]~q ),
	.datab(\data_int[0]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[0]~0_combout ),
	.cout());
defparam \data_int_selected[0]~0 .lut_mask = 16'hAACC;
defparam \data_int_selected[0]~0 .sum_lutc_input = "datac";

dffeas \data_int1[1] (
	.clk(clk),
	.d(data[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[1]~q ),
	.prn(vcc));
defparam \data_int1[1] .is_wysiwyg = "true";
defparam \data_int1[1] .power_up = "low";

dffeas \data_int[1] (
	.clk(clk),
	.d(data[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[1]~q ),
	.prn(vcc));
defparam \data_int[1] .is_wysiwyg = "true";
defparam \data_int[1] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[1]~1 (
	.dataa(\data_int1[1]~q ),
	.datab(\data_int[1]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[1]~1_combout ),
	.cout());
defparam \data_int_selected[1]~1 .lut_mask = 16'hAACC;
defparam \data_int_selected[1]~1 .sum_lutc_input = "datac";

dffeas \data_int1[2] (
	.clk(clk),
	.d(data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[2]~q ),
	.prn(vcc));
defparam \data_int1[2] .is_wysiwyg = "true";
defparam \data_int1[2] .power_up = "low";

dffeas \data_int[2] (
	.clk(clk),
	.d(data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[2]~q ),
	.prn(vcc));
defparam \data_int[2] .is_wysiwyg = "true";
defparam \data_int[2] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[2]~2 (
	.dataa(\data_int1[2]~q ),
	.datab(\data_int[2]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[2]~2_combout ),
	.cout());
defparam \data_int_selected[2]~2 .lut_mask = 16'hAACC;
defparam \data_int_selected[2]~2 .sum_lutc_input = "datac";

dffeas \data_int1[3] (
	.clk(clk),
	.d(data[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[3]~q ),
	.prn(vcc));
defparam \data_int1[3] .is_wysiwyg = "true";
defparam \data_int1[3] .power_up = "low";

dffeas \data_int[3] (
	.clk(clk),
	.d(data[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[3]~q ),
	.prn(vcc));
defparam \data_int[3] .is_wysiwyg = "true";
defparam \data_int[3] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[3]~3 (
	.dataa(\data_int1[3]~q ),
	.datab(\data_int[3]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[3]~3_combout ),
	.cout());
defparam \data_int_selected[3]~3 .lut_mask = 16'hAACC;
defparam \data_int_selected[3]~3 .sum_lutc_input = "datac";

dffeas \data_int1[4] (
	.clk(clk),
	.d(data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[4]~q ),
	.prn(vcc));
defparam \data_int1[4] .is_wysiwyg = "true";
defparam \data_int1[4] .power_up = "low";

dffeas \data_int[4] (
	.clk(clk),
	.d(data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[4]~q ),
	.prn(vcc));
defparam \data_int[4] .is_wysiwyg = "true";
defparam \data_int[4] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[4]~4 (
	.dataa(\data_int1[4]~q ),
	.datab(\data_int[4]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[4]~4_combout ),
	.cout());
defparam \data_int_selected[4]~4 .lut_mask = 16'hAACC;
defparam \data_int_selected[4]~4 .sum_lutc_input = "datac";

dffeas \data_int1[5] (
	.clk(clk),
	.d(data[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[5]~q ),
	.prn(vcc));
defparam \data_int1[5] .is_wysiwyg = "true";
defparam \data_int1[5] .power_up = "low";

dffeas \data_int[5] (
	.clk(clk),
	.d(data[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[5]~q ),
	.prn(vcc));
defparam \data_int[5] .is_wysiwyg = "true";
defparam \data_int[5] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[5]~5 (
	.dataa(\data_int1[5]~q ),
	.datab(\data_int[5]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[5]~5_combout ),
	.cout());
defparam \data_int_selected[5]~5 .lut_mask = 16'hAACC;
defparam \data_int_selected[5]~5 .sum_lutc_input = "datac";

dffeas \data_int1[22] (
	.clk(clk),
	.d(data[22]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[22]~q ),
	.prn(vcc));
defparam \data_int1[22] .is_wysiwyg = "true";
defparam \data_int1[22] .power_up = "low";

dffeas \data_int[22] (
	.clk(clk),
	.d(data[22]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[22]~q ),
	.prn(vcc));
defparam \data_int[22] .is_wysiwyg = "true";
defparam \data_int[22] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[22]~6 (
	.dataa(\data_int1[22]~q ),
	.datab(\data_int[22]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[22]~6_combout ),
	.cout());
defparam \data_int_selected[22]~6 .lut_mask = 16'hAACC;
defparam \data_int_selected[22]~6 .sum_lutc_input = "datac";

dffeas \data_int1[23] (
	.clk(clk),
	.d(data[23]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[23]~q ),
	.prn(vcc));
defparam \data_int1[23] .is_wysiwyg = "true";
defparam \data_int1[23] .power_up = "low";

dffeas \data_int[23] (
	.clk(clk),
	.d(data[23]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[23]~q ),
	.prn(vcc));
defparam \data_int[23] .is_wysiwyg = "true";
defparam \data_int[23] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[23]~7 (
	.dataa(\data_int1[23]~q ),
	.datab(\data_int[23]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[23]~7_combout ),
	.cout());
defparam \data_int_selected[23]~7 .lut_mask = 16'hAACC;
defparam \data_int_selected[23]~7 .sum_lutc_input = "datac";

dffeas \data_int1[24] (
	.clk(clk),
	.d(data[24]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[24]~q ),
	.prn(vcc));
defparam \data_int1[24] .is_wysiwyg = "true";
defparam \data_int1[24] .power_up = "low";

dffeas \data_int[24] (
	.clk(clk),
	.d(data[24]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[24]~q ),
	.prn(vcc));
defparam \data_int[24] .is_wysiwyg = "true";
defparam \data_int[24] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[24]~8 (
	.dataa(\data_int1[24]~q ),
	.datab(\data_int[24]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[24]~8_combout ),
	.cout());
defparam \data_int_selected[24]~8 .lut_mask = 16'hAACC;
defparam \data_int_selected[24]~8 .sum_lutc_input = "datac";

dffeas \data_int1[25] (
	.clk(clk),
	.d(data[25]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[25]~q ),
	.prn(vcc));
defparam \data_int1[25] .is_wysiwyg = "true";
defparam \data_int1[25] .power_up = "low";

dffeas \data_int[25] (
	.clk(clk),
	.d(data[25]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[25]~q ),
	.prn(vcc));
defparam \data_int[25] .is_wysiwyg = "true";
defparam \data_int[25] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[25]~9 (
	.dataa(\data_int1[25]~q ),
	.datab(\data_int[25]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[25]~9_combout ),
	.cout());
defparam \data_int_selected[25]~9 .lut_mask = 16'hAACC;
defparam \data_int_selected[25]~9 .sum_lutc_input = "datac";

dffeas \data_int1[26] (
	.clk(clk),
	.d(data[26]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[26]~q ),
	.prn(vcc));
defparam \data_int1[26] .is_wysiwyg = "true";
defparam \data_int1[26] .power_up = "low";

dffeas \data_int[26] (
	.clk(clk),
	.d(data[26]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[26]~q ),
	.prn(vcc));
defparam \data_int[26] .is_wysiwyg = "true";
defparam \data_int[26] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[26]~10 (
	.dataa(\data_int1[26]~q ),
	.datab(\data_int[26]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[26]~10_combout ),
	.cout());
defparam \data_int_selected[26]~10 .lut_mask = 16'hAACC;
defparam \data_int_selected[26]~10 .sum_lutc_input = "datac";

dffeas \data_int1[27] (
	.clk(clk),
	.d(data[27]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[27]~q ),
	.prn(vcc));
defparam \data_int1[27] .is_wysiwyg = "true";
defparam \data_int1[27] .power_up = "low";

dffeas \data_int[27] (
	.clk(clk),
	.d(data[27]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[27]~q ),
	.prn(vcc));
defparam \data_int[27] .is_wysiwyg = "true";
defparam \data_int[27] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[27]~11 (
	.dataa(\data_int1[27]~q ),
	.datab(\data_int[27]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[27]~11_combout ),
	.cout());
defparam \data_int_selected[27]~11 .lut_mask = 16'hAACC;
defparam \data_int_selected[27]~11 .sum_lutc_input = "datac";

dffeas \data_int1[28] (
	.clk(clk),
	.d(data[28]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[28]~q ),
	.prn(vcc));
defparam \data_int1[28] .is_wysiwyg = "true";
defparam \data_int1[28] .power_up = "low";

dffeas \data_int[28] (
	.clk(clk),
	.d(data[28]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[28]~q ),
	.prn(vcc));
defparam \data_int[28] .is_wysiwyg = "true";
defparam \data_int[28] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[28]~12 (
	.dataa(\data_int1[28]~q ),
	.datab(\data_int[28]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[28]~12_combout ),
	.cout());
defparam \data_int_selected[28]~12 .lut_mask = 16'hAACC;
defparam \data_int_selected[28]~12 .sum_lutc_input = "datac";

dffeas \data_int1[29] (
	.clk(clk),
	.d(data[29]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[29]~q ),
	.prn(vcc));
defparam \data_int1[29] .is_wysiwyg = "true";
defparam \data_int1[29] .power_up = "low";

dffeas \data_int[29] (
	.clk(clk),
	.d(data[29]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[29]~q ),
	.prn(vcc));
defparam \data_int[29] .is_wysiwyg = "true";
defparam \data_int[29] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[29]~13 (
	.dataa(\data_int1[29]~q ),
	.datab(\data_int[29]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[29]~13_combout ),
	.cout());
defparam \data_int_selected[29]~13 .lut_mask = 16'hAACC;
defparam \data_int_selected[29]~13 .sum_lutc_input = "datac";

dffeas \data_int1[30] (
	.clk(clk),
	.d(data[30]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[30]~q ),
	.prn(vcc));
defparam \data_int1[30] .is_wysiwyg = "true";
defparam \data_int1[30] .power_up = "low";

dffeas \data_int[30] (
	.clk(clk),
	.d(data[30]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[30]~q ),
	.prn(vcc));
defparam \data_int[30] .is_wysiwyg = "true";
defparam \data_int[30] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[30]~14 (
	.dataa(\data_int1[30]~q ),
	.datab(\data_int[30]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[30]~14_combout ),
	.cout());
defparam \data_int_selected[30]~14 .lut_mask = 16'hAACC;
defparam \data_int_selected[30]~14 .sum_lutc_input = "datac";

dffeas \data_int1[31] (
	.clk(clk),
	.d(data[31]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[31]~q ),
	.prn(vcc));
defparam \data_int1[31] .is_wysiwyg = "true";
defparam \data_int1[31] .power_up = "low";

dffeas \data_int[31] (
	.clk(clk),
	.d(data[31]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[31]~q ),
	.prn(vcc));
defparam \data_int[31] .is_wysiwyg = "true";
defparam \data_int[31] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[31]~15 (
	.dataa(\data_int1[31]~q ),
	.datab(\data_int[31]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[31]~15_combout ),
	.cout());
defparam \data_int_selected[31]~15 .lut_mask = 16'hAACC;
defparam \data_int_selected[31]~15 .sum_lutc_input = "datac";

dffeas \data_int1[32] (
	.clk(clk),
	.d(data[32]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[32]~q ),
	.prn(vcc));
defparam \data_int1[32] .is_wysiwyg = "true";
defparam \data_int1[32] .power_up = "low";

dffeas \data_int[32] (
	.clk(clk),
	.d(data[32]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[32]~q ),
	.prn(vcc));
defparam \data_int[32] .is_wysiwyg = "true";
defparam \data_int[32] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[32]~16 (
	.dataa(\data_int1[32]~q ),
	.datab(\data_int[32]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[32]~16_combout ),
	.cout());
defparam \data_int_selected[32]~16 .lut_mask = 16'hAACC;
defparam \data_int_selected[32]~16 .sum_lutc_input = "datac";

dffeas \data_int1[33] (
	.clk(clk),
	.d(data[33]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[33]~q ),
	.prn(vcc));
defparam \data_int1[33] .is_wysiwyg = "true";
defparam \data_int1[33] .power_up = "low";

dffeas \data_int[33] (
	.clk(clk),
	.d(data[33]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[33]~q ),
	.prn(vcc));
defparam \data_int[33] .is_wysiwyg = "true";
defparam \data_int[33] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[33]~17 (
	.dataa(\data_int1[33]~q ),
	.datab(\data_int[33]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[33]~17_combout ),
	.cout());
defparam \data_int_selected[33]~17 .lut_mask = 16'hAACC;
defparam \data_int_selected[33]~17 .sum_lutc_input = "datac";

dffeas \data_int1[34] (
	.clk(clk),
	.d(data[34]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[34]~q ),
	.prn(vcc));
defparam \data_int1[34] .is_wysiwyg = "true";
defparam \data_int1[34] .power_up = "low";

dffeas \data_int[34] (
	.clk(clk),
	.d(data[34]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[34]~q ),
	.prn(vcc));
defparam \data_int[34] .is_wysiwyg = "true";
defparam \data_int[34] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[34]~18 (
	.dataa(\data_int1[34]~q ),
	.datab(\data_int[34]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[34]~18_combout ),
	.cout());
defparam \data_int_selected[34]~18 .lut_mask = 16'hAACC;
defparam \data_int_selected[34]~18 .sum_lutc_input = "datac";

dffeas \data_int1[35] (
	.clk(clk),
	.d(data[35]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[35]~q ),
	.prn(vcc));
defparam \data_int1[35] .is_wysiwyg = "true";
defparam \data_int1[35] .power_up = "low";

dffeas \data_int[35] (
	.clk(clk),
	.d(data[35]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[35]~q ),
	.prn(vcc));
defparam \data_int[35] .is_wysiwyg = "true";
defparam \data_int[35] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[35]~19 (
	.dataa(\data_int1[35]~q ),
	.datab(\data_int[35]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[35]~19_combout ),
	.cout());
defparam \data_int_selected[35]~19 .lut_mask = 16'hAACC;
defparam \data_int_selected[35]~19 .sum_lutc_input = "datac";

dffeas \data_int1[36] (
	.clk(clk),
	.d(data[36]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[36]~q ),
	.prn(vcc));
defparam \data_int1[36] .is_wysiwyg = "true";
defparam \data_int1[36] .power_up = "low";

dffeas \data_int[36] (
	.clk(clk),
	.d(data[36]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[36]~q ),
	.prn(vcc));
defparam \data_int[36] .is_wysiwyg = "true";
defparam \data_int[36] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[36]~20 (
	.dataa(\data_int1[36]~q ),
	.datab(\data_int[36]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[36]~20_combout ),
	.cout());
defparam \data_int_selected[36]~20 .lut_mask = 16'hAACC;
defparam \data_int_selected[36]~20 .sum_lutc_input = "datac";

dffeas \data_int1[37] (
	.clk(clk),
	.d(data[37]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[37]~q ),
	.prn(vcc));
defparam \data_int1[37] .is_wysiwyg = "true";
defparam \data_int1[37] .power_up = "low";

dffeas \data_int[37] (
	.clk(clk),
	.d(data[37]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[37]~q ),
	.prn(vcc));
defparam \data_int[37] .is_wysiwyg = "true";
defparam \data_int[37] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[37]~21 (
	.dataa(\data_int1[37]~q ),
	.datab(\data_int[37]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[37]~21_combout ),
	.cout());
defparam \data_int_selected[37]~21 .lut_mask = 16'hAACC;
defparam \data_int_selected[37]~21 .sum_lutc_input = "datac";

dffeas \data_int1[6] (
	.clk(clk),
	.d(data[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[6]~q ),
	.prn(vcc));
defparam \data_int1[6] .is_wysiwyg = "true";
defparam \data_int1[6] .power_up = "low";

dffeas \data_int[6] (
	.clk(clk),
	.d(data[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[6]~q ),
	.prn(vcc));
defparam \data_int[6] .is_wysiwyg = "true";
defparam \data_int[6] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[6]~22 (
	.dataa(\data_int1[6]~q ),
	.datab(\data_int[6]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[6]~22_combout ),
	.cout());
defparam \data_int_selected[6]~22 .lut_mask = 16'hAACC;
defparam \data_int_selected[6]~22 .sum_lutc_input = "datac";

dffeas \data_int1[7] (
	.clk(clk),
	.d(data[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[7]~q ),
	.prn(vcc));
defparam \data_int1[7] .is_wysiwyg = "true";
defparam \data_int1[7] .power_up = "low";

dffeas \data_int[7] (
	.clk(clk),
	.d(data[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[7]~q ),
	.prn(vcc));
defparam \data_int[7] .is_wysiwyg = "true";
defparam \data_int[7] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[7]~23 (
	.dataa(\data_int1[7]~q ),
	.datab(\data_int[7]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[7]~23_combout ),
	.cout());
defparam \data_int_selected[7]~23 .lut_mask = 16'hAACC;
defparam \data_int_selected[7]~23 .sum_lutc_input = "datac";

dffeas \data_int1[8] (
	.clk(clk),
	.d(data[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[8]~q ),
	.prn(vcc));
defparam \data_int1[8] .is_wysiwyg = "true";
defparam \data_int1[8] .power_up = "low";

dffeas \data_int[8] (
	.clk(clk),
	.d(data[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[8]~q ),
	.prn(vcc));
defparam \data_int[8] .is_wysiwyg = "true";
defparam \data_int[8] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[8]~24 (
	.dataa(\data_int1[8]~q ),
	.datab(\data_int[8]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[8]~24_combout ),
	.cout());
defparam \data_int_selected[8]~24 .lut_mask = 16'hAACC;
defparam \data_int_selected[8]~24 .sum_lutc_input = "datac";

dffeas \data_int1[9] (
	.clk(clk),
	.d(data[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[9]~q ),
	.prn(vcc));
defparam \data_int1[9] .is_wysiwyg = "true";
defparam \data_int1[9] .power_up = "low";

dffeas \data_int[9] (
	.clk(clk),
	.d(data[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[9]~q ),
	.prn(vcc));
defparam \data_int[9] .is_wysiwyg = "true";
defparam \data_int[9] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[9]~25 (
	.dataa(\data_int1[9]~q ),
	.datab(\data_int[9]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[9]~25_combout ),
	.cout());
defparam \data_int_selected[9]~25 .lut_mask = 16'hAACC;
defparam \data_int_selected[9]~25 .sum_lutc_input = "datac";

dffeas \data_int1[10] (
	.clk(clk),
	.d(data[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[10]~q ),
	.prn(vcc));
defparam \data_int1[10] .is_wysiwyg = "true";
defparam \data_int1[10] .power_up = "low";

dffeas \data_int[10] (
	.clk(clk),
	.d(data[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[10]~q ),
	.prn(vcc));
defparam \data_int[10] .is_wysiwyg = "true";
defparam \data_int[10] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[10]~26 (
	.dataa(\data_int1[10]~q ),
	.datab(\data_int[10]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[10]~26_combout ),
	.cout());
defparam \data_int_selected[10]~26 .lut_mask = 16'hAACC;
defparam \data_int_selected[10]~26 .sum_lutc_input = "datac";

dffeas \data_int1[11] (
	.clk(clk),
	.d(data[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[11]~q ),
	.prn(vcc));
defparam \data_int1[11] .is_wysiwyg = "true";
defparam \data_int1[11] .power_up = "low";

dffeas \data_int[11] (
	.clk(clk),
	.d(data[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[11]~q ),
	.prn(vcc));
defparam \data_int[11] .is_wysiwyg = "true";
defparam \data_int[11] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[11]~27 (
	.dataa(\data_int1[11]~q ),
	.datab(\data_int[11]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[11]~27_combout ),
	.cout());
defparam \data_int_selected[11]~27 .lut_mask = 16'hAACC;
defparam \data_int_selected[11]~27 .sum_lutc_input = "datac";

dffeas \data_int1[12] (
	.clk(clk),
	.d(data[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[12]~q ),
	.prn(vcc));
defparam \data_int1[12] .is_wysiwyg = "true";
defparam \data_int1[12] .power_up = "low";

dffeas \data_int[12] (
	.clk(clk),
	.d(data[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[12]~q ),
	.prn(vcc));
defparam \data_int[12] .is_wysiwyg = "true";
defparam \data_int[12] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[12]~28 (
	.dataa(\data_int1[12]~q ),
	.datab(\data_int[12]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[12]~28_combout ),
	.cout());
defparam \data_int_selected[12]~28 .lut_mask = 16'hAACC;
defparam \data_int_selected[12]~28 .sum_lutc_input = "datac";

dffeas \data_int1[13] (
	.clk(clk),
	.d(data[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[13]~q ),
	.prn(vcc));
defparam \data_int1[13] .is_wysiwyg = "true";
defparam \data_int1[13] .power_up = "low";

dffeas \data_int[13] (
	.clk(clk),
	.d(data[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[13]~q ),
	.prn(vcc));
defparam \data_int[13] .is_wysiwyg = "true";
defparam \data_int[13] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[13]~29 (
	.dataa(\data_int1[13]~q ),
	.datab(\data_int[13]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[13]~29_combout ),
	.cout());
defparam \data_int_selected[13]~29 .lut_mask = 16'hAACC;
defparam \data_int_selected[13]~29 .sum_lutc_input = "datac";

dffeas \data_int1[14] (
	.clk(clk),
	.d(data[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[14]~q ),
	.prn(vcc));
defparam \data_int1[14] .is_wysiwyg = "true";
defparam \data_int1[14] .power_up = "low";

dffeas \data_int[14] (
	.clk(clk),
	.d(data[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[14]~q ),
	.prn(vcc));
defparam \data_int[14] .is_wysiwyg = "true";
defparam \data_int[14] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[14]~30 (
	.dataa(\data_int1[14]~q ),
	.datab(\data_int[14]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[14]~30_combout ),
	.cout());
defparam \data_int_selected[14]~30 .lut_mask = 16'hAACC;
defparam \data_int_selected[14]~30 .sum_lutc_input = "datac";

dffeas \data_int1[15] (
	.clk(clk),
	.d(data[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[15]~q ),
	.prn(vcc));
defparam \data_int1[15] .is_wysiwyg = "true";
defparam \data_int1[15] .power_up = "low";

dffeas \data_int[15] (
	.clk(clk),
	.d(data[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[15]~q ),
	.prn(vcc));
defparam \data_int[15] .is_wysiwyg = "true";
defparam \data_int[15] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[15]~31 (
	.dataa(\data_int1[15]~q ),
	.datab(\data_int[15]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[15]~31_combout ),
	.cout());
defparam \data_int_selected[15]~31 .lut_mask = 16'hAACC;
defparam \data_int_selected[15]~31 .sum_lutc_input = "datac";

dffeas \data_int1[16] (
	.clk(clk),
	.d(data[16]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[16]~q ),
	.prn(vcc));
defparam \data_int1[16] .is_wysiwyg = "true";
defparam \data_int1[16] .power_up = "low";

dffeas \data_int[16] (
	.clk(clk),
	.d(data[16]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[16]~q ),
	.prn(vcc));
defparam \data_int[16] .is_wysiwyg = "true";
defparam \data_int[16] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[16]~32 (
	.dataa(\data_int1[16]~q ),
	.datab(\data_int[16]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[16]~32_combout ),
	.cout());
defparam \data_int_selected[16]~32 .lut_mask = 16'hAACC;
defparam \data_int_selected[16]~32 .sum_lutc_input = "datac";

dffeas \data_int1[17] (
	.clk(clk),
	.d(data[17]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[17]~q ),
	.prn(vcc));
defparam \data_int1[17] .is_wysiwyg = "true";
defparam \data_int1[17] .power_up = "low";

dffeas \data_int[17] (
	.clk(clk),
	.d(data[17]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[17]~q ),
	.prn(vcc));
defparam \data_int[17] .is_wysiwyg = "true";
defparam \data_int[17] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[17]~33 (
	.dataa(\data_int1[17]~q ),
	.datab(\data_int[17]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[17]~33_combout ),
	.cout());
defparam \data_int_selected[17]~33 .lut_mask = 16'hAACC;
defparam \data_int_selected[17]~33 .sum_lutc_input = "datac";

dffeas \data_int1[18] (
	.clk(clk),
	.d(data[18]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[18]~q ),
	.prn(vcc));
defparam \data_int1[18] .is_wysiwyg = "true";
defparam \data_int1[18] .power_up = "low";

dffeas \data_int[18] (
	.clk(clk),
	.d(data[18]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[18]~q ),
	.prn(vcc));
defparam \data_int[18] .is_wysiwyg = "true";
defparam \data_int[18] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[18]~34 (
	.dataa(\data_int1[18]~q ),
	.datab(\data_int[18]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[18]~34_combout ),
	.cout());
defparam \data_int_selected[18]~34 .lut_mask = 16'hAACC;
defparam \data_int_selected[18]~34 .sum_lutc_input = "datac";

dffeas \data_int1[19] (
	.clk(clk),
	.d(data[19]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[19]~q ),
	.prn(vcc));
defparam \data_int1[19] .is_wysiwyg = "true";
defparam \data_int1[19] .power_up = "low";

dffeas \data_int[19] (
	.clk(clk),
	.d(data[19]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[19]~q ),
	.prn(vcc));
defparam \data_int[19] .is_wysiwyg = "true";
defparam \data_int[19] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[19]~35 (
	.dataa(\data_int1[19]~q ),
	.datab(\data_int[19]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[19]~35_combout ),
	.cout());
defparam \data_int_selected[19]~35 .lut_mask = 16'hAACC;
defparam \data_int_selected[19]~35 .sum_lutc_input = "datac";

dffeas \data_int1[20] (
	.clk(clk),
	.d(data[20]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[20]~q ),
	.prn(vcc));
defparam \data_int1[20] .is_wysiwyg = "true";
defparam \data_int1[20] .power_up = "low";

dffeas \data_int[20] (
	.clk(clk),
	.d(data[20]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[20]~q ),
	.prn(vcc));
defparam \data_int[20] .is_wysiwyg = "true";
defparam \data_int[20] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[20]~36 (
	.dataa(\data_int1[20]~q ),
	.datab(\data_int[20]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[20]~36_combout ),
	.cout());
defparam \data_int_selected[20]~36 .lut_mask = 16'hAACC;
defparam \data_int_selected[20]~36 .sum_lutc_input = "datac";

dffeas \data_int1[21] (
	.clk(clk),
	.d(data[21]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[21]~q ),
	.prn(vcc));
defparam \data_int1[21] .is_wysiwyg = "true";
defparam \data_int1[21] .power_up = "low";

dffeas \data_int[21] (
	.clk(clk),
	.d(data[21]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~4_combout ),
	.q(\data_int[21]~q ),
	.prn(vcc));
defparam \data_int[21] .is_wysiwyg = "true";
defparam \data_int[21] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[21]~37 (
	.dataa(\data_int1[21]~q ),
	.datab(\data_int[21]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[21]~37_combout ),
	.cout());
defparam \data_int_selected[21]~37 .lut_mask = 16'hAACC;
defparam \data_int_selected[21]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(\valid_ctrl_int1~q ),
	.datab(\first_data~q ),
	.datac(source_ready),
	.datad(at_source_valid_s1),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hFFBF;
defparam \Mux0~0 .sum_lutc_input = "datac";

endmodule
