��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$��	�LJ	l�k:�nF��v;s�ҥ�x3�J��G�۱B�+v�;��@!�̽��@�v�ƜsIM*ǫ�`�'�fc�E��-�;����`��^! 3��Y�{�kDd��b󲐪Mh�,"�ZVF�V�����O����A�镖>���J�v)�VV�m��x��- s���2mi-��V�z���@��w�: "UJ��p�6���3�r3��?ߟ��-���*�g�����_t7Nʘӡ�F)�������PEڥ$6�[�$걖�=v[�ȍs� {U�H���D~��$�	�,@����`e{���\f�����k��
�P�Ǧ���2H��uDR<L:��l�oS�;ȏ0֬`��4X��e� �?����飴��z[���TWo�EM0#]�_�Vh����S��
va�Ƀ��@�3��z�z��.��y��C)p�g.z)��\`���穫u~H��Qr��e}K�2�eL�eC�jШ�<F��ʈ[����ˤ��_��N[מ����a����k<�+�LG@j��.�C��q��ŵt���XIz)g��7��i��u�L'�Z����#�q zAŽA�� �� A�ed�<MٕU�D�����:FG�)�[�+���;�
������ ���k�8��g'�O7�_��p&�d^�M�8��W�8Gid��*;D�H�f)Jo�M1x�gTǶ2ۿ}-�>^?��@"����
>m��7P�7������
N�6��c99	��zϽr)2�"W4|O%�T��ؓBnn����x���$������꧑����T�꯲?`h���1-AphL7�n�s�@i�5�bq��7�w����0��G^�iU2��s�W������N�7�i�ia�ʝ�,��i�X�K�/8j9�쏊��0���50����œ�]�@a�is	y��f��P��z�e��P��,g�5���^N�o�'�ta<��儧��\�s��o\����M�0y��T ����7���E�?���>N�xgAs'��&�<���jgs�_���ie�O�b��t[�hn}���9�p����bMOYS�|��To.4˚���/��W�W��KMi���ʰ=@=�"k�X�n���o��v��s�A���@�	n����ѫE�`֐�b��@mc�D���.B�L�]�k�-��|���e^�/����}�|��;�� �n�iF}�ԲYÿJ�.�`���ԧF�n� A��C|��Ah��塀��@�"�?��^@�F��V��D��V�Uh����p���E�ĕdՔ+���m4Ub��%�@�F6�Y�aYB���ʩ��������/^�_��Z��R����mv? ��.�d��L{�cGm���*�R�@��l���E�<��h��w�>W�ynw�<�:hcL���N���@�vG4.b&�A��$��)����e�Zk�2�
�'�VZ�	��^}C�<q�(�Kög篱�y����L��LLq����N*2N�{�f�d�_e��$ɓ��at+���ePb�����y`Y�&�H�k�4�))|C�*o�ax|;0��\�<��+οB�|@5�d�%�oa�?f��:նs:�s�s�P�̗�4�/Ӫ�g3p/���T�����N���c��b�%�b���_:��.0�k�X������D!�Jʯ@��� �o{����hX:��!����e
)}�w�j�!�qh�e���I4eIM�4p:.�"����% H��2~^��CFu��T�k�2���cABJ#[Z��Z�~�R�#�{N �Id3I�;�D���HB����r�����%� �����u�r]��F�m0ӹS�&�E�����H��1���:�� D�-hg�	�vџ�]�$g�q/*6��f��<�Uj��4Q���_˃U�oN�#r�"������9�؝�#�Z>�J\��P[\�Kc�vQw7(���#�a�ս��4y����tv�?�q�/_�H���x;�.�y�D�k�V,������H��؞]!]~�S�8Y�+�6�0�±clR���K�=�9����Ҷ9�K�����ѳ<���i�h*���x��RZ	�;��ؤQ��*���$���cm����NjZ,R{���_SHJ���V=��u�Ւ8���a�:ҏ��)��az:�~2'�������?��g����SP����oŽ41�>7tV]:2�t�l��"�u��_��&�A*j�}k,!U���s���n�� ]��M�mkԴ��t�.8V3:Ai��I�!픎j��<��B�����hu��y�m�b�����3o��"\7�Z�}�3ɻ|,�#ժ�j�鴍��j+\�" #�0~[��g�j�NyDu�1o,FIj��*G1kGPI� ��j���w�Q�����CI�q�p���2��7qϧ�`/H��H�M�Gf�KʗL���s�џ�Ȯ�j	9AA~�J`B��L�]; Z�5m�N�%h�9����T�lh�
��r��r���h��y�Vb�S�2��iY��N3~S��3+����}�j&�j9e��k��P�x��N���b�� 1��I��4���4��b꿰���⽩�KѼ��$&�}�n_�6{J�p:?8�M9�4ѷ���}@�Ǌ��vBU��m!��R���'��xf͝�hѻ�D$�Ϲ�y$=&���4�ײ�u,;�G��
�d�*�e+��v��橫_�>�l�
�:�����w�.!�����lǉ���I7��z�"�IwǓ�.��a��|���}Qwj��jv�-����WJ��Z�ݕ��a���o�rN�ǘiq�� ��v�tϢ��)N����D�����2�lU�p��q��RH�j���F��z�S���.��̲^*ye��d��)s�M�Ak�n>��A���k���W%�=��^]c؁&tw�7�\nʤ�w��`v3|�k�P��P��X���1Z�N� L�=�Hv�и��;ř�8(�kݠl�l��2����v)���dK[L\�"2`I)��A\��o�_C�̧tD)M�<����ZN,���e�	�"�2��bŌ�G������6_9�TY"&����ߨ[�[�����	'���;���F,0p
pd%�wd�>C%_sS����6v;Q���s	[���P'N�4�·�=):~�Kv#�_~O�4�K+4]�����0����lc�F߆�3�_��j��X^�W�jUO�H�������mPK��M�D0֒n;Cs�4�Zj{�0H��J۳�6�܌��w�����o5�$��6�G�r�S�d�W@���@եd����ۧ��3��ᅾb�����th���++�Dl蛠�'ZW:�崂�����_�'d�ӫ�B�Tj��}���;�Ԍ/P����he4j� h�F�C�K�9.�������ܴ]F����'�ց��c�U��~���D|Y�9Gҝ��*�Aه>?��̿R5�fk��	�m�(��l��Wߞ\����Fر)e���q�B:e�,O��u��Fn$GZ� Rǉ��������/UwQ*b��w��4���ϔIp#}Ļo�F���8��o�/<�5�7#�*8z������|O���L�ԕb�qm�����J�3��+��Q�A~� j�mZ
b[(+]UuM�.|���<-r����?�/b*�h�8a�@�?��pb1����A�d<�G��л>��.��
��%Wmȭr��~�S�h��,p��� ��0:A%Li�o��A��,�g���N'�U�Ae��1��P{��Ĩ%�? |e �5���'�f�6���֕��f�b��x����|睌l˰��>� ����,�$��H�J�-Ƹ2�=2L+m)Hv
Y��2�� T��yz�� t�p�L�͓Ö��<�F�	�ӱG~9�`�˚B#��#xN�W��o�V�����M�<H01JI���;R��O+��y�l_�U��y/!Nt]��=�> ��D<�;�	�D���Κ�{� ��5��[���A�S�5_X�v�Zt����[��Q藍��iG&%1���l�Mx�;��{ԗ���D�/������dW�a��Q.�R�����qX��ǘ�Ln'�d!�xl��&DUǇ���h��.��&�!��
��`����&=�'�� �Kc��O3��S׋E�9��>Վ[]\���B�q�u��uf�q�&Œ&z#�������ܵ�[Eհ9�`���+��d����O����{ 	��"h�u�aڿ�`M:�S���V+ ���셵C�U�Z�4 =��L�k6Ӧw��flA�.<|O�-�(�!!MH�F�2�oZ�Z^S̼���a�V�5�>3��Ǭ���Eq���}u�G���,?0o&����v6�}�p5�²���x�A� ��C��D�F�u\��� h�f�/�_}��w"���ҵ�'쐨�p�k)�.����(��Do�����l���f��^�'0�Q[J�2�TJ�^"m�C��P����%+N!�sPm��ױcә�6�L���溻cnq��{f�8�/��c5W��UVMQ..ձ�-Թ �Ǡc&-Y�h'�W��.^)����`�#)S�=(d�	��g*�5t�Ru�(w�Q��.�;�`���Ndw�%��|J��J�/0!��@�Ƀ�|�c&��C'��5%z���ߎ��K��*�+�1YR���Vb����@o�+?�V�d��!�c;[A:��:���m��s�xE�U�׏���J'B�;����	ʓ[r�bCKH��Ӳ��;X��:P�Nt�[��l]�[o���
y%�I.�&1x�q/J��,r2�t�f	2.f����Bnr���R1j6�!�d�`j�F�b�����^zVkA��P�e|��BI�ȅ@d��-�z����W灱�֑�Ly���r�uG��-1u��\��*��i57~�ġN�*�#��`OA���_U���x@m],����3���n���u�6cX��f���R�ZL��.��i�#��3����EK�1��'�|i����B�^c�XO����?ܷ�9K��h�r�p:�K3�x
�K�W���E�rj{�uɚ/�;��E�s��0�xl=h��~]�f�s�#o|��71f�����9]O]=����s9,O)�b��DG]յ�5oF#(ؿ��J_���R�D��u
��犉Y� �[����~�y*גjK��[6 �4^����!�������e-�ɋ]h½u��jșBK�_)�Xby�ئ�BF��а�P��t�������Ȝ}>�6;!�6y"n\�%g��������� Ԏ7_�o�\T%�����zփb�u#�g�:�|T;�Q׉��G6'�"�ϼ�Y�[y0�����  �	9$}ew�o�at��(��PdkG3���B5Ѧ���eE��:,��5ܸ���[���dF̽�A;{�&������xv�S|o�#m��������G%���a���i��%��#ֿ�D#�s Jv,t�z�XO`���=5H_����D�"��Ԅ�������Ԑ�I�;̖�;],��6Zx��ξD�yH%�eE�isIz`��}`��=q�.��c9O8�Y&�#���~{իDs�,��0�U��#H��_�'	¯�/���f�F��A�a���q�"@y��H���Ҫ2/�g��D�r`�ьH\�͹�p��{�&�ozqf�"�)e�#К��rC�zZs<�I�Jg�@�/W6�j�2/W� ��8lI�i+ɮ�'�����@59��6�>���C��k�u�A�<UU2�|?*O�dh�x`����%>��?�ʘ��P����e����N7�'QV�y�{��0����]�=9�/#C���W�?M/�"�Q�O�X`�LC�Qd�+�[ϸc��C���h3��ʼ����fq��d���A�h��#y��a�yM��ᙣO�̖�8�O�v���/m@m]_E�5u3�?� �qv�=��B���2�b�������ɧ���A">�p.��1��s��̖aF��VI��sQ�j�]�uzP��{(��q�Ach�%��"�����	W��spE��D�Wv�It���y�9'`���f�:�~�2�
�&A�M��I�Vp�4��U�tx�Q�&x��C �z��3�LWU���|.錚�$8�~�Z�44Z2� @<hQt�!Ex�-B*�!h����j��ag��,��A0�"	��b	yQ,��Ҥ+���IP���G��5+w��ڢ�QR~O�3���|q�T@�%P{)��'M�6�}�:�C�Cj����
K���5��Oǀ�BHs�"��O^�4 vSGǄX��tIg�>���1%ߔ�R��JN�!J�����\7w��[nY�N�e���C��@���K�9',K��`�yȄ0"�w'����O�=�$3�9cj\T���bS�w��=8J(:X�͐gq�H������e#������p ծ��V��{�eLUƴYĽQ�L�oE�6��TwWz��x�ơ36��g��	m^��َ�%8�a�C�m�G'�^�w�1ҩy��#�㭉�1��([K�To�[3K7�aHO,�z�J�譸 �n��5nuwk�g-����>��"�W_���zfξ^N�t�r�
�z&���-	f������\�e�P��g$����@
ư�}���k~���G��ŉ
V|P{ �H�?���~��05��>�i<X�.�PB�]����Ldע�t�q�����iϏ?�����z�g�c���_�����vR.?����͆��Œ��L�0*�5�G�l����d��R2T�(.=n2D�X����sY��F������x���u]���[~�G�Us�`�)6�4L�l&��VO�
Qً����|x�7d�($)�z��k}���L�R��H��uP�˶�6b�Ct�ӻJTp�u�7����1֠�|"�ͷm���7�^�=M�Py}�^��ݙ[d^k5^��*�=��T���D�dIQ~���>&z8}��B�z���_���}X�`Th�M��n�� F��0?�%��p�/`����pB��-*��[S�D1��R���8��(k[Gm���B�H�q|���c0�8��'�&��55�r]}"��G���Q�� C����w1��D����m�� �|e�?���[��
��&Ҩ� ��eN�-fn@¢@X�Rp5C.��#��h��E�%�Z	.�,=�I�顪� 9�DEDÝҗ�$�n�Y�3�U�!��D�¾�^��)��Q�ٖi�^NŻ�n��RNp;�z�T���޷\ -���:P�xa�,�K,�C�"!��T���gl�K6��Zt
usGMǹv8�s�m:q�_��9�UM8��eK0{hǶ��3h.�W	�gA<�?1�Z����|��^�9v��*�]�T��mT��.���+��I������L
���ʲ�h��1�ĞY��M�F#%�Y��wFd�h��
��cXU�>cw���4-��;�T����ϸ�U�r�s�p�J���Ɔ�F��.Pܑ�g���Q��}�w0m	c�E�w�e�|�l�3����,�W�^�"7��8��+���"Ձ�q��$gw/*�R@4)�y:w�e�i���m�@v �G���ӟ��4��̬�;T���%�S���!�M���>�jƂ���-�o�$�C��.D1�z
�t�/�\+��kp4�۶-
,������i�x��CZ��wE�g�/ى^����
���v�4��ğL��f.�s^P.	����5�q�m�n��\��隆*
�~�ɾ^*�Vh���2@�'b��a[P�$�BJy�M���죶�D��Abx�J�l	�,���Rzj���a�<�x��8;�g-e�Բ�"�<W|'FقU�Z{O�1���"�(�� ��(^�PӍU4��7������{c5�2��ɮ�`OK���2�SL�!���7���T�J��["KD8��=��ˑ���\}/�e]�"��l�sL�3V�n����ÂLh`=�,Z��v~�*���D��Jg'�UIF�D)E�@qH��JeZ.�j��}��,�3��8�;i ���!��W��7��Y�?��_O�K�O��\f�P"Y�`���P�s2�$������:d>.�jF"��xׄ��6d�-u���.zV3�vz9<�`�,�qRWr�8�Za-y�A���_v5i)�d`����(&��^g����'Ie��m���.4��P'k��x6�t�� �*mP�����pH�g����o������7V�C2p�Kޢ����6�I����Wa-�}A�O�?H/J��P�i�r�)�"O/q~�M�.��U"�<�\˖@Y���#���\p�2�.�}����8�jL)�[sx�Y�sa���j��/�I���hϞ�� ��9s�	�l1����k����Z0�B)E����sTU�*��T ��OPv��ױ���\�˯V9���8ȫ����*q��ܫ�v� !�5`;\�r0`���FB�ga�y�W�n��iw*