��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
N�m�H2
��j�Y�?	l�Aō4�8�����>|�f[؁���
Ζ{�����0>��������'l�d�b�%#T���QOo�Rh��&42`�-�R3Ml]�Gq�]O��ל��J���('���Q�5�.����p��� 6�	J�/FM��8���b�)f�ĐI];�^�EL���j�����D�1�5�1�K%M6P�]���*"&	а��u��~ٷn$5h����k��O��L���׎D�y6"�  UD㍺���"O��ܣ2^ �4"�.��d_y&����V���k���ƭo����`���%ȯ��e��εA;�3Yй3V��l%U}��N��������aUiJ��������X(7:�_0�Ah9�[��=�2�5�����,�_���i+���C�m���K-?�qi�b<�-�a�!?@�3��w"�[^�J�������+��A��W�P���
�sYy�ŏ7j�S�����h����nK�L����E��#��-�\�9Ú��U���-|{s֒Ѩ�y0z�]�C �_@Jn b�K� ��A��a/�F�B�!�Ma��Y'�����G������]�LQ���|��gE���,\6���Պ�E?��d��򄻙���R88���Z�c��5���G��{,]n�M��������ܵ�l�{h�W�2;��+p�εn���>"q��N�G�T�����o�-�m�%�xG
�o�]n���	l��'��a��qB�d\|���Yc�Z�t�x�塳Lr��X��/'>]��59֥�'�w�ƣ����2I~ٺ}���Mw�q�ckg�<�B��<�� �b��ű�G̹�[�(�R����Dz��#hu ;��9�`6.z\��".����X*Q�dP�So�4�K��z�~�n�^�a��W��3	# ����k%��t��S0��9����N� �o�����.�Nj�z쵱�G8b�1?�v~�W��e�POOs!iъPU1��� ݀���e7��o��^�]F=c�59�s�+7�ҫv�J7=���z
��_�σ��y�\���h�_��s|��Z.����*ô�XE�@�L��:���e�P��E�U��2���Ἒj��iu�*�9*���^�y�Y��ja�3����qL%Q~����P�l8���Y����3p�V_�X��U��2�p�R�
J��p�ӥ�-�؞7�;���
����ԃC�B`)��Ђ��#�L.��FbOx�4��w�6�c��Y���ia�W�le�\�L����
NBR��@9��+����dϜBF�5��q�>��&�.{a��n��k��/|�i?ڜ��J���|�pP36���ҕޥ+�ϻC=�;7_!�g}u_�]�(��1Y׵��B��r����Z���aqB�������_��2����<�g�$��mִ�Ga��)�f�"��{(�3w>�R�5��D���t��8���A�����VkQl�"3����}�� ������z�����T�Q��@f,�V	�
�ib3-m�''�)5�4D���{�c�+&'��'�}9�5P�g8�����-;iaJl�$��W� Cǳo��zH��%N=����Iq�>n�0��| �H0�,�X�RhKM�Xۇ��tQl����Ge��j*��x�G��K.�"�b��.�o�\�����Kg+T�Z�����m�Ĺɤ�
��ó��&��)5�&�+�m,5TPY�Vw�~%8A|��=�H`(���JآD�ދ�(�K{B��ҝC:�%X�?� #�4K�������lTH�C˴�t�ԕ�(�<tۋ�$�� �?�R�o������|����O܏0qt������4����/a�+&[.b&����	�Vo�-�0�,�ɽU��-A&4�#[��u�d������y�e*��]�E�����1rGz�D�b���������?��C`�� �̲�	�Į�j�>|e@�T9�K�q-�C���7���C�kcn��DqZ����!d��su&����p��µ-�A#y6g�p|�b������^���Nf��G\�Lrs��Ure����L�b.1����w�#�����Q{�A&����Qeb�2%��>Ȇ����lsG�r#�cNr[��rHJC�4(���.Z��=���|7ⶂ�`���≶��C�n�q���?m��x\4J�������0|����_�z�Ĝ^ilCt�꛵A]��Ez����ɜ��i\��1�r����}��\��5�h]�����Q�&��x��@J7P>��E�k�f>d"�T_�>M��:��� ��qa����D������ZI:q��kJ;�XC��U&�@*0b�=�f�1��)w�j_�?��B�n�>�q��C�)$М�>��� �4e���R��c+j����ۛ�	s��/-Q�0#�;�#\��C��*�$��J�/ �4����ɨ{���D���d������F�_v&x�[��OQ�p���R�#������u���C���C%	n���oA=#�8��i�l^�K������!8c? �e��Ed���EU"��V�L
��ސB�����eP�:/�L��i���D˨��UC�m׳\�s�R��U�J�#35$�J�2Y�ro���D��k^��ܬ)	��U9l�v�έ�������Z�XX�(ٚ�ЀJQ;`��C�=2�x��m,�GWt�K��������~�Z�+�ⱎ<|�*�R�����8SI�T��A�LÎ�Q�������@���"�'�D�v��-��'����w��R��f{'o�uj�����`��"2+�/�3Ί��f�WC����m��!M7.y��/��w���,�_���"VQ*L�6���'1�+�º� Q�`6�p�6�%���%�����6�;�������_��PVd���҂���ywF��۩r�������%�H	D"���L�յ;v>d�/�6�Ge3��0�&�K����sf�l+g|�+G�}섙M|�h��\���8s��Ӣ3��r=�E���Qs"D_Ǆ�N�D���x�Uli��
@���ff�v��- ���ש��M�CHO��W_�N���
u�2[f�Ўv���íR��_���r��a���!$[KPھ�[VY�r0@��y�qM�W*�/�8�i��S�4�f�����rdL
�jldeǮ<��\-�R@����F�m�oY�MԊc>'K8�jWa�Ck�]{����/�θ6VCx`y��^�I�2���Ȥ�2���]\�pq	I	Ù�M"�삄���/�/b�:U�ϑ��%�4�8)P&)��/���l���ݺނZ��4���v&\ߔ�9R�Fp}q}TJ��M4�M�dT�;%����V��m��>y��z}���쪴I��LA����xm�0H}.�7�U"X��ʌKv��
I�$� �H�C�����Mrf�X��?��3���/�4{�B��W.@����"`/�ԟ��{o\/۵�Sm�F�i[=��ɱL1�#a�'uO�к�h�{RG�IF�ހEq�zl�Q2Ye���SɈ�&)[�շԖO��v��F. � CWyc�<  n�J�c����D�o�Чm�zo�-$y��+wL�/�����Ӡh��h=݆1��
 �����.U��.48'���]��`��E:��<��[k�晇\�X�)� ���(�����G4�U���ut�YYm��TV�h���g-�l*����Ί��c�5~:l.� w�L�:̑�ᴡ��!��@$��2�MZ}�C��M�TS����j}��L�#և����ű����l+���=�8��K�2����́��*�
�T�P���%��,1u�����JKԚS���:I��'SMw�#/���a�e���[�|h�cZw��ԪS����}�N��6��>�o�Á���@(pqA�x�I�翘��1c��0V
ŎQ��$;�.���
��Oi�ƫ�)�[W\���V@�Uy��c@_��1�����J(:�O��1D���b1��9��`�AZeo���"�`p�a����'��h�3�(g2�D����u�޿^�ƨ(s�u;�+���%��̕A)���0�E-��DbF'�E&iANu�̖4ޜ�������
V��x17,���r�z��z6��`��=\bp�׏�O�v&�(�
���:��fٲY#}�?����UBK�Ā��`�ZP��V�An�n��&E��dP�e��I]��GG�Qz;�hh�Ѓ��b�'��<�Y;�*���
�<��@�G��B��A��~����	����Z��w��)��{r��.��R\���~���3+'Ü,$lqF!�P0�'�&���]��[f�Md���?����x2[7#73aT<κ��n��1/�Gsڟ�J���=I����<-��$X;�~F�G�K;���~)���N�df��l6E)�9�A ��:X���$98���`S�qAYO�-�~~տ�:�)'����3�Q��U��z��B�vx��֪�堏w� ��Rд������W����#U��'��m�̂�(۵�1<�KT�m�:kZ�|����G�N�b�B���1�Y@�iy��a�� �!\������M�������t�n�������Q6�_0�F3�x�w���<u,*z����]��Z��*@]�w�ϖ4���{G������$0e-[�bG]��#Ci�-�X�]C"�o� jr~2L	�o�I�8�#o�[kJ�#1&��6�l'�2�m�'��Jb�;�����=�
ʔ,@�o��7��;�~��4�d�V;�>�k��8w�I�f��݇�{�KYT{𱈥x�A�;`wD[4k9Ö�o��җ�H�/eJ��i��� �M�,?� /�v�[ JEˁ��rLW3_�2p��7y��������ҲV����SM�b�1�ת���UQ�Ȃ/-^���������g V���G.8.�}�7�M��52�5X���#��؅񲢑x���#b%�GN��[b�H�B��V�ڎ��Ww��|R��}l�c�!q�1zciJ�	�X]�;!vtu�օ�'�X	͞����B����Ɉ�ݤ��G�� 3Ȱ'1��#�E	�	�Vl�Uoc���3Y��\F�2���jj��R�S��㿆M�r=y�WZpJ����p������)��eP�qS���N�9Wx���Ӻ�07%���ܛ��AO�v�Gd2w��.�_�rGe9P�M���'�+�M�[9��{��^8�o��1�<tz �M���F�{lT0�A����@*Am�������F�|�5��U�EAPZ	��c�4>ŵ��)ۏ�٫ڇd���D2,��~0c�*H��T%S��v:�P1ܺ�fI���h0���_-{�FA�"��B��Nh�;gݔ� :�F2��G�+�MTN������;1aR��}�,�߯
s��`�
��Z��@*�����l������u�>�Št�T��⩽���@��"mb_�o����	�S5+�쟎"�p/R���g�h_	�s5�i,s�%[Ӡ{dhTx�����q}R���/jҨ�c������?[�		���q�۴�kӉ�~�d���F�2��Nc�S�#ʯ��2	qE��� q�?4̿����sf�#.��O�*�����=��m ��U'R�{!tzaT�&���z7���<Y�H+�Ű�"+��_�6�*�\l }oa�,܃h�Q�&`����aU��i	�C'�m �*��MQ��������zT�eh`$G����6�P����s��Y�sǱ���a���& �C��Yퟩ����I�RN�s��P"c0�04Q��j����A������ka�[2R����\w����u^��x���[H��׷�����[U�����Z�{��2UV:'9�_�ꞈQ�v׋�9q�u����8(����,����
���UOKn;���7J����?��� �4�U�G6G6�MwR�l�`K��C��* y�e�h�7�p�u�tۍM�߇~�JRPj{O�a�B[��b2���S|�g���K�,lp������H@��J\ybvd� k��)kc�o9�^;����t���_���rH�Z�u��\�%�A���"&[ԫ�E�"stQ7vڝ�#�^��JU�KĶ��S��3�@��C���^�o���dP:k�
���t_�z7�L��؍���B�%d��QV��Q?tY�4�����(���ɣof���+��^��̘�GlD�X�a?\^��+���UV7�A� ����lԃ��!���_W��֊2������%U��~xA��΋�1�"
:Q}>�Ҹ~�����'ฬJ^��=�;h� !\ �m���L�,����,Į5�P�Wl�=�-
o�:6���BQ�2�፫:l8(-��CðΟ�g.�g�R���vK-�݊.��D݃|sK:������i��u��`����b�/re/���9��2��������-�H���*OtUQH�oa=�!�Κ�7@婱1�F�L���ޓ �	����d�yK���o��J���gBco�M���?MF�ŭ�J�����&�4��ͤ��콭gT5��d�S�3��I��}�=y�b������S��K.݆l�j���g���.Y6���J�LWO�_�e�c�DW1�����_�j
�5]�����r>���-�^T��U����T�y>�޺0�I�����)�[
�j	
��E�T�����ŶC��v�6��q�U�Y�Z����
_����H��%�\�%j��aʄ>-�q��<d��|N����2c�.�=�7�c�q+��(b�?EV6��fdN;~5M>6��. r9�D
�7�^�_󢜢��;�>i/|�;L鮖�g>��"5�-�=%H"�e��L�����̤Gs�D�.'�37�HT�N9"�*[��~��T�;���8�p��7�5�Z�C��6�t�k����/�`���)��}.Q���+rQ����\J��i�M��c���S:����zC�[�����[Y-�V*�4��_���yM.ʼ
=J�[��3f�+����*r2/5E�#F�)�O_�5Y.��77o�Ǖ�9�RV�26'��T骯M��f����6<���?I�Sb�ԥ����Z�F����<�V��P�ˑV�2���7`�k���7��]B+v|��w��W���9zl�4^0��s�Yl�Ͱ�P^��5��?�h�`h)�s�~-���A�/þ�}�{�h�Q'���aT����1
�!��{�f>t`��3������w}�r��q��f̦ځ_ )�6��x.V;��j;W�n�]�ι��H���"}hy*	�_]猛��g&�iC|��Z��b,4����)�^x��0�k�B��E͛`��.	���z3C�q��~������W��+6T��/?'>���sa�����=?CX	B~O{����6�5�şXV��OZ�a�c�u��H��	�B1vK��<�	D+�v����]V壴�n��������H$U
!	}�$��A����������'�)l!'��0���F�Wg��>c!��hd?hi>:�)��R8#��R���U3�|Ek��"TWz%"f~��1s�$��%}ٞ���G����T*l)1_^6)@`��d3d�\t�i�������Vp6遥+��G]�JB���y-<&):V#�֕
1]��FiK�灑��G�	9�:��(6��XIt�9�m�{��3�[	F?���t��e�[�����Q�'b�S���D�Ӫ?�$�`��ޒE��?~G,3��*��x¸0o�K�x��	������C�����n&�a���+�T�WR�dm8�w��N2��.�p,ˤ�����ƕ�T⛌0�����
����z� >�:h�k��E]Dm���A	0�ټ%$�Q!/J�T���W!|������g݈�\T�u~�V�@;�[(�sf�~W�h��p����������c�l���;�>�dRg�V��X���l��1Ra�F��䮲�k��f8+�����,�/�?�#��.О9�,H��E.�A���*Nhc쭏� ��P#W*�����]�1��-<&�:SNB`Q���&����!��14�˯��o}qo�n��!8y�����4׻�ȗ#m[H��^�����NFP��M�9��f���Ĥ�>Fj��m��`�K/���0�	�϶�39� D��Ŷ�w孖��k q������|/_ˊU�4�A)L��ӱ������>�M�R�'?gR���C� �����?Ƴ���!��l�ţ�R>��c��f����jVD�N�\��8r�������T��t�%�H��)�!�Y):~o*����U�q�s��x�lH�*lb��*�����s��$ޯ����j=M(ݱe�[�!p���/%5w�em.�.�J/���n5 B�a�v_�5��D����Տ�c�sN��"49�=�A@�rTCO\�= .�4f|�OQ�a��*��s��W�,�ģ��A�f4�;H����X��	���"T���E���]��&�e�����hR��֫��,!S�W�4�6���׻ 1_~�,�E����nj9�c����6.q5i�P�S�?C��h��'�ND�i�o�
����3m�P�l.�������>��?.me3�P��Fn������Ә��jM��:=��&lw��H��w����)���	�����v�������z6�����3�V���T��H�?�t�y�1�l]1|'��sD!�`�/8<%�Rߎi��%���c1,����q�ގ�Q���ȡ���	���7�=G^�}���@":@��H�1�˵�\�C*F%�{���s b�8a��<ȴ�8-��A)3U�����$"���'� �J�4d���V��^1�ɵ�`X�����,��?j�zHL����\/�0����u[��f�6�!2���m�M]/ZҵTh~�#��I@��c�sY�(���&*�;��2o���6X�OGsc\a�r�f	���rc�	�w�ؔ���<@1�N���8A9�=2}�V%����aEW�1w�{!�Ĕΐ����舰��>��!�6�갧B	o톷��u��<����ҥ�y��2���j�獨a�$����M�ϑ��aհ�q۸�޶�A^�#y�*�S�E����)� 6ja�A}�����n�m{U�v�â&�1�x��<��sR.b���$ڤ���z��s�)H����<���C� [j��V7E�{f�����$���/U�[@�~y�͗\G�I��d�n;NWӴ�Z��q���(	r
փ�J�;�u�jd��b�q��˫�sA���qu���Ԛ������7	�T���GCT\U�kT��)�u���EHm��#�X6ԸN��E�ɋ�:��;��Sw��Trj��V�"�̢^�8�_\�w�<�CqU�hm� ��|�Fԡ�D]�Ȗ�����}���~�Pĉ7T?1�"��$�������5���:�����Ny���l�q�nB7�JkY�Β"w{�(��H��[岊Qq5�/����`�Fͳ󸾬ӥx�Cs��ن�> Bg{�W �SS"cG~i'�,�{/��E�E��߲N�a����˗�0�xW��1>�@���O	��(�K��ۛX�uel��r)�G���誃-��7���U6}�͈A"A�FQ��D��}�}	7����D^����S�^�\�54���
)��KZ�5|RX	�1�F��`��	,��s8Ȓ��^���n@��rC�h<���P��t���Ņ2�u��ޕ��՞89��x^�y�ތ[O�����۠C�Pn�|��Nzҡ���`+-b�F��{�@�8 _YY�����[��j�C����/O;'��%�-��$���U�&��u�їn�ᗃ1$���MQznv��D!�{o����U��[�V���sEF���`��P�{��$�6�>?��=OP@������>'���N-�����:�AO![�4�M^���)V����n5Z�\%�
����	�f%�bG[�{c����¯����IH]�I��?x\�Y��ۦ�݇��e$8Yof5J�z�������xD���pPQ��`��k�^���B�tW�z�r�r26	�$ľ�Y���*Ē��� ��͂��o*:�E�[!D�Q���j�
�5S�m��#<Z� i:t:D�y�i2�i���E���6�F���}K�����)�u��n���3 �[�)>@0���#��EQ��m�b�����CA�Z%Cs9�����!�-%<8$ŭZTK�ͼ�C�S��ȶ[_/ R=G�Ϣ�����kk�|���6V �D�l�z��uNe��@�u� �u�خR4�y�@�\�CdČ��!��j/b��q�8����%�������*�ا;�u�Mٻ)��Vއ~J��z�u��.�.{���9�{�.��7E��c~��lr�O،Z��B����<�S?U	�����6((��Z_�xf��}c�������kzL �6�PfH4i���*l��<+��I@��P��l��Ȃ���X�Sr���Y� �N���UN�&,{�f?��`�&�K��"��,��Ȥ-N#p�'߭�XS}��Y[�f	���y�g�3h�zfӓ����9��tߔ2�!�2'p�;��W��;��ɔf�d$dRˣ�^�:/�{ �L<4�Wpϣ".Cs�މ�C��z}��Iz��x��ct��(��d3T]k|G<n�b�8-��I}D��'�{ �#�տo�V���[V-�EJӵ��٘xŻyX�f�H���#k �!Ƹ�7��F���Yi�F?����cP�����PZQ��0�R��$+��F'�<�~m������';�5��
=w˥��"
������:�F9���������� ���y�0G#����W����������qc�z�k���]b`β�5�n}���AN찗�m�X#b�qU���|��S�]��_��M��3Gݧ{�_a�v���=ʫ��9~��le#�h��iZ���p*�Duk�2!��������hh6� �g$�� �,�|p+����hgzWa[��w����_,�xa� �C<W ��'?��o���88���i�*q��������@���5�r�ĭ�P��;��B��o(�5a�c��K�1N���{?`��	8�ϫ���I=v)W��~�"�g˹Ԧ�+�*��}B�'�`�����)@���N��ҎB'�y�+#�S�A�؝�<Qm��h圣����_�UUo5�#8�$v2p�O5���-]h|,ۍ�b�*#'�)�O�7�E��p��l��k{��
5@�,��:��Mr}0�ۅ����dųڔ���\������	r�O�U��v_γ�{M,�Z�K5�R~3�L3��U�!�RȪ<@P�S�7Լ�}��o�L���ջ�yZRXۅ�W�1T��߹he[N%0 �N�5y�9Y���G��һ�=Nʽ�v�/ؔ��l�i56.:���}Z�-Q�Q��T�:���^M�y�KVB�}(��C�*��\�(�|��̲�p� _�Ź�9���y=_⏲��d�o�"���>��	�^��j ��2�+�}k���b����@��Ӗ��?BT4E4���
�͛�a-ο|�܅ԓ
��*��/i
�����Ч�"�I)�����o�ؼ8�R�r!�F.+�Tʥ��H��H)����a�δ�Ti\��*uZo�!@���-�nH��v�d���H�R��]Ε��
@�0k#l�:��Q��{�J>��E�ݒD|h��|ns 0�VX!�v��HF<y+��+dW�i�z�
���P���0���uɽ��>�6䨣ԝ#�OvN)]��dL�e��)�N�_.���KU�{,9m���K��.񆛡��u�ی^�m0'���l���$o��RjQgLƃM�ΣIr�}��o�ow�����/�A��苇I��:B�wWFt��|�p���0ݼG�	�,���t�A�j�p��ߚ��=x��T��T��x�O�,��O��'VP��kj�H�=qs=�|�g:�u�(a�r�Qb��8�\���!%'�X��&��4��hn������d����3�Z{W)uY�>�Y�m@�z�"v�y����Th}�j����CI���!���W|Jm�֒�b���`�֘�;,� �<؊w��>�K��#�_��X��'�����`�[�Y/`��5rG�ӶD�_���j��;���:L�b����<���,���Y�QɪR��օg���kj���b�#a,(����!HLoa�P�54�n�Rl�4 �Y�h��XG��=�3ɳ��U��6Z�������
B<:z�I��#!���r���c���Q���Q��"|*f�j�\�j֞��ƙ��N|HC���;��!�m�mabn�� �vd 9S3 ���/*�Q�_Z�7r�F0�&�ťD��8++���,�rg�GFYX���=����K�Z/�<�Z0Y�	�1V��Ya����BR�� ���& �2�g_Ӱ�d�z��'F&�v���SR�T�����	�\c5X���V+�nQ��t�9z���.���%\��㣖�k��3�+=�	ƀ�%v��}p��5�s��RU�f��Q薗��F:���[{B����f��o?���%ٚ����h3T~��k���ps�S-��K�\$3�pJP4�0F��ԥՇ&H����o���YOj�������~�J6���B���^��/�����1]Ѓ4�����~&�15,�0 �C���d\��:&���K�E��͞�Q�c%QǕ��O��F!�i[½��" ��1�uע7E��.�)�<��C��Ȯrz�Cl��ڞO8w�}�0Z���(��3��B���D�v	��"�Ň��P̢�{�A��i��4����9Zv���ʥ��l�z�%���~���y�X�f�]�hx�IK��J�I����v�nCh��5d8��qǹ�,����A�Bx%{�;B�U���K��4w��~�h}5� ��F�����l���-�D�s�
�-Wz�G%��O������~�soCt�uf��R0Gt�r������ �!O�a�pؾj{98d�#Ҿ��\��.Ԣ����?�o'}hM���;���/���ϼ!=L�C��F�q��#!�8�:yo&:�Ai��N^D��D2U�H�������'X�����4i�%J�j�j�ҍu1��ej�� ���5����/K���C%�@�C�<W�f!Vj�g��.m}���@�8W��;�!)f�����#BT��+��Н2�c�n�ǘ[?k7�@P!���(ʂ�ij,�SN;��Rr��� �@;�;���(�-]*̌��!=�e�*Q�?�%�Ȇ��gz���z�;w_��?Xӓզ��獽%����<sƊ1�)��^��;�� ��&*� ���]^z�z�M��SI����v����G�4�2Y����4��_�zU �Z�gB�"�����fƹs_�b𡗸8`Omr4J���2�<�Gf�V�^�I*7�W(vw�Q&���p7�e]� �bF$��;���|�B�S��y�ZG!Ƒ�𐐥����#��;��>�0*k��d����]�gEÈ%I��d��^��y%�;��=��c�����t��+�:y�!�ԛ�!qF���O��Yf,)�B�h ��Od$���,l�<R�#�$KG^�6hŤF�����l�C����������w��.G0M[�4D+E�Y`��Z�t�Ү��HWނ��B[���2��U�ŋ��~��ُ�s�kB����jc�x�ƀ�p�Sr0M�{��;tɼ�ʮb�ꢀ ׾=
��7��t���dbҬ��O�n�����^��k���_����jJ����	�U�]�(p]g���rR0���w����|��f��k��7��=�n�mH�E�h'F�)
(Ǯs���r�y� �������M�|C���'���`r5\_��?�HgѼZ��
a�����.S��a��.�1���~Du�9�}��u+=�u�����0�q��D��}������s0i��a�,Y?2^ ����� g�`{�<$�@k7�B�[n��5g�0m�B�=\��P��.�f��J�^�IeS��?[L�{�7���C�l~���̎U����n�7/;u<i�a���(z�X"�PS���<RR�wi�w 9�Ny���u^q{�=Ӕ�e���FaFWB|�3�sk�9��M�,[���郉0JzK,���iY��D����bG#S��� [�=����UU��+&�[�q�
.����E�y!+�9�u�Ϳև�-j���8�6�m�(I'�3p��颂���[x}���I��$���%f[�����J��v��7�#?
�	����-g�%d�j�,
�����%�"�sO��a�P)�W��҇_m�F�/m���$ѾZW��p0�d����}BO�,b�l�6|8{�`	T;�S;S:3bP�c�^��C����20�mq.Bծo�[�n�S�� ���b��h���L���6'�� ���oA��z��ا�?���|1הf$[%�&�&d`��L�S�����S��u�!,6ԌzG%:P��vb�d⎭b�(�L����?br1��
��I�'�c����n���x�<���Ϧ�bvѕť �U�NTQ�"��%��z���Pm+<�����_�����%x����]a�,�¯�����W�zn�\�Lh����X���� �so{$_�,���$��OA��K�G�n��aB�[U�VAJT�%�E�ޙJ.�DH3�p�#�IG]+b����Y/M�?�!���,9�oX�.q���q�+�Ů�\�s���ݣ:/���ɺ�P��F�}U��Y�K�����neo���9Fl��É��O����Pȇq��*���n�V�o��A���m�i?����!�VD$�O����I�\���we[�s�(MGC����9�������F�_&�L=7h��`	�^*��W��E���o%ۤM��o�c�Տ��C�<��5}_g�CxR]���N�&�{pC7PFX�m�4<ʁs'r�c���¨��_B8��C��7sH���>�y���$ޙ�X5>,��L���Pj��-�]�1�~��a6���ͣ��A���(I��'��D�V1`�
N5+s�x��
S��^��C+)v��0�g|k�g�Ԇ�m'll�oD@�,�����C2�8p�_����?��ϊW�m\��n���Q\��C˽��!���w"� j���*Wb�}��7n�{ύb�\��΀� WW����eSfp_�0�����Dt�"�6a�0�M�r�`�0��~c}���1�_df,_��y��X�8�H�b�����-�2~�<f׭�;:��W���(��޶�d�dq �yR�̌���<F���S[�r��\�����V.��ER���l��ˠ��ܴ����/�Cp^��ϯ,�-�o=4Ȃ1�w�8ܥ(�a��_�S�����f��g�&j�qߐ}	#���Ӽ˄J����3�TJ�V�qD����k�}��>
M��_�=)�-�Z���)�H,ڶ����0+Lg�u�����a&��b?oS$R�$a�$�DD蓳sÏME�H?TYs���e���1ƹ���Y�*�Ǎ}��;9��/��<�aT��_ b!��i�X�)����=�}��П�h�i�ob�>f��@��s�����ߕ�D�<����l��fo<��oܳ��hB�̟�3�E�C+\���������0�"�k����𵊇S���Bَr @zO7S�ø`��x��޸1F3��K�P�������rSl,م���8g��ս	G$3w�_�M��Il89@`��*.�Off��#gKm�Q������<�+:��A\F����'�%�S��;�L7�<�`��y�f�ɂ
�\2\��@	鲃�3�4���Q�O�����O=hU�~���ÙZ-e�l�	F�O^u��1�;l�-�����_�>8	4vä���^c`x]z}�����A�~Kuk��a�_�a���!<�U(��G"�o~H&-`-��zt�B��O��O�Ȯ�?��c!�xkUu�3�_߉a-�a<p�i��3�[��Ŋ�my4@1��VP�,�5�2G-�)�e'Q��>{���$�6��|D��.��Od�\�r0�6bz��[S˩�;���*�=g�|�N;]A����������q~y�	 o�3�H�,��߮�[x}��Y)ǞY �f�a��(��9�>Լ���5��j����x�m�C�{�:��4�
�����Yi|�q���ր����5���Q���S���si ��~�󲖩`���9@/�0d�L&>�֝��{[���k��u�_���k��^����H�c���Q?��&��lt�F �o�̛���*n��cl��j�C��'=GA�O9�7_�c!<��6���3����*C�|D�FGr�窨.��|Ȅ��l�1��-���գ����W=���s�4��kݝ���Fl�,�]��^ %�7ܼ�/��H��?3�����S3�Vщ�^�>vn	�a�YP� GY<ުMM9�E"ϸ˝��M�+��/�x�O�g	�QPt�!7ҽ�d��J�,�q�Q��głP�#��+��Y�;��Ƃ�B��}�"�r|���o�e�鞄]ݼ(����u�a��;�O�^�/hǅ��$@�N@��dqA.Po�OK���3]���Wp!��pp���`�!ٓI�->���ªlG�����Ew��_|�>;�[H�i��i���pyU��`�el�q��J�����>;�5��R ��>js��76z���S�n4��1�����_L�@��|�̖QsqK.C��<�~%�/�����*{��r�N$*[��eSqؘ����/����+�+֣�<���!����Z�]��/�����~
�n�(��D�����B��>e=IS���7�p���35.�Wk�zaU�l�u��\�(x�����e"�z����*`��Xq
��<?������~���%A�r� /45@W0�����(ޤ�3�䊩�aה��y$�о<�5��͎$���NOnkQ�*;qe�i��?�b�4��1��{��|j��⁳~���1q)"��e�SP��������av6`8A��9i��皫G�9s͆k�.K��{�j���8��~�#��E}m�di�E��c6��M��ct��&�%�ܕ(N��Y��>���N*���~��R��M�Aw��	Ү7��[t���ļ��N^��n��5ޏ�o�9�UJ*��.iR��i.B(���r�����GZ�����DT�}
e��ٌƽ�פ�=�V�T*o���Fs���:��AZ�_�� �e���f�`�����$z��C�����9�����V]�V$��C�+�<!d�-P��	����E��������C�����Bu<?�(�{6�=�Z���6���867�OX�k��2ˠ�|���6q��n�"��G����q����K�����$)! �ᙅ�
�C�!�5��$-v�ԝ��i�ob�q�`�}�]��S���N���8fd��H���&Gk 7o��QC�27Ot/�p�Z�	��%�u�ך�c٪�8�I�>h��*N�z&T1O#��ݢ��+�Z��߲�0?���Ąz�g���OX�p��t2oڌ�B�67\&��|`%u�<���_��w*lU=wY�^�iH������?���^(�Ӭ�Y�@���B=D��# �~�p�v�#!���4{'���vvE�kٮ���9���Q@�=�4�m$W�a.��ܙ=����W���y�� W_���P��9׆+�Qƚ�&�G��pT��jt��T(�������k#�~�7�ӒJyq+ĖQ���ͱc�������,:�|��rM\~h�NC+ �畦�1|�ob���h{6qn�r�_�x�z�w��F�z��]��aE�m%{�l��W7�Cz�eFj
kGa����a
�	��7`�M�D%.2�Vx�3�p�?Tx�֕x��oJw��`3"�Hr�֙�n8�������JP��f�	p�F�/���|���V���p��/��Yh|	5l�u��
� �u��� ���+v�� �O��$nⳉf���>N�&�R�8��M��A-^�Mt���u*�_��;(N`~�ç�e�~�W�w�p��/�3ئ�5����Çj��Ű�m�I?�,�����pm-eb�`�j�p�0��->_��s����t'�Q�^��t��am����J}9;ϲ�۾cD�4����&� 4a��<�K��ґ?���\�ː^'�l/�^#��-����������ޒ�%H3=�juG]M��'�D�U��b^q�TR��I6��	� �SC��$bF�# ������Rs�%ϱS~f�	{x
E}s"9��gA���|�{����J���nI�{�R�}��)�zP�׹� S����6N�y8��\-��L�=��
�����1Hj{��@��k^ w��<~�y[)�P�㘯Mߍ�Хh�����&��w����_HH�QC�kE�_�T��4�po\����S���0PZ�U�?�Ĉ������~�:Y�\��2�'?s���V
�_�XoT�R��P%aRx ��ϝ����@�Ӿ>l�Sb�;L|B��-��FH�֚JC�^�,�*%FzpƦe�	�� ���Ēw|����1{�"X��Qׄ�[B�B�|z�FU��P]����R�lA��>�V1!��>t�?=u206�]0d��+.�D'J�����D/��,%��YUq`��/� ��F���]�%w[Im@�Yj����\7�6e��es1P�֣�e��Ln�\[�?@��D�k���l<��k�su��og�m9Ɠ�Uџv�ڛޛ��G���$���
�1������#��c\�R� ��NZ�X��_���|���u�}[(������Oc�S�6���,��m\�0�c^W4|pL��g"�z��	/���'�m�^F�$>�b��G(�3l���Q6}'���]���t�[㇈���p��8�{�GV/t9Z�k6�>FQ
|�Z���9���6AA���)��#&Ӗv����D�΢?<b�u̞��P�=.�1=IxU�yF9�n`���� 0�(�(h���ھM�p���D����؊��Lz�,��n崑��ف�xGL-lG�^_���ȘJ���[�5�"�'��rkE��������ƹ��/
"�����r�$��g�|�z�n�����|����Q�&&�䠽Xfx�X�/�2ڶ�Bl��T�p��T\��0�a��1Yzi\�&�ۄ��N�^�l�I���G��:P��T�2બ`�r 
�%�c�KJP|-H�]��;KJN?1-_|Z�%[$'_��Q�U����n� �@uŖ�`vm����	Ë� Kg����&Z�,� �"�׌�|���DiZ���'�L��=#�����6���AMt�v.+�BrÛ�& ͏��π��{d>�ӎ��g+d�����J��K'$<��ӊ�f����������1娾�n7�`=�L�V�X7���e��������!T��\/٠
��H𻄻��`g]���a¾K?ŗ�g>��Hj�ӊ��:���~H���,�Z�~$�u�a�^��d�g��Q'�
;V�.������\�e^@t���L�)l%;�e¢8k�-��� VA����F���B�О*	3
��G�\�k�jji{
�O]��
V�uXecj��ú���?�/�e������e���D�dK6DZ swT������/�ڥ�?���93��3�j��nX�������6���M��^P<�f��o�PV��;M��B���fD8�o�6��4{��b^��;m�5`�g�����Rd�B�/�������i�	�|�7�,YD��k��)!0!�E�auڥw��j��L��15�M��#徚
آ㖬�Tބ�j%f�+	�}�����S��~���Z�+p04�S�@����C��~Xr��Pu��:UveJ%���h޿�V>�-�P�{_ ip|��p��꺨F�O�j.e�Q9�Eq ?���Ju�7��,m�6zi�˂,��� ��RR���5c�{qg_Mv%0����$�������!,@�𚵁tz��,Y@[I��u"3�d`؜�W�R�O��N�V�	���eܝ��*��wĝi�`0�Q_� �Fu��~�k@jH|_5��y����v�%��&�>%=��t*>�7MIAVz�
�1>>����vT�����e�o�.�� ��}���~�_���V�2�g�]�p3Q �hʗ���ݽv�c���b�����X�h-�)����~Y��m�I��dc_z-H3/�-ǝ�@/0'�2���0dRև_�"@�G�r9�L���g ��a8ں����:}�o�Â�/���B�\����0�F<5���o�S7���7���`�諆u��}�*�j�5�v'��紳<a�7�կ�ǁuxP����'21�Y���%ku�=��D�+M��L~�M�Csfx�04k��Oa�ؒ����wa��ɮ��Y���߸��7�Z�Z�� �8�G�����T	�V�J3��Ń3!'�AӪ����hs�w����wcX��2�t[[X�$��tW��)�<��M$�7׽��?^Ƌ���"(�Ϯ�o����'���ŃG�*��o �Y�>ü��ypLΟ���u�J�e1s�"^z�>|4�� ���mq[��A��"R74̧���i����C¨˱�~ᕍ�7�!�D?]��91PQ���eufU������0{`���kV���U�N+�m�6t���P#���:*"6F8٪��9���Lg�h`89'�ш��S^�y۝��?��X���@���R5\�-����֊���t�5��F6*ɯ~JɁ�Ml�κ��f)�7|*��;d�k��7��!K���A�.��k<=��k(E^�����9�%�7��I���OoT58}����K�L�uu�FzE���y�$=��O3�}����84]������2��1)>F7�|̍|Z��r�1v�e���̆N��}wG S����9�`�Gg�
�� �m����nl�O���7:BkF��s}�!��A�����9(�-<�����kַԡ�<?��]M���4`S��� �ΰ�Uj�$K�Z���B�#(�$!�{�;�B�������hf�m�"�D�6.B$���uo�$���N,n��>;�_\��~"͸Ȥ��t ��ݶղ��M��;�v�K���G��օ�<i\�?��I�x��dJ����G�����'� �QI������S�ύ�r'ʊ�A"If혙a:20�I��$���ي�L��
F�D���#��X�Q������i.��5�A�^�ǒ��j�U"��aY�>d��@d��2�yQT���UX��#����T�������Bk4	�=Q��H��됄<���⧥l��Lr[�V�A�oA���ES�gQ&����~�M�2 ����ؘ;Gn��p�*��"
��?��
,�~�\�jK�|����m�z@Ʒ���*��tG�Z��so�Pp��R� �I��f��]kj+8��!7�U�np~����O�j��c?>��%d��
��`�f��m�Q�y����2���:oO�����Y�ߺ��� ��胵��X�%�OZ����V�׼mY��Oޭjj(��Y"Q���̏l�6S��Ⱦ\��g��n����ɸ�
5�A� Xh��.C���<��;N�8Qo�e�M�k�rk�rn�f���n����(��h���	��K�/�j� qL�랰���B��i#L�\��!��mbZ�� �YM�8l̾_�	x.���*����A�<��h\�n�`�4�$g6Ν'�	8R�+�ǂL�t	��+ؘr7�'��~���m���kO�a�o;xp�[�қ�з�i^�|���Vz����r��7������p��I|�s�����~��)����N�a09��e�
8��b���2��Ԩ�.q���L��J"4X��O�B�>�=?>1�{7BY
~=���*'��gTh7���Ȃ�wF��ZERW�ѹ31����Kg}�����@���w�SS��5�u9��̒Lɲtj�t>i�G.����Ѓ��-���JH�~��W�*��0�N%a㣥�$�	d��B��3��;�w.m���R��m��"�,�2gG���;e�v,�5}�P	�6� ��kR�
M8��1�
�����Z	-b�*�2Pj>Xa����l��	��T��Y_9�L��f9F�U@�G,�@rHW�g햧��_�G�,c����d�� ~oC���<�Ȋ�a��_�C̟�7:c��n�@bK/���ַ3�\b��Z��y�g��ϼD����1B�LW�a�)� �C�w�P�Z ^��bG/v�K!�[:7�	���L�j���%��4��T%�e��]�@U:��
MmAg���I��<���D�'���~Y���@3	�y�+�nI�Y�?�n,&���!