��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|8���e5�I��d8<��.�l~GjqG�F������ӷi�FՑ�!aX8l��s=I�* �3J��y/��D�)�}�űv���D*�_a?��!L2�nN�L�4(�p�-��M�h�B�~f/�S����@�������cpd�+q���:`�D1�~�$�4[?�vw>��A����8�N��	>kN�R�FLxs���t~Ʃ��0�°]k:+TۭG�vb���U��b����Y�jWz�F�\ړ���D����S��Ǐi�sd�I�*��
-�kdu=�e���x{!c53���a�^�d㎄j\��X���]�ߞ�v]~�3��YuD�W� �C$Z���Jj���XfҼ	�fr��@\$���)HA�7��۴��<�!�>pB �\1wt%�3O[imؼ�ɪ����;w��4�QPl�>�,`���Sq��j��xm�d�?ٖ���M�2,�B�>����|����n���E9I�W�1����,qj\�K"V�q����M��=_�̠ja?��<�\٣�^j�g��\#�]Y{	<����poNVH�4;W�gr���ϗ�f�o���x<!=XI�˅���<N����O���HV0�ʕ�}�&���!>�6�&�f���uYP��������oQ�ե����P� W��1�#9�֖4�[�M�*�븻�����Kwp�2��sާ�G��#�-�2�$�!�,qD��cJK�3������F��vLG�Z��x#���+���dmy���f���Q�'���b��٠�X�c�r��������Ҡ����1�����.���F�h�?ìz|�dc�z<S����A�K�P��)O�/�Tv:�_|F�-�� \'ܮ̈́��k���L�Y�z��LK�_/X�s<` w�ձ{�ƍ/|�&N�HƤ0�(��I�V�kfx��XDZ!�%�7�:��qiw��2j�s@lB�2�,ٖR����}�e �ۊ���R�&���jH��C��%�Gw=�Y�C#�t��=��p
�x`��?v݊X�G8|پ�������.f��%5�U3D/wG��d��C�����bmM<B
���5��L����/M�B2Hq��%l����k��P��$&�9f3��M���T��� �0X���i�x���@Ud�i�/q�T��a�"`_�=�{j�֥�:�wD���%�~��4$����_���T�g�eȓ�1�V<��V�t�@�~!*H�����(Q��7�p6\�4�|4`M�3>? ݀�!%�S��v/\�Fi�c�D�k3����b�׉HH���7��Qc���u=W�o�;��c2(��Jo����.���[~,�\l �D���O��rD�����F��/���H͡x�&<��E���㜡ŏװߣ��Q_g�r�m9�Yq�m���8k���P������/j��9���=�pj��o�������h� ���/��0p�63x� �|�����v
-�x`nNS��w�/D3lJ���'u��:���ڬ���>�܈<8vL�l���$��/>A�qgW��Q��N ���\�`yp����'򦖭J�6r擓�O�ϓ�L
[ ")�_ �{�Ok�*;��Տ�Q>�v�]����j?���kVV�E�3�K�y�MM�_~1�������y���8'��l���6����K���!��*�S��7WJ+�-4��FhF�d��ǌ�@����,���x�~����C�n��b�����1v �R���8�+ä�i����PZp���U���^��c�_�~���C�9BFc/fw���L�f~���f�EȨ�����^~�G@!��غ�G��Ȅ�Oz�&N\n���V��|3�>�����W�lN��^L�F�+���9����ո��By 5�S:��&�LY��"�N�b����!aC�<e��K=�A�&>�`�V��X�#E���܍~P��(��g5�p8{"���}��'ƥ\rP%�'}2����E�t��t�Y�}h+~#W��9]ı�Hn�x���	f���a��h�-�&�>�Z�w?4�� �0f����̕l6Z?.cX����`a�����T��k.�ܣ�����ᥦ@k�Q��w
��T��i�&��?zO��0�*�}�G�ѕ�p���6*V�S�urr;NN��D����e ������dS��[{��~����+���|gA�h�Mp��/�� 4��R}�@x��-Mn-�F�W�ř��N0�F�x<g��%Be&ո��A����7�w�M��/g��p��8�p,([�q�tR$y�N˗j5.�P�z{p����USa�����)V�̲˕��q�-1�:�d�|-���eަ�ҁ���*Hm� �A��Zr��>���.7r�5��]a} ���qp�j��!�頗�������-F>�{�s�{,��@#a��>
]"�?S�MI�%k�����'
�}bؠڸ
���ꮹ&�0����hld�!>�������}���;]���	�	�q�W1��x�D	\����t�{%{Ԧ��)��"	9v(3U��s�A.���&x^�n�B7��su���B��A�����Q5�x��2�އ�����B��jky!/T_}�ގ�^R&#��PU�P��5@:,=��AU[�[`1������ 穸ܡy�O��y7������y'�.�_0�v��s@Ω��.D�Ŋf7�PD�L&�N[P���%vl�%�I�w;
�M�ۣ��|���Y-O�ث�G�5>�"(�x`�[���ճҗ�4v�q�Hl��)�����Gc��2���:����ZP4����5+��l�­��s%��r�dt<����҈,����'�:fP�)C�ѣ�$:aJ�`G�xH�:DLb���('n�Ysq��G�>���&�XH���s��������)@sW	W�w��� x[H����D5h��P����էs��=��e6ыԀ�	�O<~AȎn�>��H�#/b�o �X���}�����4t'��j8��������wO�o�I1,�eΧT�(�pFj���E]��[�v�~�R�#k�w�Ea�o|w���f9��S#}�3�P����'��Q���sٵ�:�XB�v���o�ӟ�Boh����9�Mp���6�!�1~��I��(���Khԕ�T��ٓ��ա �2If�}O%�����m�`�^=��&1��a+f����nA9��L>��ۄU����av;�X���?*���Z߳4Y���K_hW.���|9	���D�	p�6ʁ~�R�s/��n�F#X�g�Կ���I(�I|�s�Ԣ�.���#��m�K�cꮀ��P��Gx����!=�?�VsM���9?�"��iVĳ��!�z�z#�"�
lOO�;���TS�#x�wr��Z�7
1�]�U����0�G	Ƥ
�m"���x�*���e&;m��)�B�h��u�#��y���̗���ȅ[���*��_N�:׀p�Aqt��7>b��De	���`������2��f��w"�*j�n�i'��1�Bl���ˊ���^_ě�cZ��HT&BZ�$v��)��SuP�,'	��{�X7!j��lb����[H���>�/���ģZHw#Y�o=O�L䏘��V*�R �����x���"	�䁊ئ�6CG���P�k���t>	:u�N+&'�V�&"o���X���{L2�� ��ʝ�ǥ��"MH��4�8���8�2���T�P��%��/��$�����FH�m���]G�K���_�j�Z�]��R�r�&�=�A,�	��SnT^����>	��G�l�A�I��7�+�����2E�^q�L�T�T��T�w� pp��Ӓ�
I[����0�=�)9އM�96*�W��vń�0{�t<�ߓ�q,�g⛔�2��'��a���iK��@8-=���?}�c������T���t��`�
!��;��xE�Ԗ�ɦJ�G���n�1���N
�P��"�gmN���x� �@0;t�
�Iӆ��Η�9�\Pg$��[0��n�~�����#+��b��[g�^�#d�J���4�����V��~"��Rlŗ'p	Rq��Z��H��~o����n|�e�zc�Bb��	j$�@���+X���GV &��LRR�w�����݊��9FLV�l/��E��ح�y����A�O��$�Ů{Р��љp���ݙ�������}��]AE��^��T,ݹh���U�Ww��1H�A��-����ס�>D}4��X�1L�*�G:�A)�z��b�E�1`������6ڨ+�Dͩ�`*�a�d�q�4G�chX��[�q�C����ȗY'b7�g���o�h՝�@Q��B���K���OX��5�¾�v5RC�
��7��m&��K�eB�`�.���Z �������g�&��6�+�ak�]b'��P��P=!I$�����(tQdϸ�81d��F�it�ܶU_�������)�ȶ�A�x(� ����Q�����{�>��[��ɗ_Օ����Z]�gţҥ*��ݣ�pq�h�o�C����rC���gQ��#�� ��4�%�|�B+����cC�򊜦��o$���H��¶�E��W��RS�Ϥ��.�F���vN���T��"�̯�;�^q=�2��ި����Վ��ȸBN|'Je�*�PW8Z��d�������p���O�<�~|cݯRh���B����z��&|�yXC�bF`e���@6��M�W�4���1	�
�R��`Tq�����",$����?&�W{��̑�*��ݚ
��fQ)	g�ȦЄp����f���į��fb�D=V�W�'��d�~A�<
�E�8> nbڥ_\��H� �H�V]��q[d�X# ���B0/�t����2�{4�˖l��T�'�{4ny�X��>���S��^8|=s��^W�J�����NSM���G��!����[��EZu=���O�F�K�8H�n�f�&Xn Ꚛ��?Ծ*oSL�O#���g9U�e�����"%g�I��@�ra_>o��7�Ryi1��\�Z�{���(��[ϡI�@�~�Ά��4�!I&B�����&4+�T�Qe���� 3�t-�<�w��m"+����9p��tZEe��iD8M�n\O��BF8�hJ����qzE�IZ��H-{�3��Աvf�.5���I��z�(��гEHqW�kd��7�����o����O�:�A�t7�gsǈȶL|�`ڴ�<K2��Z�.��h��ױŀ��]�X������L����1����1
r����*�$Z&d���+I������ͩ�J#l���"s@>@�$���I���8 �cП�������.�;c;P��M�jp.}��K;��f>�ź�E�^�T�xwE�͊���+�Mi�m��qW�� ����R���H��Q,��2DK��\D�H˞��_
7�4�iE,{�d�%rl�b��aؗWJ�0X~�
����",3��Yj�����F���������0�5���?����*��&X��]fX g�;��L	N��2I��ດ\�ǝ�����NM�z��W[ �i9�j�,�����~�A@����%5ޑk�}��a�Hx�tģ��9yS[���<�p#BO}jNq����C���7i�D�\Og`1�?�Y��a0�5^dmx�@�JD��'s��Aa�6y�_����sp |���HGtE�R��P|���@t��Jeɹ���,��pݽއ�<}�e��>ۍ�o� {���yO��q�uj�n�x�_�#7�n+�m�EԂ�G\稩��������l���Ȱ���~9uHK�ݥ��e�{��4aE���b�y����
�L�,j$ҔS���t2Щ�w d�Zy~�+�g�Y2q����ز�S#�)�Ɨ��[�Y���������W�ir/�/F�U�O��/8�r��x��$Ƹk}���ㄎ��t7�6n�JZ+�-B���MXp2�9w<�>^?رWeO��T����HB��M�q
�;�����e2ryX�����6Q>���[���!y�!DIXS��ܿB��&�V�>�g�Y�˃�6�GϦ&h�(h]���E���T�/stQ���H�$I�峔�q�m~:G�[p[�d��>�V6��7��?{�3"<;����}�P����E��lܰ��X\���T#��#��|L��d�{;ц�m։�N; �*�����lB:�G���#�]�ư�⒂e=��h?��eT����Z���Zd���c�f5J����ܿ�`i�7��{��>^���BS�,$eV׮���b?wN�5鶏�R�W
Z��h�2[�7I3r�ۖ"�p��j��tF�3����[%n�+�1��w*��hZ|QC��F��+U�J���������t�U���Ұw�\S@�`��ŭÏ�"�4��p1�L%��֮�7;��*��'��B'c2dҁЎ��.�EÊ.�C�rcn(��f0���Qg��#��td�Ŀ����(��ӝi�Y�hU����"�%9�~7J|�7:�A�	;��� P�E]c�óf@s�����mO׫c��4�}��]������ūd{oZ��)�\fjM�?)������ښ&��=	�����>�b%h��i�������?�qKXUN8����6Y��g�h���:1���Vue����Y��dC�C-�WRm|��eQ)�A����b���ch��\�3�'��3!>]nT��ha��_	}1z��?���f�x������z���4��S����B�Z{�_G�I�nO���@�(T�
$�V?,o��#n��<9lB�q���-�`kT���ڽ@Q�O�UN $}q����'�ϓV 3�<�8u�wiZ��P��ͺu$��ԡw��O��Zjcu���qU������T�\���_��V3l�~YZ�bwXP�K�����:�G�͒>�ŭؙ12A6�s�k����������oZm+<�I���
h/&Q~�%h[�Kl��t��FZ�n����|���!¢i�oȖ����oD���%$�m��N��$E`X�s��vϸ��ǥk�Ѳz6�DƸ��?U��{]���u�O˴�,��y6n�ܴKb�ʪB-�A�p��x4��n��E��օܞ	ڛGYK������^�/1鐑QW�!.`ۻ�bx@���D	*��7��1�:P��F�b�6��μ�!�PV���S$hoN���σ��tc���؟'�q9�#��Ͳߑ� ����RA4G�|��r�) R����o��ұmZ$C@{�v��L�Ƌ�t�>_ ��/O? �]
�`��^o�9�S�TԾ���fS�ᘏ��s��}��!��?�i��;�f�]}�%�%���{g�"j�q�)�5? ����ޜ�����ј��ހ��jF�5�,am��ٺ����9�B���<�q}�6
�
�NV�ǣ?�?D��W�h���l���ԛ� �3�?+��2� 
�1Mb�,�'�SPO��3�z��_r�[f1���:��U���jۉÄ钜�$�U�yn*U>�8�^�����ؿ�Φ��E��`K4%:�t�x�H9f��ITG[L� �{�Q�8�6.qO����H͆��Q��z��~	�al=X��w���.��U�U�0��ت�ц��~�����vFX�'��/��* �::���v�Xg=P\��=Q;7��¥�K�DOU��)��w�n��} �Y��}E
o�x}���+Z��Y�(=�#�����U���7B��Æ���rN�=�4�Y�Wu3���9I�6�7��@�d������qp��O�qV���(ۙB����ť��e�l�k���"_ܸӛ~o��? `��Nԗ�"��m&�`�|���$;�ɺ!�F�&k�q�آ{�V��W"��d�w�_UڢrǙR�I�
Q�B3�/�5�Ԩ����@�[�vFpq�&�#�*y9��Vѯ���r���r��3��>�eߌȳ`��z�ٽ�WL`�\�Gy:s�npr��֩x�#���|�nvŚ�����U[ (V�D	C��d�,�P�k�F>S�B�0qҋ�(�ZhѴ�2����Ű�b��Ŧ�Ⳁ��TbN!��%wu?m���lP��C���A���Ӿϛ70Ţd:w3
r��Ā�@p\R���g��N"TQ�Z���	qa�z��/PG�'�-Cʦ�<���E�w��}x�T��Sd~ۈaHLh���v;�4�\'1����%1�Ӏ�^�;�w�#�:��j�ώ�-ZsP��z��~��N*-IsN��0�jV�.�2QC��r�'r�0E�!> `I��2.3(�e�2���$������Z��?�\{T�im�P��+(_�ff�[V��N���4ĲGϘ��D�Q?�y���yf�u�ljS�������T�7H��0��)T�O�w�/D ���1��i��~v�Ze��wk�	^�����Yh��hqA�ՁŚ��%o����pƁ���kj��TZ}�k1�5�Y�$v9m���,��Wj$��euxʒ:��'6�(K��>O���lZ����O]Σ0";da����j*�\��sfܼf������B3�Ec"\�ޏ=��.��;Ѵ�n,��o)�V�Q��a�'�#�í�6X�P��k��iď�������>逵+c��(�8/��;�#BL�'0���@�ď�)�ҙ.���ϙ�DxQ�=mOx<'�Va��nO�2���?�R�Ӝ���zhW��F�o��;*,Ƨ��������Ĝ,?�.�����C�sZ�^�Oܠ������/=��,�orbu����L x�@qvh+*xzxo�ކz��rZ��R�n�|��b��%��F���6�J�Ub��m_1�陎����a�m����t�!2L(���Q����Q>g��FYFF!U���˲�4�h�mz`{!Մ.�P���,�A8�Է�﶑�n�IoS���'0���!Y�s/�"���y���{%E�΁̦�1��gĲ�7���9'�W4�G�d*T�@h?�~{)��)>&?Ni%+\OK�Oʺ��")i��T��ښ�����n�n,W�բ���
��Sb��
��8PCg��횴��^�@�&�`��8��<�S+T�OJ&�V�ίCL�KeȊй7�T�&�R2�\���Gd�� ��_D����������jZ.�5PwK5�vVz!e��>��DŻb_`�_R8�L$REԶ���T�	��#�J*�l~|���)p�d ��ZM��=� ǿ���rs�S����R���hN�]��CU���6u\0w�.�o��u�pv�s٢�H���>��A$�ȟa��J��`!���\FJ���?���[o4c�LgB�K
2����9��6�c?V߂���n3p�y��N�CZ��Ɣ��2��S��ꖷ����n�<5����iW���Z�4�0��1��<��>�3��V�������Z~���0E޻%�M�x�̤|�=ul���ɐ��������؜%�b�J{����.�m��-Z�e�?��F7��en�f� #l�uU4?s�gFW&V��2n�Mz�)>�zI]Kh^������X%�����0���c���\����O�Y���`\�n������ �Fēq��eV��1��CВH������n��^^�k/��(�����U<��f,Z{�$�BZkg��?�2�2�������I(�{O���}؜_4a�9�%6Fҭ5�HG6&l��J�fqj4|�_��ae��	�7џ�����S�DV�A}D=��8 ~Le��!����[���W[y��.�B�^;�Q�i&h�ns��d�|�r7����{����N }C���,9=�=Ӎ>�:y�4���D��]e���]���.�{v�8JB��1i������k�v
��S�@���$nI	��[~C<(�et�A��@��~�v)-�'�&�i���l�}CN%Nr�]�8��d2�c[`���5R2�=�
G�Ѳ4�����7 �q��5T�lO �}�\.zt��`O}-+�������P!�SbI�fՇ.�@�%���TI*�ꄑ��z�Ȋy������Gzp_#�>�Sq��}��o^�nx�h:z�>��9?S�1��ŊX�`ɀlA܊f�.yC֮��Z� �N�PAiH� �&�.��Y��-���f5�يB>fO]0n ����F��2C�R�۴<�"���1L��֟[؟ꇉ��Q�D���y���Y���C����¿��n�گ�!X:������5��ϋ��X��͜s(=�i_�N���r3��MGv3�/�xq,l�)��$ۤ8d��`���u&��@�=Ӈ��<��5;�O	�~�,g#ƻV����[!�l�l���^6�X�^��G,S4����Z'�d�yx�x�9�i�
���"O���8��_c�p)I��<����Ol�����8�Q-�����v��t���`s}u�? J�R���lzo>R�î�t�a(%1����*�t��uV�D���݂���,�yW|%��E��k3,�����iJ�Ϣʍ�q�	!�\ym��\�6�,�7�]
>���Y4����.sx\�;]��{`�%& l:X�L�b+kȏ����@����Sm�;䌥TͫoQ3]ٖ�j�������'�1���]Qbͪ�M�F�GV�Q�����t��}|/Q���<ۛ䈑N�a��_�������!5�FǏ8+��u۠n����Zq.�k_od�
g��b�ۓ�d�7�X}#=t~`��k�B�e��!�xؼ�b�x�r.��)���@�sQٺ~^�{c�*�g��j�ˍ0?gafŘ�I�_g�Ԟ`�>jX�%(Z��w����OqqĎ��@>[ Py�P;�ן9#�Su��Km(��D�7ώ፛�ϖZٗ�*��;b��� �c�u<�Q{ny�-e�f+z�X�,))[ Y�f|�v�$�c�:6$����@8���z��;4�� BZ��X�>
I`��b�<�b9l�~	#	
|�(���Q�bu�c��p�^Z�ɸ��~-����,s���hOwS�88f�P�/-�'��G ő���i�̛-��t[�J=��u�)j�J��CX�ʓ�H(�����Xt58܍�J\|�+Z�@���o.w��g:��#.l���a?�tFO'��O�� �\��1�����AP��1XI�+�!1֐"�K129з�8<�-�Z�W*�MM۱WW������Ze���ܷ~@uj�ȭKj)���v{�����t ���D����Ӥi�<��m�k�n|�}j�p�q@�XFNk�&����@	�K���B�D?�o��G�O��u�+	�Z����?x%�r�3Y:�(4��d���[F2��Z��@7|��t��Ԏ�;_�M��^]Q�2�%���W�L���K�k3/�BZ0�nD���5[G�Z�:���&�1�v��w,��:�K�r6����+�o_$�7���za�=�p�ڐ�x��6�����<�@�LS������-%���Q:X;w��4�&T3Ӗ�qR�n(�O�m�g�&�_�~�n�I.)}�^��*�J�3���p�U��d�p�:��c�E�:@"X���z��0%��t��w#^�j�J�ü�dzYT��:�̉R����{X)9�I���	���f���az/�NX��kWX�0�H�~ذw��C_p����4Ы<�V�%����)��`�,p��V��ǎ9�/�g�����+��l+k�_t%`��;�R���.eN��]_�4V����Eh ��j5~�����
�PD�4s���a��8��!ȢϦ&�
1�c�6��P$ʘz��s�28xVR��#�7�U��a���G��̥2���}�삅q�b#V�S;��_+�O��	4|����
ܨ�(�?�Ȥmܾ��oE�n]��
%���+��=b�t)��{���r�C��Shi՜�����I3���E;!�A|�	pg�>�-�b��^�*AHe!ӣ=�)�\�@�E,Z;A�Y��aq�����x�I;ih���y��ع(R:0aw��"7��7�\5�z��T5퐺!�mq/�w��`B<A�$1��B�z����ϫRl��P�w'1�j�52|�����X��Vϩ1�� RPM�	]'��1��]_�T%�mʾ=ܓ�=T�&���sj��5�NT�;���-���	���ނ�6��Vov��-��8�ۓyK�S�'Q�k�~��pq��g��^	�!�f�]I��N~�'���g�h~�#���WV�8�|�/�`���$I��(?���$��4ٽr4����biU^	[�xi��`��c��#x-�K����E�'���z�G�~�d�؞ܼPkR�M2�K�(�"�F��Q�|!b��O��BPr4�� PO�����y�ZJ遃�7-O�ϳ��ː�<�Ih0-���FJ�T���� ���N]B��m>�*s#����sW��<�2��N��fA~N�M�6.Z��P�k���o���V��|����tw!Oɾ���ra�^P�ƒiq7C����߹cT4o���jQLA�f�n:mN٩{�jT��-��<��o�b�����ͼ ٥Ń���`n�"����7��F7b���������D������-v����ʝj��#��@����Hp��@�������[��ME���'���M�����ef���ޖq���v�Q���r�@�S�1/9L���J������jc���#�����/�ԡ�,��������ᘑ҈9�
�r�*���{�Y�B�g45l�%9����i�r Ð������B.�z�)��e�6�vz}� Mޙw̛A�G�sf�������#粚S��֖��Y�w@On�xƕAl�i~Q
�Kz��&���$�y�	ӕ�ٯҥ�[L��dYE��: ��ٞYxP��M��%)?h��rU~��r+ƾ>����VG�m�%��n���ωJ<�x1m`�S���g!�鏉���1�h\g���V��37�	A�-ů}�&f�q����H��Q5�H��3 ��Ñ\���yp�5� �7��Վ�,Om��ޜ���)�-=˄��%�P-�d�g�y�H�#�	��ӝ��6\Ռ����ҿX�Fd4﫿S�����-��;��:c=n�tL!������jL*	��`�H�ڑ���@1�%�	���`��ӔFJdn�&�t�-%�m�v�����^$�'Ćה�K*��!�p��M�P��Z�r;̠_%a]D�Ur���i�J(Vd-G� ��u���c	 54z�$���yA�;NvO��A���t��6�l.�q����_�y�Z�9�9�7���L�5���Cڰ\����>�]�N��p�M�;~W��-u�?.�>�d�F�-&�V���JT(�DX���Eif��=�7���&����Q���F���I�;+�"n�Sd���Y=������
��i>���oC��.�X�GP%��Z��	�̆�!W�ɜ8��3[kB�]������V#�b�<{��
c]�t6/G��9�U�)a��Mf��K���	;���,�{s��@v���d����/��v�P�5��m�\G$��R»c�f�F��Y�5V�"��Iz�k��χY��+H����V�D�جӑx1B�ÂGC���^��m �&�hZ�V���+�9�ޥ�f�U��4v,�9�b2�hց�5��MO ��--G��'i~���0\��i3������¶���y����m���B�ma�=yr~��4>o˺���_Ag��;����҄X�H�HX�2єpE
~�	�5C��Ko%�wZP�qs#"!�*�����4c(8�m�G�����pX���9T��k���]�Y#g�D����㫯�+e�fTPKe6�$��{>l�z):�f�cR������W��W��ؾ�t��͚x���SE����H�@h�b T��:�q@G�b;��wg,�L�̡��})2`i�E�!@pػ�����Uѫ�_W�
��W���d�#��jҳ9�,� j/�8����c��ux�q��JB�t|w.uF_ ��w��ʛ�s<[��6�U�u�A <�`Xz^�?�\li��*������K�4N9�7eV�;T�$�P�ǛD4�^�a\18CJ�E�TE��fv��WC�C��<�m��Ü��x$P��%ŵl��Bw6��`q!�.O)��M��ɨ�N+MJuy3�L��[p��r���=~2t�>��� 2FP�vhz�08����'�\�i!��uɡ��\qh�t�Y.�αq���g��9�)?-1G�`i��%���:���BZ���]��	:��]0ǾA��޽;�5�X�<X���!#��L��lDO�gÓ^ӷ���g#iІ������r,�d�r��u�|�(و�5���q�HDK���1��V�g�i� ��r�7*��� g�~�J��@�2������=^o�F�٫�fZ%"h� ;gjl"ZLE��A���+T�-�U�Yh�d04��K�iܦ�ym�C�5����T���{S�*g���G�f lQ'h��H���5P�����ET|�E��Ta'���;nPa5���e	}0��Y�O�� �[�W�'
���f�Η,����Dg��,����b�F�4fd>s<���Q�(&��-=酑 ��׫������t�;�<��D����4�&![|kKK�,��曝U���f+!��ɲ!�ָ�xZ?IQ-�<+���٣ �^��Mn�,���@<�AQ����������?Ndb�-�s�xN�������-z�������"�q��=�ΰ���oCvF'�w�S]:�iu�U*>o�<��Y_��̵Ĵ;$��A$���� K��'�s���%�Gݦj>�_�����sS�6�t��#�t;�Y4SBIr2������	��o�Hj&�,���^u��V?�uV;�bk��5�7���'(����2k����j�ה�y���p:��;Ȩ�Yh�l\I��r�Y�	��>�#t�\�6��
(7�Fx t�紁&2$�=C�u���_��ݢ�f�I:��⌉68�uE��C�Ũ-��6э��#��Nn���,��v U�/����kd6A�O@_�&wϰ[>�SJ��R��VYk�Lʢ�?[���}�%z~D��v��>u`�����b�l5��j�l��#z�o��-[����M���H5>��+�ӧ��*C�36��-`"fK$�N�ʗ�4�.s���No(,`O����sBqpu��`�`?������`
�T>;��.Xƀ��
Q�<�c����1T�;��WWH�Q��YW�>���:��I��S<l����c݌���ւÛ(�6|��!���l+���2��q���?K�^�a��+?/�0��5A'}_��0*nm�$��%�7��ҕ�s6��yuѐ��kԘ� ���9�
��E�c�Komd|Ǒ�/��h �� :���1j8���8�)��d����x�2�O՛(k�`9�����jS�N��Ƴ$9ZF:?qY��;}A�t>���r���l��?�E��l$�2  v��A]R�2G�<�6���	��4���-�����&Ж�_/@/Tܸq\]����{E��.�6$���ݎ��O�y��М%%o�,Z�
:u`�4�Dx��\�o�Icf��y�a�zL�ɥ&`$�TPN~(HYX�H;^���Xz��-�[���-�!�V���`!���4���7GX�~��J�����Py�86l�dĮ�+$!��f�A6<
:��g.�>U��s���i��s��S������m3�j-���h|��`�E>�tܳ�,v��ڢ%q����*�����CR;[��Q�!�葜�в y��e`I��(�Y�I(�����D�d���;� c��g� `�G�!2xG��x��%\5���|���W�a�c	�����o�[I:IQ�(����|�z8��<�x�[�62�dO��_jhS��U�h���?1���i=�gQ��d�Y)t�+F�o5D]�O#�q�P�/���]z�(6�Uˣ�R�^��1Q��Y��<G���(�1�:��
W�P�G��;�L��Vr�k�hok���iD�8���벳G*����cТg�[@���cA�Ϧ~	wk|�ս�@�Х�x�-~�֝�[x�X_����W��W����F�A���@d^��_Cb��Uێ���c<NI':�PT�ƘD-�����5����E9�۶@C�d�28>���
Y��W�x�� �Ѕ<s/�����(eI������>N}{����VIl����on�oS�Z������H)"�w~��Ϧ���j$q�U�_���]<,;C�S��������52��Z ��kH�j�&j�DY��Vu���W��$�09c�O�)���1/$�;fPj����i��$�Un�"��p1�}�թ�&l�\0�$?��Stlk_��Y
��n��f�6�z^�������	anH߃_�����0q��k`k����޾�99?�z��m���z�;'u�+�'H��*�,�l�������=��'�;w'�E�	�t�����!TR�1��NNT8�)dJ�vvn���肯H�/�&���b��*�)ڄ�j��`ʷ�X��_�iy�,g\>����%�<�ٵ-���:mz6�#��sF}0���#� ٔ7�κMITH �a���+e�U�D��������>?#����߮|��$�{G�cnac�X<ք$��se�/I�B>�l�mJ��}6n�&A�F�%z	�b���9����=��ǜ\C[8���7�5�lR �V�u�c�PN�$s����R�%I��U#�J4^6Yna�FK�ܥ�i�$х���4 X�����ݫ�.�Q*^_H@�B��<��leC��~�Њ��n3Δ�т6W��	�;�5���u�Ҡ��A�L��	xƅ�)�bIԮ��`~��W.���	`@8w�ȧ]�u�Ɇ��R���ȃ����GݩJ�='�����x�p�H����YA��FD�^o"����L��8!3OA?}��;|P�}IT�����}�]�kq���sW+wՏW�Hpn�u�����LB2PK⛔��$�6;�snOl��d.�������I��g��C�?�"w���E
�-P_" �������˕vZ�ӷ�f��^[���8�t
zpzRѴ-{(���D* `gwi"� <�;�l�
�+u�
��z�p}�.|9��ԱII�p��9Z�jxG�ּ��s���J\�͑OPm��'�p��[~���-�͹i�.IX����L�E[��+ˑ˼�\;@���\��� ��7a�Cw�@I@����خe%���\+;�;b!�v���G'g���{��B��n�;���@�A�U�s�Z["!s����@��ܾL��Pv#U�ٞ��8��^UbTA��y��}SS��|ðR��͇"T���£�lQ5SA�'���/��J�)ȋ��hB]�cf�����d.ё�8�UE�zf��£i�:��j�h�(��O9�BA��]ug 6t��z��Ƶ��6 �u�#SM��
�Tegi�� ]�-Go����%is��+U�w|����8�9��h:Ǚ�*�X��ŗ�͜�>݈N�@-l�-�T#�,;�A�����<�/�N����B�����.R ��->�e�0a����,7��D�y���\X�,׫3v�Ͽ��I�+��,�V�9/�8��9GC>��}�r=)�y��IB�s�$���yxG'jozCx7ƞ��n৿���#jw���bNm�Mq럕.r�Y��v�D��S�O�~1����Ws
Q�Y����a�;R���{@�_�t�]�sS����(���iI!U�<�R�xy0VݢO���0���;�������R.�P�fVb�hKjZ���s�h1��KJ�>*��L���q�u��+���o�=j���\fFG�3Ay*� �Lֲ��؜�*|K18�3I�5�d����$/M:�A���h�A:��\�M�L�����	�?������������55�� i(\}f٫R�"e0q���z�_�Y��8��еʃ�-0�hy��؜N��[���:7��AdU��S��Y�����&�O���_���D��Դ2XR��ĵ0[&!'/� XS6m�w;9!���n_�)��$y�a��{���}���#;�.�+ ��2)&�n�+аfJ~-0�����d�R���F�哣�����N��U��Ӿ��������a~�A��Ҁ�1sѶ��c��D#_/IY+$��S�<?~���B�n�����xm��a�bq]�m7�<\�J{�3Qn�8)~�]�g��A��*~?�X3�̒���m�U2���a��>CzvywU�����oi��EV�1���Ӫ2W��3s�_����6LA�*�J�ƪ#^��[�Æ�bh�م�H����z�U�[ClU� \�S�ϗ@Y%�|��ǹJ�� �����i�ltr��9?\	Q�qћ��8)�@�hy��-m�!����\�Z��- ͕�ڽ�?�K��P���y+����)���?\���#��C�*3fe���m����<�^<�hK�.d�ļ�_}U�L@�;�Ƨ��=������V1�X��9�+J�*�1Q<�?ͻ����-k�˷M�\�L۩���,�~B3�â��x`m�,�fF��R��\�Σ-�R��{U�|[A*.U<�@�ڿ�2�}�do��S��~����-Y�ŏ��5d�y`��� �ͼg�j���#מ3�%*��k�7L)�靘>+$�G�z���+�}peK���k[�8�؉�$�^ T��^3�z��-��5�ڊX{TΨ�x~�TM���~�C�� �wKQC^�;�n2B��PB�'\������>�Oi�c��r%ؑq�4��=�_��)^�:�����h�FB�n�,y!S��XԿr@4����3)٬3��<��9��6@H��t�	�P O�&�p9nT�Ţ%�Tokb!����;"��T2yI������I�ځ�N�,ڠ򋑘`�9�Ěrl�{y�E׿d�t��B�������/j���qS��dr%:��'vU?��d�����R�EU�5�:F���o�}MD�u�b�Zg�0G����@��"Q#��|�$x9���WKi�����+���n����t��n%y!X����S�������k���9D�g�8���1�&��k����D�b�J�)��p����Ѿ�7罓�i�IGM���W���bҿ�e����躐&��|2�L��
��������Lq4�5by�9.�4�>v�FOc����q���O�����Â�б��{�J��2k��gX9���Zx�b)8��-],AWͲ�|�N.���؀���"dw/iNw�Z%�B̌���w�����bLγ1���B����5����'vV]O�|�ъ�4���X��q�}4Ř�B�kf>���sO|??DƐyg�M=ַA�g�z�ߝo/����b��N6�%�[���E�uq�6ߑV���,�͝L?��s�U���@5ޙ�����߈ �6K/��D���âB-2���^��JK�����p8�~�F�,� ��0���(U��^���tO�ġ�2��7���Ed��U9�$���l�fFx2��a�EOZ�e��ymȿ��܊%������Pu77��S��+�c	i��yR  G�]�:�Qub�n~�w�)�J��*UNw�m[������Oʾҫ���0R�苦H�
 aE�gӍ�+�@+M�=��A�3c�jn
��]�[��ͧmd9J�	�#I�yYh�eM�Y���]
('�p�1�M!��Mf�����pG,�Z�[�:)t�'��2�P�"��#.���w�'��;�-�1���,.�^�Q�%c��b=/'}W0�tO�BuF��d}׽	�}�M4<2a�ϻ�?�4���eѪ�Âz�rwcK��ӡm\ސ_������*���<�0q0Af��Rm�7��p�mέ  Z i�LC�}�1;["����*OW ���Mm1��ŉ�-�ŵ�0`6����"���q��A��!d�-�;� _ᒂ�u������jS��g��J��F:��|~������I��"\��N���aݷH5�\bS�#�L�Ʋ�&Z�F��dͫ<답ԇ$z��`Ӧv3�@�Y��*�����I�{E�|����,�7�<���RېҐ4�|�|9=ۘɓ*�qx+��뤏m�Qf�UD%}l�O5,��.�s��{��rq��bZO�S!�ꁨ�3�"YBYI��E�7s< �.e���_L�ˇ507���_t�U�y1��Ib���������E�BD�tǉ7O��\�x�[8���g�w����.��w����_k�ܜ�t�� �H�(`P�B���@5�s.[Cx�6�䅘���N��_gg�r�TR�'nˌLA	z��'�2�K��w�/&]T~Gw>�\f·��  c�
}���ɀ���7:�
��H�a��,/���`�u.`��4�\��,$�i9��' �#ng��@*����u�I
 f��j���8�'�������ѣrS_(%�<��l�e��c�w
��?���'������smy��/yHDD8K��� ����U5q�t�P7+8���H��R�#1d+�<��z�ڙ��pO�6�ST�0j���2���e���RPb%,��z�ZLۏT/�-��7�s��ɝr@�$�7T1�������f����+�[�j�,7���K9�c�@�[�nj��g�ez�%��[��a��&(p{LrR���h�>�V�N��_�9�0��&_�4yyx���L���ؗ;��&�%_}ez��~�js�D��Nj�X��L"�;�@�7�F��X3d����(w�:uC_�Jt�AqQ_cN���8G#����~������� �V)��I���M��%�
7�y޲U� ��`�3��0E8㳆'��%M��I�\����bvT�7���M"Ș�ni����ܬW�Dj�%;9�Lj���T���ҡ��	W�4D�=�2�yL����T��Ǣ�1��NYj��E��C�u�����w���Å=�� �8X���P:��\��p]�"wS��A��rQ�>��~���!WO��h��V�ns����0�̃IY�E}hU��:1���i�=�}�A��C�O�	8"M�C�ex�X�Y����?|����5�(5�p�:��Pk!2��ZyJGO-�1��(�FKp�s8���;��A�C6��a�y����2�d!mb��μT�i�Wr^=*�S�'����4�6�~�GD��ct���{��AR�%� �ԇ۟eA	��@�Q�Q}ɠq$�	���!���L���9Sf@�+���U۠~��1���a�	,@�]X��,)�ȶ��P���&���,"e�Hiq����V +7��~=�j�8��Bo��+< ���R���o�+�04�D��
|�X�y۸=R�T1��'O�r)����f��ũ���pĉ{���2	�VJ�?��2X�o�c�zp
�ȫA�]��C�P?'�֚���ݏ(a��������2�����oD��n�85K.�ܲ�`:��
��As�n�8�@=��8�	:e�|��_�7B��d��9���E	:�f����Cp�G�!���°�$�����+�yC:�_�7#ҝ"���'J���2��<�X�C�7Y��0�ן�#�*��]}���>Jk��Ƭ��fᗃN`=;�|�����"�ˊ,QBmsW C���=	v?�H|��+����8�ʇ��He{Z~���D��]z�3�\���͡%3X��;T���n��N�uV�q�yJ&-�j�]��߽����D���{JL=�@�^ �/��Q�d|����r�rT�j��>`�'� �74�g,�}I���;�����w����LF�J�V��j���v�2G�R�Ό�ا����ɞ������-x}�-�@��Ԓ]ц��D����P��u�c1�Tq�>�UG�4m���:-xO���O�7>��B�ț\��>d���`�m'�.�����Z7�Ol����;�u�r�U3����}SqŪG	�k�6�e�;���!�1"3g���2��[k��0�@,�����N����P�e$Y*�G�_�.j��@c�G"�&�t�OY�c��\�]C�{O�<�(�L����%<c�؀�iU���'BR:�������l�	��\k,#�]��BOkԸi���_3�.��%S��j�j�z���o ��E���\����V�RA��Hs'��ӂ�ɢ3;��.x`j�أB�c�)��T�,{�D��O�͝�w���؅4���4N�컲x ;�0�����h�W��^�@�	ꏘ��K�J�[��������U�~���a�z ���Kl��]�шz'�8qa�M�0��<�yC��
�J�o{e꽞�����tJZ�H�-|J���I�ZA��%����%�|��,�U_��x`^�$u�C�6h���"��aV����D��̈g��C&${��DiJ��O76Z�a��"/_>Q��6�MQ������,S�P?k-iI��M�Df���qׁ-�m�尲Rg��A��x�l�nyH�1�������9Ƣ
�z*��2~M���:x<p��f��os��jt���d+�0v�b�R"��� +|5����rLtw�j���+H�&f�����_m����34��m^ǎէ V������Nf��'�dˡ���j�����b��Jf�K��VIR�Կ�Ko-(6Z��P��4>⵩p���$������e*�%�`׈{<�o Y�������J��0fQ�:��{h�)�yǯ�N���;X	B�:����s$b�[ǫgl��� ?���X��K}�����6�sV��i��*�S�FhmD9|rf�u|�-c'��D\7ׅ� 1	I�8�z����/m�atU�l��bOOW������.is���=���A���*�Zec�$�5�g��.(H��� 5ό�W�@G<�hU�vFM��Q�p>�Ir��FD �fu�{gi�� ܣ	H[��aN��t$9W�E�kH�cɽ����Ç|�4�7J�+�0�$M�����vSܽ��j�2� �)���$﵋��ԝ�㣖�Ej�?]/	���9-
��Cƫ*<����^���wO��+-�rg*
�*�Wo_VS`~SV �ސ| �ubh7��f�n��<n/�1� _�5�U��c�+���q>A��I�4��DZɴ*���d��$���2%|�Y�2��1�C/I��@�{��g�?;j�W�K��̍*>�B����v�u�޸�F��3_��t$<@��8U��?��w�ߐ1`��'�������b=_���c^X�=��F�Wn'4�뱛6ۯ�B5�:�k!���$�Jp�ؚ��W���~Ǡ&����x(vO�������05l���0s�ñf�tP�6Y��ў��6�r@.ꏔ�]q7e��ю��q�R>�4^�o8�1.Bm��1�+��|�Ud]�!���֎�<*:"B�EYsY�yC\��qk��+R�0 {��*��]��z�����w;�v	ҽԌU�N��r�g��]�9m��@
���H?�MĘ�c���nvӃ�!���]ؾ�O[$F� �;��X#�k������b�<�d嚄�q
wB˔Gc�c�W��^ ��D���ԋ��N�D���ڂ���$���W��1�������2�������7䵣�\�ú�Kط��%�Ef�]���wOA�bw�la�����[y�=�Èd�֩�3��`| �䚢�w����pD<��bv�*f{2d�7��;�X�`�u0�r	�)�nU#��KJ&Ɔ\kߣ�x-���~�j�QN�(+[�x�$�)H�ޒm��Q�R
Ǹ���6�$'lL튯&0ANP��{�.F��s���mP�w���`�,2���\�u�l��9��G$�Ѽ"�>��'G�*wV3Y]�$���:��I��;����&	K;Su1w#\�������x��'Ǚ��ᘙæ���S����{��*���1y߱@�c^۠�:. ��.�	ˈ*8�0y rۃ;)��0��
ԗ��Q�N�aR��jmF��	mw�I�t�j�oy�S�z��g�y�v:S<�,��� .{{<SJ�1!4�)����Ov�����mu�A�E�91��sny��p����4��,����'I�N�Mԇx�pD/ヘ[��.�g�/���̢����%��|�uY��me������TWm)� Pi��g�sC��l7�^(P�t�]�Ꚍ�]��y����@��L}~��>Q��,Ƣ�A��)��Z*������	�	�K׌�㧊5�G�a}�0�wvع�5B�-��BJU�]m�D7�V����,,&V����]���8�m� �?�~�F�+s�T h�D�ܗ1P�鏌�1��z�V�f:֔��f�{��E��O���@-�'�I��A���|��K�Y6��~*z����S�vJɝE�r�����{�A�S���2���N�b��R��E*�ϖ�vU�BJ�znZ��b9��q����@��NgV�S|�f�ѵf�a�ɩ���_���q��E��V�M	�8`l�`��|0⹑}�qm��Tj��:`ZS��,�4��>s�Q(����B���W���/k��~��U�\IK��;��M����f�&Y�sX�k��E��A�����u���f���镮5�}����O���0s_�\�\��1S�ϝo��[����gD��}D$8	� a-M}\V��ރL�� @�N�۲�"pm�r'=�r?H9��<��"��+��+�yԀ����g�Rv�Q��B�H�6�w�K��s�	}a���}	�E<��a<�OY��+t� ͯC�.ݽ��Jge�h.ZL�FJZ�6u�'�˫��b$ ���:����|�f�g����\�O7���AE��8�`��(�T{됴�џ�;Mf�T�\���I�I�]���=@m?C���v}".w{��SE�h���*�K��4s$�8d@��$Rw*=�ק@�)�_Q�mH���CIZ���y��(�%��C����ڃ0��J��4�a)�M+�|;�j��JŀW���UTF�✝���N����N$��GM_1D�$U�f�y!m �t��'��H����	�lG�xW��:,"v�j����͘�v�?��Դ�*ʙ�YΘ
,��ض�'}L��t���_ O ������AB���Mk�.SW{JQ؄�Z̴�L
����M��M��X�8���Yh[�e��7��6lJ|�0�� B�WRpW�b�pǿIލYN��}�]Ӧ��e|;�4��gF^o��N�����,�d��"Z��{��y5?��>}d�w
�JH���Z��=69�ES��=��h�M�s�1�B�4K2�e rı�q�-��t�r-`܈�q��m���hl�1ԧ�w�n�h�2t{Va���2ώ̻}��uߊ�tT�S�J�!C��&6������5��	~ �	5o�H��,����_�"��I�K� js l�G+_�rؼS�u�R���7�>��k��"�s%�y
��ڢ��Ț	S���_��d��,:=�����5�������)~��:U�+��i����t�@&
�#w��b�:8��|̱��L�, L�f��r'�+���~,�MU��n��nE��w�M��A���k���*��~^��us��'Y�^��|��ܓs�ԍ�p岪�t�5Gb�*��g��!�_v%Õ`-�{�!���_�1�Ь�5�t��i�e�:t�zmR���[	���㐅��۩@���6$T�C���A��`�y���>\��#����'e�r@��D(z�ȁD"�ϕ��d�.g�Yu�ƫ�Գ<��q!e�z�Sx����Z��"wSO�\+�½J�R�)hP/b9N��@<$)ߘě�s��>����_�ɣ+��|���db�Oi��X��W�����~Tn>ُ!�����aι�8Kќt���.`��J�����Ո��18"����b��#%�[�~��nW�������Np����B?��	1�O�z����@�8�j=%3V�c|��҇��G�O�y)x�H7�\����P�(��8/ܼu��9����v_��G;��~	�o�55�o��sy�zB��-`��
�$��4{2�jf��6=���~��ɜs��q^�BU��g�
<�ǉ��}�g��w?~��+J3�o����/]��HR+��ܙԫ�-"$m�﮵@��T���0|O����2k)	y�r�f�u����:���X��J�̟5���,�kv��u@LGG�QX�ɍ�v�lV�p�˟ư}�`�$<�w�G�@�؆�qL�)q�̵׵��(b�Ҏ\���)�_���*"|:{ۯ�7/$2s��4A�EWg�=��F�o�kF.����UE�����m٨t�kޘpN�t�Y�S���ʐ���Dȶq�/�d�|�V�5�����
ׁ�����s�g߲�p�3�%F���Q]V����J�#�r^֕�TDK�X�iKgc}J�j$5�}5�NX�i�MrQc��3�z�?�xA�����F�׏�XZe��H2]_�/��I����Ƞx[�DȔc?����?����2�ސ�����	rφXږ �]꒠�3b��;`�+��Q�=H�rE�����h=>