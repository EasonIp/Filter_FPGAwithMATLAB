��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��ע9�!�"��F�Wnb� �i��a��c��v�Ϗo@��Z2�[�Sh�+����,��ơ� ���
-�2�4�˰�=���#�B��Si���絬J�A�Ry�G��!�w��ķaB�� ~"t#��#��������L9�-Db����-�[����f� b/Q>�B�K'
*�j/O��9CB���0V �<q8x���f������8AX&�uN���jx�|k���<mೌ]�N-4[��F��	��oV9)ӻb?xq.��A��4���zbu������^�,�c��/�5�䡡�"ټ����)4o� Ĉ����OH���`,��Ƿ-�^�_	xr3��~�i~�MJ!́�<%pM�m�nRvޝ��<�)�l�;5Fǘ�T�نa}�P���S �F{���>����%���y�ԅ�RG�e-����`��L�9,�͙΂�O����Z���#q�X�H���3_��˽���09ܘrp � �e��;
�#j�h~���%��8;��긒��r�[sm�"HmA�zQ�1s���Z0�
��m�:>>��[=k���x��}cI�u�(�w3�l�u\D�o[�HE�����\�-��;\:d\���NA�j�l�^�KV�<.�����Z�1���%�E�b8�_7��T�t~m9Y��Ħš��H���BIBEE6́�c�����9��T+Sl�b^�h����@�odhL�w��1�f�Df��D�[g�ר� q{�{�i�C�~��U7Zh,�/k"2Ɍf�>����*R���\�X�/H=2��)�;�!Nb��fG��	���b���*�/�o���֨����oԅ�3��pA��L�����v\�=���k�3�	S�g�B3�Y���q�{U���a�O���}^u�mt�f6uҤ��nd���:>� ��X�����Υ����<*��rE�D�}c#�=�c���X�@������Q~���y���A�v�ƹ��I�@�]-%s�O��&U�H��yR�"�6�%-�f��/���ţ�qF����M��l�ż����׏�sa˛C̃�M1,�����靥�l=��r�Є26o�R�F����
H�q<�)�r2���F��7J��!��U�屛���יzV"�abq��9�) �W��	�k����q�ܭ��`�����-���^�a�\���|���e�S����՟�Re��8T��,^�ю�]���H���H�>�Y!���0����g&����UBs���$����ґ�PH���j{�ѰQ���K��̱�°zN1Eqjz:���lJiH���9O1x��a�.�G5�blt��!d^	��Y8��,�m^]�a�DV�[��@����Iw-�����{�R��J-��I�Y;� l$�GZ��B\�fhtOچ�s/��Ń����Q�ϵO�D�2�d`��%0�(j��~����nع�}	����#�����6<���P�>�BuS��q�����^��Z���Z<�u�XnM.ö��N��:����@誜�6/�N��No)%'��Ʒ$����dHz'�i�L|v���ZQ���-��Jz��/��4s�9� ��(T���fV:��ah�s*��\$J̱떡uh4C@�փ��Ƣ���3��R�tO_��xF[���P����9�w�w8�Z�N^�J�z7�����y���D��k[��J�+�X��[,e�i�WO�sʱ����ͫ"gu't#�/�j�ιu �Wh�������to�y5�侺զS�ř&(��^���a)�>�<Bv��~��5�%p�L]artM���;����6U�%�|^��d��'���7Z��`I$�i�0�H?����p!p�gK�R{��;��[l��i���S
�� ���BX���<�%'��[��~��ӫ��9-t�{�]�%�}Bϻ�m�!M�����-)y����7W5�u��S\x[Iƅ��d7�l+���N���
��d$ƀ��#D-x;V�R�8D����-o�xAT҉�f��a�\���Y��q��Ef	���c�|L�8\<��N����o7S�ˠ�7w6 ���v��Qu� �S����
w��Z�;��7��i�a�������i2ݒ�,�C\F+�JWR�mؓQ>[��B��g��R�� w�`\��(���ޠ��p�.~i�u�'{Ƀ&
�h\���Ꭱ�H��|� �((ÑV��;�`ΎXެ���?���EQ�)ڞ�X��A��	����{����G��0�5�gy=��c�V �7]S�-������"���NBM+o"�Wc)�~��4''b�zu����y�k��%q5��,�ѫ����,����PiR��nѤ�Z�gp����ڶ~+|T�Mw���[�E�����xC�r2�o�R��`n���B�8�JY�c;7���J|�~��ŉ�+r���_�xH.��6��������vSm���:��+?�V��~�"cl?���r�0*�"Ӳ+��a-b�ɲ�]�k��`�u��8�g�yf6K~�a���&Hrۂ�-��A�6�)�A%!_Nb��J䝃8I�yGn�Oy�I����P겧���-������G�C�yϿ�f��R��z�fjEሁ�e5��;��i����J@rm��j���M�g��ڪ���ٮ?����jE��&uY��X��_Kē� ��^!v!|�@�f�����n��s3�w�A_��&Wl��L�:��a�%W=�h�O�l9-��,�xteb��6�W@���f�rM�똸�=
��]AɆ��('��ૅ�T�B٭�1�O@w!�xi}����lU��,+_E�d>��W��Y֯Ik�f�~}`f�K�w'�� �)�1���v�����l���Um���]��ʄ�G~^��ӥpHBp\��X$�6�������.�-;��F�-�=Dd7.��d��Pn�ap+Q0��U6�rV�Y�4 �F�(���2fƜ�G��Z�	�H�O���ܒ�oP)^�	�����Z�q�$�}��݁���j;�1�����[�>/*�tA�T��!��>�b�#s&���>`0I�xO�A��8��	��mr���/U]��+�~��M�
}�<������MS�,v�v�&��jn
��ɍ�gzw^���@ҸԀ+�܏��W�2Gn��`�l ��+�@%��E�`��1��� P�Zcu�A�]2�46�P���Yu�ڍ�� ����Ɂ�i�(�w"�]/��g<�"�:�n�8����t���2^�,��{|T�� �)���K��c���V]y:�R{�օ^3Ϙ��.�ܾ8�D���+-�Xռ�
?��S��z\�'v�IpT~l��N��WO5�ҝ���Ӡyҍ�ʣ�~�����x������\ֆh���.2���~���]Ȩ-�����&yk�dSłp����ÄQ�E"����:ȗ���5S*{�����	u��/^dn@Of�"$��m$Aa�'�	נ�����"#t�"����If�O����-;1$��	�Zm<�,�	�8��_6���랞ܒ���}�x#08�a3�����̰N�p(svFGHo m�
)�ݿ�|�� Ap��af����-�s�1^Z��*���]-���3�&�}%�;ۂ��N=f��^X�w؆@+)�Є��V%W��Lhz^��\C}�,:b�����r�r��\qao� Y>x��>jMm��V�
O�0�n�`����tE��|;gONڎ����)���J���K#��-)M�#��]�B�|����sB�Je@���*�%Xt�5`�Q�p:��խ��5���2�z���e�ð�t��J#�9�Ƿ"���S�A{@-b	�����GMF��|�T����� ��6����៾�:����LP�MT��cV=���E��(��T��;���̨>L4�'�+)?�wD����FR�2�iXx z|1Hg���
tIIG������*��󜸐F�t~�����l�e���a��	���V��BB2��/