��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��5K�z��!��[��S}Σ{$Gx^����c��Ʊ�U�I��h��T�(6k%a��S�o���MW�>��:�m��]i�t���a���שBT��M���7+�
=���CmT�vъ��  ��?Ta�C�S��9����3�E���rq|K�>���.��|4���CR���UUaYQE敆�ft�P��W0	��(0�޾��Ac�� [jC�f9	�#����T�ݩk��BKoR"g|�lN���RB|�mr~m��j�Zo&�r��C�+K%u�"��V�K[�7 1��m������dx��s"y�[Љe��<x_8k,�=�# �!GJD�]7���t?���c1�ċ��U�X���,�xL�.
��o���1R��Aݧ�e��:wey>ה��H��!*��h,c�2��LS�L�fǢ֮��2)��d��:��|	dJ��U���eڝ�
5�yϳ]$�J�Oq�Y�l���V;�2�/ŀe*�Fs�^�=�Es�tG�f���B@c�b֏�M ��p��G.��#�W�;vhO`"xSZv*oA���ԡgD.&���D�_"���"y��qX2��@f��J:MY�!c��)��Į����a��q5)�S[�~v�,����(p·�$�޸m!G�@���$D�#a�·rrp�v����S��It�l]�LAX�y�dN��]8i�p���'�D�:XZ�7T9�6_Y���b��XC���4�Z�NU�������Yߩ�1^�톯���.�[g
��8p���,��f��B섯��S���W�� �l%7�S p`���O�x6����8K9}��Xzѝ��O��@�,�+Fn
�?���C���e�،�.'��#L���#��'k�&!/�s.��s��z,��.0�5��W$�ܓc��Y�i�ý��~t�lm����S��V��%��;� �����ɦl���h4���+K�,P�Y�A&���h��T"���WxV�#�2mj]4&�Z$W��x�{�n�>Ww]�l�j��y�h&�Z1}�)ZSc��Tx2��&B睃���g��
H��[��Q~��{ F��ZMi,&ò$����Lm�Y�+V�ĸ=A2��0� �c�7;�� ���R$ip�A�
{p2�B:��h��]�}���S(-����#<�k�ݦ�����p�P��I�h+�V��њ�?��8�x��)5��z�c�lY��i�`�M�e
�	;��F�jK�<	��_hӧc�X�BC��E>ݰǃ��ʣ���y����la��c}F�q�3�L��23s�~�T���fC�X�Ϟ��k! ��*�ʷ�H'`�i���E%mv�������̺�9�f85`}���bI\�,�@������|�L��}�V05�@'S֤nEu�,�\*c���Q=��3����Ĥ%fG�	��x�ְ���?��~q3�>�8${ �)I�6