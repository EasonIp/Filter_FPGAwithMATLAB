��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ��S��#f;�E&�o��X-��MQ���a�1�̧�^�"��0GO����IS�#8Q���+�%��i�︡���1�ڞ�<}g?�֨����1p�u?�%��ؼX}B@��{)�z���Az;S0r�V6�fi��&�ypó#}�!f��p��/�*x�wye�}�6C2��V���d<���\.��V���OA���l4�?�pڅs��n��I�=iΎ��P���v�aBS|�iw"K�
�d�x]��HFe�<�L�xf�oFo�)Z�*�k|�a���i�y�t{�i�[���g'��BL��|I5��=8��]���F/V�Y�|�l1�Cb?�~��[�QC��kΒ~�[J@��Ld��� �q�,�݄}噵�V;����3�FbJ����L�'�O;�I���I7@�E�~|'���8ZՄb[8�d�_�����Q!�^���_tf����̽I�����M��04�Ь,�R�W�ǯZ!��f	�t��c9�@W�{���-��|yt���N�F�Ӣ�����3A��>)�(�kj�D�?&���h�adO�}�߱;�Hz�"x�ďZ09���ѸB[w�\����*�������5<��4h�-Cw; {-T�.�	���d��}��AE6'"4���2N��������E� �F]a� ;�u$�aݶt������ɻ������`qRC�H�GF�f��>ă��js��n�� �tzէݛ�n?�jh���W��Px��]���aTO	�;H{��1
#�_�a��Fsu�԰t�%��5�ѱRS����v���8���wqfƍ~�!˸�i&��fI�8���Jα M�'~��L^�P�����#�����m�?{����K���oe�iv;���=�7G'bL���;�>��P19��:�vh���?KI�{��������,��_8,2��4`�b}/�˲u��>�������N"�HGµ�r�B㺴�ߢ0B㲙��/="��s�R8��)�KD�A�a�����rx�	k���AiO���]����5� ��j���^�}z���;ϫNY��zx8����[]S��F�(w��c���%������#��s���=�4𬞝���F�m�x��	�d<P�q�����4-偰�2���x�=!̉K�"--�yւ��n����tB��֨+=�?��ZT?�ٷ�-�uџ�Q���|�t&��i�Z54p�/�����B/[���@y��仕k�rr���I}@s�'�9W��gE/zaߢ�n�rkՈ����EK�imU�<�"!�DN<8���`�h~����KɃZ�D=�WN�6d�?� ��SVM�'����7<��B�s��aƚ�-_}x�20-[�}������w������t~u���c��	�k�`g�x|�A�$ �Ux�5��]a �Yf����u9�ܒ��a��� ֵ���+��C���Ê�B
���V��Gm��i�E�����v6����~�7Ӈ��xe��V�����o%^�<|�W��b`�t:�h%�[3S(�!
���k�+a�+���+8ZL���ͫ���M�+��Z`�F�YavǼO�T֏�p����K���5���z8�(8b<d*ʃ����a����$;,�x�HDz{�qW� �}> ��jn��gg.߰�u�a�YKA��VҶC�!b�U��/�qg������YЭ���-=�2�����K�l�Lk\��ea���M'�5��'����g��{L����Av&p1I	zL��_)j�s����c*�>�����w�;,���7'Ln�Q�:K|�߻�����xn��"F�.�3��R��55�wXGTzh[S ci��i$�B&R���kypJKL-�����1�}���h)d1�wa9�f�V_������W+M���Lh<�V���ĺD!��Y���J�7sr��xk�.Sl�6���DIKR����3W?v�&�þ{���������烃�l[����F�Ϫkkg/#�!&��������b�j�v�Ts�����]S�HV�2jZN�����B4S.4dJ��ё�6��Y���J.��Kc��eαfEӣq]C:��2���%�����q�T\˥v�Ɍ<=�5��G�;������$��jG�[�%[#6Y���=>�/t�%b�0�"
p�˹`7�M��D��w�{�,�϶(	,�̏o�4���'��ϲ���RYLl�����`"�TC�+�,%�"�tda�{�ؖ$��<	L�YY�B�a���z?B�z����o��)C��Q�V/#�%������_�U)�yiWC�}�C"��b�W�Hrũ�˟��~Z���,R�Ƕ�@��5Dd9�
�wܼ��qE��������H���m밆�����jn6*8$>t����A�a����� ��U��T�<*�Ѽ'
E�ó}]�[K�6 (&�8Hy�8��C���<jk[������5� �[�H\jt��� ��p,�jQ�����6S	��^�(:D`d��r�J�w#y��E�ö�Q���C�b�?0�kڎ�D;�&�a�G}�t���%��>4��[z������F� I�%���p�q�d��+�_p%��& ;�]�)����#1�'�걜�p���p�ҙ���D3Ϗ~L&�]���+*o,C�)d� `�o��w��g+�s&�H�[�1�0��_�I�q]�(�C<���:���Lա�Ӯ�����2k�����W����8�B[1U�e�"'�s�C<�HIu�fD3 1�؟�5;=�3-M��a�pA�*Kڗ^�jd�y5瀦Ɯ�,��L�ҹ��Y� !wY��^{�U��GT㶁�.����
' ݊�Y�}�6tB#k����o��3���L��{���U�_g��N��EhqSť�@Y�=�M�5[��Xr�N��RQ�����ɶ"��q�1�-Z)i��4�cD&�>]���о	�ɶT�XG��x��|�l'"�i�0�{�#E�g�x�b�l"�R�lƷ�;PVTv�M_$ ����%gN� ��_����	7(?�'0h�J+�{�|�-�2
w���/��-pU��i!aa��p��iOis��(�+�y�x�����d�5�?�R@�#�;ק��&����v���*�`�����^��^y�b'���ܷ�Ѝ�������xM��6�g�fޖ
�̋"�Hws�)���tl}��9]X�:�E��KV���w��e\sp�������g0)�`��Ґ��9�����_NJg����f|���n���8;"^�u7��������1����=��@,ʒC�ۢ�${[�WN�u1��O�$H�?��k�g�6�/�C)b�7�����Ԭq��ըΧ��j+}����*��PRe	�	�$��s�(�c��� ��W-�|.ҡ"H��2JW��~DR����O�1�(�[<��j�i�����Ȼ��<���G���/�q����n������?�H����;��9�C*���G���)߉�d(�������HH���D/�����ƹ��_���ٖBxk'V���bK�He������n�઒�d����$a�?��J�����
	~S��yH4'⁩\\V���g�G�DZX~(ރ���ׅy��&~�Q���T��K���I����R%�է��y��q�r;��C�Fn����-N;ʧ�3@��$�Ѯ�l*�Ͳ�ҝ��A�`F�x���4�e�{��}z^�m���1h�~~�3���:���H`����V�$�8�F��u�c�qK���f~n�⬄�"o)�\ĳ�˄�+�Ux!�h|�%�f��E�B^E\���ňbX>N���[\�j�

�lxQ]���-f�TcTra�iK^s8t�酓.C+�M!nPɲ	t;�3����΍/4nNW�L�:�CZO1o����pHi�ݛ�LPQ�sk��Ɂ���"9����@�������EO$	`����Od�%��iss�=L���R��S��<�d�U�,7�;��[G'B�^e\\�a���B�o����ʮ"��n�X��,�z�`�å�f��M�H���(z���Lg�g��#���
z|UQNH&q�j��y�P7�6r�عGt�7	9>vJ��X���e��
n0L����g�%�%(��h�yEl��a�{�lK��
,јH�JUq�L�!k���Lc�	8zHo�v5l�ZH̉>��@(��t\<���i~��c�O�6��e�=G��-� �ԩ��H/�jq
q�#䣈�<� ~�����<ͨ�jC���|P{jן�BH ^C�/���ԦNȭV9��#-�����pc�جǬ�T��Rl��#�[��A��^WBH7�Ю7�
hY҆�̞KՌ��|[Vd�Ɔg�<��X=��D������u��S�jݮ1����6�]��UF}�.q�MԒ>̙8����{���cÉS+i��!1��ݪ���3���Ɔ�cZ�~o�@``��
�:����s���6Ѓ����\�������3:�DUC��2|�u���%����I�r���Spk2��H8��2e��/�?A�7ڊ�4`�١I�`v����KN��ڳ�Ε��[�M?�|�_0ry�'�b���i���q��+�<��	�x<-�@��<�۞8rL��8H�k>��~	e�x��U��c��55�{B����7�f���KLF��X,��SQ�;�P�O)h�9�Ѹ��ZJaK|�l�(`���	u���!�t��/�L��zܒX40��o�#�㠻A�t�A˳��]Μq.?��)��ɘ�28$�M߆܊�Y�Nu����D��I���7��r�����}rO��r����e��\Os�Eb��F���X�]��������?
���\�Dп���0�ƿ�*A�gJf�=f��]�rl��]��W��/��kK͛�HG�\i$�p��9�v�;�z�����O[�o�g��=N"|.����4�ML]H;���\��&���Q�ڀ^�|�j�LyH �q��X+����p�^��a�A�o��k��n�k�g�.��_����xŃU��cۣ��:�+�L_��٤t@��Y�{>o9j�a?�cn.�O��ʼ���͠3U*��"�ܢ���B����x�P:�G�r�	4/����ƃ���n�+�|���Q�P'�D�A��v�?|a�-t朢#}Q�<��ք����ܛvj��/�@�F_�-�Y	L��N@�p�-#�i�T���)!Q1��E>����MM�_?u��ߨ�{�[9x�x��[���S7��uU�o�-�%�>���8䏒����ȴ1�X�Ҵ����P�h�a������}� �!����f�pawM�g�h՛��AY dv���[0��xMa�l~a�!��]J�k٬ ���ta��+���_k���ZI�?�=𸃲�!��ȜX�=r(�|O5ԘE��ڃտ��7�S�� a@?�qYF��t����Q��_I[�v��^���Ey�g����Db�Q�"V5N���S&�:�����Fk��b���X@�3�E��=�]D�"��d����028�Z�Ĩ�E@@�YB��'��rK�ò�mci��'��\W�k�Q
�
��g�e$�ݞF Nv��C�&���8�uQ{8*�{�D0Ȟ)���\���!���Tƫ�B���.��4�)Ԉ��nM�veq��y��v��ܩ"���-��o��Хo�lى������M#?;C�q:"�j�l�ח�ˤ�6J�t�Ē�ϼ7+�:�W�ST/VM!��)sW�b�*}�$^i��d���/��Q�a�ش`$�{\�0�K9o"B��aKtw���Kl��_Lb,W�S�l���'ͳ�^#>�1*JwM��>�
�b!�p"�TS&�q֛��W&��u(��D�:��Uxh<]]~�X����� �%�@h2}�}���i֌�m#�L��
��lzU%�
��!�W�V�~ �\ٻ������3�`������2#� ���𾙶���}l�~���t��$-A�:������i5C�!�ȡpn�szH7��O1���Hb!��/H)BW��~nD��i�!Lo�~3��'S�{A0/%+��Y�L�;>b����4�y4d�Z�Y>����}"cb9�e�s�53ش�j�͹���k�:%�c�ؿ9wk�����sb�8~Jvop�w��>֬�kp,����H
�}��MX�A@䩟�Jh���:����I�2���QKm����x�`ˣm�J���J��M�?n�gn-�xǌ����EދO�K��\��nOVqZ�yg<���*� �2�z%�_�S��*��x���GS�F�Ց����Y�x��t����9�����7N���qzrJ+�W�GC���n��C������J3���23}C�G�X�6Y�Rݝ�/n�מ�I����F�^�d�{p�G�C �lnqB������D%��C�CfT'��SH�״�����0�=Lܗ�ӯ4T�*��G�(���?�0�3��)?�E\�A�~%O#���G���:6�K|i��8�	�#@(�Uz�v䧭Q���B;�<�j�ђ��+s�cO��}�[0�����Ѳꆜ�SWL��0Iu��=���%޲P_�Wث�����qC�������m��1��a.���&�L��O��jZ��O��jzhm��&ku�S������RLEO�W�R Q�pQ%�Q���Cb�#2��ف���[6�5)�w��A�|�y����nӲ^�8��-���w(�}�_�� f�I1�,� ��"��
��2� H*��<섦�)�89������x˧~�D������'��4�Ӻp>�Y�k9��9*���/m�XW���JAշ:qx��7ԏ�.��*(�0���kE���v%� c�|`ܭ;��{'�7�oz�e�ֵ.�h��}E?j��!��l$��h@��ϐ���k�*�=P�t%��@����������L[��đ>�d��6��Q����&�.��XK����S�6��eډ��	�p|�%[^����?��A&�\�)'io��������)�K1o���������Ij����P��}H��H�"(ͧ���?��v�	�v1e���}&���԰�-o��<�����졡�Y�G? �����/�� ��Vތ��L�ߨ�F�`�e/L5p����FŚڻW�k+>�#��;: ���r=P�ѳ堈�l����:ﲞO,�DR�>	�]�q^��2��h���F���8�]K�ۻ�[1 �΋�oi��0}�5���9�{��|s=�}���;z� sA̦^B"[-zM��s��{o+�z��4i^c���.P��G��Ჲ���i�ii��zD�R8�6�<~d��*��K�sq 	���:H"�.2�sH_��m��{~���k#�Rq�q�����[��1�?���e�Ф���fԼ��A��l@��~�E���n]�e[��M�hIs�m��ƥ�K���f9�x|t����]���
 �X6��E�\��S���DR~���!n�y9����zؗ���\I8��n�VcH���`o�b�!�9>2�}� K=b��Z�h���C ��ۓ��L�&���I�h�� �y��+-�(�<�Zǣ1sb��0�)����ea��d ����Ơ��R�Ǖ���yY��{�	��O}��eb�:��H�a�a�����~�ߍ�;���dQH���mh�g����mBe�P&y�����M���G�3������7��ro��Q~�aI�ޢy��6#�$N��&������m���]�<���s�}k�zJg����Rk[��0xS6{x��څ�%JM9����Y�}L49Պ�Y��SZ�W�k߻�����*{ƽ;2�_ĘCdS����R'T�M��_�UN?`����z1��a�	�,�iE։<�&TV�D"U�|~s�UZ��`�Т�.U5박��	@�����}��QCK�C]{wOz��-ZL��LW����Ň��#
b���TS�h��X0��5�-�2"�%�v��������?8���af�+D��>������1̑�R�,�GWv��v��&>Gwz5#վQ [�Zx�M^�&���������q��:gڸ���(Y���0|M�[�-"n�N�����2����ٔ�����S���F���n��T�F#�0�m��~�>�?"(���}�(�F�Kc[�sH"�+U�B=����P�7m0�HXK߬D�'bz��Ob7U�̧��	�<m�n��S�H[$D�n� ���֥���G� M���%�q�RY�~�,#Ueէ�$�A�m���) 8�g�RI#�h�������D�ג��C9ʫ��,[μ�Ǝ��P��B��QKm���rk��Q����}��۲T��B�(�6�h�p�=�~�5,2/�o&p�!�_�������+7Z3_��e�5�c�ZoM>����ex�������e3����7��Sm%���0������Q�E�3�b�`F�����BkG�F/�>�F%�=!4�\�M:��:��g����j�{�V�J�9]�	M�4ّ��zN#Dj8e�����̃@�ZB��34rH�7�?�+/#��j��֠���P���/*�.�Fa�\��6%�^�<W#����m�HTkl�u���~aj޳kN�P���Aw������,p�@"��?1f�J�����M^��R�7��m��Ɵ�X�9ݕ�E���sa��!�#!Nk^�@+�}�C�� ���:$zh��W��9�{?�?�IR*L��o��?*R����b*�i7.-�����'�xW�!4W�y)�l�����قԱ�)�9���J��'��շ ��j���朞�����/k���Wśc��֬'ڪ#�r�^Uk);�`v�lNwdB��e��e0)�IQ*~<�d7�*o&:Š�l!�-;X������e�� ��^���8O�$��:6 �|�o�6�Z�`Ƴ����i�[r�,l��F`^wt�şƳ����]�#�0{�Q7E��=,���հ���1)�o��2�/n�U�1�c�Ds1j������2�	���Ɯ��/(��IQy���bF�YX�o7����Fn��5�oC��꼲z���!����B��^D��)�����*�1}H~�|�����@�Q�s"�m<B׋l���1����u�]j�Z���wiYa�����M�^����Z{IF�	6��%�,���L��� ��O��i�:.�CUx`e:
����+�0��~�xol��pq_�
�������P*��ή�*M�jG���R0
���-#�=�'H����������<��y��L&������Zzj�����t�dxXo�/�W���
��yC�|
��G��+���>�x���|�j=;Fl��:��ז�	�E�ݗ5cU� sF��Qmz|�Ү'�'�)_���P���L,�/i!��<~3o��˼�~����>$�E�1�ö��I؝�t}9O�L�u�F�J�b!�O��A���蠹�a+� �B���ã��˗H�V�Rּ5�����$'�P���`,�d���*�)&2tlOg�Z�×�`�8)h$��c�:�w�-�t\����}#� ZP"FGY?���j�g��N-ɨ�q��}0���b��f[	\ �6�7�*�1V�
�ֵw����Z���>��Dp����l��:�D\���g�ue$u�i������KDR9G8�#��r�P���.Ma��lDlb�,+n�m�{�{�_��
�K�C��J������Y��6ܐ����K�S���Es�GU;� �$�w�-�(�λ��5ZH�h;���=O��'��C���@�6Q>���@�:(���C,p�űu':���K�1�q�{Uv�Io�t�	���� ����ʍ�o9�����'WN>�Pgw�8UD� ��F=����޷�K�cY� ک�a��'l���QW}?j5�z� �P�ey1��l��w�"6��#���I��3�x��쉜��T|?(m�T4֋��V�C�G�H���r7s�/�%մ�?4�b�B9�r��0Ivv+G��],x�W3��ԃ�K�UW �'��6e�-� ��h�E��_�:HJ��̿�y@��7y��$B���-�i�������!2 �87q#�Xz�2�K����N�q�@�E0�r����p5�qat�b^n-��F!R$2��m͋ղ����X}/�m	I_lKP�]Q���n��LD��V�/��G�D�npv<��~�RLN�{�C��$�l#�赅������\A��5���:��h�J�N���H��E��J�b����F*d~<eVei���67��^麕��P�L?�X~+��l��+\��|��P�f�b�Ҡ�b�+����BH/��:��%vI��aC��> wU��q@Kh�V髸�J��8�v ��_,�>DD�����wK�R
b�p��"�2��g��eD����)�}[T�'����qY,��k�5�A��|��tA��"��ϲ��f�^^d�waO�>BrO�}|��'fg��z�G�r� �{���X���TD�$8�p��S,	l�j��bgd�����4x�5��¢��xxŐp�\��� ��?�˯�e9HO]X��C��x$!��fF��t�Vg�"	������]��1�l�l$7 ��b�9�"A��nA�J���o��bX�ȋu����)yxߧ�m����%׀ۀo'��R�}@�?+��v�h7��A�R4���B}8��Y�*�����@/~�U �ڜ��N*i�3��宓����N���k��a���4
X�k�����w��Y����ܽ����ϗ(��5Ӑ/��@G ���i��or���A���0�Դ)-*���e��(7ʹ-$��͞8�J��B�8q����j�9TjI'����V�y}��tfv\EW����݀B�M�G���{�;;�$�[K�O,z��jDI
u���|�?]��WV���۠"����̋�]����ļr/ݒ��G��	C"�cZ�˜FV�H,=���
��kIrVj�g�G^:-I�#�����}g"<R� ��$q��Ȳ�Mm,=K���C}["��j�� �j�V�n��b����5-�;޶