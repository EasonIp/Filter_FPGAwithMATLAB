��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$��-�z}��w�˩�R��E�o�ox �L���47��7ӊ��h�$v�|F�c0���������?T4��ѿ���f�������d]�:�3����4DV�LN,�,,s�0����<�]�j|"f�r��j��k�5ala�t���c%fA�.���d����-�� �@��T|�<#���ս,��Va�xj4-E�^xRj��J��hG{�3Yh0B{��2":I�����ʞ�
5�+�w��g"���mc���<�V\�*��" ��s�I��읱��	3+��/D=�e�� �V C����*8P������JacORϙ���D�a�8���/>��=���
� ��Jrn���Di_�k��+B�٪����|�jc�����x(%���U���6q�?�L��rV"a��l�褄���"(�ã��S��/z���d\F����{3�^-R�<��dQ_1W�^�Y�J��sl3�^w��.��#��L�9J��0�l�z@�{�?>�re+�!	D�{ ��a�__Xn�>ו#9H>'�Q5�\��3���.�cm��f����
SK�M��#�yM���Ӑ	.��b4��p)�{�:2�c���9��=��ߌ�#ȸ������YTQ|����;�Z����t�e����ΊA��1��<����K*l(2׈!&rK"U�o'M.[[eG~w�=�=S���iC�\�5�2 ��)�
`L��Q�;S���~j�5��}�����W�	����� w���s�[��R��G7�_C�� ��k�WϬ4���G���������t�<��e��k)f���I�-�>ycl\e�n�{"�0�U%uJ��^��ɩS�T�Vd�}��|Y\�t۴�}�(��ZG�Σ�}�ڪ�Z�:���*�[g؎]���
�@���+�¸��&���n�|��o�����*����ȨU�6��k�4e�=쫴��G�+��f��BJeO�4{�Xr�1���~�S,�"�	�Y���M����>��w\+ <n���V�I�m^�6�#��>��	�/e�Zd�C�ݲ���a�v2�|Q���k��B�V�㍇9+�^��J�b���Drp@*��=�]bV�.��2#�m��1Ⱥ�<�����Gz����9����wJ�.���O�"f��,t��a}�έN�n/W���;j	J���_�	� R3�k���D��k��P���&�Oeb��m��u�kE�J�$/���:0c�K3#~#oZ��p�@�7<Q�9��뚮���d0��#hQ~@�0F63G%hC�E���"��omx����9�I��̓�S��~!C^��T�3�
K�-�A�~3��p6�".<)����,_��v�ov-[uрd$	��U;�eu�aU���x*���3[����%h���^̹�3's��6���X|��X��IX�F��  v�@R>_zRv?�Z��C�o.��[h"��+�|����߬�����*+�C��Ta_��}�Ĭ>�����d�s���QoQ�ba1��&��L���8K ��H���p�%OB�s�ɘ��/a�$�����̴�I��=�������c"G���Xa0f�@�<UT
�Tý)�'�%nGI���{|C�Ʈ�U�>_��0�����˼�
&������*A-�`C�0�^�;E�1�Ѹϼ����J"Ro�2������z�S��2lg?��1L����f�:-!<�t�ծ�ԍ���ih*��w���o ��a���ț>H�o� 
���J܄-BQ_�_����^�.@�Ax�ט�ژ��B&��l3��:#ق���(����r�o�r٩CO����/XcT}�vL�Jp9˰���󭏳��Α	��w>	{ܘ��اLޠh�u�3�������XB���2@s�ǖ	N��/��5��)ω�>��]~�M��ݜ�{sU�*{�v�Ϲ�s�>�>�v�}��B�^��8�Ƀ���st��ԛx3�	���DxXRI�tao�>��oI�c�o(#�Гq]\�XI�މ��]��Gރ6%m�qk���yL��x��)h^�C��S�ă���a�ƕ*o���e�Nqs8��G��X|W�k�VA��x�#�^2��t�
+�6��>�f�l7??[=rc�3�����41��j}��������}?��,eŐ���(�L�{�B��v/PQ_o�B <_�9Ӏ�q$V^�����;uT9��QI|��^)���a���ѩ�n��C��<��Kx!o�p�t~ >IqUV�O�Bķ
�%x�گ0ȗtt�jR��%�X�c�������l����4��?#�;��T<��A��R��ۤc�" �����(x��vvE+��5�&t��<��.9�)��чî���qwT	̶I��4�T��?�0�����d�.,mg�����u��	�S�>��u[?�=źfq��Esj�E�,�a-F�N8k��?�_?���� j�1��kf��E%W��ڊ�L�
H���	Gn�^���R�1�0�A����m�C� WV���k5���x�|�̄yD�`�:b�;^� O��g,N"?�n�B��~�a�g�K�I�����F���=�V����b�� MUwVG}V3U�f�oW����! Hὄ!7_��f:E�ԧ8�Lw�4�_	mb֕g:�AS~�\(��p�L�E�[�Z���ph����F��g�<�^u:qs�%�S�x�,A�x( �݁���������̜�cƴ��e�����aF����HaM���4�6q-�N��n^���_ʟ�pγ�.��\�_WY4a����q�L(����V��a���L����0W��d�(�{i7
߱��.�7�^�\�d~iV�}�uu�~��O�-�F~&���I�8����es��n1x������K�/���9�8���/p�o����'��b��!!c]hbfO��i�7C�S�*�b|�6�L~��ۭ.� �
����>�����3@W(¶,kC��F]L B���e*�@@\�6�W�e��re�����dhy�DԘ[q���9і�"��0͘@����W>\�9|��e��� �G��i*T�W��kJ�,���y�9͝u�r��&0��2�>Q�Ae�E�g�Tظ)�\x���?K�}kq�a�Xi(��	���%��d�Wl��(ֲ8U�r���V���Ok���Jߏ��Ibv^B�C�:#���U	oPh::[�{�;�ԁ(nF�1��dh��ΧD��ڧ�Y�]h!wJ�-�#R��	���N*�f��=n�Q����d�Q�!��-P�(�O]e��M2�m�1
d<�<+�9���֏#hil����� �=�&J�Wc�'�d������W,�-tuӞ��Se����_��+]1�_���u� )�Υ�i�X�^o�
��|�u�_���^�:o�Ɖ,�?<`��V��Y��U��\��p�r:�8���,<�'�ݏ0�q��AL��|���}��%�
e����;���OD3)[��R�3����ڕ���LO�`듘�hޙ=��q��|�$0F��8�s�o��4c�}�����_

#�0L!��W�?-*����C�NM�P����U�8NC�k�n�I�egI�qx�An��O9�����|���2�gK)%���{�� �n�p�$5�V�pmƳwz�q`��^����T쇎x��f�(W7�	&���z4ó8ԆCԴ�QB�Ek������!�"=��ϋ/K�#�yVG��!��q�r�UW�jH�!��2�?E�?"��X�6|�^j�Ťm�3�݂k�	�)LzQ�:Kf��s����\��8]�,Q����D�',���Q�q���unk��pIg�~�t�WE����ݬW0�m�u@��ҍ���IZ�Y�[l�s�����JfRσ$�vt�)��`M#`��,S`w��
�2�4��Ӄ�vA>�#'�D�d}�n�g;I��Gn%lrS��y*AaD����F�Vt��^���C��ƹ����m��S����ß	���Ճ��~�%�Ѣ��J�۸e�nkr<����-@���l�j)����hm�BM�ɝ�`8g�fC_v;e���7�ޓJL�`T�@��m�ߥ���׍��>�1^`�%�����	�ߏ"sI߯��PR�y,`F��'�P��ɾU/�a�ЭvD�H������w�Ws%D��b��x<YF�i�G�5�,�Ƽڤs�Q۵ �H�A_O� IB��%ܩ	����@�`��!n쎙����ǃ?��:��Zc�i}%�v�5��
Pj��]~���� �`4����I}��S ��iӆx�.�$�Dw˞dQR�Rϼƍ�N$���*1�X�o;���T��,8�cWǸ	<�Q]�P�?#�!�B'h4���PA_Z�L�l�J�e(��	#����"���8�Jj.��  ���PYil ���z$_�V�ӟ#	�������|%q�[BşhU��]�9�@���k
uv�^Z͸�M;/0P*�%2e��6�䚫���]ɹtw�x�B9��w�J�]n���ي4�Ok�._ܗ���W��/��wEe����t���C�J[%>�O5�8�.� �%�?ex��U˖�����l �zu�/�l�V^�T �|��7��]��W�Լ��싢$<o���DK�w�mj�s�x"!8;�#�_�� ��P桰��� x!��3�F�Hީ2�Τ^}���w+�c;P��FZ#�T��KfM�<�u�&��{�g�l�U�w�q���Ac[bz�4���eT�,�g����n7'�nAd�
�h�<�N|��0�b��ĘK�C@����&RbH�$�&�h�|]R��)�6�r�?�jh�AXI8}:1�]%rP��YL�9��%}�o���?�x��S�J� �\�M� �ԫ��=�2��A�+�\=���v>���8t��r&Ǽ�=�!��I��Rt���ѵ4%���\=%��甧�UB�j:��V���P�I��)�k����6��6t���o�TL������~x��"�k�3>�?/�����2�4�+���2t���z��O%��Ai�sc��B�L�(v1U�lHg_�JLğ�N�=��l�鸒����8��Y��wz�$�x���g~����Lf���;Ńܛ�RԘ����NQt"N"Ę4L�|�X>��U�2R�	�Ѩq=K��8i�퓪��4xek"lyJ����yl~�R���R Q4�b���!���o�=�CP	�.dS)'}����|p��9S!�˹(�f��Z`m�@º,��)�����g^t7?�pl���|�d�kH?q�ݲwS�?��_􊈫Q�>A�/�MQ� 3�d*�V�",��/���1f�\G�*z���\�����<�Y�KW�Hi�aEL��X9�WO������c�)���}��J}�¹�G[J�_@��m�9���H�]U-ԛ��Hx���p����W�ռI�\�ƧsA�� �Â;t��	~�Qʤ�]���r.�S��,����8r"�R͚��D��R�iyglo�hp�p��g*��v���giG荬�W�F�-.�lm���^nf�2�Or�g-�Ƭ d�����=��;8��-�祓��G�p�d9n��>��xG�Ao��6wG���ٲ6�P�g�,;�������n0׷�;oɯ�h�WYG�X��E՘�Q�Tn�Y�+-J�t��:6�v.c	4�R�^�|j,B�������5�g"�z�+��H
�6��y�i�qS���-$:*��|7C��Q�K[.(�M��^K��Uw�;����j*zip5$���H��Cκ�5�[�S��|ve)�P�Q6��LFr�>�7�ʳ�q�K�&���D�5^����暶�=��&�9?~�P~�JUYB	Z��A�}E��������vAq�C��$�S��i�L�v��U�`����(c,VD��� �Té��������%`H�k�?�Z�����L���=#�5�ϫ�����
��Q1"�
� � &���*A)5�cM���jx&������s8;%��?.�t�k�ztT̝���G�r���[��mt�y�h�4�a~�F���&5�����Y� �AΫ�Q���K9;EX�s8{�u/�M<V��)ƾ�4�Lo��`��-��%��j��{��;B��ܠ��O���y�P:��^����$�$�C�F���7�8:���������-.@�s�4�>�0��oO�hs=-��R�,��g�.�����s��P*����1�����UQ���hn+�LM���A�&���v]�p����!��Y�E������F�z�b]��>�&�|k�KJ/�^��\�* �&���s�y��:�	9����'�O8i����������Ss�u�4��ҵ8D���R�X��?�'�Ƈ /wG�a���8�&�"x)��G�&�I��n���R{�Gql��?q��=�W`��MX��W��BA3�T����b��Vѡ��R�
Ro�T�f���
y'%hD�'2�[��%_Q�f�s-'�aH�y��.U������?x���)�n�!���a�s�����dŝ;�i�Q�W\i����Dg�h[y����^q>�S�F�Qk�5�U�L��Z_{�t�e�g�u���?9�!��w��(��+}
�Ơh������¼�"Ns���i�Ԩ"z������J�u;�=G�rt�9']�Ζ~�GU&�~���tXN-(���KO� �X��X'^OK���ͯG|i��W@��NA.��WWxQ4D���Ir=���|4s=P�z�uQPa�6>͘��X���$G��9R���5��߼s$��nz��J�.����߶��8?Nќ��������a5E:ҡR�$wY��H.��]����מ�0Ю�����7�XD���j1�b��$�,����W�r�X~jt\:{;���m�������`z�)rK�Gv�������z���.5C_)�]��bi�����W�5$ݛ�̻�*��UtG
R��k޾~��2��@;��d*#���J���`�.�:id��T��)����Cs3p����T���k�1�,�����;��q� %��}Mrb��҇s4�q

�~Ʋ�랑Ɍ0ų~~*�6$�k��9�{�Cv�ŏ�At�䎛t�'�GӞg��� �@������]|C�aF�j"Ŷ_����ݸ������U�U���"���vy!u)uO�&1���k�y�隹b���b���ր���ڝ��i8�N�g�nW~��.(�<��E�D�ۑ��`���Z�HB��e����À�� ��R�m��ԫ��?��6u���s�V��;�O%��e�A�r���d{1|(+�V@�9:�#%}Ӣ�7ܠ{(�Ƞxn�(��Iz9�7$�[���Qׁ���px��Zs<U3F7;�{{�3},Vٛ��⌜M��
D	r\�c���.<Z�:;Þ}cYhǱ�S��T���#�����w�`�y���=�jT𝩠�v;i��C��̸�F�iOͅ�2�s��nY�O��X i�6�k��P�cH��v]��9/���%���a�>#�S������r��懶X��� ���$>����é��L�+�����*NO�n�r y7�H�":�Ƽ�f��@�WF�u%�e���]����譮U8(�)K�����) �x�n�l����g� d�9g�u�T('����t4��u ���ui�~�7t�=�Y��	�G�o;5�F»�^Xh�|~�S��e@xaǬ�J���u?G�jr�Ւ�������۬O�-o�R�]\�N]��.�.H�ؿJ�����9�CI�^�`&�meZ�:}8���B"��?wί�J� jg�bu���4-wW"^0�4�l��o��BZ�>�1�ioF��WW��%���m����	s/t��\����m�j	@���5��ݸ,���Z����to�|^o�C��"����m��RH,���16i� pUt�;�<�!ϥ�ݘ���e�t�J|�"x�/;]7�e�$Քo�"�E_P�}&Q���F|a�#��ޱ��"m0�v*��M�ٿfB��̳QKF�d�j8����׋�#��`T�����Z��ns�w��3ڄ@
s}.��A�H�=<���f�EeϠ�3�2n|�U�(��nO�y�)���@th�?Ю������~��.3p?U��2n��H[�Xkw |�cG{�p�S����lO0[N��v���Y5���3p#)�[��Y��r��|̤���T���b���>�cp�Bi�{��;ax7v��0�V����>�Ǐs��֧|�r94$��o��]搄�7�`�/E]�$՚�!�)W����.č�)� �>Xv�~�z`�
��������0M����y;�4���|����0�y`�҄v���p�Z���EE��=���x���!H�4-;���*�������P!�R^H	J�,ݘ�f�k��L��h�;5,:E�Pǐ�VT�Ũ�=L�YK��\��c1�Hq�
O1�@R,�ﯭ����X��=��h�A�K�M?�%����肕��cfC��
����۴�
ft�=��E����
ƔafUZ'f��WiEo�`Q���t ����tJ��ފ��q2�]�WMW��|7}���Ir���z
"
>�}�ސ3^�.cR�%��O#�T�l$��#������+�M��Х���F�Xi�X�/�r��]���;$�,"���~��{�8��s�X"�Ccnh}�X�r�o!s�_�,E��*�]���uq�ϙsԷt&l�+��P��#P�&���f[���k���|�M/���7T$0r����cC����T�-�f�
����wXa(9r���to/��8��� Q�}�5L����n� ���u��0g��8���/);��^�$;��`�f���,T�r@���Q o�H���+��׎o����Hv}!������24�W1�=$����������tL��P+������?I]۸��z~���I��������y�K�|��r]�UGцdb;$�L�6K���?�DS`�ty#�x!�¬F��Bߪ�;Ӷ6�h��F���{;>Y&T%���Ynh(��7��� П8 �Ɵ�&�ԫ�=�}���� ��^�Z݈'ҏ�JԷ��v�sa?�T�Z�f_5��02��ˏ�So��S�v��4�y|�M�Y�>I��&'�W����M)���`G�P.��tV������n���[`��I��"KN��?C��vsa�U�+��v#�������4�Z ~���,�[8�\�q#����� ��N��3y�[�H�
F;�����O�{���{mr^��jZ�n���x��¢�i�f���3����K��r�^0y��
c��|g&�4{\�j��{������@ڎ��S�`�}G`���1ùjM������mUi��J������1g��r�VyO{�L���J�������$\Ep޳1{5pґ��I�@�8���V" m�4�2��0H#�c&x����֪Z��_�3���g��^
]��S�}iQPg<�u/�����o�ߨ��ݒ����^l2o�z��ڝ�C���� �Q����-�v�̔D�\���MH�	�����W���B64d~�&��%���t������D�?���;��"DÓ��*Y��^����v��-\�܏K��l=�5�3��5�';�����
+2�ULw�@�M�`�ˆ�V�="�L�8Ϊ+L� �|�.�����+=سۯ�2ė�G_�i��i����<��vE��������O�`��ɱH����H���� [��;;��FF���ۇ�Y��.~�6���,ON2��|���.�p� ����-���/��a���`z����T���?){����y����������Щ��Ʉ��K�H�|���QЭ�pXxRn1j�5��e Q�:݄K�������c��x�w=���k����C-0�Rd�m��3K�������on����1";ߞ�7�
K����4�ņ�}	�}c{.�vX�^�v\�
 ��Ks�6$���b��f:� k���2o�&>B�X�l|"Uq��pj��+�X��	�)�Wc=��4�|� !^u�rU��ʆ[�vޤ<Z�y�d:t�M;O��􅽣�p�4��xLv���j�IY H����&����|�e���a�-�QR/�̍P�aV��A�mS�Mί(�9���t�x��t��&G`����	qT*6n=��
Md�S���-&��0]� `t�|�x;�q����vB����Ҋ	䟣���K�h��7`̛;��y�'a��7C�����.�Њ{�b!G,/T�0��]���ѹ�8-�1��;�ם�c|�h�W}5
5�_fu�I��^7��r�fY6ξ��l,9�'�:з�=I#�qmT4s�0!�9�j�޴ԭfH�,jCk{X�h�J�T�<�\��w����l� a�ʴ0�@Yo�~X'�ث6����cU��_cC>o�k��3M��4��}�>��AH ��"0�Ѯ�yO��ύ������a��P0u�0뿉n@
�r{��S��b82q.�A��W�`O_��T�x��Y����{n��*-8BE"\zT�Ǧ��+F&Wk�y�����`3P��O��J������̖�y�����ҳM+X��X��8ɽ�a�W���;��%�Y��ʋ��I�-Ӗ���{c_��E�� �_�W� $}K��x!�ҩ�-+�g�_�W:�k �b��#0��̈��XA}��7��V'�;�ԂA�|i����y�m��}H�q�&�oy�E3)e�I�T�ۋq��T��9���ӝ�z�i=��k,�P� ��1�+-�Pӊ�g�}/�c�f�I̍2f�l�0jR����q���돑��kk�����Ч{�}e�,1+W�(i����%���e+�V�h��M�٤��`Y9,�ɁeU̺�/,7=f��sϒmI��6P"��ۊ<��e�5[8��|M��F��A.�L�B�Lc���բEg��Ѩ�)d1a��y��X�zߦ�$�e6}Ir�M�~���A�S�VA@.�nj���)l���_s��[1�F�XwE%OX.����4�=_�ӌ�<%4SZ��Q��(4�O��=EQ&�}�M�y�����������j o����(���,��~�w�~L�#Rw	c�MG�Q�=�o�ml����OqP�י�0���H��Uq�S[F��V@��)�r<ע'9�)o)�yxhX��xV���s{u;E�����CӋ{)��%��Jҙ�)��J�XL���eZX{�N�����*i$�t�8i6S�U�El��Z�#+��uni���X�����>c���׵�V��\�/b˗$*��=.;M���4�k��*�:k�3���lxmT~�K�+֔引�
4���p%��zO]}b/Vc�	Y��b��m�\e5*�zE+=�B~�x!A�|�^#�k�{>�'���)��k���+J����>oj��u5L�QbÙ{�]G�[�H-����ޮx L�M$N��4�����V�e|!�7a��n퀂ģ��P�°{��I_�� �(���P_��*��,�_F��z��}��
2��:0��;~1��f$ծ�K�/��L��}�������A.Qx+���0�E�K�!��^��LJ����Z�(�d��_����� ~E�ď>�K��iV��+�Ύ�3>�M[j��f�d�-����X��X���.������(EZFP��g2tr�ٱde W5���<�5�S�U/F�H��-��
�l_\��Q��m���
�	�^�Ɩ={�c��b��e��������эq�R*#���e ��Ȳ '�iذB��ڙ�M��j�m1�zG�^y�a������²���_BX=�bV�j'e4W*h?U���'	t�O�y:NUۉ{׫�@�('�u��f���H�m�����(�U������ۤ��� �p�ͣG���b��l���Y��T%R�/F�Ҙ�鲉�B��aI����}�^\�zIY�Z�^W�t���΃�,��پt��)�s-2W�)�*$�}ٞ�=^�"'����19�j��rg)��f�U��f�?�y���1�^t)��0{������ܤ��k�n��
��h�iA)]�R�t���`���J��i��Hp[��.ߋ胪�������ì�J]ҾS���O�ь��~��2��Jْ�n'���wN��}� k���K��n�sx�d�-��W�^<d����/ݾ��� V-#	��K<LlJ
�F�}���[S�S�O~��P���6�E�B"����r'���0�/U6X���t����O���LB�*��A���iW3����u����L�zkrf��9ynb�q-�5�c��u����;����E��w�V�R�PP�
��4T��]t��lJٳ��7Lz^ct��C=$���#�U�,�40�T���7[7g���9���L��C���޳O!�3v�r��nA���&̻K�A�Yp6N��Dn$ֺM�� �T��^g �/���F�V���K���-��4��oU��^�eL���x�6L#����Z���_r<��&���6Pz��DٷS�~�~.\�>��]r�n�8~ϣ@4�>�Ko�5ܱc�^y�Li��r+�9�UXs��\������"���6���=�?�m��C^�/��19n�����_h'ޝ��}0*)�ݢ�ĬZq+��"�TO���R�x���R|ر�]L�v�g�5�J܎�9#`�S�/��D�ݡ.\[R(蚡� ��.Kӝ�0��F��o[��Oh�C�Q>�Xj8��ۻ-�{�A�s#r�U����,�m��\"�g���YT��5�#�7�S)U�XfT�C��i��#�T��)�T/�ԑ��A�h��e;�_���ӭ(�C7z�C1W���Y���>�F����#6��d
U��j\_�^��8~��GE����\��4�xB�h�ѓ���C���mK����D�P�ղ�mh5�cka�'"L8xf���G��ϦW"�&��WaPVX��>q���޵��hW�}&v3�Ԑ*宯�����l���.}�����0�s�t�m��D�,������ v����v!����*X'ApL���'@m�Q0�X�[�`�U��^l �ט��k �@sy���{�~�kfn��K�qH�q1b1���7l�H���\
0."�h+1��	���4g �nNY�yA�]��K��\���K��fx�%�Ｅ�v�G�b�����Sd̩�q�j��
������.�?e�:�
�Aޫ0���xOP~�%�1V�g��(�Q>sLz��U ��l�I�r�rG��6�yvb��+&[�f����J\�C�m�Ra��c�yC>�OQ
�0r~���8�*x��Qh�<0L��P��T~�qhj�����P��Δ�B��ݷ�K܋P�6�/����ӵ��_e��<V��wi5_�F�q����'�^q���eՁ��k��w$��s���{���G�]{�$��]|���WW�/*�R��z���gE/�D�n���UJ�(GCe"��~�iv�e�����v��b��@s �#�r��<7O�>M���il�»0����_B4�UM�l냆Y鵛=$�t8�H����]��;	#J޷6:2#|�[��P�^'ﻧ�*�DSS7�:�/4�3���Zn �cl�Q�zPЙWS"Õ�<��Z�Mu�xM
x *h��kM5�wm�;�D}E���Q-\[^�g7X]��]���<!���C/ֱYlk\Q9�"2d�O��J���Ѧ�e냞�hHLh|�;a�50�@ �n�´<5�A:q��Kͷ�V�O]��i��Ši�x�]���J|��,i�ZC~��旝`X�����P&�����-���T��`��c��/E#�T�h�gW R�20����/���6�YIb���M7�3_H��tB/z�ZS�p��n�aV_��fW�����}e����1����&�K�"��cLc*�ō}2�a���B��l@Z�4F~��l�sP�OU�nVO��QA��LOj�bV~�����4G����PLB�a3b�![��c��<@�W(�0�&���F�t*�R�pM��ޫ��1���U���v��RW��E��$�Ή|�_B��U�u��6�|	Fj��r���_"9M���HR����xR`�P�מr�)�����u�C�s��9.�^o��bdɌ5�Aï���2�!���n�V$Q�GY4��4��2������܍Lm�"���֐LĴ��]�.dx��@�
�B�)H�FC���ș�o���%B��W%)})wT���3 �䠰�3�EB�B4����}�&��+�V������=l@�5�[&�*�=|��i�/`�TP-#����/ϼ`B�㖎�y�Y��0�����K0,�|�`e�m�0,�Z�M^$��������m���bF,��0�U�fBb�L��{+�[���H��0��)���/��m���\"���Z���X�����]<(����k�E�_E2DU��2���~��u��5��0IV�J�B<<L�P��� X�TR%i
��t��B�"(�<��F�e+����M�sj -��(��(��e�
g�h�pS�����8������ºY��B�u���^v��|Cێ��ny� ��Q��)Ƹ~\<��Gd�����_�!��n��K��pGO9�
��~�N�I�g����8�,v	V��6}��R0	!�!��!��)n���� �,ήX�qҧ3��3L���[�"-=�۪�DG�ըm}��q}cB4���G�(���Ҭ�Ch%먨d<��g�|�tړ;��-�r��C1IX�������zA���"X|t��/j4(u������Ǿw��_	��P�,�˳���E ��	���i7N�J���?���(�"������5���D���\�OVV��|�+�'�'��}��w�M�;�Z��p�Ro�h�hPY��uN��ed�,��,hSD����)�� �o1�K�J�\�:o^=}�}Ew�µ�<M���W���Y����I�nqN:�AH1x�7/��?PNhi; ��uM	URۇGC�u��:�|�������5A�|Km�^k��d���t69�Y�;���+�y�K ;z
���k9[�6����������e`&@�˪��	��#_��ů/�F7���.l1��W>їK����Z�i�ƭ���y�B)��@��vgo�TTL�Q��Q��Wl�(@O�� �� sga���x��oV�8��T�c'�����}�~Y��R�`�:Y��'�bt�/d�J7����S���[e�s|	$!�wP���@�?�K"�$E�uD��K�����Å!|ݐ�Sq���BɻupsҥfüJ?7���ާFjA�+��ᄔa�<C�
��e�����^�)�a~�un�����^�A3��z�:�L�*xbI�9��$�a��b%%��S�=�>W����Ud�ꦗT4MR�!G�?���?�jn�:p'NV�����&0�����h<F��s���~�#��I�Я� ����ଏ|�4&J�G�U���&l�Z�q ��� D++����%ZO؊5I�gՎ�;�*
־��$^+X�x���b���,͌ {�8�����mc�%f���/�Cw�q�Qڕ���I��Hg��T�����uU�PZ�Z�Z`�,�W�vQ��J��E#g�Y�$6�}�����ո ��=��t{M
��~�_����L���H�w���~�ТU�J��Irv(�k�����)��)>��n>41"��j%���ϧ��[Gq
�y:y۩�;l�jp#=�o�l��q2��2����p��[vU�ס>�4�{��u���F�:�bz1oI��&�����`�(��j�f�@hJ%���;�����g[A��I�&̮1<�r���u�8`��*m�� v�����k�Z8�&����t��հᗴ�����ic7���S����'�e�1��֧�f��x�(��F�ŗ��wp��I�{��F��,wNM���'mN�8������ID�;������+�o�����٤k%�;�Am��fCF�ϐ.s]�߯ 4��K
_/jE�߉ʥP����e�ltB���3) �9(�(�Dђ���fY��g�������q/d�z����d���mOm��d3�!�p����+�xXGz_����
�oW��g6H2�O�Cti�㷨k�l�~{uێNJ�#]����[��0z ��V���?�囏�P͗TuO�����4 ��h�@�6ZAP��H��.���ˮ��^ˮ�*��YD�AUl�.�at�ղ��E����(�w���o@��>�p�e�瓍���x�A6���=��Q눨?F�C)n���ܓX�zI%����4<�&&"o::� ��!�Rg��i[0�Y̺�W�'^j������-ɕ\�]w�	T�w��<2�0
�W�����Av����[��4*z
n������̒e{�"4O�Į�L4v��(sOH�厵!S�\�=!Z:�{UVk���OZ��*�,�|;*t���,�5՚��]B����Vr*g��#T?�05�ϳY�~����,��&����J���K:薾��6�_m6�R`��Et�Z��N�	�~�@-��<c���>��P��j�/���Wg�N%c@�p�?�
z/�l7\��p}fL���X��/��^�"�e����8s.G�]s�e���,ù�j���pw����AE�Y�4̷F�}q�~��]���K��Ӥ	�7����5 ����a��ʫ�׷Յ������-|�_C��6�H�@f��W�߭,���.��zb.E��a��Yt�]ʷ2���(�~���&�Ա}����j��I��<޸����Ϣ�o��]�^��`�g{# xJ�J$;ѽF��Td̮R��%��� ��@'���,Ć�yg���!�W�_�Ð
��_HI��"�mrk�)Q���_��S�)��#��ǎ�,�"��*qJ�$���SH�>p�ֶ�{X���)ߪؕ�j����Ef��F wS~6�%9�i�B�4���wxk�b-z��L�JGJ������k��>�P����Fq�"�s	��;2z���8++d�NuC/P�����y�����Һ�	�[���>�T�R�<�Ю�lX��"�U����<C�s�U�F����֩U`χ��"@����8�����KCSI�r�	3�Qg��$uZ�+�ْy�|����%��)�EP/�x��Q
��jY-��>3�2];\^��J�W�0S���<(����m�Y��Z�cZ�C��${t�D[��CM�r��P޴��Rݟ*��wLG�I��X�gß|x��_��w�N�×�$�:<��U�ҡ����(i9�/yh@��3ȨD �?�M0e�2�H�+P�,�T� �ǺyA�r��#`ܸlA�r�K1p�-:��ho�Z^��|@�P.uӜ�6I���KvJ�So�
���R����� �]��Ie�mI��������`P@a��)�"@?�SH��$�� �+fk�����eoM;��3���r�����Y�5m	n�f�zFm(�+�9�:���_���VBFU�]��܏�х��g_F\9D�������*V��j��ڨVW£�Q�ٛ�GM�v�썮�YV��)(�PzcS��M�U�MJY�&}���pz��F�Կ=�|�5����5$��e�fP�O�',5E��<c%"T�ƏD��ek@��~3+��p꓎���!ܺ?���� ?�O(<K��of���J]��q�-Qd@�o����f.�e �����ֹv����J���"�Y�lB�z�F���e{���,=�]���w��~�J�)Yx�$X:'>� �/n�Ϻ�,�`b��9J��Q�:���-�k���*����˴�X,!��$��vZ	�6~������eI͈�c&�V*"�b����m�,�M!��f	R�vK��y&s���� /�>Rt��G�ög5l��`� ����cB7�G���a�j���3xh9L}Cgl$���P���� �9��ힴ�R��H����b}.�v7��H����k�x����~����q��nh�P�ķ2v/�8������)�z�[��W��a`OfJG��x�y��7*�|�Q�����Y�]K�2�:��0��kr�퐨'��h�lDK��F���W`Ft�*ߕ��x��"�87�5FS���{��<7)������]_�;%��[	�HOm�Uh�Rk��I�%�c�aWC<F�W�DI�Rs r��h�OQ,#�U|�n�n������l�_Ռ��4������	&�H ڰڡ{j��Q���l�v9�M8�e�2L��W��o�U�uW\�I��RxA�X�cn
���q��u/;� R�E:*6���A3:uc#��:����<��_mOk��"֔��_�Co�+`�K��f��F�[�>�[2w���2c��i�Ӽ��.���iw{����S=������`-#������<�*��X&�u*RN��rW��?.��=j��2p?�{ ����~8� ��O�x-��9uh�&󅩯�<�Mٲ�YK���[��<?�:|EO��5�g����6	8j�L�K�,�҈A=z4'�ņ�YJ����_�\�ԋQ?D���H��
�Dܣ	+��Y� ׌[JȏQɰ�Eq7��50Qu�kڵh�������eU��pS�A���Eؗ�Z��^���<$�0�9�ý�?xg�#N�fdW�-�4͐Z�V����&������/�����d.<��;�{V��	�X!�M�%�\@GV5�;a1)ZV	}�M�[+=p�����>+RG$���h��p6zx����J\i�\�TF�C;fܺN�S��Z4��Ayl:w���l�O�ϑ��3B�˲�G�ԅUn���=��&�m�oZ��J�]nU�������*갠L�r_�^"��'`���D%��?����f��+�������.)�u��J��Y������4(s�q���=��)`6r�����R��`�k���e(����p�,����+xZk7�v�aݙ�CS���C���.��"4V�L��������D���\�����6O�8��*N�V^��!m�	HAw6�@3�aO�6֩�����~�6X�e��yR7�G��p^�W�r���Q爳��	>�\[,��0�7S1ܢÏcO�bq��t�����*���Ë&Ze��Ig[���PZ�:�&��<~n�J�����=*d�UX���('��P}��\{Z'���JG��d�`���B���u�	�J�+��i�k-��ԕ��A��D�1O̊�~�8`�XOk�����2��}:�ʗÞ��5Z������-�57��'�5&V��.���Wr��)������T)u�5��<#vƈ&����8�oʨ��@/�g��1���0Z.f��m�I����*jJ�r�	NQf�55��>�	�bV[��$5�:Q�j�,���Tm��}��l��=�j����Zn2�������-�@�h�N�xcB'Z�?�?�,���<rl^���:�2��]���aߛ�5{{阫���QL�t߹UVw����謩�Bqq�3��`��V�����x��O~���u��d��B�Ԉ�~�:�7̃o�g�Ի�����*�J�ot���� y���Tb�,���x��>�Y@d�H$]�*�h��<N��Ji�zMT�F�����n�֧~W�CTL���x�z�1LW��GձQ���5��Εl�����iK�[ x4_S_�\#��Z
�6E3�	YW�Iي}�iB���G�����3_���.e��N���q���=倨ك�,v�k�Q�a��<K��G�H�w��c�lk�#Aư�N�l�lYp��?���Uv>�-��$�lb���-]6C�x�Cht�:Ͳٸ��.�5����7�[�R��׆�q]�堞���x�E�;z�R�6~o���x!����ȅ�����Щ�Aޚ�������M*:�^\�ح����s����$LI��9���4��I��-dR��E_s�H��dS#�:.r�i���8��vv���a��[J WZKd?�Cb3X�צ�[�閂g�#ގ4�ņ��O�����g��ۦWi�AR��S�8����'@��,�����x=�wz���!"G�eg�t��Q����>���-P�|��.d�U��*`�Li����I����BC�AGX�Q�d(f`��e��]+NjWr"4��\����b�F��C
h���p�A�>�ز�xn����u�T՚��	����	Y��>�㫘P�p��Oz|ǖ�V)ۏ��]����xUd$H�S$F��`�8�Fqz�Zu�8~��Tt�@�Cc�!���tB0�j��G�7��i�p�����/��DIw�[�|s�yg
eXN%e��W!��8j��.��$��&&�U�+�"̗�^���ڳu��D6���F�EB�Z���]C�^�ch��\W��d,xcs�a_��H�4��g���"��׼66D������흶�h��M�K��f/[��x�^��U��ַ�����3z%�{t��B8/&�e֥L���[&��B}�����"%�9�&��_j��5�'��9o���������P�ʳseaw촻Ai�k5�E��r���>H�$��TWϖ�g�'��F������CX���GQ�ո�[�j��8Y1#Ϊ��ޓ�<��W�/�<okQOb�iF����9�.w���]�?tsܪQ�c+@sӶ�'z�O�?ѻ�I�����p�䙭Y��h��^���zj�%C�5� / 7��E �s��}Z�a�����ͭ����9�騷�r���qt�,<����6�p��p�H��y�M�kѤ����`�hӑ��Mfo�絣l@\��WI���|���cot�sB:ޛ�Z�C�e���d�
m.^������ڳ���AI�6�c�i\&}}�4���S����&tN�5�Ӧ;�\z�m�##�pPl5���N��2<&'�S����VE���(4�J��E�a�O��t���-'�9�H�Qn�S�h�p���+x[�=���ge'���;����w�	*?��1��W2x�6�v��?�=�v��m<w�c��s�
��I�-�F_ZYA>�^ �b�6��2�D�_�41��'�;���'�ttP�*F��L_eo/~��pdTk<���'�~���H�86�+��
l�19����7~�z��SM����6�h���qO��)-�D�M��}����཮�Xu&�0�7MK_ׂ���Uz�sԥ�l�D�g=?� ���p�rh(�b�~w�sJ�k~^������ޔr�����SR%���t	�N���j�*Gꍞ:K��|x��4&.�+���A��i37�����X�:�b�Do��2�����q�N��M%o�K.��}��ui���G7���$��莰����*���.n�MJJ�fMi�<�!	����rH���v1(%�"���j7g�Rj�`�����7P0��uGW���/�Q�3f�Ķ������l=�hdb��&�.#���,�'a~�����]J��xd����F����2CJM����&�������8Ͱ���L��fɌ��T����0�;DŜ�к�~����T l!����
���ɤ_jʗxr��=\�Q�;� ��3�wY�5�U4���Q��q���j�ڝ�P/i��IIo>�L#�k��	��g�҃ǫ�]���}�#�9���2�a�rܗ���s�B��#K%�w��H�[�TA�5�I��s�A$F�©�ag�6,��x9@�lF]5�����|XQ�;yM^^��L �.�7�X;���VKf�%��uZ	�82��b
R����R$���|t�XO9�<�	�5k���t"�i	��)������瀴}WP��M���8�b�o��x����#����7�b9��{�[� s���E@Z�_����g���C��	o��~ݾ��8O���CU�����%�-[��=Aqg7147��=Ͱ�c<��G���@����"��Jҙ�`��?�"S%���I�t�r$�@���gP"�Ϻ���>�����d�{�I��1>�DO-�b?;�M]�W��
��Z����k������T��ܬ���	?�)�7��tN�u�3E���V����
t�+|8��4E�rD�
��lݔXdW�|<خ���l�29,��p�Z°�A�`p{uk�7�r�md��F��Tn�[Q8& �c�v�35>\E9F].�#3��[�せ�m��r��G�����p�S���S��e]�.cv{�d�Ԛ��6)ƄExv9w��q}����g��tB���Ԁ������B�u�~�&��H�S���f��v|� ����̈��v߅��@*��O���fCn�!:b����g��):/ib�$*X@[�<K�(���`E��N�o4�)Ԕ0lik0�N>0	f%E�g��~�-��+j̏��B�� ͊���&0V3|h�v�^��p�C�c���K.(W"��2*.'̔�n����L���Ԗ���r�Әe
�0��a�B!����z��wa��Y��I�d(c�)ᢁ�����s�E�x���`��-��}��i�Hl�}�H��ll�}��=Ur���&|�_6�X.����#	YZPh� \{�ۨa8~�q�j�L
:0�4x�i�y����Z������ӑ��`�:����@�4܅�#S'�Ѥ��]��MLo4��%~L��~�޸�ֻP��a�;�
$��Q8����&���u8��41��0VJ�I-Ozpl�s}��$������^*��l�Hq��G�tU��K<�̍Q��j�w&R|��ij�v貍�w�{�݊
�E���������we�}��4�/]�4w�JI��ԉ9ׇp�ם�p��-�U�{�Y*;#+��5ܻ2U���݆�&o�ت2cj���F���z�~ɘ��\=K)���ۛ���$\�Lo�w��aI����g3D/�Lj�i^��>�-*e?w����.�&��r�_� �z';"�o�<�A���gX��Qត~��n�l�a��]A;��פ��p�FDډ���7��ǇDlȔ!'.��	� ��m�x� ���4��� ��۔�F�F5����d�j-���t�Z	Ua���킗H�Z��J\񫵼�I937'���V蟜��Z7$�����
��:�2����薿M \a�4
�w�NV��d~�9?<mG���L�a�P�i�.v��o��
+��RvsJB��d�����j@��J��N|!Н��5�FT�7h�k*&��k��K�O"�gF]�<
6�}��l�p�-���v�J�����en5>L�?��:�6Sl'9(�덛�	�1�T㈿�R@�C}�#���>7Z�B��-f���-(��k�[��x��%�3���3�AdeGV��u�J}�Dx2��s͐s�8�z��D�ޚ�e����˔�a��wP���S�:�x����z�ǧ���J�Ø�GYǆ>�b^ꮱ��>+/�������f
��0�?m6&M�,��+�B�q!wpRw�;�˱Խj����O�0����rgoX<`=I�P��B9�`���P4��7�}��h�B������	��>�+0ŮO�KK�p���u�"��u�eư����4����Ca
CY͞T����)�xu'����ĔFs�`��a6m7��U�E�j�-�.{�̅����p�l�:�

��I���u��lA�X����W=|�W�������7(�$R	.
-�� ��ߦ'y6���NE׀H���f�������2���8���?6t�~�<ċ�`K�{[ [�i<�[��ɚ�_{�����Z�bQO��-~�2Uz�w��)@� Xo����3'���#�|�3�x�s��O:j����3֦
m��	p����P��ˊ�����8�D�ةZ�c�����,?69N���z�
ӽJ	�A����|�xn��l���A�4#1[�{�c+�2�:	XӋ[�'[�e�-1��WR���\�}�� �2s�ÜN�M�9��C�۽t�H[ߗê �C�HU}6�x�7�����2�uE�=HC�����@�hH����)6�������Br�@4%lm9�rY��� �wi�q�ُQ߂���;���=��f>���V`��o���(�m��N֨��QI�쐟��$ŲY�4K�ޡ�d;�y���a��{�Xf��^(
�����R�Ƞ!�I�K�A�濻���Y��/'���v��敷���c*a���)�)���v#�%?�v�ώbq#�M�)Wïײ�vn�w/y�"���j]�H�����O,�c�/Y[1ݜ�MR�&��1�6� ��p:�Ad@�*��^|M��#�n��8Ƭ>��_��C�8��ł������S~�9S���8Q[��V�|���%�U4��m%5�]4�4�W��"Hg.���
S),/D�e�E*ΉAg���B$.���v�R�aҏ��cT�=����V��R���2MU"��~���˴pt����S�L��2��;��C3�_�87g���#�&)i�ƶϔ�a.�nB�񮫶�����킹E�M�:5@���<�xA�Щ��T8���<\��v��7�z��F��AN>^��p�6{���9��d0���|k�}�d�w��E�c�&\F��	��	(�t2�Dnւr_@�����(��:E�����nod\͘;���"�|P�7a�?fG}�����y�Z|t�=u�,�5��sW���-���[�Ӭfh�q�W�U���|����I�
t>�_2�6�4E���(��ehMYuqԔ��?�L�wX�_K��nR�Y��p;r��+��
P!��~�/%��n�H�%���/傊y�eXo��d�5�(���
�5Y5%E�m�Q�ߦ����v����� �=��v'P��>D�M�N�����@"�okI��f!��'�a�U���ن@�@0J$�1�c�Q=�T��xn��QL;�cg��f#�.���`��]VR�w������P<��!�k\��L��s��/2�{U�,��Z�7}<@W>_T�N�^�� �	�t�3C���wP�=�.�}(2-�&P�Z�x��X_��F������mN�@�=u��\�R�Eoę�鿀M!��F�JY �2�,�l\�ƭ���(=�j�������!6=�֋�R�`H�n����8�GC�H�k.p#���"9+W���6��)W7~`�˸� ���O��d|	���ѵ���G�Փ�Wl*V"�9�I)��;y�ڗ!��
�[�Н�O�+�gKB\��Bb�g�ѭ  M1&?%���>;Iar�J=����<Dߚ�;�Y�U�=�_��p�!��-s�:*; �k娓�j������9����Dc(��)�����z5�
�����*��X>��R{#�q�8ĩ��j��9���\�~;�
�iNZj�@ P�Y�����Cz ����B���Q0�ZX�޶�"�� $���}G�S��Q��,�Jp�K��_m[�g�I����]^^��W����G
�z4	ڕ�_'a����Iȍ�򩊠�'*��(�C{��|ً//��gήG� �X� 1��ܿ�)0��`�u\�NhZI�P{���Ru
�i����Ѡ��֐�ћζ��<|�Q�r��\��C��e�
`N2�l�c�ϕEe���_�\��]{3�*�T��D�O0��L>��9R˒M�ef��XW�FE���b��8���;a�v��oqF�XHMv^C�S}MɞK�{K��!�������U~F��ئ��x�SҼL᝸������o�-��LH�Ҥ�u�Ǘ��@#g,�:�Ț���̞1��2��mg�޴�~c�Q���{7���5�T��F$��$	-��;*�̧?�:������牖�*�S� <�P�ȥ�e[��b_S[��<#��Q���LL�K�H\R%Y�0R�~n��J4+�3����@��Y�Y�S��BFR��[>���<�]��+���2�ʒ�Z�����1\.ڛ�
g��K߃;� �)⍕��*�1�B�w���U�t̜�>[)�q�g�҇�>�Qݴm���K%��_�I&��4�ʝ���pk~�]d�e�5�LDzj4�k�9,1Oz{:q��t�>��yA "�x^+�6>:D s�9���M
&��[�Z����Q����SbZo]��{0��mWd�*��я��+�f�E�ּX7z�#t͞�m�U�b����a쬜�lAy�R����W�M�.��	|�H���Y~*��0w�q�;�$�Is�#����N��_�9����Bޕ��rq�Ѵ�i�Ӱn���
.�)pI�	��p�%_��=e��k��\� ە�E -[�ti���0Ȧ���k�rGsJ��*o00c4�4@��d���S���z��i�L�@����l����`\#Ԣyq���&�p�{�$o�Q� ����ff��d�x�y	�����T�Cq�����p�@�赟��=�Z&��0�0KxFo���o��v�_w�R>0��˺]9d���Rf/����z��� _�Q@�P�B���S� b[.���.?S�����Zy��CB�o�!k�-ύC���[�m��o��X��s�Ƞ��,b�;]�rJ�hE8Q~[�D�ok�D�:�{���Tl2y��B�Z=�F4�ء����2��r=r�p�:M&<sKAo�����gz"i����(1�� ܸ�ϧ��ށ�j�����R�=���'g���F�4�l�G�h�m@��4�s���Y�{	��<�����9a�^��31
-�A����2����U�Q�ale��w��U��'Ƒ_S�#уP�h�wY>��f�Q;,g4l�0�{����(����E �֣؂�}�Q�&|����-�Rq�����eo��n ���0	~��Tyk���۩OE{��'��>8��-��	��Fn s��9֗�M��b
 �q<(q�8�<���<d�rL��ǡ�9_�eI��<?�Y+'�1�O���JCDǖ=�������n�[����e��a���N��*BVW�*�o�����C�X*.�{�%(�s�Z�G>5G��#@7�Gɸ�V>{���T|~�l�&0���&f���e&�ַ�e._�)� 8����TG��*�t9��N�����8�x����Fu����'�s}�>s���T���P#���權���O�{�����I(�S�69��lR��H�Lk�Y�qx{�$[o_/e���}x�X��E�<�AAwf��y�4d�Y��zё�b qޙ�(@�s�n����߶'d��]��Ax��I���;򬰑W�﹗T��/#,�9�j�sT����(�b<���[~wYs����;���S�*��|:(�$�3D3Ǆ��W����_��f~�]J�:��ٝ(^4�^����&,I�lZ�<��G�N�<Ňk��*��C)���bJ_&�������p�~ 4�1��m����B�A��<m\e��#u��^���&?4��3�3D��p`��C����y:Đ1P�m��B$F&�>�t/Y�0_��rbKfE�q�Jv��e�g�mh��*�/��;�>��O��ҺXl����$�T�͛iJ�f�6���_��zu���4�dK��8��0.��&y!뭔�ͱxy��D21ĄF�ޔ�N��ae�V?j��鴟�75{�\���s>���"��}k�x����ן_(�H �����Xn[D�� �cK�����F��d���xcc��R���Y�/�DǜZ(��ݶ��&�J2#�ϿΜ�KR*#�Ns�8�lV���Z�\�����⌉���Cբf�';ö��R����\��ԛƗHO���}�aTQEob)�G���I4>M�;i��=�J���]���d騯��ZŨ$�§O�r�Go��y�6��V���5����-9G:tL> �iN�i��l$[�T/��M����`���{��Ѳ������,|�ˬ�+���*�P��(�~�'�!p0���T>�Ӑ�5�wH��_����#������5�5DXD*yV�!�ݑw�Ј�`��I�&���hc�S �,�G 8x1�F���������8?Ş}�����"�!������x=\<�����`��=��!7�I�F�Mr[
&켃)֥(�'����3�����M)u�@�E*5��󨉴�3`-ٞ�ʜ���A^�E����&;��_%n�ݹ�}��i��p���ؼ�hU����jD�Mw���<Z�k�ݸ��t���)�)/�jv�HЇ���N"�$�SE�]����b�&R>^R.Ntj4嚇�MV1�e�A����Fw����^����֑�aVYf.���^R�#&G�����7�i	��{q$6!��|��77n�?�U_�VE9NŹ�Jr��;�^	��z*��ҧfj].&���}���/M.x�*�:�N0�V�����A;@
�Ld8����:M�Kps(�s������.Y�5��� J�3 ��W����~ޕ+�����mR����m�4���9��fVOA����,Z$����G�����_�M:�˧��C#�s���$���i����Nܒ`��&<U&\¾����{���e���a���jk�X�t� ���e�5p��`2Ϣ ؠ�7��Ǚ��R�Q�$�/��g�b��r���Nt��E�S=T&��vT�{q�����0%�ݿZ������d�3�*�Ŗ+w6����_ ޥ������>�:In�oļ)X�D�����d�a��?PH$���(e���W���qv|7��49�c�W�׏�+���\�q�n���P�hW
�K��__h�� 6L���D∣� rM#ļ�[��(��a�4��ēn97f��ɲd�d�DVjhb����	����f���=��d���W�Iӛ��y�{���F�PpR�ob%g��֜	n(9�/�7�&hL��$] ���N�Z[�a5W|�ƠA$?�_/˸��y���V�q�}������ @/�0x�쟐�� �%j��FQ�AKR>W��%$�id�5�N��"ȿS]N���h�2�����+�^]���*,���r�'�����5����GO���4���n�WgjYG	u�ӧr����֘����4mFg4��1��+8��5�0�T�a���:���X�����q�����3��[��mH���)��@�gh�ֲ�d4���L��H���{؆��&D)g��>W�5��_4���\i��I��
[I�D��,��7	͌�0����dI�y�/�#G�u�Τp�\|�2P��j��,_3�v���8�^�?�t��8~��+�0��k�G�'qJ��%峖M��O�?nUx%tsf��������<��]\0'+��W�1�_a���obD��;���7Y�rj �%x�|��u)I�:~L��lǗ�b�C�,�<3��vAR�������QS��=6�5?̞��
3�&$忇)�����kG_?�)Z|�	:íes�nQ�Uyw8��
\�M'�ҭrs�)�!?�z�4���7I��D�B�E�x��<��I���x��.����DX��m$S��e<_�rũW���8+�v�Լ��"_,����ѸF�,]�]��[M�o ���LO�O�3Ǝk8�G������E*�JV��L�-p��J�JI�I��58�ӗ��']��2��{��/��\IgC�XJ�N����s!՝Sg�֕*
��>�PT!�F�Z�~��NB 2e�
����ɍ)%��N�>��R�}���<	�;~^I��T�8���S�ٽ�7�f�r~6��@�
���H	ǨS�t^2mK����k��m&9 Ͽ*���~!O�rW;^��5}�(���{�+F��x&Y93�*T�녡垾6�jB)v���Tn��=�C�H�WVMV��t���&�Es�]{�Տ-%Ѷ�{5?F�+ y��S�P(�p��H������o9�٠�ل���pX��I���:�[_�����T�h��q�:c�Bt�pJ�ؑ�0�UN	�����7�Ь]�C��F��;�Ѷ�1��@`P4�ǉ��CHoal&�3�9h��i;�`���G���a���{�&�\l�Z~�V:Ā��U[��I���W5�Şb��*旡��o,���b^1����#}�f^���s�r��sN ���m �Y h=�zoD�~t?���@Ʋ�."�h'��R��Hz&=W]�Q�z�"%q�O�mL��dc2��������?;�:AG�Qn�.g�w_ط"��dkQ�3�P6�%����(�!��b����ډ�I1�9d`{?E�z�!�P'*�*n�>�����Ś��z�����[��\	Gvk�3sOR��f��V$p�l$쨆��>	8O�C�Dۇ2@R��{z��t��XK�����p�S�y"R.��P��P�`�h���9�
o(�>��,�'+���:��+aة�������9z.Z��������6Ge���|�]q�KY�3�p���!�Y�M=[:���Ce��5M�Z���$3<:�!�#tq�f\�	0'(��;�����/
��RA�ΟJ߀�C�������_���7�`�F#k~����>/��������c�(�������0N�\/ޏ�YOs菶j�Lτj�8B���Wnn9�Pat�j�����&����$4A�T�5�
��);��57<ը�g�-	�J���X�|��	��'U����M���[?��������H�b'�z4��XNuT�zB	�R(����V��q����ݹX!&SvPa$���W]�A�ߴmԄr��>�nf����u�ްn7��u�\�6�K���@��tM%(*.�GC�@%ٔ�wX���e�ϧڛ�<goϙ�~�1�f�BH�kH؍tx)����cMڍd.��@_MZw
��`\����x�^��M���H��^�N�SN�Ԩ ��M�S͕��~'��d|\j��3pN���[����*|���4�K��=xH�̑�5��O�,�9��#�0��d�C]�y�H�|}`zա�di.��}Xh功��)4��f��F^�-<4�1%���}�1ރ�B��F �4&�TU��YUњ��S<䍞�*4��zP)��ÇKq��I��+�keL�ΐ��%+Xu�Ϲ`)�Yٙ6�2X�l�>�|π�CA��%a���7զh���a����ܪ��|=�;`�������[�-ɔ��%�r���ݲ8Q���p(�-���Vo+�:v� ̺����6!��p`ت2����P����"���q�B�稿���K�OA$m�K���V,� H(*`VR��>�t�ºb��N���T"���*�o<�Iʹ)tLI�I3.��˛F"%��w ��ƌ�#wUH�n ���B��9J���,c�勗
{��y��_�(��ɜ01f��q�����#%�ȼ��Y`0������A�oqr���y�(��G�쌴��w2�/
�K�Jr)~��X�oM��͕qN9Wܸ�)%��+���7M�N�$& �dp\Vs-F���� �h]����GYrj:��o
l/'/������Bq�i&i��H.ի��C�dK�S�9H��.�(ȣ=��j��	�_���� vg�&�����E�թr{^M��@��Y���"�Zqx�ւ\m��@�4��<������${�zK�����&<�!��+fe�{쵇?6���S�iLW8^��a	ʂ�G���&V�� le�O��\	�b�k��m�����@5L����|h��� *��߄���V'��Q�x{(��=Ah�妉tLZM��b�I���ܤ.��%�����q-O������QF�2�V8��G-�{��p�y�+����[E���(����Ԅ�)<�������}�oEv���X�D���I�W,��oqǱ�/��Jb�%����k%x�0E��M�*,�Ļ����k�OȺ���_�i2#р��v>ix|Q��R?nn�&FgB8����#�_���C����%��dUճ��K�����(���������R��J���"U�i�����"�N�$O0X�P��k�+�xp�OK�u�8pWl��Ĳh�q����;�����=}�[�=������b<m�JZպ!�.֖Řu�َ?K�x�6o���9�ג-�
Ʋ�؉���_=+�P�`�\4&;���¡4�2��q*�Z̆�h���A�(�5��/�c0	b��
�g.BϾ
�N�1׫&t#j��s�C�ؙ�빮iPX?��rqj3M��x�!�e.b~�uk�V�T��O����]�!
� yV�^r�6\���c犊����!s���]�hg��[��j(Q�\����<�Q��4��<�F�.Y��-b����f4.�'�-�z��^L9��B�ɹf�HFT�^�s#EjI+.����'(����՚�/(��`�OGD� 3]FM�?RRJҹ����!9�/���(�1󵥼�Ou�̈.��&Fr���9������B�<���$�s���"��E\(e�tu�Dۋ>Y�\�Ol�Z��_G�cp/废�L��&��[���.x��:Ģ��u"zv�ә!V�,+�ʎ�j�0��쇰]��]Fa����\�On ٣I�q�A;��O�DWS�Y�K��]Y��I��1���bw�"x/��q�v6�h�n��c�#�o�����x��:���V��.RY�-�8_T�	�G��-�Hb�U�h�]�fN�ѹ�.��u�PN��[��yÔ��������/)bJ�Py��G�rqrlJ���㍔�_Q��L|S�
��؎k%e;G�:������#)�]!���j�qx,��ކ?K��uE�`�#2׈��H
Ms�&oD�~6��>7��V8�RC6�;d�9��K���x�U�_�S�����Z�v)�� ����$���R������1� 7����S�v��Y/�aݙiVhAE�(ũ�?���a��EW�� �{��9vx�`��,&�B!��^���j���^\8��������d[��ٜ�}����?8q!ޥn��l���]��W4�bsP
�Sr�5*k	�y�_�[�0���0UI��W�bmC�������h��s�O�q�cʗ����(�ѝ{a�n��
w $�6'c6v.�0<���r��	]}���f�����Vw%io�TQ������i���[W�CA����f�D�n\.�'|��%:�8B��d����E�R��Aˊ[Ϥ¡�r��1�\H�1n���þ`���4 kI>r�E��h5�,g��p����+�A����2OӇ�/�l*���@��� ���p@v��+��QV���A�$]�������*���ȧT��k�~l?��}��q���Q͸���;�E��P���ǻ9yca�������{�Z��U�Pi�L1]JHtx݌0}'�Ÿ���>��ށ����)U\&(��#�a) 6�f*ʔj+�!Ċ�*����&u{�5��	%!|(��Z@��ym�0�?��韕�`	[`���}%ٶ`��8��h];?�멱EI��I��"���P����N|ŐOЁ�K��c���qPH`�!�7���w&�������ώ�+}���d�7}X���ʜ|�H�^����:oI�t�_�A?��
E;���R��roo������
���.�C��Ե
d�h6$C/nt��m����r۪��+z�>,�F+C��Gr$��%yYD���7�cbW�\!VK�f���-��7D��!�:��l�FA�����R�#F����m��ҷ�a�e�1�����}!bM���{����w�&
R����*�^ȥ�Lh�w���[ن<���U>QƳ!�Ӝ=r>�NC Q�����>A��l�[�c��t��4x�W�Q�Y��5���C�$�-X�������(LV��>��������F)�%X���'�6r\ƅIעL������d����g��0����{Ӫ|���չ�}{�ZS�}�N�xp��`*�`}"wS���0�e���mh������MO?���?-z,��V��M0j.K�B)�~{t����PK�����nB��4�<��^6�n][�##�������d�i�{Sx��_���Ck��a��mE�2�Θ�����p� �W���*O`ca�T�
�;��~}H����:7���`��P�o�>���Z�Wz����^���Å��e�e�|��8T����^�d����?`ϸj�I �I���?d�Hܔ1��ya�$m������V�T��#�݊F��I�[���I+��Wl�闝���)9�3Z�3����3�2�Btz�[@�/�D-�N�P���l^@Pt�Ш6*�)ɦ[�Q�a���D�)�x_�az������A/j~��� ]���^�+v��Tf���c񴠃g��\�*	H���e�a`�.�:G�&}�`�"�(�:��6��";u���[��z	6>a^�P�C�{d`;�B���&�Q�z�Ԇ�'6W�����L�'_�ǰ!iel_����㟳�j��R��@��K��h����ڲ�����S_r[7�<�%WQ~�㲵Z ��Z�'T���2u��Jͥ~};�s�[[k� )�@Q&�$��U��U�pW6@�,������Q���zS.X����;j a��:�=��I�	�/הN�X���(�3�v��N L;(��{_	��2�-�ê�.�$c:/��77
%���:Ҍ�|�I���ߝ��}�vq���J�-��CX���H���`?��C�<�f�N	G�P�"��l���g G��)W�M�p���0�S�7;��!J��Tj�x�����	y@mi�d8i�,�;�:T7�ľSrKv�>�W��x�J�-����h,�òP�Cć�A����\�Y�ݧ�۔uv��B""W8�n�:�e�M�KB{�Qmj-�eCA[�)�_���'���[`�C���S���.�Tb���S:)��۝|@5+G鄩	lU!9!����iV�5ݵ�����Y�j��]j��� ����)8�jz>M@l�����vî��y��,������LZ׳M���r���i[��vpИ 	zO�{I�ƅ�s��^�UـUr����]��r�
q�K.aW'�"ė�����6�#��
mTyӗ'0��7�.���K0��%�g�r�gun�a�	lI�Z�f��E�‼c	�@ ���މ���:pF�\*��￶+蕒 ���R�Y�b�K��4pU�,�^͌���C{�؝��o����H����aAZ�<���A]p��x
�o�c�8�e����m�D���T@�=?�)ph����y
Tu#"I�K�cLri��#6;�@h�����g����'e�U^u�����t�.�T�&1ǭ�'��s�2	�킿�^ϱ��/��Ǳ���� ���Jq�\[�?�[4��'�wr�E:UN�ؕL��W>�V@;���9�+�h�>"����	k�e�}XUR�s�%h�˜�&�L.���?K���N�D62��l&z�B
C��|�%(��Ǚ��F�S�D��$c�G]�^~k~s��cOL%G�/?V�O� t';���UZ�~E����.��N=�L�����\����N^$
ə
ʆ*<�l2�N�{x�n/m^'�Bӱ:9�����������P;��#bN]���lAf(.8r�V�˄�aڵ���E{�l���<Z��|l@0�{@���!�����4�ş��YN���14�Abr@��-�5$���>v<�c�^��!�b�Œd�或k?�V*�%�D�)<���mq�h�	�7L>lg:Q���CZ��DJnQFym	V���vA�~l�}H� n��Z��gA�z��3��P.=�L�VRM����u��ٖ2�Q��lt-�J�8���p�M���ɍ��M6��Ĭ�P�2�������{�uoI��&!�Zt e�C?hx�wS���2�o�G�/�=#%1<f+Z��hVbu�9�?;#q��+1b$��Ul�q��hzBGzߑh �9�2��H��Ņ�`�i���q���m�-p-^������A��s��w��|���D:�[��)��T�^~��U�y��~�����X���,�~�j讨Ғ�S_�����:�^fN�L̩�6����v|��@���w)cS�tD�$����L�;�@
ív�'��e�3
6�5,���k�P?
��b�PK¦3��3��-�4/�{$��"�Ӧpi����b���!�HϿ�F�@/����ZP'��,D���\a�e'n+Ս��#��~���0��l�s��%��4���_B�����*ޘc�x� '\�q�slk��p�WAL#H�^hzפQ7��� z�T$WƖ�PX	y&����p̭$�ڰպ櫸w������� �#�9�iƀ��B���;��Ɛ�H�J�w�H[t �Խ�u�m�zi������{�2t����,��[b��7$��a%ؼ����CX>G����prnaҎ-�߰�_#����q�>m��	����M6_��ě�|��ǈ�V�D�<���*�
�����*�h-o��?������c�R�T�?����*�A�Q�Q�ǉ	��od���~�̕�[I"���w�N�>�=��L�9D+t_7����ST�%��Z� P�4�ܪ��m�V��\>������"���NCap`7�5�s�xhϖ:�����I����ӺӘ��|���Õ���W��&�
My�5�,�����c�����#GS`t�&�h%v0��)��#\;���ؔ���tD �W=1��d@�qV ��%�s�M���$ 2,�H�Z�����^@-1���V�Ta��!��,i�� ������M��Ŧ�����Iف�`�����<�w�}�՘�I��9Vŵ/�X2!�X���6��B��n�q��H�0��j�}҂"���w�/H$*�E� �;�'�w ��?3��1��An�un��b�j��h=KS&�;tI�1t��pWA�!��Oy����w2u��o�aEyE��Î|��Y��?����?��i������6��8� ]��N	��{��_k�9,�G���0�Hg�������>3	�.!�(�`����[��:;R������S/���_D*:��+�-A.�N�w(/�F>��>b�Ǯ}���zEk@�rrc�[��[�k����Q��+La �����K>�y��>��=���_X���؆~�I�(x��3g�V�ί�$���%d�	��@��"���dU%I��V�j]��;{�07w�Sy�G�[}o�b��9}�)6�ܿ�9Ar�#��M�C��TW��'��YM����ף����h��OV�)-� �N-����j�3d
Rʂ�
��ΝӐ�N�H�������y�m�*���(̃��E؟s�W��D#��9�����k��;0��v���}���?��=�E9���ψ0���_���B�wW�|��]4vT�@�L��A�nO�"uJ�E����W33��>����"������$'r��T[Dϡh�`���
_c������1g�*����K�����k+������e� f�΂#s�k_���J�l����'K��<�(]xU����Mp��g�z0�G�@U;FxY:|�
��c�5<�L�| �<)��$� ���V�&�x�����f���:���>X�Pb;
�W����� �����T�f7���>b�?s!�1�>���4���� ���_ΕM��c������D�3�g��6h���S.uC}��.D�/AJ'��+8��2�RjɿQQe�����Nɝ?j^�$Ն���	�ɝQ�����]���^{p^vJT@�`�៳��I�ɤC,��J9�3+����e�G~`��P`B�&������b�D��G��K�=툋f�[��fW���\RS���p�Y�B��T��k�X�V
�m��×4��,̣-�a�3��A�Ə�z~�)�!� ���Ǫ��z��HH�`��`��O�n�^�}�#)�w3��HOj�Ml?�x�S4G�De$`�R���ݽ��6&�������Y��>����#���̗��P��(��EA������{�v�z���K~�I _�p�3�To�c�!�n�f��`�.��)����t��`
}�Uf�
��hfe����j7���Rnv�b��X��<i��ρJW��0����I*|O�'_���0�kF��ȊU&��y�,�㮹�,����G��a�����+��k��M�F�u��Xǅ`��AQ
Mz8�(�~-\G'�%AE��-S�S&�$bW,Ώ�W���+,=�[{��[_�Q�z�5u,���r���s��ý�[�.��9 �K<�C2�=�������8G�ܠ���JAD<;.C���a�(bR��M���?7�-�K�)��%��^���~��
�VU��ĸ�W���+B#��3����
z&����Y��N�,����FA2i[Wsq��6&��I�X���W�v�z����!W���{L�Cc{=�Әi���wb	*_���_�lu�N9yp��^��M�y��AKɃ�!�A�q��y8�"�Q�%%o��I���EɈ$�#���F������?�Ŝ������\��Ymv�w� Ny�EB�aVp�s=\j8��6�1�h���XcV���م�м�Ƌb~�&�]	H�g(x:�\M���@4fP$��OW`�=�.�\�j�������a��~�O&.pn�2r����Vt�
�F�Y���!q�
�q�� �.AG������B,�T�B껀� T%Iy��)���3b<���/D'Q�l�nJ��q�a���SL,'&30ʳ����^:�"�?�#�c��E��&���|��Ԁ���a��0ݎ��AC�@)��sC#kƨ�B�`���;�?��v��x���0/���7���ȯ(��`�q�&9#6QMΘr�w�n���[�MC���L�"F��%��z�4_W���$[���bD:�U�R�����;�]�1 �l���?�&O @�*l�i���j�K�9�uX
$���/�{^/#'�d�c{u`2'��jţ�@^u�k�h�&M��)5ϧ�`�������~=�.�þJ5Dd��N�41y�r�WV�R���E2�:�\)���c5��a�Z;���cYư�I���|���Žg�[M{e�ҁr��,:�׃��E����@Wqb�Ӎ�]����'x&���'�^�hG��ª��A�*����&0�=<��1t�% $o��G '3��Y���P �Z��������W����VB},)����E����Q�B���J�n|�A<��e>H)B�|.T٠�d��� �C���<c����j'n�BNŝ���-��]H$�e�I��+@.�W�8)}<�	��*��`Q��.�4L���݊X���8l�E���K0��ܛ�~�yw��i�ȭs)2̞����[�J"��K�l���z�.f7M�C��搘�y$X�����ZmڣV�U�W�0��I��sMZqCi��-�1>Ŕw�±�Ҽy�z�#�)��6�[䱹q��(9�Z��i��K�}�d����
�J)�u�<� S�@3[D� �<�\��(^;�q�֚�ǋ�!�_�6��SG�X�X����W<,��;��A�٨��0���L�<�i�a������Zir3���Xs*�=����6���D��z��MV�����2�l�8��2l,��/�>u@��H޾�
��6;��)�*�Kk�g�SQ�=dnO�`�~�b�dx���q�yQr8��rY]�ՠ��~�=Ռ4A��Y �0��^�J{�8SWrM|#$�HguS�WUIl�l%��6�o���#{7AR�J������l}l5.;aҋ�F����e[��[$3+�MW�f7����ReM�y�(��M�v��4Pa�#?�c8@U#a�B'�u|�9�9�:9����"Ns.j+�K֟@M��aYAmL����~�������j�ӽ�k\�<�����b�]�mS����I�ub������SW���ŻS�1�TpYtM-`��9��_9&��U_����
��I
�廚���X�n�D~T��W�=��Ԥ�Ļ�H�j ��h��Z ��T�m�S���T�`��P7��H^"�uSoW�.�.:�zg�}Wg�R��PnJ�ա���U6�~�}����T��K1b��o�|%����NRر�4�xG�v��ڍ���s�'��=����C\��y0�!o�ƴ�����3��xv*�bv��� ,Һ:��!�]�|/碻�������!��(s<r�5Ϫ�+bۅ�/?J����hau�S��F�8F����72��t9V9ơ1��=ST{̜�S��hC=���$��H~�d�%�9�����n���z|�2��#U:���T'e���$���Whirq_8�nqO�
��n �O:h�M�A`��kB���}5¿���B�e��!�82�~�N�#(��,$��n�C�`a �22����T�3�T��E���7-�R?6�����K� �(���'��X�ԛ���^}Vߑjn�]1M�"[mޞS���M���J;���"�z�D�O<�,`�y�jb�`@5�F)T��q��dk�C�ڍ���&�H֣1�@�)e�A�Vt�Ƃ��h�q��ʉ��X�5�Y����a;��8ɶ!��p�q��W�n�3�m�M���:1!�����'@d��n��F/C�K�l[#��K���
��V=�z`Q|�dZ_Ǻ�M"��.N_*�<�*{߉u�?�~{�qX)ng|��DbH�{�gRL�!�v��2��S :N�Z����mՇ�(�V�Wx���-�ݲ��Y	�Kr�Fi�m(IV��δ����!Q�K����0ǂn_\��P������k�X{`O}j5夅G9��=�>�1�����i�A��/H�$�?�9�x�L�J�-2��PpvX���& �2�HeT=�z,�}@(��H��r[fJ7��\�ݥ��U2����;&L�I%�1M0�tb���z��Femlv��`0 ��<� �0�Y{$9yq��މ��eD��B��C��?���L���i.��*�!e&�'�z��Ɂ�T5+`sZ3�v�7C������ǁ^w�A�`��4P����<bȈ�n�,sy@��dj3�,s���:nS:3Yy�6����(.~�����ư�i���q���	�	R�����
�SL#�ي~�;ڿ��JN
Z�n��O��m���%�O0·*���jݎ����w�tTa�]��;^ѣ���=9f=�:�	����%*�(nP�H�;�7	��������0��K��`�\��.g�'5,io�9�ى�1.�M��hû���XB�Pg�#�54PpИb�N^#2h镈~,bZ��T	\�P~˓����A�$%�J����㭒��������[c�i1pQ�O��L-��q��v����:4�����Lb�9� �h�s�m]��`�J��ڠ\!�[T����L-��2O&1�������+���f�8�V)��"&sPlQ��k�j /+]�\֬��vr�7��쥪ǵ,�T0��a��!_�(����Bٞ�Fv%�]�2�}S&1�>:.K������'xy~����1T�7~a �O�5��V�k_�N5�@)|-O��@�fH��N3��兪���0�Q22���<��N�zZ
p�e�B�����1�B�|ulk7�;uRH��t ��HxW5����N����n�z��H�Na�㧍���q5H�˕����U�V�I:�9�6:W�X�Ж1��k��{�W�HŽM���u�Uk���L���|���c_�mw#Q�-y���'�����H��*��f��\�1��Nq��Fo�K���Foo����y7��~لe~J�%�������z%����DI�	؂�]����w����y���M�Zv�`)?���/J���%�G>��ŷ9rw�C�~�m���?K�?]?��ɟ �Ak�Y2��ʋ�Պ�5}��畒Dd��;W=5+�oByS74�a������W�U��~H��t�5W�-����|i�����O`�xc���T����e���v�u��*Gk$6�&z��A�����4CဠN���
����;#�}��g���
#�����>��TV8�}&�B]j�2D���ko�����h�Ń1�׉�����1y q���U��kd2�}���EƗ~	�9��)b�x)��$u����7�@�$�g��'G�{��{t�&mq[G��TH*9k��멨Mc996ᘕR*���~�5m�F	?� 3�>݋dP��Ѳ���w�0�cK1ږ�W���:�[!���?�04�g{��#�R�u݌���ws@����q�Pk*���p�H���4U�h�LVG��0�Eۖ����l����?t��Iml�Z-z!����"��TFt��:^�,a,}.����}�f�(-�WP,Zζ5�^JN�z��R�E�r�6��l�z.&���g�U���롫&�测��*�<���N��PҤ�J�A-k�w"�b%;�~���dRb6�\��i燱-�#���rMQ?��1�y��Qx�/Cv�iQ�&�i#�i����x�Q7 ��^@���x����>���ome���D���r��;5� ���)��n:�|�\�u
� z��N��>�=Gz/8��+�N�r�~�J�Yt�
��j��0��c7/$���;������}@=&�g�A�ݩR,��q��S.�+��@�d!�ƍOw�׿������Zt�����:�m.9��?=>�zIOZ���
"�Cs��-�.��u��->-�|����*�	&f*�t��HN�-�N��O�ĉO)Ao{�ջ`����0�:�v��r6��\����7��hc'}�����[ �\����7��g�P�.V �2��$3i��\{�o�=admr�n���j -K&lk�}�Q��g��z�K��Ԃ�MI���Fܢ^Bt���k��01![�]�N��Y،���~��g���Yw�J�)��n�e�	����"�@�A6�Տ�^#ȷ0{����j��
����>�^�����O�]�Mi)��W��|�A3Y���h��/E[��~�;_�2Oe�)�j�J���,�.�Ì!��m  mcuZ��T-���r)�֚;�CV m����]z Fy�I%#���)����'�)Q��X4n�5���U��&�o�|R��{�В�;��m��<��zd&������g��+�eCL��L2j�U��w�����]�Y\�a^�鰵�!]�j�es������7��9�(����fH�0��0�o�H��hp5p�� �=�gi�x�oY���$�MM�-4=5����$�r������jԚ}s81-�b���eB�XƤ�M�ez7:��Fb���8m'�9�b���z��,��+W_�J;pvNn�]�I�$����5�����h�[�	-�k�B��`t�(CUa��kDO���m�5��P_}݄8�?6�������pil��O���C�Q�����d�,����'��N��B����d�m�Jc�ޛ�7v���Gٷ�1Gv�<��rF�m����dX���[QO#��7���ãt�_�=�ס�����k�m�_u�[��K��]�Q_��?��΢5��RE���)h@�7��uԮ�zR>�}�4�| 蹮��]ڜ����N|='��]D�?c��8�.X��
H�]�{��l{o$ׯ��U5��@ǥe%��st3��5�[H�sT�TR�;�Q@�pC:���Eh�uԹz�k奮����C��=�����0���Hɠ��6�2GFxf难����Z��2�z�W-��(�Gf�vRM����i��qy�G x<?�ʣQ������{�W9������;�Y��~/:��m�#�(�u� ~�Q�&βej=����l;�cZ��"�fm��,~r �j���&����	"O�?I �Z��4�(R�F�:z꿱h��ɇ���#�Q9%�IէCz|��i,�P81�������Z�/�'E�R"�H�: �4�x񎛟��x�j�I�V(��<�?af�[HL5����2��F�?��#�̅bj���U�������TsMJ}�z��Ⱥ�����WA������i�FnbYx-����XߏJ�Eρ�-��ݑ"���.�Q��iy촷��t�i��\���Gۀ�s2�H��>Cr�2�_I���V��j#����ò�`��"V�哕
�/ʫ�հ�J0�`����ʼ�i:��A�W�4>j�1m����U�P)Լ[�. �\���aC{��`6m�u��2��]��n�Bheg���~�b�^�hPEv�,����uN�q4�Jm��' m)l��㢒����������|���|������ľ�u��5�f��[ �x�� �	-0�����[�{�ȑ��\��q�/��̿Ӑ�4��	�d����Q.�wwoAH"�7�}���_7L��[^i��"��D�s�(odz����d�X��Nz!�<6�9z�F�K�k�b�'�V�}!���B��u�[%�3�.�߿D=uc�<�q�Y��=Nb:�j�l�:˟OD�?J���4R� 0)�\�/f�����������\B�RP4�z�O��1z;{ƾ�2v�d�$����j���$Y�.8X��<_S��z�T#����;`*2���=v�G�9vSa���y���K�ӕ$-*�]6jq�5�"C����G���%��_���Kqį+,�z�3�зQ�>(�@.4�]`L�{|��"xUrؖ��	���֟C�A�Z��̓h�Cy'�)��P+�F�6���:ϋ�/L6�v�]��!�4 �h�uƥ~eԽ��Ĳ5+�ޗ�3;<Q�tEYx�z�/��|����� �Ս;U�<���eD�PwT�xsM-��#�g��]��ONلd��e�m�{�d�	1��S��z+!/r^KIC�*n����@���Yj� lJ�X�����V����
����ٲ{�\��Ka�'q�q����uD_yp?�s�q��U�i�S�_�vugǌ
��ߜ�"����u���(��o�L�a1�P& 0�na�@5e�"ӟ`�KRڞ�'�f��Xu�^��PJS=���YoH�ԿTÇTP䳙����y�2`ב�+[
���	���[
c+3��U笍y����6����]vY�n�^��%0�a�f�l=gf9x E���p���3�P��1iy,Dr6�$ =m��IN>�YZ+��~�<y�����e��wF�o1�y����d�^������v�N,sG+��u� {wUƁ��ؗ�.4C�x����s��)���O!}��Ȉ�ӎ b75lb�V  -G{�4y����6T�*~d,�%d��`M�����X�J��|KJ_�7�# ��P}q����XQNQ����
�7�#7�S�����B\�vw+�,�j=���#��2�)I2Yі��b_Qs�%sqMh֋(�ۗ Ճ��3N���� %���4�a%Iv�I � ������"љۜ�e��6�ǆc��K��K�}?^2�'�5Wh?G��v^%��`�c��6��l�H��F~t��,'�Ag��v�bS��Ems�o���d�OK�h4�z��Va3B֑D�D�x�u�jE�oI�zz�!M�~����C�s}8�~I��,� �/ST�z[�zF�
]��+���u?���)=��"ܑ�G�I~��'�˞��(�M6�*��d�jك���U��#|x�^�Ăl3�6����B����C@�!�%<{�L%1����	u+C�]7��Gg��**b~��ёe�Tm��CT/��,��͸q���bQht{�ӏ}n�G�'�}h�M�������1� 魑���b�&��@����@�5]`y�*e�v���ɤd����6�<^��I�c�����uS�F�2u��1�^�p9�/L�
�4L��{Ƶ���h��59��յ�K�]�"�QX�_@؁ r�F��D'��2W��áNiS0b�*�u��o�������+�1��Ă�TuO��:��H�t��EX��GBM��o��n�lJ�k�3�E�@eg"EI���� %=G�h�S\*)�l�=�����
��f���O��`^,�5�K���/�Ĕ9HU��f&�x'h�Y�wƧ�K�x�n7��K����_!�K�8[���D��:�z��J�Lن?��|�S�;�V�&\��/�!�zĖK��
�%J�A�F�^e�w��%��T����g$7|�Y]vl�ī�^�D����`����-\��D�q�4m��v�+�3}�e:�8��	|��G�������و�� *ˉ���}��Ԅ%�����$EE�Ϗޮ����cD�F���\�F�:�q\�!p1�؍�R�h�	�1j, @��WDh]�@�Gn4;�0Z�vBD⺽v�f������3���Dj8		�faӉ�3�h&S��5�/�V����M^:�R�Oxc�8'�ɿ�u��)���w$p3\î���T����S�"\&���
 f4e=5$�Sw��B�>�U)bJ"�a��F0m8�6�.�F��vv�nәj4,�-���g�~�m�mq�7Į��͐�U��_(�e��%>�Ǆ��S'��Y첛�gΧ��_�h��!wU8G&�`�.�~�C�_��W��E�����W�H�Fb�2���j�sZ�4��ĔZw�̍�K����.e��N��~�	��(?�0���<�,����[L�	�u3�� ˔��O�_DW&'�/a�>��2V��M�dU�e�盛]{��]ͫe��T�Ҝn�uP���g�9��>�s{,3LX���vV �"�	UM���e>fˏ��-,�D� �B�׬}��	���Tx&���-X�b�3�m�1�)l�6yݺSF���&��bGf�YV�믍����K<�i]����e���#�t߷���ݛ��y﯄��I�D�G_�28�P�JiF���0�?\���	���0 ~��h��-Fn��څ��\�Ll4F,؁]?�|�>����/�~"ȏ~�bA^u�m�K� �:�8���畧8#)��o$XN!H�F����q��9@��^�W�qv�<�c�W.�$\���vK�y�HS���0P�����8��-�a�i��?��/9cp���T�>@|�u�4����<� �gT�hIE�b�Z���6�1p�١����62�car��롷�N���4�g�a�h�9����7�}���7՗.w�,�KMuP�Ӡ���,J�q����\�Ԁ��s�.���l� H�](�O��xH�\�-��H�W�^L���3!�>�	˞EO-g�Ң_��a4� '�-YU9o�
�&��rI�wW�������O�,t�4G����ܨ�Vw\�*9=��ø)�$�W����)T�s��gϲ��i�x�@�Ƭ)Yu���;I�b�Ȱ�M����vޔTf�ik  ���=%;�4L�l�Սo7'�=�f�"��;�;oX��qT�C� �+���`� \�*nmH�B���6��9`M�-�)����p
Z���#�x����|뛷�wA��l�rD^��l�����Wƺ{�?����}�)k�;K�=��MP&��;%5щ�<\�fsV��E�"-��iM:����M|3�C��iWy)Z�e�ӾQ2�2?�/Y#��B!�Z"D�
����\�?xI�lN$+�0l�m�F�$���:^!�ߗM3ȗ���.0u4��ľѐ%er�#"���K0�W�ð�ڂ��o�5����^�d����54�����P?:�H��(�̪�{���#r̖֞�/H~�J??�i@5�y���q3tNڛ�N���A4z�qt�@���� �����r�>(8v|޳5�D$���Q��O(�AiĮj�F�ȗ�P��&�������?D�;܆E)��Ksq�P|����2��i#y#�q۱=mή�*2`��$[�����'�p[�0Ɛ��
Q���@�WTe��7�R1 ��e�;0�神ǩ1�5R�wL���Y�q����� ��짘�s��J�~�I�!-�A;�-a�A#c廙�!��j�����|Ư����!	�^k"L��n�Ŀ�V�c?�٪��d}]@�"w1�$q��V�=�@S��^�p���]��MS�V���ek2&y]��AǚԿ���;	Jb8��#�l�W�g�1B��͇x64�ٮ��H_g�U� �Ȧ{h��x{h���+#r�.9}��Lw:8����'��}�@Ǆ�{=���I~���q6m����ߐ���7��{5G��E���(n'�j�g�*^3c��ʉW�	3�]��# �V ���������H;֝����M���a�w���G���ժ�䋜h1����N��P��� -K^g��į|��;+Kp���1nqU��2��N�d ��Z.�J�Z�y��p·����+[�Q�|�	��_�׎w�����{֔�
�����z�¯E�o��}�"Ô�4�����S�S�M�O�Gs�eP
��ԠR�g+&�*�S=y`NxW^:+t�A�K��5Mjm���U ЇPK�"�ZסN�w�K���ȣk;Ϣ/��5��2���!�_j/�����5��Xy��ld�T�ܗ�q�?_/���+gÏmU��:,�5u��{��،VS7܃�28B�]Փ���E��<�5��)0h��(�����-�ƥn�?"P��2(>���c�+��u��g3UopFQh�m���$Y��U��_J���
F���)��NK� CD����c��8{��� ��O��aV�t�<�ʳ�~}Йw���s;�Dq�׌��c	�dC���OA�M��������]�4���]@�-s�W���x��@'I�.K�!(��O���d��*����U�O=�l�8�� ��J�Va�HhG�Z��2�{�x�%��)�F��/���[�L𐒯�{"�Ż!�K��"@��o����<W��m9��^��q�C1�n��"���m[#`XP�$p;/��@J��R�������'�0��'�g�ؼL�n4�[,N�>c���Δ?Vp}�K���(�����-݋����/WIP�6�UI�٠�Lg9PE�#�5�u�����F��o�_�/�#r�:浂��Qb��#� z|����J��Jf�� ��o�pZ-1Q�B��Ϣ���ﺝ׌Z3��#<�����7��u�Q��}r�˫G Y�&�V4�K��kt绥��.7u�
,8����������/��y����⟼׳�n���:�RH/��V��ΠD���4b��M��@�d�s�|�h-&2�W�˨�h	G�R��X�p�5Q���dM-pb�i�ڲM�������t�r�K�g���#E��� ��
�VŴ���"�^D��_c�F��7����7�"�C�kbol8�����r_&�(3����+�x����H� �Q-��X�Ӟ��
�euQ�^�G'@,�ml�#0�$��у���k�(js���-ʹ�Ach�e�|�q�����d��#4p��<��G��p�zob���4�L,rgm�Ij^y���p0v�(_�{�2�]�A8X�'K�Á���5�����'��E�/�ƚ.n�mK��<s9�Lc��?K&DlŢ$
eh�:D}����64���05�q�%��i��8�ٴ+�JM���]r�̍��Qz֙{�_S�Yq�J�H�s��W2���o��h��� �I����^4Z`A�պe���7�t�x�DT�09<��礤ݳ������V���R�� �W&�S�ٚ:G�,"��s�F�e<��OjM����k,K�~�}$�b�/��5�wCƍ�u
l��>_N�o˺~2����;�z�G��~�1��t�zi��1�f�c�pg�K�� �}o�zv�W��Ё��yt���̷�9+�;tW)4�=�RGǤ�<.�@���[�U��g��<�\�c�s�^�e��jVe[�$�y�낾xp:X�TV!��l�� mX�b�� R�T�Wԛ��h�Ƶ��p���S��Y���@j�}���������_����5M
{����ŉݦ�9�-�lpP���_ɑ��ɫ���S�l'���m�FģEv�^��}�]͑�������@[m%=�X�k/2L��8�����U*��+���\WM`/�!G���b�q	(x&�h�y�N}�(P�ͤ�6A��l�bdΉ����tj�b���R�GR�K��	�ĺ������D�^�W�i��
�mu�򣆨�t.���Be����2�Tu�����h��x,����O�?�)j5���q��sA	̎ʫ�Ժo�b��ke�v��䭴Jt� .Hd� �詏���o)&9������|s�>�6\�.t}}��t�[�9U-Td�,��"���<;����\��][�}�5��l� �l��CBB#��e���:J��8���6��(�w�(�GV=N�8əy��»t�8�\QWLq���'�d
o��%�v1�� \������\�vch�U�*�*s�{Px�����I����M�H����d?�������KT�	$x#��ü��P��K�^4���mP��P^��$��1�4(�xiq���VA�B>R҆%�RDS��e�5�g�l��5��$�t����7XD��p��?�q*�6c"�Θ�-�����\��l�D�j^�>�Jx�0��s�7��+��D�!�;��-Ϯ�w������Hȣ_��Y�f�����"�5��+Ź��E4-�,�)���r�����4W4eael<j�Z��c`]��j��d�NJ���F|5��Sg�ZI`���0Z<��j��:{�;��ؒQ�4����w}[$՛i�^۩Mg�(���E'!��a"ds�ŃvO���yJ�Q3K�04t	w�|�������6ﳲ��o���@w��/Ws�v��K�"�P�/@�F&)l)�߶��U�|!�Z:ƫ?�T��V�b�P6:�=�נ�FkA���t!x�h<�ה�-\�S�3b�%�L���#E�Qm��r��)XS�����xp�J��<���w:!<`�"e����ؔ���"�4��I�:\�ģ&��ζ����᪽<��`�ʖ�rkW��V`3@L�ׅ��{����PfH��U���{���@�_݇���e�Dy�/�<���_���C�p��?R��RP�]�0�9�r����5<�1g��Ҩ��_�a
���ZV����e�r��t�X�O��i��F@Y�=bD�hj�G�#u��0ꖺ(�T�<���*Z}��#�/m���������|iM���F٣P~v�� �qx��We�Fr�l{;g/K�'�U߀�yzvF�2�r( 	�S���2k
n݂@/9O���Ύ�T���;�zSe��&����!RV����A��uV8 <�V��a�0)G"v����u%�u����az����,���}�q���&}|��}R�23��lN<���~���q���d�����^�yK,UwՓ�l� ���\ޘ݋���l0h���d���(zx��� ���ڣ�e�ɣ���J[`�!�C!.���g�=l9C���,%��Y�zU���Z���F&��{�'���FND�f@k7C Є�ȭ�h���.	r�xA���F��g�O�1ROP�߭gGvF�������#���s�P�MU�Q��S���`�B `�z~�
@�(�	'�:�ە�ل؊m$��0A��*�L����3^��v.l�Sf�)��q�;�n<i����������W�H��Dtz��
�W���/��e��PΩs��||�+��}� .����[�4�j��N?q�ݕ|U��Z��e��
0-�A��,!3n�|�y,XǄ)�vq0m�n���5��zU2`�
&�8�c"RjO�a�7�$08Fe���>Q�D���֬i�߰J��׈̤���=A�8�~N��4���:��b��1���Is��r,v��%d���}��-L�u��%���S�ǽ��@��?�ঘ<�t��fςgG)}2��]���� �uH�����/v���`�:g����o�_� �̯�>0F�m.�3��5����K�O��v`kY�j��k�V�mWK�1�,"�����$͙�7�83��9�����Rd�"9�'ph9��^JP�+��՞�%l�:����d�E����y<��V�zY]8����̘cE^��;n࢑�����An���)��,�Gpz�TE�����`e ������zK��0ʾ
jd�Q�Ȁ�/�3�[�hG������/z���R�$��K���2W2�㑰���~�h�dzH�������w/8����Q�-�Հq���䶈��n�ڏ���/_J>�
�ip *v�[|ܩ�N
�;vm��Z2۷H����l��rW�EN����� jm��B&�&{mGXGא�;�ԩ{$�2S��倮�͖H�mC����T^ю-��pA|�?ލh(�6����\X����˦6?�|���
f����#h��N^5�F���=�F��t�+�錴"�����0�8Il~�9Z�jS¢z'�φ�lEKS")�����.:�1�_V4&"R��~
L:�����O���^��s����� h�M������>�/w�i�_�����(�8��� �y�6�-��� ���puR5��ii/����>:��lt��M��}S�FR�V	?��y ~3����3�2��J���qa�Zu�L�0	ް5٪9x�!]�~q*�!RĻ��_�rlQ������]�kgD�vʠ[���lt3��@�A��c� K~%a�Q�Y$�F��z"RT��6���c[`y�}yB���QC�����'��lcc�k�Xb%r��F.�ߢ�<zZ*UW
e�U��"����N�P�GTݩ��H�V�����y9� ��ΟVA�~(>(bW�÷��A5��k�n..��n��	��q�����lZ���r�m,�G�����UW�F����騹�0܅VC�Hp�Q'EN�h��.oJK^�z���Q���;5��`>g�]#[�N��~���ng���,{;���U���d8���Q��:d^Ԫ۝\�l�ZD��!�8��i�Z�������DL��5��-1P��Mİ=�Ih�tЍ շ	���}x���\��+|����BN}�������$a�'���1Պ�I���Y�Ĉ@�K.YkH�(��z'@1�
�m�������LQ�MS��{"�L丼-��B�# �f��K���5u\H�a���d��֦�l�d#͵>A<�*�˺V�|M(�%:S����饻��9H���?�bU�Ϫ�(��E�B��g�$Շ����Y�|&),z0�������Q�1�k����+�+��x�
'�y��Ky��l<�-w(��7i(�f��z��=���M��z��	�Xd�9q�R"�4�n�xw��)Ւ��扰�g(q+b�M�^�i����cn�↬���ph��MYVx+�P����u����Y'X��R���ޡ�zHr&z���UW��k
5L���~�!\�$x�9$T���w���iq K�C��s<�yz�6	��F���M��8���9P�Hq�G`&&V��=Өb�>�� �� �@�L>b�q63�-� �=!�V�d&`�G�U�� �m-!��m
��^�6���O�Ņ�9E�=��[�N��p�$���!�R*��%���6<�Ԡ��-s]�K�I��5 `f���AY}Q$4Ŀ�x?:�r�^1փ_�G�BЉ�	�4�TS0��=�Th��� c��
�Y�U#�k����
.�����xf�K:O|����}�����,'�&�N�b����J�����ܒu��=&7*tDAt+�C�DU63���������e�M5�¯��Z�.���-HT�����_��p�iZ�dҍ|���l�Gg�ɛe�/}FP�>F�%ɶTG��#h�F��q�SMdw�j��h"�?�������S��G�/5®+�V�
��a��`��7:�����Y���z<��p�0�X"R �bl~A}�L�C{:_f��͞&�C�w�M�&��
�*��<�~��,K�5Ю�D�~�f��iuF鯝���l�yg�Ϸ�]b��81�cp8o���e��W����d5�d����-�l���z�=�0�����,�OR��f3��f�[h*�g�[ԯ����H�N>='l�~��}���kHtn��v��@�)�Q�����/Ȥ=����8���nE�3p�RB��BK��G9��>@��ů�Yr��E��I���*-u��Za�?w��D&�~�4ul���� ��?X��lr�Z�+C=�#z�T��Mw��a���^����|��ˈ�$��$�����'>b}�Rv�Q�:<ė��f���["�~���#]�c�C)a�-U@g�t!9�O(�v4��P��~9j���k|�qN᨜.�8 ��*��@(�ы���V���A�;F�V�E�[Ms�fB9ϰ�0:Lo'�w ����|�$j�&�YB�k����V���O��NЬ�eF�����M���c��&�ɭ-�F'�KF�x��s��-#����̒e���݌yӫ����z:Q�m�w��f�mRH�o�N?b����yؼ���Ƿ�H��S3�ڻ񠴊�y�I��]���$��"2��!��>6:{����38 Z��G�!�I��R.p�%Q�)�_{���CZ�~f����w ���uݪЪ����y����xzn5x�FFE"ڽ��`
���|��Z_*yLPJ��ǧ =ۙ���#V�(>�e�\U5�E_|��۫WPObb�S�����������N3�@�<s��:���۝+��7>�W�
z���R�I��IYax�C�+7򭧨����eR�ۍK1��k�k&�E:��LL�Q���S?A�G�3e4˟m�~N�^�ob�� aE��A�*�A�N��(Z��������4#��]��Lܭ��?K��L���V�yeL&�O�+&�VdWTں�/#��l��֯h���w	����-u��[�>B��l��Z����utp2H�tv|���cp?��Z�z7m���)>�wJ���G�41
��9��;��r��Ia�X("U��@,���V�c�وA:���7��k�E����I��]�n�\�;�4��//wN��k�ۨmgIg�3�솀�٦���Y��-c�pw2�_��s	��8z6����R9rnŊ��}��z�&I��Sɩ}��oSO�@�3Xl㢠���{��ۥ�n��d9~�(���ɘ�dN�z���\ɦ��jY��s�-�cb��� �����fn��BĀ*�3~cǗ�R"�����m ;#ڱ"2����˨�KD�}X�/�U"ax��sb1�K\�����D��I�nPt��hx%+�ċ	�)N,U3PZ�Qf2�,_X~J�WE�KVh�+�ymd4DI�;���~P(���!�;��d��s�h���A#���nĉ�r�݃�Ĩ��rL�V|�����z*�
�Jv��X��e^3ӡ�n���k����k>�Ri��N���RF�O���N)Y�611L�����f>�<�]�%6q��nC�t������Ba��Y�������^u��^E�oy����F����.DP���nM�6��f.�*��]��C�p����X��ZB���b�V(0�F�Q�v��7�w��^pפe��b�\r���	hRt�ʁ�G���1���� V����x��yǫ���K��lRP��U]��ib[~ﱑ�+��E�z|�(�,U��e_PVV��yH���~!*嶶����+,N-�K�4J����V�r�Bv�mݙ_	\#z�/p�N��oWtk � �:� ��"��J�K�7Ly�n�ۥ�@X.`5�ӟ�3F�X^u"qB<�
ښH�#&�p�ւMD7f¦���1}�o2��\�a�W��v�%y|�X�uX�z�2�ej������.��5*5f�ܞb�H�8=�R.g�?��B�F�In����GJ�@����g�N?����(�X0�\]�`�*-��O�Q.9\���;�U���fR��|�-8(�Xw�U�M�!Qޚ��Z����@+�� ׳�Ӫl��͂~�0����Q�v��M��ʭ����ힱZ��H�n��p��%2�ƀ�AZ���ʯ�{��zQ"!d=]�*=ami���	i���޿N�����8�����~��a���P���t>���9Q�����5�4����9�I <��\Am%�h�8����D8<B�K�nb���b��ŃЪ@���/:|��ѽ�Z>���������QqL�"�p�ik �>�?[�����ݷ��`}�	]��62��8�Y�ō�T�o�T~,e�ZзqèD��7%C@x�۸CI�m�wrչ�E�������v��ݣ%�RϬ��Ԥ���ѕ�tЫ�ס`"�Aw�1��� 컐h��-M�Xb��bN���}�z�k�/ns��k;H�nm��iNch
�N�w/���l7e͖kԉY��	���@��R��\"�����ٌ4��
|؛�#��.���{�uGB�C�O���Ѓ�����[�����,K��.�?�;��C��24i�_��$ g��$4Į�W;+�����И��|���/"������Ʈ�pvs ���=�:�G$w�V5+
�k�r/�a�����p�6���j�%�f��ң]A%��?�%9Ƶ.@.rl���Ŧ�4����Z����h;�;%Z����.��o|�9]����d��n)��\L�`b�i��6�Z����U���g�SR�`��\����"��O��+�S��c{��;�nD9���������F�����~�j"�G�r��P��i<-B?���L|���\��A$'� sp�����g�^�5��CO�"3�3+?���'T|Dac��Nr]��G�r5(���j>j���^N��+Tb�T�q��)��Q�h��&�{��x��?@
b�J��J��}T��Ç��7H��N;gH�"Vc��9�xCt,�ks)1�&<"3���j��M�~�L8�Z*���K��Ŀo����2�J��"�ޡA�Z�h��'�jfPH�Mu]4~�,�����
� T;�V٣���H�76
�5.а�;��fP:�n'��g�zgw۟���C���Kaq@\L���M��į�(��"ň��8��^-,# �O7>.��K�z�>p/4��,�r["��g�Q�3$v�#���$���E6�����7��UD�Qg�&�x��$�	�v�����.	�������`]� �E�m�0�VIs�V {j1�ӲЉ?���v�4�s���j�Ep�m�3e���E�=�z(��ښ]�cӀ�)�Kx�xc7M�|T�!��f���m0��pW�H��պ1[��}���6�Cj���_ Y�y��i�����G��-(��է�.�酮�#q�:�����d?I�x/��:GP��)�`-���e�AvʆE�߭)�h��g.��o�"�2;�{I���\���?R<���wi�~j3F<���-&���1ڲ�B!���q\F,
��'f�#[V���YE^�$� ��o�U�B2sl��( �e���_��ۼ�e�P�qӾ���3%�K��#�������5�q&W�����a���)#<��*Q�L� z�{�3�������'��<���w-��ߙ���jc���K���9�"�j���7{F���sw�K�<ƯXA�anL)#��>*���PP]Vա��9�Y��)�h]�s<$Lu�p��I$eY��w�A��N�m�3�����nS2��\�/Ąt�AJ��b>�(��%$���m���V�)����ZŅ��HꇑsЭ�T \�����^�D���pd�Q�"�Ȅ��h;O�9uƨ�9�k3��7Tq�u׹�GjlP���/��o�~ ȫ���:2�ɨU7=��!�� �A[],��F��ǼvV��,ԿZp��Ƭ��\��xx�5���9#ݟ�{a��P�&k,E��AA���D �V�l��)���.�JpQVso�w�9���槲�o�D"Glf�����^�d�Q`kV�G��6E�@���li��
[��"��_)�<��Q�j��Q��07�`�*��(\�����j�z����7�x��pg����z�)э����w�u
����#	9�c�@bF'Ttqά]8q�&�����5f�E:��_��Y�䘵|%eQ.L�^ܔ ���g{MN�=6�G`Eqh����=�="<�x�x���L� }y�Dv�Ě�\���\)��
-��:n3O${&b#��* Wr�r�ɋ���-�ډ��Yb�OtsJX^����Y���=�i�6���� ����+�8r�wQ���#ƴ�KE�V$p�?�x�\�A�)Z�Y�w+5�d5��[GD�e��v��%g�u�<�?���9gÝ����4~���*�q��4�[	��K�:�n]z�gxWc�na�/����"釱^z2�v����� B��Ūx�SڹA�խ�.yxHo����������������N����9?:#]�fw�ey3�{��]:�aaOIS<q�"�_x��Q��vuE��
 !��9��a����;u�?]�6T����sV4�U�Z������)U��y�5�_@ ʻ��=�&[�NpZ��Q�:��
��|�>����f�O�����F/����pvd�I���@k7���+$p���I��?�S"�[�r�QHD#=�䡴��t{~[��	�A�۷��Bߋ���-p�xܔ���_5�E2�^c]K[�Cv� �z(�VƱױ�Գ�~�k�~�$�x��'I_Eg�!����92��R�i���f�q�gG^�֤3j�k��p��H�� ����憑����=~�c|7�c���7~5�[�@�;%��\(k�j�V.We��X<}��v鱑��;��iq����g����WjJ|ϫ9mɢ���*Ʌ����{*��-j�~���u*z�7�G���R�^r�4ƾ��sܭK�s>��(�V�"*�{����g�?~1�^obja+(#2ZVm=��J4���(}�0IZn2V����	"�W�Z��F�ʢ0ʭԆK�8-�[p�ۗE��
4��%���
����y�jQx��IB
V�	�F����2�:e� ��.���d^}��~a�}F4V��?�~HI�Bq�I|8�	<s�/�X�{r� C�Z�4�J��ڼO"�"�Eg�SB�+F�^:M�ގe�nHQ=Y�ZIiY�Y/�4��S[	��t�E��&F�y�γh�LI� 
@T �?aQP27�R���$����ќԦw��� �[ANWv��mQ�!�Ú�R�a��z+WKS,3-�Ͽ��S#8�:0
�'� �H�]����Qs`��FE��}<���r>��=@��;�z@YOH�K-�/�ÿ s�n=���� ��8~��3��u�_d��Z��U0�����z뇰w[�QZ�
���@����'�n�#�A���X�A�E��o��	�j�#Q��95:�#��
�G�ڱ�
�=eӶ�,u}a���ƪ��U>;A1��`����K6��y{yt"�1o��L�fF��<R"�tJrr8��F��)06t��2�Y����A]'�'"��ZhC*������2u!g+KK�և\����A��W]i��:���nE���4�\��QpkU�ޭAy|�A�R��	?�l�#�^�J�q+x+jc�� �����.Q�ױL_��v�MF���bo�U�\� �cC��Z樃T��i��܀R�;����kq����ܳ��בDgb����T�ۦ��{?
O�Y��+�@�cy�	 U�z	ۗW��i���^���4�ۆ�T0/5Ɍ����n�!WP�61�Y�]�v�Z� ٔD��ִ�-������f�?��E�'`:t'�( �m� Cå�RR�8�m���{�7;)yQ�׷6*���۔�؇C2ZdT\Ah~��7�^�,0I�O�b��^9��$  �Ճ.?{�o!�_�춉}Y��>�5	�N�9�f�P�� X�>@nW ��w?�᧷����#t<��W@ �h��X��{wgt2���(n�I2�5�R�X։A�3f�J7�R����Q'�=A?�c��g��)okؿ�cꈆ ��.����mz-=i���_lrx�`Z���+�ůqȞ�1�v���D�s_��J�b� c2�5���gF@�vW��jO�	���f����c؎���Deqdg
L�/�	�M(W/��,��&V��J�w�T�[k�Pr�
ׅ��4t��KT����]i����
�mb^r�F�,�9�ZS[��9��ԃ �&�<v.~��#�_�3�xu���m�U�"T3� N�`p3	��שt1�ߙ�ꭀ��_�=��4�لR���;��L����[;���ZH�ZW�D����yu�c��b�wH�Ci4
06P_�=b��}h�C�jѵ(��3�A�X�91��|��u_����`�	�Em�K��	߳���@1f�ܐ�]\phhNw"����q ���ַ�X�֓���ҙM7���\�x�p�$3�n]�U����ƚ�=�{d����M߳z�{�I �2@�>yu�N�!T1��h�{�����oyd����d�2"أeX^ҋ��ƽ90ˠ��":{���t���U��XhT�V��nIdҢ73L�U�?E4Z^�i�Z�?�Iп�C|�w(
%��!K�|v���)��F��>�MT:�\��-IZ�%T%��t}��Q����UCep`��Y,�(��7P8�.i !�S&�~��@����#��!u�R*)��:��f�	�~,�݅̾�jr�p����Cr���]I�a�XՔ��mR��9�<M��:=��j�m7��@���CT$�����mvd�M�x��H���K>�Du��Io3��v[�A/<���vT�{L��E:�������p��}ˉ�̓:@g��ǉ:5S�����Q�����OԶJ*Nz�o֞u^AR�}���:�I��DvL��mi�h*�!�8�_@��m[gh`���$�.:�������f���h��S�c&�nw0�@���N�)��0����9!#���7м=�D9HǠN�;�P�A(��=,'�k�r�c���Yz�����Y%�YQS�ܪHr��֜z �O�u��q���Z��6�Py�ʈ�pՁ�_/&&�n��cc+�E%�&7㮀����7d����`����.f����1s+$����k��n�aG��Y0�D�ɛ�Y>M~����H�F�3F�q+��6�%ޡ�},����
q�Ő.K�^`�)e���SX��s�i�7m�q �6k�kz�ͅA#�xw|T`9(TU��P��\�Q[�����P��b�Ȓ�\O.����0����z��p|L-�B|����7��~��62L��3�S�
�b�$[��H�x��z;��G9�PG�����7�O"�'���!�C ��,�͜z}T;��eo�?ˎ�s��7b^��Ff6��-U�Q_D�q��1�$۸��t\�����H��ɿ��'�˞���Z6�Jm��{^�e��q�1��!/n�4G5������Щh�|n�5C���t%4��ryam9^Y�:?Q��$����b��;Di��d	h�^b�>���Ib7]���� �H���ɝ(pR|��]U7t>�|"�W}#�EC������F�����W����3y�ƙ
�C����W�6~��]yj����u�c����!9^2��BCk�д�9�a��Q�O���`o@� �g��-���m��ܨ�1�R����s�sR:�t�?<Vx���&���B*;��;d��U��U��[��A4�q�"��jT�c�6<����Q�X�K9ZQ�)/j#q��¾�diT۾��_-?�7x���|D��� �������n�ә�Y.PҪ�pU���5���Ȕ8#da�n��Vh��r�	� �v�u]Ά�#�:P�ROƈ�!��P{��1�FÑ!��J�Pݮ��m����⟜����](�.�]k���(H�K%��\����A��"]ߥ��~����oӈ�W.j�̗<���Q	����f;q��q�f��U�1Ѕ.���+��v����Фd���fqr���ee��8g<=��XP� V��zt���V�W�2]��@q�ڊ;�  KR�,��'���I���@H�Q��b�R
�7�A�ގLR��RS_����#}�{�6��cWޕ�+��8���zd4�$c��53�X]s����uI(��Lݞ�<tq�cѢ�.pJ� ODIEf<)��H8"0>މ����Ei���MCP�%	���B��j(E�l�W�sb�JB�2�]c2����ug�����y��t�b}^���%���0Ϲ��f���0Y(�4�����4�k���h�j���@�'�!Mb>+䊧�!(�v��$_l!���J���`��"�)�Ǹ��of�&��s������<���-�G�7痶-���`_� �K��s6����
�|���'��+UN��5�b�Ѫ����F������U���Ra�I��h2S[`39Jq����)�(�OΏ`�h�O)�̧KM�kK%y *��ˌ��-������܇�Đ��D��G���g>Z��KVH��tP�u@�e��my�J$aj ��JJ ��uj��W�����v���LH{R7���q�� �o~D��Q��D̓�=#�&�D�q�s}�/��5�������oUT�ϸ*s�"�1�AD�x ��"�Mr�ս��<���!�ٟD<�}�E�_H���ud�0����`��,�Ib8�4�wf�Bpb�R^�#�F��t��x���*����N��[�j��CzLs������I-��{̻�IЫX�f��.��B�
hS�Fg��`(�xds����"��)i������9W�M����J�c�yw�jX2��Ď�fFqUr�k�6��)�:Br5V$K��<��(.:�,�w)��Qܵ��Sz�M܇R���@�I�B`���g��)����>A�����8�
6?y������/8$�9	���x	s/�@��;Q�(� �2���_��䈩��n~�����=��b��\P��d"y��"%������ps2E�XV�q ���A���/�s/��&�=fG�`��w��27G���	(Us�r���z�$���g��,\o�XȦ�"��>x6�7'y�:�NK6����SJ�Ǣ<B�t�����s����P?$�&
��*�u�mɱ�)��lx4���S�gBF�3��>F1G��B�˪�W�܋���0��fŤ���v>���|���#�24����5q����H:U>x诘w�Z]��\�顟�BϹ���@/&�0SF�z�ݭ�����7lve�`g��IZ�Ot3�t&E����$:����,4v��vI�G�|����(�ӗ��P�X��<(d�e�������n);Ȗ��9��
hSL
���=2�R��f�{	�_4�����hT������)�.�P�B}��������<�s0�E/S�N�։J#?޵	�5��_��"(l��yx1����J,~��&1�u���L�4�R���F'�G�ռ��W��Ƀ��ھI�C���'ٹ� <�a��u�� ��[{,�#a�r��,,���CR<d{y[��6��.ڽ*~�,�H��n$��l�V���&��d����q�Z�r�R�t�{�Pv$qZbA���w]5?P�2�;,��|1���?V�wif�*��;Y�ә�qw��4W�{Lq�sT8����	�����ƾ!�X��`n��*ݷu�ޏ�h�]=�es�S�Q	x��J�����Z6�"wW�i�e(5{������I��o>r���`�2p+zS*�3�*�b��t�U4z��$�Vw��f9�!jy��{T��.�z����n��8�����֛�Y�]�Q�/T;-5`4����'zcv��^_tp��� �C�&����X�?�z�\��ѾO��	�Qy�d��Ԭ�ǵ/'��13&IwQ���μ���jHen@���I���6�E��~vPE0��xuc�T\䜖�|�u
�*�z�)æ����lL��q�O3�e��~��9�"��E��/�H��?��d�x(��EL�m�f���zlGo�VH�G��?ý�f6��^�+�6!MG ��Y7|��ӎ#�7Fd\����;W�-����0�`�sq�ߜQ�jl����(�r�#��\�j�QV����g�y+����L��1�d;ʄ������B�������w��p����]��T�NC�N(�A]��w-�hg{R�2���-�G��τ?E�}��'�f)�QLf�[�A�%�KH�g���x.:��zw��F�}���M˨��`�)�sQ�U�'&ȉ���C��ђeZ��m~(�K�Ғ�g�"��Y���V�
����v��߃�� ��u���^�PVY�M��Z�j��7����n��&э��~N���a���!���I�����s��/r࣮5�u�(��\���`G!�$��?�q[�rܛ�3��V̬��'j���l�!#��ׇ�P�	=T�!���B�+�Jϖ_5��fzc6�v�e!����gl GS��߽����@�3m6�(P���Maj�H��1Cy�Ƕ�L��Z�`F5�೸�$D�Ԉ5���&���5�AИ:������	�%�쐮VR��aÀ��U��<���o"iڡ�M��)[�%��ȕ���k"ȇϗl������ʅ�:RwR ����w�Tr7����Mu�>���q����ڼc���h�����$��^�-3@����M��y��m*�x21��:�~��qr2��U���t ��@K� ��ue�G��<5��Q� ��܄Hi.1���C�c�u���
���[W8V�3�`ԂA ����RT�CD,8�x��S�ϥj@G""�j��/z�u�t�~l�=>ጳ3��������T����J��),p�sc'��ڦ���&{��~�j5R>`�h5��>L�@�U6߼�x'��1���$<7���I��4~މjj
��4�ņEC���%O9L!\��~�^��3��d��t���kE�~�O�K���N��I��&��l�Eһ2~rǻ��^��^{�dY��]=������|{8(s�S�تKB㏟UM����!�]��)ټ_cԅ�:�N��]�:*�\N���%��PŲ���W�U�|5p��p���Ȗ����3��x���
e;��E�c��՘8�`�M���#:�e�Ӛ��g�>݇ |MBY����8	vJ��d�较z���9��B��^�]^�\pʛ>9��Tj��>��������CX��n��jq����W�X����0����H��[�PX���"�~��m~��n�J�d�G���t�o�0B��Tw^�Zmܐ�eS���!i&z7�@��&1h�MCC5��?��u`��!�+ێ��7��8�B��V�2��F (A@F��y$,�]~8�þ��,��Lx\ìUP�SH틽G�|
��Ů�*g;�ڰ�P{<Q����ef��]�7�on��#���t�d�/�q:ºV��h��jˇoŖ#{�N���#|z}!zP<^��/a~<,�%F���Z���j�3)w �Y�B�J�4�k�9�N{+*.lڄ�|>Mdb{5�MN�с�����BPH'�)vE�`�5`x͹������vg����"�rw�Ԓ=�����;[m��𵮼�<�i��Hk
`������z��͵bے_ܸ��َ��w*��$نy�n2 �7c����Ran$_�"�TP�8��������gV�Y��YQ��}�K�n����������R�!F�ĩ#�:�SY؀&A���ܹ�/���O!�Y�{�Z9/%����
�& P�Ʌ��8n�ϮC�z)Y������	]�w�J������f�#�
��bW��E��d�(E&�XwD��ݦ)8>���Dr�(�j�-Zx�����#�Qр��h��H]��z��)(��	��������3��ȳ7�=��ٹ1�(��.;�3e-��|���5��{)�������k�w
�Wy�31���<�-��>��,`��!��}�sL�.�����3Sr�J�i�!����
L^f���Cڰ&	U8a�����B �YX��ª9�ۢ-�P)sM����;����t�$�	m8����P�m���J�q��wDyP���ql4�n�]Km9����D���`GR������4��Ƚ���L{�>�(nI?��]�g��j��&dY�lP�7v�n��r ���1Ѧ\�N�&4k�����<�`��-a��F�>�/4��P��8�?�B��;���Y����:�������6'@\���L��C������攚���aTXg����Q�eR��R�r������6��6��������?�`*���/�Ӧٗ���H��"w�������`�Zo'�N��[굱'Ps[��Z[�*���O�*�tߐ��/1 4����t���9l7��E7;�/���X{�3T�=X{�\-�����SPi	� �	bN.�%�3��2(B"�g�a�+��{����@@R���Oe�Έ�2K���?�h[u7��;����0N��?�ÿB� �;���;���CIƐ�o�R�
�
Κ���-�R4��|��'�L���	<ec�du�}����&�v�i*����-�"6:�}ZΚ�+��'�_�j�P@Y�&��N��>��x��_�z�2Sf����}A��o?�~����ǂl��n���Q@l�$����rBD�%4X�a�p�vsZR<x)y����C���&��a�xD�Yg�H9��7}a��q{�4p,���Ί�>SoL֪,��G۹c�
�{τ�h��H	Y��ؘ��t��jVro�M/@^�Ϫ.1����Ǜ)�{M�oYo�,C�%mq�$�K'��Y!>/��s�Q۸��7���2J�0��v͂�<.aM�Zd���&�%���M��$� ��8��kZo�E�+�6`��n�{-w�R��=gn����ҳU�7��q}�T��Ec�֎�v�q7s%�0/���fT����d���z�ٍK¾�b���B��RȨ��h���s����E�B�#�����a������Щ������03j�h�)���=�ތ���ĪMb��}qʷ#53<0 Φ��I���=ξ^W��V��D����� Fܡ8$��13(�`�)�A;� ����9S}�\b��+���U��ʫ�.i�+��d� sV�T�A�Jz�F`0���d�� :�A�Tz��Z�����qr�(��.b��y(������`H���p�K/�7��(|%S���p �>�����Z�n;w%1�֛C"��a�O�6���p��3�x�&1�=��9SQ���ә�y���%���2��s������I�qB��Ki���<1}-ry^�>f��}�������| � {�i�|��b&��}�;4c���i���ib#w1�[���
G��q2w�����GdH�,Mw�ȝ��4�e9�J^�������"L�F����o�/�)� 
��F��G�K�8�bRTam�7�K˨�@����4_����:��T�����I-t�P��=����g�+�`>��-��i�p%Eh��	�|%e�e��)�k0`���?K�6!J��Kko��x�Ӎx1���]&ZQ�{@�I˕J��UlR�GX#޸��]v�v�ٴ�u�H�ZB'h�pJ��Z`Y�K�ぞ�f�L6�=3���ލ{�A�6���d\ES���n��h�#D2���%�#��:��%��2}�A@��<hTw�
�_s�篛,���>��x�\eR��T��Av�7lԬ��R��3�=�2����zB��m�T�����w�4�ՁS����)c�~���M�x�������s���P�8��`�5CK�s���.+~ֲI�`�G(|��0n`��S+�s�o�[@���ǰ��, n:����B�	��t���B�{���|R#h��١�ՈP�����`B��5ŗ�Q׵�ſ�6~�.^��GD;�x��_���	F��on�s�#��_��S{N����/uZ��F������BZћ���U��>��< TT�b��B��Uwp�:��Jm!�(v���^�<[�ĩ�0���].C�ى^%��}�bdP�'�Ĩ���9��iX���Ya����P�0��3�K�G�}�w��$����@���w��'42�²����k7�/!eB�P�v�S�����Oš�|C���K���2	���;��dȸ]:��(���  ���SYuwj�\��A� `���$�J���(|������^�QU��Al�ˏȑ����%;5N��	��AӅ�Z���
��N~�j�������eh�z�ξ�8v��I >��80�VbL��G�/h:�ۺ�K�5$��0�]���<w�B]�r֧ԙˆT �����QW�O�Y5��>��>�l�bE�s�n��&�SG��R�s�ŝF������ED�=]R.�X�|��)��(��OU.��jj�#l���#vK['��=��	�3Y��bpՀ�a��̡�j-kh�A
� �J�b�I5�g��z%�Yf�U��%η��Ƃeb���|jY�����$����TD{Zh���!��Ra��"��ʚ�xh���e��
�?*�|�E�B�*���|.�UZ��9�jHK��&؁�>�ȘS�=$������U�8J������|��<#HpF>�Ɖ�ˤ�]����;�\Y��\��$���(��'�F���aաK]Y��p5n��̯;���WA�D���}�:j�F	j�\�d+���IG=�)]���y��A�i(2^�
�N�|�;��yL]��"k�4&q�,JӸS��7$��(l���I�Z��E�[z��p%��u<�wʹ�ț��rKoy�
�}W�&$�rS.�9�0>�ٱ�tֹ_T^E�~�0�q�ⱂR<�FN��x?nC�LL��\ 
aE��QӸ��^�G\,u��[o�;1*0��E�=)���(+���(hq2.�dbv|��:-�Km�(�6���+�$\aH�?Ǯ!c�{^��Fj  ɧ4=�b@kLl*h_љ�3:��'�4nN�5� ���n���^~?��f�`�Kn�R	�-Ce��8/�, qu���N%��_�hb��2|��1�S�"����C�hp4(���o,�r^��fm�'s�)�<+�^���iR#nK��6,������~�FHyI?���+a��SE�h�E�f�v��u���_\q��cQ��	U%�֒�z+����|�t�IF>��SgW�*d� .^p�q�2�,V� ���=U�D�&��OSM���	���3�(�bP�B��GNY65�|�� ���y6�m:�IP+2�ߑ�E�wx���6��Q�.:�ǤV��VU�ghB c �|�t;/��wyR~ps��OU����
���S�s�����G���{����N�^:	�*�ta�����q�>$?x A/7��l��t�n���������U�Ǵ�O�\Eӌ�����B��ڹC<�Q|�^����ch&��Vx��N�]&dcP0�H���m�Wa�؃��F/�E�m��ƺn�_T/`1�>Ʊ �-�0<�ծz��m�z���<�dW�c^���.��
l]	�w���Z�hOI�F�o� ����q��x��c�Z��%�r�M���c�|��|�	'��[30�Z��KԄ�������J��QrF{)F��f�^@�~:�{9^�&*&������3�D��uER�	����V�8gBΎב��ڹ����g��)�co�/��O�? �9�.e��wdv�H���g�i��y��\��Ċ�����q7î��˚��v���~c\�p�����|���d�wpO�pto�G�[��@�:������m�(5��o �d����E0��n�"Y۵{�l��O��2\����g�(��q�b�3���7G��q-J����e��yWk���E(ϼ�J+�w%= �����P=�~0�
d���\�=�����yp�*'��,ȨdR�Z#]�^Km'.2�6(���;t�J�i�+@Փ��S�.V�:29��c�O�Ez�"�F�$��TYsy�d	d`~�^(s��dqGl��(��#M��{c��r��N��q�C�5�蜕��K�t������[B��3�1��ř���,j���� �X�X0#j�q�;���K�92��u(7s2��w�[���=�����g��JZ��uF�%�K8���D��G�$"�v��v�))X��i2H��XF;+vױ��q#O�D���|H}�.!GJ`8yy�Rd��b����ϩ���ad��1ԖH�������r��ѷ��6��:FxRROHƂ���,�_(�4z�<�5����`�.�j�Sfi��z��|��]/\���C�	Ɏ�
t�E�{�; R�f�Ix0�ym�z���:��j�yZ�?��&��q<� #Ԉ]Y���Ql׿?��P�Ol�-�	S����q��0��I[��H� KqA��Ú"E���=V	�ыVy��R@HK��-=�m�g,��챗s���Ǡ���군6á��(U�r}�h��j�X~R��>��|H����cMr��^I�o���`�?E�Ĕ�����	�v���|E�b`'��($څ��G�Q��p��s�x�~������9�@@��Kɀ��hf&<���	����%�X��]��s���o�y|~���i�h�0J��Le<��b�InN��Q&�E9b��'Q�C�E˼r�q[SSg��ۢ�3ԪC]����?��;���u�7�jٸ/"��p�:d��\-lA��AuĘB��<��U!�M�r+ӻR��:4�"nv�=�`�r�
��QUj5�.���k�A�9�����|��7�9��������L�dazʢ;g��梯�gNF���.3�=
��\�2����I<Є�����Д�U��ΐ3����Q�g��NO$	�y��sc�yTa�jWh�ЍVV��8d�F�ˑ�뤴����Y�p�G��� ���ct:�"���J�7��t���ڵ��B=GZ���n[+��'�n��Su�'�?ߏ�I�n�M�=96����镢B�U%��Ͱ�6+!'��v0
�d�:�}�������zT\��]\��9�u,^��B���jc/oz��=�l'D�=�5c_�n�i�����K�tT)j�dE�F���4��D+Kae;U���q�����&,E��F���qy$�U���7��EuO��BNG>g�JM+U��-��,=Lu�$���Y��h8ZEh��߅�|c�w;�sl<���p���_�{r�m��[�#��I|��Bc��������i�~�4���xf|E��	Z���&�a��W�'��a?�Pb̷(@�7 �C7���z��Ϙ ��e/	�D���A�`��4AK����dŊ�<�Z�=�Xå�i8i�E���>1���DT��3�̒i�>��E����D �"�Si��P���B�O �W��u�C��_�T%�ѹ�ݞ��,�~�^0��\�A62��Y�����.�{p����&st��"�f����H
}��w�`@�`�z�0�I�tr�	27Z�1.|H�%{n��k;�x�-F���Ρ\���N���;꽊������Q���U{=�r�}Y�J?K枑%}��Si]�&Ό/���w�=��" <e.�k���A0�_W�W���񼸺�֚"JVSU��.b%��Y�Ʌ����e����ܽ'A)��.�J�u����M�Pj��}O��a��nhv6���a8G�BlW����g�D%�e�V�;_��5�ʼ|���ud~�Ђj�s�=_�-Ӽ=b�t�K��<�;Δ�6'�A��݊���B�P%I!����d��W�	�n����l�QlÑ�*Pc5O��KA�<	�r
]QDeD��x�������$��1K�u���;���|�)%�Ls�����N�؛CyI�&6�dnK�C;\>�%���������f��]�>�w'��\��<Ȫ^������@%3��闲n���,�)�e�Y�\�{���).���L5ZG֬���zl2��{�Ɵ(��o�ߨ} 맦�c'��2
�bQ��z��j�L>�!U��fRA��9M�"��8�_I;H��c|"�!H�8�����5��~�8�����$t��V�y�;mG��A5�=�"ǭ�S�:Fjٽ�+��H�hE���]�H�"��a�Y�F���dI����QʴT���'N����;�ϻ���,�����o-%�	�W��/���h`�{H��%�F�Yޒ���)^L/�ܥSt�N=��Ղ�Z;)��S�l�>n���qIw�H?�� P��t��D픮��ւ��]��O���(�\jB�E��м5���Lz��-ת�}�/�ǲ/��'���݁+������&�m�p�{0P�j4��t�ҶG���/A� �1^�?���8�D�U�v���?��8V���;�y~��}�;�K����D!|���]H����3l􉏎�9��?e��#��y����瑰PA�&�xGL�)x��oL���oQ�)�/1%iϼ����z�_���x�?Z�J|�9�Њ������5d��r���~=t��Y�Ab`�6\�����!ä��N�yӶ���>)(ӫ=���=�!�I�>Ӊ�v��9��0�t�y�0�Yih�P7`�Μ�5���*�'�[6Z(d�L�,�L���d9U�>sr��� mp�IM�.��:�߈�(�C�g_Q���?֖������Վ���Rֿ�灋�[j��	8�aCQB�4�$i�
�Z�}򠥟���CZ�Ӫ�~!��L�G\���t_ڼ']������/(UV�f ���n|R���E);��j �K�؝���9���9��;�i���u�w�H2g~�,������/�Z���p�uxX�g�<G��Ax��;8E�^�jO8S�Xm���Cմ٥��mkN"0¨0ԍ7�{�8Slǳ!���W�OCa�7U��.�pi�i4�,ג�U�HKyT&W� D�t�PI��YXN������XcCb�(���Z�^&��U���z��k�J�Q�e��=KL���D����Ս,�$d�1%����y_~����+����{sk)��@�g�GD��u~F�	�?�Q��#y��da��X �j��W~��EkVk�ݬF�-����@�gϋ1xQ�R/�A���?j�ʀ��Gn+��N���-̚3Ԗ�m�B�x�vz�&���7O�y�� ͜j刢M�]ꏁ�b�ꯅ,Y���<�ңA/[h8 v��9�����,�/�U�6�^�W�����E_-�F���������n ̓F�Ǆ�|���ad�\�>3.����<u{�M���=��>�����X��c�]�?	٨�˝��d"����������%��fM�w�~�%���\¦pȏ� �0���L�F�[�gAp��ڣ�ճ<�]��m����;������Qw�d��J��2S�D �{4<�>4 A�/�S��_O=��IZĩ��JTZ�dU����>تS��*�ダ��������E�-��<�3���ra;�J#���=��*�l �ʻ�b�AJ�F���&��ӹ]�g�Od����#`�}Y6 ��;
~t�~�.5��A�-ypW6w���չEM�6�1W��0����0��r7�\.
�II���^���������B�K���3᫳m��l��.g�Y�A"����ה/7���h}j+��*�~A����.P ��f���M4��.ɠTo�H/W��/���ȩ��M��s��L��X铹Xr���i�>����S�֏�@ֿLc��-�/y:K�����^��h!����J@4�T]�zv���/�-&G��^�K�+�!�\�rh�)a���xi��W/S������((<�*yy�sR2$����F!r��&�tlW�հ��k�����#�L��)X�P�\��7�n(�<����;�����}IB�iȴ0��P���QL����U�VK��?S��֨�xyn���￑F-���;V�]G K��U\�y�Z� �}]<�ߌa�0(R��1�
�R͔�����\ՠ�5�{����/����(�g��_
�/�Ĳ���t8>�@{a����u������7�_�.mG������8�d�	¸�$ �O/��y�a#E�yḨL�	�l�y�����)� �a= <�M��TBؒ�����T�'��q�yzXh���x=�ɪ���tV��H�Z� ��$�#	�UaM���3^V{0wHw.���U}_�<�ԇ�3)���Y{�;Т����^L�>F<��I��N�������ߟ��Iɇg} ���/�:����_'z�7y*��=xG��\L���-d�n�p��^~�n�&L��K��i��-�	�S�K)�^�{�mG���� aY�wS`f�q_Wu�*��#-B}��>x��m2����;oJs�drѬH�d�v�+M��:40�[t���3�wܩ��M�Hm2�@ˆ�!�U��/71����Q���m�qfx�u��{��d����)�T�f�£�	��9�M�G��	R�sʞ�W�5B�T@�.�*隆�������G���g؜�>G����/!���!�9�5�;/vV����)V�Z؁�k�G"F&r�}�E�$�����nD>��j#�+s�b����Kn;5�9A�
�tPϊ�[�'|X!L$�kǮӂ?䯢t�|- �)FMD�T�����I�������<�@@x���}k����*�z7oc.���w�#{��uSx������~��4�		رaf�ﵹ�3D;����o^�#>��~�'/����D������^A�)��R�ݻ�Ғ�w�u(Q|R�0��͒�1|��8�k'�p��,��~v�58��򠊷���_��Yj�7F*�'c�A�pK��*1o��烰L%��*K�9������������k�K�DM>���@TۜfcA�����踢�r�8o�%�<UR�s�Ϟ���#V�^��P�6���L�"كg����[�'9,G�	�e��g�__��<	U+Qt����,��-���J�� /�R0ft� a���;������>��^�y���k�-�و����s��Qh42���0v��ҀXW�|�9��s'�8]���`�l\�/c����Ң�zɯ�?�o�7*����KZ�N~��&��dAYn5��qg��e����.�.�Y�w/��Y�`�qb�\�!Y2��Np��,Ip�1G�Up���շ{�ώ.��^M�ʬ��i�/��H<�u�
'ߏ@m���(�u����h|�#[?��08��fӄ����VԜ�M� ,�dޠn��2A'�؃v0h�ΑǬ��v��+��E�3!m���w���RZz���������p���a}^}��r�������Mȧ�$H܉��*d��:!�q����qFrh��H��E��̪�E�ra��	�#'v�Pk�faX���XS� 
5��POkV����-ϯW�2�KD�Ft����Ǉ 4F>דᏼHY��hs��ŀ-���5���a�6���"w[���=b��l����s�}&k�WP���m��KU΁,�ٖG�P��סP�ா�I1�V��$�\X�m8Z+H�� h��;�oY��+h��"]:�2���T��F���k��C�����2K�my��|j�1��z:g�>Ƃa�mM`$:��o��Gp=���1A�M�1J(��̡�d�џ���z�G{�T���5<���TT�fC�nVP�b�r�JuO��4�̛w�(ACbFE�sK�#���`}B�	iz�'t�)�qi<����u�3�]q�A����ӹ.r67��������%*���m�%z��;g�%)[�F�V'��w��w�^�eC����ŗ�	J�jaq󒲺H�
X��
K����c�|�\��XLם��r��/Ol�V�6N�D�ŀ{yeg��O��x�@O�iR�&�擵�'M[���g1���u��9G����%�|�����O��TX��8_�g@h�h\��V2\�n����?��<y�-x�{1C�.Z)������_BJ��'�$w��l���QB�?h������t��!y���&�D�}w�g+!쐾	�C�"#�4��9�}�Ժ_ѡJdz��"� ���7��:c"D���V���=Վ��M5 1fX�hFEABT��b���O�v���fr;��a�h(G}��xw�9��/A�A��\�'q<�{ QX ʃ�� Xu_GE��/�1�Us{i��8���I��8��ᣡ�?S����`�G�����m�|�Q�����Vո��S�7L5Ft&�O�uݤF(��UpgI��W�{@�^>޳��( 2dZ�֣u�%�L� ���S�m��gIN �t�D�S�҂6�B˿M�k���x�=*�Ns�4��If1X}z��!y���M�~v&��J8�U��=T�_�^���?��T��20�w�G��������TŽ��r�N�em��mr��h:x����"hä�g�R��(�x�22aY����=��C�W�r��`?�g^>����_��'��=�v�pQ\*��� BBu�*h���bm��%N�|�|��{�{$L��>Ů�H�څ�� ���i�N+]��n�h�j�	8�%�ϻ�?�nѹ.�})P�C��CCy�7����H�{�y`���C�0�b��IA��	XH�,�Mıv���+�����X�"B�T����]χ�l���wu�%��e-�� ��|���[��>Hva�mC|�b�ft���6>�X��os#}Crh��K?j�=��+�yɄ��|�%sW#���|hb���mZ��P�&)�_������OMe�� ��⦎��k�i@J˹�C��;�U�Sxy���-�
�W�
�
3�rB��M0�4��L��@�iߘQ��y���5�w�e=ɨ\���R:ha����+i������u������k`�ڤ[n�uٳq���׎�?ٜsdRy���bwFqU7ꎒ�֕a[}ڸ����915�q�:�xIŷ�*[�8a��2��d�	P������r�M�:,D�������h�,����Fi���-�C���\M8E�f|o���4����GE��)��):D� �D�M�Ƥ���Z:��&SoTE0IR�s��"/}L�a�hZtehP���y�)�(��[�<�~�J\�jٙ+Y�p��$�"���šx�f9]&��Y��w|5��{TD��'z.����7?�ܤ+���?������&&��a�2�lt�h�k��ovv�� �~������߄]Z4y���A-8fg#�bD�R;�l�L:���t��(�A2�boM2��Hf�h�S �q	}Q�;�Q��`�meC��lanc�	�}������x��@��)� r��}6��͊�~�bf�)P2���^5�GT�(�Ӫ�%ܡ�<�`�^��S��8(BB+]��*�(�0�otrw�v�� Z�93��/������jj��Еi1$[>�a�t�<����%
�*F��I|,�B5Ė�xލ��_n��)]��Q���q�͸��uƳ�{7�� ��x�d#��J��C��^6�U�-XǪ��gu�0�����#����	�����p�5һ��.���F�͓�e��F�h��i��`���� ��/:P�����a���Σ����fH@,�<g����r/㏩����D���Ԣ�x�u��J���\`|<����] ׬�N��u$1�DưB7b�����0�N���>׏Y*o31��,���5~����MazQ�z�C,C�9 @�}&��8����6�ΏzH���/hc�`�<:H�K%�ʜ�$y䱳eK��O�f�6rIo�7�9f(&c"Bc;͢i�B��/ܮ�:;������qz�J���#{��L�+�w0�J���!�p��y�����V���#�׳{�j�˄1n'd2j'�7�!�b�C��Q��o���Λ0/��XpG$�р�pՐm���,/�~w;|�Y"�Q)���7��߇��d�;�Q⯓�(�/��P��m����4:�ե��hI(�'[ '����$	�#
���ax����C��(E�WVի����N(=���DQ���xI0��-��OD8xMa6�n������������4�+
��Y(����[L#� I� �����h�o�� |rV����O�h�bI��A������R�?p�qh8#�y�Юڅ�Wr�W+h�qd	h�s�<Eْ},�S��<�w�!�����d	
P��6���g����<���&�7m�����f��RU�,���q�̀e K��"��"�4��%��'�����r�)�?�̓I࿭��z��N�W���toʹ����6Gg�>g?4}S�.t�pד�J���Ь�#�Z�_1��{;�l��)"@C�Q5\0��D��9Dֶ�.���!������pP)$e�Gn�zN<��0O����3��>(�����E��Ct�Eh�6"ZN\�[�A�%���6�K��eB;�v;6�m�+�v�D�V����CK�MFK��Çs.Zx3|��H	�����R�5����yzo6�1��zr��☹}v]zT2Ed��<�-�HS��H���j�Ƌã�1�����5���V��Ub��R�q���_pr1g ���\�r�4R6ċw1ض��%�J�L/u��������h�a���f&�x�����nd��l*b����� ��)��S��F�ƅG٩���ݠ��S�6�j�&��F4�
+��\΍�0�	Ej�F���mAp��x#<�%z'��ņc�eI_�O5�"
	k^���������e���sc��&S�=�v�p@o'=6�};v#��$^^��	&m���ޞ�AM}w�p �l��l�h�33\�m���?>>�R��q�)��+������Eڥ5��R���I�lT�F��p\0�l%��No�_�KqGɿ���Q^}+7NW��+	�ʃ@��~X��������z&Op"���>���ƣ�����l a��r�"LS<'3����4u?q��HPZ�9�e��u��ѣw"�<�ƫ��ov�(�F��e�Ђ�N�l�7��e���Xf�*���bxg��q��T&�Lb��OQ���l����F�6����(I�-tF=?v ��E�blML$�v���-_s�u�:��k�o|	��|3���/cȒ`�@ZrS���4�	�h9g�j���w�K\���ӳ�Y��6K�+y�Qg�[�e�;�x�24LS>f'��ah+�����m�_.v��RG=��@BM��U��5e�U��������_��!u�LY�\���N�ߕ`G��ԯ�z�b6���o��v�����f~]&x/gu2ۅ����#�Y"�P��b���Ɋ��� k-C ���f:w^S�dp���.`�M�."?��m_f�v_)�E�?�v��ί>k$�i��O��_�]5G��^Z��=B~��1�u�W�o��pn{�74
����)�I�=e}�����Sb�f�_t�&l�&��o���eO�n��4��r��5��Ʀk�+j��$3��*��:����"�N�k`�(�&j�l<Ը�P�mA�N�kV�殛jE�M2,:��WNvf;ҙ][��`�'�Sb�w����)D���TD�J�༳y�dY]���[�?�gI3��0���.�L����P���k�R�8�Z�˝�j7�A�[F�m6%N�d|��zvbh��=�.�����1cKڣ��M�<�\�4�W�B��9/Y���qQ��#x����=����J��S�X���[M*���ȜO�o�;ő.��*єE���v�%���A.�3�hש}^.�Es�3�n6(��'a��bQ�ɡ�ś��V�TP�vʖ�>W搼E���.&Ѓf��EpX1��A�T�A�?�_5�Fn��X��K�i�����:��g���ќδ�v
$�*ْ�ľ
�ܼM�"-��83�����X��:2��XϘ��t��K���F�i��5��@�SW�6�p��9{T.'lLF[ �l.�Q��)1j�`��'�js�>gW�k���:����B◿t�*g[��X��ҹR7_|�\A�0�>T >0�k,�uթD9S�0y�"Lw��Lpj>��L%4��x4�W[��:���"��-oO)0&S��}�J�+6�z!�LH��%��8��a�x�!��eKڕ<�rzu���a�zj}�J �%kd�h����d�u�����\I��u[�<Q���A��<v���	��s�z�X.��g$Q�f�qP׸H�ƍ�I��Bm���>,�LU� ��ƥr�?��S$
��kMrmBXۤ�Q8�n$�DN>9ဿ�p����7E �x^a�hhYN(qL�F}��#�`YhG��0!��2�L8�ۿ�x�jV�0=�U0�y]��-͛�O�42�YiX��D4��9�7;�aΚp�kL?U�8�O��pvȕW��X#"6�I��K��\��X���%���1Q�8a�]��fpb�`��r:��CfC��f�J'��ণ7ߓy�2'��E�(�P�C��Јd>�
򂬑�1ٟy�E�B8Z�+n@[�G�sI�%H��a��6�*ú��k6L��.���\��d�+xz�P�5l'J�'~&WU&����c$ޞ7S ��@ktŉ��$3� ބV1e�w% _��y}̛��93Z�iN&=�k�.�E�ru��^t=+�T&.��(�Y'��(;N�$��QIY� U��D0�L�:���,;v�7������g]��v�+�W�5�-tϮ�/Tb�6詣}�|��H�Q+Rwd,��4��� }t&�`:�����-l����79�g�e���c��<h�Z2�䜷�׹3�=~�zA��B�~���[��C��������y���Y�{iߤ	�K��U�!8�SSN�6�/>��!�C�EK/�}�ӯ[�J�l`Y�X[ߕ���S*?p�x�o"�뱺N�F��ެ���ZD@@��6���������Y�=�-�hv ��мUB�(��p�T��#�-�q��W+��z��"���_F�t��6�G��P��t4e�O� !���ގ�x��SI����+ӈ����b/�e4����|��c�.�/ժ�_UUk�6��*�����|��q�#�#R��JK1*m���!k�;}�t; X.8�U�.l�G[�~��'�������W��&�����8�(��d���c˕�N��4������}d��V�nn;)x�����`�=e���5[ݨD���VA�Fchm�J.�]�=���%��W��Aȋ�l�lG��a*��PXR�����n��|c7x����^������L���{y��buo3*��n�����LW�]����WG!�iQ%Ӝ����I�.����r!3�t�f]�����V�vw�{��+�I��^ ?"�y����i��N�5
����g6��g��%Iþ��j���>�:v|��Ei�4�_'}}����<H�S��,�`gQ��:�S�ٟy�j�>�����]�<�K�mԲYf�}0�����]DAKɆ��緆>0%wfy+�}�7d���^Yy����*I�W���ǅ�R��r/j.��u�����	f��S=�ɰ�v�^�����*�ۑ�j�g��^�[f�HI� �ηG�5���L�8��Q [�a\C g_@+S��#4�H6�8%�k7r�{�p�|���u�8x�E���A�V��M�ٱmq�&S���	%�F�Rfڭ��V!����a˭M�`���)(U8۞� ��(�1ĭ�O��Gݒ7;w��C�kwV�J��>MD�0�A`>q��ؑr�+�1bۂ˚8�_Ƕ>�s8���r���'x2.�RMS�1Y�ĊWL�x�n�,9�m���ʓ_� Eh���>Du�R��	lIQ��w���ǒ���%�g���$v�/�Y'�BË3��x'�p�h�c�H�����n��y���T��ݱ�(�va���� J��x��٢XoЮ���S�h> �diƬݹG.rm �Ql�d�Sr����B;h^d�_�[����1Y�C`�aCHhکK�t�
��E�4�C��vsּ,`�p��N�Cq�D5�~����)Y��r;Y]��i>�����?�z(hb[z`�Y�Q*�F�R[>aȆ�|Ar@���O��$�i��W�}�#�}�j��Yiʥl�E�����0B��j�AC̑8�`�W�>7v5������k���*G�B7�;� �Li�wZ����ā��c��>yܘgZ���aw��)gMw�YD����|���������0�0�	3�`7�I�q���ߥ{�U�?Ee��P���)l$v�5�ğ2��C��P�7*���TcY�Fx��`��g&mR�����8�[��_�-A�q�1��j�U(B��[�z�xIf�4�o}D����'�DŽ��ɝ����׌��O����3����c��wd�Xߤ0�S��Р�����O�6�ddF����q9� +�D�z��]���'4���#X
��[�â:�Q�����~����c��#���?����)���]�q��W��WT*����y�H���"fA��$�U}h�2�yR�0R�kI����Y3���n��\) ��#L2���v!-��=��Gw�QZ�"�g%�����HEo.y�����r�8̩4q���O,/2j�&��yp�|+��2��j�e� \���/r��a����뗂r�gcM�93*(5;We[�I�g ���a��	 )�j�7�`sỼ#a���]��1���k. =�
���~C�n��6�4�	}7]gzR��~)قn�ga�-�'Q
G$���$�xAe�bR	q=�$��������~J\yn�餦�j������=�$��ʥfĢ�2�m�q�f��VOⱕ7$�,LbN�Ό{����ūI}���}Z���-U���W\'��;?��m+Uo]��2&�{!�q'��Gq�Z��y9��PQ5=���ʝ�&)%4,��7�  ��y�(=����2�����׎�([�6ZX"��ﯔ:�MѬq ѽ�TX�;j�	�v&�=o��T��]�5{P�������kE����AbY���Ϥ��@&�=��Td��vc�������2�݉��S�_ǭJXۿp�u���zNoW�%�Keb�"��+A9�v�1��4lp��1M�����j�eC�[	m��+z��䁅^2���zz�h��[u��r|�#�M�u�C��K芺e��޲��&t�a�X`%�V8��U��������}��v�NͼO�YI�a�l���%�R<y/��t����uϸ|̥]�}�k`>&�O��6U�M+��1+�Q!0���T;+Sd��XV�n����v������-c15�S��'�3d���a2�P � �>�/���i�07m̊҉E�I��L���(�B�.�㵹�D)lԖ��PHPhF����=��S5�
'}Ȇ<��s��}k��A��3!<W�"�X_)��@�Ӆc����Nٓ�[�z/N�ͽ/c�ǻQދ���4��>��.�!3#�e�A�!N`���u���I�x�\���d��[���K��t-z:�F`)�v�����0�$	9.�A�A���Y��XR��1	��[�(���LfYO>!���J˞�ۄ�<�?϶J�=ճ��O��O���lFkh��5��"�)b�8Eux�;�� 
$��M-���7Ɔc-]�R���n#�l,i�Q���_P��_#���d�
��
�UU�ܚ������>��t��B�:�{�I��l�
`��
�f��'�R���5B@:��r�������֬�RnB�*�n�bJ��%f-����F��/h9"[ʫ�$��wU������S/@�yJh{�Xÿ���6O5�^A(q �/0�� �8��cH��t�lQM&��^Қ0sG.jn?@�:Wu��#˰BH/a<����0Y�'$N��Be���k�7�x��U%ŋJZr�Wz$|����U{�lU[O\�1���@br�'��`���!#9O���F˙:��`Kt �8���pSU��sŪb(IIc��С�!�q���U�io]��!�6'�*�ؤEx��� ���F��gI3Y�Xs�e���
z�L`#~��t	ȇ�M�[�!���s�N�8٢xS�m��p9̫HE22{��+���N��i�fF�Ѐ�/�b۲����g�|���Z�k3H`�~����G���&��e �I�7 Ԓα=eIb���)�� ~.\5���g���h�Jhvnl�2pZPH�4m���ߩ�@��\�ƻ�#ĤSW�ؐc�AR�Fs"|��M��U�i4�:�s���mj3@�5�l��fT'���^�b��*���ƺT�^���aᑐE�������Wc'i4HwF���BLO�>��%���U#�?5r����a������Y{j���8����|Gk
6��댘�n��x�{y����uO
�����NdC�ڻעяX �5��[�ɰI��a
��s�+�Zh�Oӧ��P�dE
��L�� }Ou0�	�#d�ӱ��o;(pJ<QyU�1�Ү��*6=�����P:��%t7Y3���hyG�y�ێI�Y!���/��l�<���N�k �w�x��g��3��6��,>#!�{-ש=N�� h�2�.]j<Թl��YJiƸ8�Q��Z�xX?3�B�M��+��>۟����U��r0ZC����;8���_�2����`����|.���j6�
]Oa��E҆��̬��K3�f��4K �P��L�%�]J�	,ň??a��v�,V|��?�-�&�.�r8��\J��P3ql盢-H��������Ly9r2C��:AX�D��	�ְ8)l`:�{�*b&�b�w�@�����WІ�,<z��ɑ�jOM�w{	�΢C �2�֣��mpš�)�3qD�J�*i�ꖆ���_�)��PR���	����rր�;�V��d���|ĩc����3�iٽb�j\����ѹXZ�9qt!�zLI��#�Rc1¥� �?��e�R3oUMn��Jg5閷��T˄O��3l7#���^D��hY�+v��P>ğU�hU0'N[�l7��ݟ1Aό���5U�o��&��bw�������3��}&`�����VAC34i�U)2:p�[��^R�'���~�qV�������͙)��bJ���{g�B��*1tp�
t�������(�ĝ���L�\�._�guuƖ�u�^3��LqY��1��'*�k�p�rr�>N���ȱh�Gy©�g���1�}2�Mw��ݍ�y ��6����3������F�_����AD�Ia*Y�^��HIp;���E:�� �R��0,Ur���S�qG�Iu��Y�U�3��V	
^AS�>�����wK7ky�믪p�}(Ee�0<�S^�RH	��t8��h GH����F;`6IM���2�F_{���꽒� �������b1�(�)1��aE/�mO�b�~)����<�[U?lM	KAR�h��L�Η*b�$�$F����Z��B��e�F.�IE��gSmjy�O8�0�*�#���\�h=��ݬ��CC* ��/��`��K��j{�@�BԦ���Ϭ׏"H+ݑ�?�+]oSw2ٔ�%W�a��L�k��UZ�!�ǃ�E G	Y;u��B��8�9�8h���k5˂x
�nMO�O�i���1 ��>G�1A�Ҷ�i�#�<�*7�|��u��^��b�*j����w.��_��"8w�{N����B����L��9J-aF1Z��{�id�-*5qE�Cͭ�;<FTp��}"�*t�	w��DGڰ#j)�B�Ŏz��Rdϩq����_�rpo�����X�N�+�$�l�m�?0����P�Wu�����#����%�y�e9�p��8�?�ݩ��7��B�u����`$�HTL$���9��0R}�QFo$����~�Τ2�]$肏�� ��oAX�F�0��|�8,�d��xk�\� ���f��ih�����o���\�f���c���O\�� D�~�]��3S�J5u}�6�
�����i�P#����l��#U\��>�������a�����Q%���n�0�-��Y�1�i��χ�7۫cx���}�A�����ʚP���ER]� ���iKI��;T��m�������:Od����z�x��W5�R$�OO"�
���%��Sm`EUyڊ~�������A,�C�O�Fʤ��k��u	������R��H�p�K]8�p�p��|B��Z
,�sT�F�D~�^j�.윽.�߸���3�Y�Q{�ow�[�9�ⓒ�>����k��&���N�ӱ��B�j{Y,E�y�bEa��s���_��3GY�t���Yy�C�n�!��6+�c���_`O�S�6���HQ���p�͋T,DW!~���3�]�Lq��Ų6�C�g"�ƍ��n[g놅FH�꫕��}x-�g�8Q����r��SZ���� j�Ay��?���}�o�p:�IV��҂���t=M�oU�7�6��w����4T�]�E?:	����N�u�����[�l���d:�
rڗ������ќ��v[to_����� * =_�����C���Ţ�q��-�ڈv�̺��p+D���%[	��{��#賧�ؠb��hp�Ǽa������s��K�Ni� ��ɡ��jLU�����f	Z%2���������h��5�WK��mS*#��fG��\��L�& m|���M<��|u�B$��FӸ�}TVL)��2���i3�m ���m^B�|u������ƂӤ{��U1.Mf�,�I��F�9��&��&EΔK�[�^�-��ל��r�ČkY�F%��q�h5er�C9�V���f�!���j�����"�)f�Z�E�a�Z��_V��sP�	w�V.�?�ͅ�3h<����L8|�����c	����_�6��"�q��<-b������M��%H|�(��c" �Թ5|(�(��:Q/�s��-TL@;y˂C2�M��������QS	�,T�2f��$�������^�i�bғZ��7�_h�
iv!|�ٯ)�A{�3�&���J�w�Z_�h�5_K�p��A^��HG��
�p�ޗ��<{"S��s����F��� S�f8��1z+�:N��-`Mo>k��>UZ⋴c[�4�
�!���V��v�x�W��	�V�So�v���J����m�C<)� ��1�@gm9�*dDe$x�y�����ib�0��q~&�T@��VJ]��F���^ӻ,��O�r���yi9��� P�������({#�*�"-��OO[Yg8ِ��&e��0<��0��Z#��~��)w� ��{����/3obے��yD�Dky�*��'�g�O%��Bwt�W>_\Vj������2h��#]ڸ�=���1��3?@��-���:H��Y����u��I��%����V��˒���wb�.�ݦD�dM�]ۑӗ ��N�}��P60ƾ�+�A)�@�(��z�ۇǅf��Y�F�&�.�<T��4�re��Jǿ�7�)�u����]�%�8�m���)8썡y��6�L�5 h��(�µ�T
b��7:	��<��%����6vQM���r\��*��&a"K�,�SJX�������uDr��|C���j��C����G��I��&�ψ�<\zUrX}bɨڋ��L���NO��}!�~�3Gj5Cd�D����xOk��M'� �Hj�P�Y�x���|���h���7S{s*DV>'���X"���'?�9sی�x��"�����8���b���C�6E���p�����z�ɷ�u�������	os��[���J��1�3�����I�C�Qő�'��A�a�NX�-h�!H��-\��>��'d!��y���!��OE�G$�l1���T�	��9�]�3�e>�l�>�U�K�,�[�z��0�� Ŷm6o�L u)T�O������)�]zwd��~��z�j��0v
�6P�G/Tv.4�A����ׇ|hm>˃�M�,�0}�L?�.'d�}~mÀNIf��Zꎱ��zA���=f�ߘ�xlo�^�!����s�[s�$\��Mn�ň�f�w���6�;+l��<����q;3&uh�I3��5��6 �k7�3({!5�Q%'<�{%�f|��i��zP��3@,,����Kʌ�WVL9��>�s���}2���+�-�ǡ���: [4�����`��E0����dBə���uA��I���t��(t�3�Ya��s�;K�L�0N͵�<�aW�"�	N� ��I��u�(֥}b�Qxً.w�cҿͿ'^���b ��<�x�����4���XW{�:B�eM�_�B�mL�#������]��&nJ���CF^�Q��`fM.��֔��8�w8g��3 �r��V�A�ϯn�<��Ԧ`�/3!)07��c�DY9i�/�z���;�L�t�7�H0�� E<B�<�Q�W�Й�󂵤M�F�6�P�g<��f�P�I�cPb����`��<�܀<q#^�Z Hׁ���Κ�K+���`��P��aEޭ �[�/$�6�j�N.I�?��Z��$�ȬY�]*]{�@=�z��h�!�i���~�i_��Ȏ������}��R%#���q���� ��G)yKr}�`T6�y����&�v���	����Y㓝c���8��^ fi��at=6�
U󚚷��"���@޿�4}U��U��S��X�m@m�Ã�7ǥ�Ċ�ֆg26��+xl�	����**�Q :1��f��D�v����Qk����.����s��hz�/�VB������s ���Y���l9���;^�dH�j�LXfV��Q��%�O����=ŕ=��/�.��0`��`zR��H�,S3�i6��>Թ����~<l4��,꽜��L�n%�k^�wI(47�k��b�=Y�}�k*�p�/�˱�H���=D���~��8*���@s^�x<�q�g(\[��
������}^cx��Pg�繅m��7'�i��� ex�l���i�O!/���{��\N�I�" I¼�����J;[�{�n�x3� yf���\9�O3@Q�~fX��;~5l�(G�c0L ���kd�z�#���
W^��Y�fҠ���"j��{�eM�	��%w�l���#`���{�O��O?^ռnC�A0q����!m���S���E����@rAzA���T�\e�'��%,v�e^�R�K25�6@!�">7Vԁބ��ġ#X0���ē�7qH��>U�Œ�=��}��5V�Z2��'��J�Z�2�ˎ�z���Xw
ͦ�3)9��r��P��$�5ʋt;�\�pM֒��'��Wb�Nf����a	��]�S��'��a��F�����=#dȠ��rTW��d;q��N��w��$�[�>?k٘:3�!��bB�ਪm��<��k"��t!����a+l�>��4U�/���J�O*C]ݠt�Thر:�����v]�����Q�;�㗉 p�����Oș'
g�0{M��DzǢ+B��R2�}����+n(�q��>+0�NQ��	��y�p1��m�����uG�f��-|�?� ��Rl2�����*�t0�ϲn�oO�]���b�Z��-�+G��fk�� Yu�n2��0��7�g����bx�y�оP�|�)�h �A��F6L�$�i׼+�:
��/�����bi�7~��$��nicnL�&����*W"�yk^��1#K`���/M7.�;X�3
aĻ�K� �dE��K(S&.L&b7Z��̙��n�?�E�7lG�Ւ�����=��!)��ï�yx�����M���Иp���@�U�MY��ӆ�������LK��1�V����5ȓm^�5�0K��/��Q�/�E皎�Hb��)ט�8�t�U�$��T�c N����~�/I'�%9%�G�+U6�1at��t��(�ꉎ��(�8$�A�z��_^DyãN0t����|�	3?�΢�^ےk������1���#�����1��������M6{8��7j�W�?���P��*	z o"���멾�C7��lB)ZG-�I\�z�e�jr���n�?�q9���Q���<��h(��-�X?6�:�CW'�e���$��_T��<׶�/b���+[J��Jm��T�T�}�W��2+]�3�'�� �g8c)Ҹ	N�����8�q�N;�3� �+����S�$0�+Qc���)h��!_��E�'��=)͓��7/0h�A?��Q
�,�P�0�q��c�~���h�C��ú�Yݠ�^)8��a����z̊hHH8��(�&D�qJC�B(�W�}�Vt�I�S.���Q��G���]�ȏ;���A����B� ��i��K�S��a�x�{�n�FIT����^���n�<Dw�ʲ�y]��:�zs<���ݐ���.2���*ŗf0�긘 b���;��;��W�'�ܐF�Q��q)�>�]�O]-j�N��ZK���C���ݭ��7���]G���l_���^��#!���J��p��6���S㑉R)��V�W�P��s��Ή
E�+�N���J���uL��EΧ�՗�!e�Z�;ܨõ���!��5Q
PV���X�'Ilޅ�un ���CJӃ�G��F䎤���7=:!��h�|�f�FE�89,6�A�Atƞh8BS��`���r�4^���c��#I�-6t�(<�VG�0���:F� ����~�j��l-���GJ�S�D����uv}��}����d+ц@l�CC/�5��%��t�2��bvK�M�h�$�B�J|ڨO��đ��i�+U��T�2�����]P�\jaQ[
%B��B�Ѫ�+�"J~wq:6��
�{�
�Q��{Q�4��6/�X����3H��癛v\�YJh>Gg�X,�S�*��O}�˰r���p��.������&���d��f܇��¸��}������t)k�:�n鮊3�^����Y91���4��I!���3j�ԫ
v~�K�F7��V�����!�b�;��=)���i<^��-��wD/�rk��G�ZJ�$�N�>(@�ݠ6��He �����mh}O�X�)U�rbK��(K���l��&���2pP�Ӯ�ɟb����"���I�z�AL���;���<�4�D.,�վ�.rE��O�i�&�:/>J��knp,ꕗg"蒽�uR�������Q��9O_�z�(H��N�4qړ��e#*��H(�F�!�5 �ť�KQ����r���.\��z���/n�՚�x�P�\��h�s�̣�[��bW�*�(�ɗ�Ͼ*���z�а�$�	K���7ѐ8w�	E;��<���-WyI�0�L�C����K�N�B6\f�-�B(�Tl�hh���Z���>�M�c�T!j�dЅDi�A,��;S�Cj�Yd�}�!ʏ�k�P����Q/�n��|��ˤV~�1j8˥Ϥ2����%Nx�-�zFD�"��w�o�Am��b�?r��_��MA����`�o���$[
,G��8M��c�ݶ��9KJb����O���~c܌�����S� w�᫁�k��Dij��.��{����2_3�0~�K�wϦ`�lp�3H��B��Z)�'�C-�mE�*	@���)Z=7�.����|��zg�+I�c���`U�=,$d�`��R�G7�0�����[��/m_��4����6(o���	�>}����z�T��%�u.�@���Bx����ְ�3&����w'3��A-��SgE<��Az4��=8��7X�-�\^�
$�[	�ٔ�b�L��1�d,P����+��6��L_Q�&��'9��iF<D
�q��2�`ɏu�IIyӠ|��Ȓ���^mAN_��Լ>F������2��{�R�1��>~@e0�$wtEhtK�o�Dm�����(#��;��^J�Ç�4�`Y��:���¾𪪰H��:k>��g�����=Ρ����;ņU�&Q#2G��������ެ�n��RȬ�@��h'Et�n.���Axj�Q�ds�{�:�A� �[tVz&dn goȪ.i����W��m�D�zϘ]�0i�`�،NJ��ٯ��q[tQ���?`IaM7��Ҟ�u4��t-��4i=V�렒��cb��F���x���-o7їԗ&�>��舼_O
EL$ܼs	���L�����:�r��h�\w�*�^P��)���������p�^;�!=[Z/������=P�/wߋ�&�W�X:$9}�Y�mD\���������[�hK��tb$dz��ЅTWb�Ｓ?�O('q��;�_��
�(��k�jf�ޣQ�2Z�|�� ��9�Џ�j7���Ã��ۆ��y�T�dE�:�.�/ȷ^���Z���S� ��jH-����Ж@&�&s�˼����v���h���훐h)��*BgV*���G=���P�Pq-!2�Ԯ��r��9a�4��J��"o#l�@��rI/����e�E:�=l`쀰>��C�.	��+�D,�ex�]5���+�S`�r@���-;A�t*���n��7t�U��gj�r��0b�-M�n�w�G,\���'[�����a���o��ym��t}?�_Ȱ�P�%��b0�I|�F���yTԑ���rW����\�Kx�[W
J-�����D���vb
�^y��ng,�H_6%���W���A�Sj��{E~L����D��2\A���f�w9�2)��|(�mr�'8-f�(xj�z� S�8����y�&+:��X����1�#�<�̘
����^F�*`6�P����,ӧe��+?O���[J^᱙��_]3r�fU����(���~�wق��(w��RA�ĸaP
m��~�u�m^M��a4���}]��E��������|V�>o_J�Inʢ�0#]�X��6:{$��8�1h�P�s����^�f�dB��c�$Ԑ ���~�%#�m22��6����-q����u����;�!AH���i3!�cU�Wb�(��H�s��{u��p�4M	-L=�k��Ԅ\5��{����ZR֜aU}��Iش��P72�2��|�!$>Nne�!�<3�h ���@&#��~?�Rb����Og������v�I�[��f���8�|��AG�q������D8���L�J�^�2+'����O��Ȑ(�=���N�E��8�H4_(CE�N��`�;Ta��o���yz�7�ډ�q.Y��JM0����E�3Ra�(}T_
~���3�uv�%zSt����SE��j��烦��R��@	��� ����Ἶ�`9������k1���bl�e���I��@]g����k�w��![��u.��/��>�Ú��f�}���G$����ᴠ��6��G¾�WԒLa���Z��߬�<���W�H�$2r]tt����7��d?����`�������]�b���ho�|�L���L��cGr{�ғi���}pj�^,X�;~ޛ���3ߍ�M�a�|;�%�Yؿ�UP�O}]�oG y�y�C'H㯌��z$ȻME5΅|���<g�ZJn����ii&�@��qt�3��p$�)��D
��������:�<#ѧ-1�j�=<�
~U����f��ݙ�����^&}����߼5e|���úb��7���H���a`��|L��3�B������)w�}D�u�uj7�5��۳���-AB9y�5s�1�qy��G�Z�e��l��+K��?�� ��� �<teN���b_�͎Y�M�|�MKT���߅���B�bő�V�;�y63}��L���NR� ��C��JB-�Aq�}A� +m{Op���S��(.���-��3� ���p�UCb@䗸p��ZӮ�g��|�eX����PR��v]��V�Ed�\h��.-��i���'�/DL�nũx���G�~�&����	Zx)��d�V�C���U ]�	pk�m5渑_^��B�4�J�/W��P��4FjA�GE�`\��F