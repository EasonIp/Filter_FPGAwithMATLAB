��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A��#��Hb�а~�g����o�+5FL�cu�ȗ$��ƃdY=�7Ў.�;;yfP�)o��#�u:�E+Pd��U�(}M&�#�ນ"��:'{�x��v~�rG=��t\�O~��Vά�q$H�ɦ�| ��4�W�V�sh�Χ1U��wGpV��5�cKL�r*���۳(�^�:;�ϐ��<�K��l�ޕF�Vpԅ��e�)�h�.;B	t�o�Q"&����b|���H����I<O �y��d
�4�.5t;��|Yx&����d�c�KF��1�	�j�A���d.�8#�m\�*�u>�kIB76�������\����o=H˹\����?<�DM/n_�R���U��!&l0��~I�R��!��_��4sw�7`�P�
��f;���FzT�
��g_41�H`�D�|�g*� 5'ٛ6WPΛ�xՄh�����T���
���N��'"���Z�-��9��B��Σ�O|�꧍썹=ŉ�ΘNtc�)�I��.z�ئ䪁LRT�'p�l�a�p��UF�-�x�U2?j©�ڳ].m*��8Xa��5�0KM�/P��>I�x�X"r��U���߯4)�ۍ�naN@�A6}�_s�O�X[��i:ӽ�@�$�:#7�
I��H$�M���~ A�;��b��=��0�:���G�&�A�]����#g���mA�b�^D��&LJm� ��HH&�1;ګ=��
٧�oK�L7E�B���� 7�@����K��B��5�*���V��^-�a�*3�������z
�AN�?�3�n�T��:��ˣ�VG��`��	1p�j�0i���yS�<�w߹�ށl_��&��� sw�W��J���>$�������b޺����0d�]S�F�,V���o�fRI����/�@�5�T���[�`�˯�^"��D�O�SP��,��|pJ�J=D �[�@#��e����fa���$<=���b�ڟ�$���G.��Q�X?��=KW�//�2�d�5�A"��NT ��D������=-vLh�K���j��9�t�*������Pw`<O6ʆ?�[��7$ڍ����%�'瑾�����¿2Ԏ���* Ԫ�)�I�����@�ҡ�d����J�w�߿n�mM&�0���+dz�G��IS����PD�e��]�ł�$���F����.&�C�G��Ɗ��5��i�uGUc,%aw��5`�G���}��-��d˺�(Y*j�n� �m��ݲ����6�oħ,�xQ�9}j�B1_�'��zPC������zD��m��]��D�V��Ɇ8�T�Ô?G�C0DU�$�
Q�q�D��r���D�R�?K�ۄ5�D�������0yУo˨�Z�1𞄰mX���,��=� �_�K��������Ic�$������2m��:Q�:j?x�'s��G�_y�#_rJt̈��R�����������1�>�N6��K}�G�����D
f�_�����!���b�W�=�_s�+�V�g���)e�'���ʳ�y�� ���@s����:Y���T7^�~��o=������TOS"N�2�a���p���<�+q�p��6!���yދN��k_��K��ކ�x:�2�.���U�P�e�!1k���EEKaS��OJX`xP�2�xqm��ڹ.�Z|����j���qH�5��Q!-L�B;hSAxe"
D�\]�0�����yt�N���-��Zym��*[~�?�|'�g<0�$1�(��|h�������ְ<��d�.�� �i=�C���xE��	�TD�evL>��`Aܟ��		m��E;�	�Pv����_ab���2����'u���{�6��G�����oG�l��$<�(�o.�׼�킩2UlOS�M�l�̼��&^%e�hʎ<�Eʖ���`��(�1�8���z�o���1rAU���YMp'�Cݙ�j%!~�5l�Hp?�V�`}`߫4J����<��&㈑S��D�T@}�H���"H�C��8�nļ{�	Y���o~~��w��i�?9�c�+��n�xύN��h���:ί��O�kAq�^����L*�43�7��wkf����q�n��/PKr�yq4��lۓr���;��鷁���Ƣ��J�g��"��ρ��>�W>@8j�.,Y�H �_`��˭1!��Ko.�H���I�3�xj�N�yC"��ӱ�}��ɯn��Rr7�C����!ڄO}\8O��ه�(ó��e[������%�I�Q�����A�PO����13���Am:�Sa%�[p���RT�s/9JIb�V����ܬ�;;�.7z�H��n�aWỵ7p�V�������7�䍹�g�A2����e�J~*�Q"ޒT���'��(�k9�j삝 ��r�[�x��?;��o>�v��+�`[^���f7O�j�i]<��q(Ü^�p����ѝ�gǬ���h9�F$�U����,��gJ9���������y'_T��Կ�QEY,�)��nVPe�)Bh���*y+d@�1
)~�V��Kl�ų��%lc����v?h*c�1x��O���e�K�_�NB�[Q�)ī��tGW�j�m5�A`�ѐV�j&���%��:ȰYZ��MP��B:W1b,����٩Kϼ�	i����\T�n(���}��3L���ɸtL�<n�	�Ǉ<*�������C��C��2��è����=g�W�}5�.�{T�[6Q�=�\j�D��9�r|n�����l
����#��ޓCv���#�I�lVr �n���C��`߀��D�^��?'Cׁ��'���ʵW��ެM� �y��}�[z_+�^����;T��������Ob�>�ƻ�r�g?�O�b5m	7MǮFP�nK�゙�j�x������ *��4�CrL�i	e��#�&�\ѽ_���LI�� DG�x�JM%�y41HΚ����D�>fZ���D�<ীb�Af�z�D�	J0��c'	̼���5�\x+�=W3~(6�H|4���Q|`�u�"�U�J��3aN���o�&1,�=��hE��N:���\^W�m�&����h!XH���.�|��L����e�c��0�C���LP�V/�D��|뤯�����>PZ6�5���2�>j��Bjp��9�#X�z	��z�0T|���hJO����}\;XH�ǟb�Ni��G\�t�(��`��W6��f7�|9,IЕu�J������d���e0����yQ�Na8���*�4��9L��(Dfn�*_% Ų,^���{s�$B���+��|��S�i��|�(�F��H^
���"�a:x42�R��v?&B�9��W��!a�;��_S���]P�v{����f����-��fi�)���M!��b ���yK�Գ��-��1IsN-�qL�/��Q�ڼ�,D�Mb���*�<BF�~�(� ��2��D"�b�� ��P(�3��f��nI|����H��n`7EO�̏���o�畈��y�f`"[m$�Ǧ�IF�2�F�c}�O 4�@ʸ�U�F��Y��X�$y�6���zO��M@ ��g��5��sђ�pEG�o�(����=0��Z�h�a���h��PG�3��N��ܩ�9�9�f�sF�D���ͳ�0�z�<oǛ`�2�M��y�(��:",D�a|���FcS��?Y�Ѝ����L���Gg�D'��3P N�]�PP��U��`���oT����@���ڥ�M�l�ҕc����=���.���Jz��ŉjH�y�ю&4E2�ᶃAI�kӍtK�7�ǈQ_6�r\��7UG�|��Y"o�$��Z�C9���b���`�0j��rª��3`ރi<,|⅍��9%)�fhm''#�������ל�<"��c�ю���="dS\���KR�gr�`m�8��&�c����Sᕉ�Gm�e����/��ź���#�	�|e�||p����1gCSd�v��k?b�{\���SHvɝ�!���~!Y��"k2~��H�������Qx���f�n,�3}M J5;�Et]�I����~���h<b`�����g�&�Z��U�L�Ss��ejU%�`J]9'�/ث����1[�6<hl��9���� F��[0X\�ũykZ%B��P���y�*���'���q���)��|I�9���
��0���.��sS�L�ª6���Ld�	�n������<v�<�٪b9a�ȭǢ(�Y|u����߹�	������;-�UdX���=A�+�rwK�O������:�Bq9S�Y��T D�0a��r�ָK�KΧ�{9��E�T��5�h^�3�^���:r�`��fo�_E������%���	�. �ܣH��ьJ4!M�B�!�j��P:Aٳ�y��X�5��$����V�F�z�� 7�k���9���(�0h�g��)�W��������� �h.�΢R�.��a�,v��G�ҩ�^"�]��FQ�eUj�B�r'�@O~�S&��v����6)a�Y��Yq7z�ݞ]�_�0�TK��G�/Q��� b���~�W'��;\OޠRmE;�mbΛ�V�vP�d��&f���{ �!,�H`f]��(0�)�F6�J��O��P]6��d�����vF�YI�0��Ö����M���;^^na��w�;�!�A���U��$4��