��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������"0F��}�h'��8��<���9���-�j����,W�_/�H: 2���x���CH�^�g߹+�F��0�tw:�j��{�)�0��H.�'�[��'0���ck�D����L�Lq�&��IzV�G;]V0~ݭQ�����)�47�gP�ILO�"���tAf�?V��-8�/b������$�9~�
�l])V�"q��&=��b]��[��rL<�\��+��1:����Q_��!>5
9�͖RT���/��Ől��W�f,���th��sC|�o�lԾ���3I�*�)���l�넢�}�����'�x�nM�Y
8SE0����K�!��I�C3m�G]�3�����v���:���fT�~��g��ͅQ���o�M|eL�|��|!�)+s՘*��έ��b�E.LMi�.�*���Xh��c�NV�R��W�N������x���H>����e��!w|�%%'fE��d�__}{,Nj��I��"+����[�	��L�QhZs #�b�n�(L�Һc�C��Q�6��l�Wl��2�m�
����1�@Эn���\�^��@�*&�85^�Qmwݰa�,�C�]�k%~�$z�U�;7�Cǽ���A�B �T7�C����El�
e��wl����(���>X^vQ:�&>:'�>�I�xMK�����<C���^:�ȹ�*�P	 �k��R��\�q�G)��<�@�듻�*�=�5���s&�μӮ�����uR�S�ɱ�n��f�l3\���)�oH!��c�ޖ�� �*N�s�)��r���ʯXo�k/ZQYDD�C*�S��1"�q��KS�[��M?���91_](2	ԄKJ����%�g���(_T�[$�K�R�isq�R�0�U{Fȭ��+;�N��o<�$�e)2��+��ړw8C\T��/� y/���,�f�F*�e��M6�u/|��P1�k��O�NMq��	�Q_8H�Z0! �z��[�c�+�'�:��h+L�ᘬ勎GQL�|{�P3�G2�<�0�R���c���tW ����=s�Ve����z+�S�7�#��N��^|p���N"�M>!�c��`����:��#�}!��䜵�ǂ[����8{?��L�un�2�DL�=X;�e���ɔ�Lh�� Μ�����YU���������S;sn�$�r��ɓ�[��~�4)�_��|iM��9���l���U@�sf������f��н|dBs��J�r̍� ��R4,g��5j���ԦK ��&8$�E��T��=4����l��^S�~�j|-wq(���m�r�f��Vm�ACH|�S�F���.��Ç'5-]��t����7�
ݺ�N��y�"X���C_�ߤ>a#[��1Q����z�Qq8K��HIc�k6h$�����*���Dxwt�b���Ti����W{:�>8:m1�>����<e��z����,c����M_x7<�O�'�4,ƒ�F�E�=��{@�����۬Y�S��]�78���0�"�'�q[�I�dN�Oa�X�SE~�'�b�6�ףv��Q�[��<�&����)iMք���������%�y�ko9Uf�b"��^��� E�~ݧ�c��|���c-��K�W�z���c�.�	&��j N�Y��м�ا�������r��l�`���C$H4>��^�I���ј�h�l��P���o(��-im�σ;��ml�h}?��S//1���Y����'0K�+8^����A"�L�����aށ�k.���$/����5Q� �,��5��:8>9	@�J��T� �\��G��q��/Zo���p��v��ǌ�"�껰�y��ۥ�[g�>=�e�m�2���^^_��l�Mjn)��u������)��<-ݤ���sU�Id����1�G�b���`4P-w���2 �@�WF	74uƐ� ]���to�"��p�!�����q#Ϋ�m:7�&TT�)(
Oe��f`|�ȺV��l��u�%�Tʁ*]��[K#�v�ܧ5�[M=�D>*��S�V�=�
�H�1he�{U�cl>��h9�u��d�Q�8+�C5��7i�\��1�m߈vz��xi�=`��r'f�Q�th<�>�h ���ye�JXa�}�Y���R	�n_�c��% ����C�3.}����iY�&����,9再P��Au�Ü��+!=�"|$z�(��qd� �s�v_�M�y�0�6.�a5�.R��ժ68q=b�Rʏ"Z/��(��B�e���h�D7+�,��Fb���7;��u�����<,��2�c��@%�a g7��M���6�;hЫ�^���[h�U�� �8�*�z�Q���#�J����0��|w�X����>ۓdƷ��mENz�M�S���v��Sa�����ApH^A�^2�f+�ͺ�9!��}���Ӡ���^o:��";�� ��Ƙ��B��݄��6ux�U�5��t�>�.�ф�^���p�]���H�H�cy�E�T��q�k�>Ω�ɉ���8���O�����[.4�)hp9�E���k�"m
�~�Ȟ�Cx�Ꙍ��3�E\��l�Ҩ���QtD#���o��{�[Ɨ;
%�������X�2�&Wg�I8"�M�n�U<b��s@�h)�Eq�1%vqI3�>�s����Ig��_ӻ,#������9\�xU�s/�n~<)WK���kI"Te�K6�V�P%�k�f��z�A�P�1�ZĐˏfTB���ikx�� �5L����%'��d��Trz3�RU�fX���!�6F�)���l���9��3��p�E�V�{l�4��4�I�S�^���L_+��i:�`䗗)��!�j������K�z���}=1M�"V�@�pb^�c~�I�@��-�'�� ���;h!�w��%�=2s'�"�!L@�Ŷ^��a�=ޯ�����[C~E�S��FfyG�j�k�@�*#<e���P���ʰ�}�ρ~�IƹbX��","�Õ&�v��I�|�n�6���w�4�����Zզ- 4���]T�;A�ݡ7R������
�qԺ�>^���L+E{��a2�\�6,�����.Pr�G��ȯ>��LPeK_���4{�@}e�ïrzL-�Η.v�6��|��fi����!����y��ى��24�`��˝Y^u�S�f���t�z�Þ>o���'�\SC����d�.�]����&û蜠izF+DO���0L�����ɉW��_.�U�r�لJhޖ�����oŖₛ�P��UW޻c���N���O5���k���'_I|���$�sʠ���΋�sl�VM#�$F^�+���Y��Tu�jN8|QTM
��rXỠ����H���.a��&��������'�sT��Eh5�4�-�\;9��x�ғ� /���BcE�.+$ш�@���y�z2pŁ�P@�;���g3��]j�H�mf�����=Ats�6Zx�6�kvj�����Se'C$�_ ��;�Tz��g �.��q6�O�L���6�������MI���O��b��D��ea���9��:�nƪ��� �*�c��^�рx�[�>Ҿ�}
J_lӭ��|�}�wl����*^~��t�N����Ð4t�+vrW�G�s��4�)������}.���fgf�֕ex�x�C��\0׺��fKd�B�߹��8×y�q��o��1���iT�,�%�#�	�v=�5��F�xo۝ZX<Q�YwW��pR$E�Tґ���m�W��z�T����A�N�Z|A~�?�����'f���)w�H��}��kOLdO�e.3�G����cLq�W�s��Z��w�(�dP�.�/�8�+M~]�M��t_�fS�-�UI����b�F�����Y�j�0�����L��<����f߿���:j���$>��p͍)�^$����o`��}_eo��g����g������"I>7vP}Ἕ�t�Ѯ(�Kt
�s<p���RRZ�!Ǣ�S�H{����"�p`�<��!^u�q�o�{���K$�rk��K?����Ȍ�ku�]�D�ܳ���V�N	
g�25����gDΞI�k�he��Ɲ�q1�q��1M�b�(uF�`�M&S�+��4^d"��ؠ�����UT@����Xf�A>��R�Z��2�ܓHؕh�� ��H�I��d�J�V=�@���bT�֧V{z�H���H�=�m��:���RI�t�$#3�� R�YWZ��O���<�R����:K���<��R�GbV�H��+|
sM��Ik�����Y{�L��2MY���UqD�AH@K�nSP���ȒQ�_���7:
MGZ����V�Y�D4�=1A!,���"{^zY���g/�¯�L��[�U�ׇ��b��aO�C%�.yu��~�a1]A4�7̄��{�[�uE��p)�j�WC�l@��2���^�цh���/�ύ's�_����=�:5\��������nSXx'�n�A{�������5����[/^��b�z�%|�I%��2.����n���*t�>�C�=�Vìd��rPpdm-S�b���\����[�_<�����`;����|���P�FtT�'z����~����Tk�#����&dy��c��A:�i���w�\rϛ�>�(�*�IYhw7�y%	͸�Wc���[
��#6����>�R<J�Ț�Ɏ�gS�P-��uNr�2Y�����e{]�0"!%��i�-SGL��ar��ik���g�ݸ=�*��Dy2|�5��!�Ž���`>�d����������Sz-5m6����Pu�9�Uc�+��L��H�k��#.�`��E}{�#_�C!�FNJ�n��J5�QF<F��e:'�!;WB�$k7]jG��r7���oCoZ��'�Z��ifX��Yp����TUX}ZBMFE��YaU�Lx5EHy#"$�ϳS�Z�p0*%E7��6����j�4����ͪ�iy@�Kl�#r쵕�;=r^w��R�CN�Bt�i���V�¯:��������	TB�p��սn��x�de�¥;ә޼�@���h�3$7�] l�e�[z?��. Ř�BJ�D+��%��]�����b>�,5��I����^o;n�k�;-���BF�_,!Q
9u�ߌt0�m������*tbO�:IքN��#��E Q����8�,���R��	C]2\zÕ�l.����)tYʜk���H�qU� V���9�Jb�I�~N"7~3��ק����&�7[��Tc��l1�5��Y�('��QAW	�h�or�l�v�S��i���O�.���@C���>�]���b҂u��a[8MR�%_�e��B���q���&)��'����U��S�ԲU��φ�m�q'wS�K ]f7B`�|vT�������Ux��A���&P�ժ�u�Q���q_��D�o�e/�x�7ه*�.�eRw�!_�殬�{Dy��dt�ߍ���Fsw�v�����o¹��tf���z���A� �:"`:i�3�QEQ��N�7;l��������L��� ��uP�ۂ
���.�*-E��!Y�'�U�_A`��ы��AԠ����[����4�^1����ڠ���|�ݽD�w�=��
Ux��k�[��	���� S�b���}P���}5�c�>�p>�^Ulș/(Q.h  jֵ��{�R؊�0���5�.'ْ�g�dQ����!�g��+ɪ4�~[r�$�mn��3���E[<�9p����˼��ā{6s�&��c�h� gg� ��㻈+F���e�����nW�ۘ���d�k�o`<6x���lj��F��(�Rr��G.)��ޛu��Q��P��&����2��EY'��:��{A�H�Yg�mkW�iWY��"f�aZA�B#4�r��?'d��YZ ibav�/ʏ��T�Vq*φ�#�V&�Gn�k�"M�k��\e�<���N���m��U�CLv��� �b�ΗB���.N�u48�L*d����������E8^��I�?���Ǔ����L(�=Vi����܇/N�X��*�93y��KHo{F,M��T�i�E�6edU��{�������w|vt����y�>��7�`A�ELf1�[��M�\��:�"�7�iWnj��b�R�D!!:-x��¿ʨ�Au'Dq;����\���@#�<>�KĊL�h�Z��14਱����IeU0�<Ǘ��*
oS;���T��+;�Wz�?��1Xm�*�v���dթ@֡�GJ|��u��񽮄#�7�u7T�f�N[+��a��Vm��p�{i9�w����ې���n~�p��7n6�hF0(.0p �����*H=n��<Ist�2z�>�c��U��,�����M�W7ܚ9�\��?!C��x/�'#wl/��r28{.�+�9�U�,�`mVP7�qO�@Q(|�뫳�ӑ˭9?O��˴�ڝ��cdKo����cD�j� �8B:γN��7\f���x�T�$��ۺ�v�v}�`vlЎ�W�8![�<{�˸ߑQ![���_��� ,��/u�a��r1"�$�t�`l�v)��;"֚w��S��G�6�ih�Je)jmh^/�ϺY�7Q��I�J��L�c���j��@0S�v3 �.�q�;���;J"��j���
9r#�DP�-��
^��8�j���'�I.2qh��t	�-��{�������{��������Dn{$]����a�˶��GIA�t)��7J􈤷�|�ѝ��3!�R�S)�rj୦] %�e��~�7��|�̳=�`I�3K�X�И"8\-h�'^A�/�y�-���!<���n��0�ކ���Z��Q�s9��/�(}��>���{�<��?1-�wR�ᔙ��ɝ^�ok���-I{�t�(��������j4y�e����>��Z4�"K�$���0�m�s�MY��`eO���Q���A?�{O|�CwY��~�q���[? �J�1����6�����@�K�d��R���?��^EG�=X(�5`W�v.�8��"�u�%�,t�1���L�ܥ�+�Á������L���̭|T��>���b]cfy�4,[�j#��޻�m#�_�[;1ۗ�e�k��&3�=���٣φ� 4t��lq�gE���﷪�b�x�JK�k"δ���I =m���PJ"I;+X��qv&E��%�yYG�<��F;��K�T���0��L$(��@�`M�H��,(t��崁�ب�n�� !5�[��G��e�c�P�D��B׫Q�n���������4Z _�K����C�hwx�#E���*�˹~���  *��J3`*T�Or��"��@���s����J�)s��4�\�90z�f�;7^=��e���z�:B�"�I�<:���i��h�9"���C>?�}���`Gu+�5� {d���wb�
)&'S��`4q�д�Pn���k���r��x�-����a�b��Fg�����p�H���wt�u�]���ːv����U���]N�X�H�r,G��A��)r��Htv!�v���]��� � [���;��Fo�>�[LA��SZ��vYN�V1y�'�bÌ�CQCqb���6�7���R���t�ԛC���l/�a5�Ɍ1��k$��ݼÄ0��`��9ܸY2��K\�A^��[����a��"�ýE?׳5 �6�O���D�b%����{Y�����|RE�au��C�p<�)�m7چ׶Z�~�;=oN�.+�(���q2�;e��֎i$t����뉵8��qR#]�N�U	Vq��+%������b6Q_�hp>�����4<�88���Z�RӨ�4��8y0F�+e#r���g� C&��@M� rXN@��	M���$(f͹�f�>Lٳ,|YÊ��C!�^F�T��B��6�4�ԭe�8E��[�ʺ������MTJO�c�l����!�ʪD7���V~r��vq�}I�r���ǠI�M�#�fh�$"��؟8�Dq"�.�6l?����ׂ�X�!KNŧ~y5�~DE>շ#��C3ա��IE_k0�L��&fSx]�\�o��ξnŉ�o���H֊i����j-����O\HaE'�u�v8�4e����^|�t@/Og"��kU�AH��5�qx��8V��.�W���q?:?��μ����3)/*�Kk�n��84����������_Eu!�Y�x"C��[0��A�qh"~�Z�5G�i��D �cp��P�p>?��|<�ٛ��} �e�F�'	\2d�X�B=a۞Tto>7��F�>pX��P�eA8�5�:Z�_b;��;�U%��v/��e������v���"7�/�p_8�J��m���;v'i��5^��J��3?�ݏ��LV�b�t��e4Qu(���f�m�����&Ǯ�␐ʿ� dǯ{�.�
�{Ө뙮�G���K`��1ָ�X�`�j�
i��0�Ζ:Ɓ 0	C���x��,��� ���_C��?�sᾹ6@���-֋��[A'
�A�;� �ǆ�`���L�|�gקrǒ21, )n������yL�d�.��eJt����_��.���� �_�����Ci��ˠ�fNO+�:"������'A?�\=���®�iK�P61snƮVz�g�o[ͫ�����֨��L�t�؆+�ҺB��u��c��ŋ��ɽF�+�0a�	w���_�p�j~�
r#�"��0�+ۖ9n�$%���/㥊r��S�D��ߑ�O�����.�_���h*���m2I;����IATK���6�SiG �`FH+�p�^ʫ��������1���t���IN;���]�X_^!~׭�VrG�L�IJ�^ZS��b�0ZCX�H/�@|ܜ����~rw��jSa![��W A����h���Kp�J��M�  &��O���I��=�o:�Y�傞����aYm޽5�ù��Ʉ��	,�����Ee��f�`���]a�O"ԢI�\6��jƂ��}���z���_�X��K�{jb�u�B��a��������րR4j��s���"��7��QZ�$#�dUGv�3��y�_&	�y�F��P�����zw�W[�wnE��l�qr"��G�ؽ�dw#���0��go(����"��`�v�Ιv&��G8��[Ԑ5�?'�V;m����~�њ��6&*6�>�|h!��7���OO���{���#������O���T�cE)2���14@o]��&�eO��r�ꊆbd���Ts�v@�ރI_LT�)���2����]Fm
JY��� +4}�*���cm�HhjM�������hg�^�Q�D�.��9l�&{�]�����e���au��:l
�4i,�֍�����I}P��������:������A��ku���
������6?@�iL�*@��"�PP��u�qAw����c&(�e�5r�Fש����).�{o]��˽��7��P�����u�c����#���C��#��]Nz�Gѯ��]A�Qod���nD~��8g�ġ�~�>�N�@�l�{kY¢gA�5=�5�����eG��K��~��w�������;r7�=��ֽ��b"��闢$'c�;�(}�D>�6��_H��M�R����t�B�����|5�17�JB���H��ř��l�Z/gЏ<�@m��6�v�uzʟ����}qP&�~�]Ռ$2��p؛�e�4�S;���P��tǢ|cQ�;x0�H.K�쎜s�vo�����z����Y�2��d��Eɞ$Ss�k�X��{�H	x�	�2�]SY� �Jr����M}[��j#Z���K�žO1q�'�:CH������d~E��ظ����W�'C���T���^�K�;�z�����P`
�l���:��!�3�l�8ʒtyeiu����<�<�U�FVXa�^[x_<˖��:5�lE��;��;dԠA���
�G�C��dHX�8W�c�Z�"9�;�� Ռ� ���3�#!(y(p"CR�yˊ��;O���Tp�w� �2P�u�;9�#�V$~N�q�#*R���P<b������4�A����Vt0'#�C诈J`^��:q�zvя�-�� ���$�դŷ.q=����Ҥi����QKu�!�nx���>v�־����^)���rp[�U��ܛ$��1hǶ�3�O�.�6��'߂_�l;������W�B[	��h��.� �u�]���-�c�5�fo���3#��=Y�G�/&���d:!�[�W�U�Sۿu��\������{.t�V���r�kh�����Q9�ҌP%�S��: y �[:�t��x���xqj~�
���ޖ����sF ����*bV���ZE�AǺ�'��o���f��49�$8�^�e<iOW�#��'x��q��z�4|cPG��v�������:��\��9Z�]��<D��X�(����� g׼?����VVN�&��Ky���?��ai�\�lF�6���*��_׻q��Pz�|�� ��vb��&`g�����O��@�:��cY� zqV�-�rc�=�4��PB1x6��#j0p��b������uȦ��7��N�k�ٰ%+ح���҅&.^�s���~=��b���!��+���KW�j����{�U����ܖT3d	�F|mog�Cn����-a}��pz�[jNϹ*d��E�a�u�H�gJ3Kx��L �Dp��\O���=b�Kp�lg������R��1���^��jq��3�g�`[l�u8_�us���TC.b��FIR�<S�`� �s����!�q�z^�Z�� �Jr��W��\��{V#N�V8���%�d	Ϛ���6�^��W�7e�ɐp�9m9��zlG:�?1��}��yK�G�i0~�]�d�;��ݡ�7�Qo��g>�0H�O���tX?L[[�Gz�qvǨm�7��uӔ�W�Sc*��=�l��"y�^���>xM51@�;л�~�D	�~�t�EPf�n��N�k��#@-9���:��ŝc�{t1RЙ)X��~�����cMŽ�:�4y�
�}�E쁁�ś?c�ȯ��)$�_�U�K=��=X�d�G�ߗ�t1ķ|WԘޭ@}wG%,��@��wr'+y���������� �a�=���D�,k�G�c��v�y�6����9����{��G�i�E��.���b��M	�鎠˅��0�Id;�0����[��{jɉ �f����vk$ /��}�Aȝݘ��(&>�GG�1~V��%� Ηo&KX��nV���&鏏�7^��6���L���|�97��<-�pf�I�];�Ks�K�I�@�Ld]K	_�ĸs]����P;��a`v�<sfj��	�j�p�?����|d�pZ�ԀY���B����q/ �_L���Ğn!������=�m��-�Д:�{K,r�}�y�է��{<�	 g���=�dHό���f�s~� �%�v/��7�|��W{��]�)������Pb���>0��H���&�1�5=ܑv��A��c�^l�C�ċ1���� ��g�5�+@� ���r2W��	�c��$�ؒk���wd�,���<ք	$\ 6V8�e�bb����_��@1+�ڱU������k>&vz������ ����~bz�U�Α*���5��6A�Gi
o= ����D%����o��c���j��F�f�:�x^��i�P���R�jG��5h�/^��,�pwC�D��k�{N%��A�݁Ϊot�w_���zG���-��X� �k �vPBͼ]���:���)6�]| "<2����@	w���"��
��̛��٨�B�`�wWT��랏pƬl*M݌�/h�m�q?N�WzaBaפyEN�1� =gO�>���-�3`'��i2�'��Ibf�lд4p _q��Ȕ	m'�2�gF���Nى�Cn�fP�