��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$���G�S*��ʃ��6blg<���15M��ps��O��1�>{����ĩj�{nLDD��5�����!�i�X���ec�uK��.q���l �I�����2� =* �-m�k$g��(׸��:[���-��M1I?�3���wԠ	�H�l�N\��R�_���F�r�2(�.v뫭	�M�GO��JM�N_LX[O炋9u���ϪM�XHܻ�@��"CMx��m���Ծ�&�����e�0����Ћ�U���k��D�^��|�H�¿\���DH/� b��h
���l�X��ٞFr4l��A���v�+�NN�5�M�g{�J�)�=��ë0t���>f'�t"���}ִ8�DBF�'��ήDŬb=��q�� V�!��@�BZG;����@O��K0�Qj{Cbs�耀��m���l]W"2HO[�i��.wH�&�b!,*7�%� r�
�}`�̃����n��J��P����Y����rl��ΝĈ��Y�"��	���1�&$�0���"|�Yl�����7�͎9�@��C��ӟ�o�r��K,"�n��B��E�Y\[��S*�M�����>ҞRv�������8N+��̪��4���������-P@Bƫ�g_-F�\�����;���1����3R�1?�Q^�$�Y]�x��9�=w�ԕq<t[n�Mݗpܼ;��E��&<��*���b�����8N]�.jSQ5#w��M�A�QR�����_�@����qt� ee�`9��� ~����9�<#t?tfm�^�F�@t=�Mw����̖�BL1�>aAِ�lݯ�B�3�-W�>h,�X�~��^�F�Ua�,��L����^Ez�\��Rx��+n�'L�To�ԍeM�7} ���buJG��qy�jvۗ�b]��=��oAg;i	r�"?7��I[���� y�����L.������tI<}���Kј��9i�
M�dx���ɨT����%���Ľ�W�T]��/�|x9{�OOe��\j
�(�=XO�뾪3���EMB����q�Q]��T3P5A��8:өEp�E @9�*�i��񝪅������1�z�ݬ�U%=kVe�V&b~&��E��������.��H>).
�O�/��Ԉ�}X��g e�E���*>m�/ea^�ʨg�3Q/ni�)Tmv^:Y��_#(�O�͎M�y�*ю1y�3݃�y7��iPs�	`DE�̌f�����uW���<D��dꓱ0O&{а�坾��-�.�*���sG��œ����U����J*��XPԠ �z6����d���{�������W��H��@p�<+8�8�D�)O�����	��G+^l3p9�D���(1���8A��,�m#C4඘"�ڝh틈�֎4�7OA�K:��T��׊e������Iyt�nIӡ�
Δ4����B�on����~�������w��ئ��u�����)�'ʜ���Q^�0u)7D��]28p}�W>xt{"���E�p�sȐV����d�)I�2�