��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ��nͳ�R[�ظ�_����Qq���G�]~��\�^�W.Z��ke��X�?�I\�zA@���Y"���a`MBl��$���X���/~%�cg��OU#,��;o�w�F�~�wy�0�Sa��qC�$�_됲��ݗ� ���D��.����v��C��k���<�$J��3��I
����<[�P�}&ʁ_m3�P{�
A���-X'�H4Eml�}-���i���[�f�c�:p�D�oU�5�"&�
+�W� �\�� �Fe�V��nv�|�����X�e�(l=�u�gz���^�O�`�y��ѣ����^���ܘ��7����l�"�p�l*�P�.Yb��7E���C��!.�����GSo9<�],�+���%�o�"�/!��&�&��͜�X{o�`����Px\��L!��2��.�<��p�Nj��Ξ��[� ����I"�O�K�k���z4�f:�ޠ霩�їr���"�&M'Y���|����n���׃��s�	�\Fe��L��b�ʸ5zM(6���0�.��)�"�#p�$N��b����d:�t�g��Į1����#IP���PM�C��$�e��6}����`)܃C�Пs�]U�]�O���kۏ�D"�"�G�܀[~U���2V��:SX%�����o�7Wt�,vv��T*�qDHD�0�'e�M��? ˍD�?�5��I`L�aXn�G�>o,P�%�胺?�̱�d��<���Z+ǨO�y��]2�4����Q^���bXl�J�2����C�+��ݟ۔�lU�r|1�:qC&��6��l�hӦyf���dx���P�����6����6�1�6&Jh�VO�M��J�.�y��R٥jR1��}F`Vn��`px��W�,rCG�h��n�h��`�o����*'d���I߿�ή^�}��`X&��8�Fz<�U��9��g���.�A)��yV)j�O��^�n�@�<_�0�:���ߨ^��t�u
�1��{�,y��9�Fo�����}(W����H�&Yz
A��y�%�H��x^"����� U kl���ֻ�s�mO.+�(ZH�:��B*ϋ`��X�Y��z$�}����=���}��>��r0� �@��s�˽�um�[�ye,w�73��y�;��j���.�,}�a��__Χ=�l�RQ��* D�3��X�z�u�gG"�����/v"r˟���)�+ʷZF$�O>�b�H�O[��6Lxeq��h�N-�3�ė˳;9*֣�>�"t@a����@���Լ7�W°��Z.���A�M_�6a6�s��2�׸��)�b�b��%8�s�X���VqB����Y��З�^�}·��5��`��/�qv�G3G�"U ����i�9?��ԓg���D�6/��+^�q��.��n�Pz�F�d/�!��l�
;�Y��-\�
��}_�!q���|����/|��[;q ���:�/ű!�5*��O��w���W�_��my�iJ=�ɗ�͒�G�A7;jB>�{M7�R����Ϻm��Dl6���s�����j� �?d�	*np ɴV�Q0�+�˔ȕ��?#*�r�$��$�l+H����� �FY��������\4��9p�<5/�OB�j2�TF1G���N\g>��l3��	�6rz	���M���%��f;x4�[�Gʝwrl�BF�f�7�,�?eM��q��X�--z�h�/�W��Op�s�?t�kb|�>�E&������I:w��j�h�y �+#���X�p��A_�Ѥ��T�����G��F���H��=���Uq(N���s�a��ﾊ�\�w��t�E���_��G�a��=E����̞��m��X����R���,Y0x
`5L�]�2����Q�An[�#�0̋1���/�3ΫM��L��W��+7�IG�r�\�f��(�:8͌0�4$u�<�;Z�qv��ڙBF/����)�!��:\K~p��˔)���a&�e�Ǎ��� ;B��ƅ�s�$U�}7���q9��,尀-�{_6M�#���b��[dW���=,����p�KC-d�d*���Pbo�mYMGՆ%B�qZ���T8�엍>�^c�Ɣ 	���_(՜�T��h��ev6.�<���E�@�����9H�}@����p����I��@Y��h[��~a(�ǡT¶�_Z��V�5��7��`t`�� ��� �0ئa�rY��ݟ̂�Ü�jW��ʽD[���$�t�ND@)��d�d6%�L��g����7���&�J�U[���� ��cXrE����~fk�UP4��8b�#V�N.uIՎ�cM�YT'd����:�uH����9��O
�`J�Ϭ�ȿ����k~-�6�S�Co�\s�hk3�}�A@������be?4w��t�b�My����L��Y��$P"���
��n��:�+L�R�ad��~N��\��I.g��r�ذAioV4V�V��0m�6��Ej�p�߰�ot��oF�A��ɣt6B��(8�����(�ua��~҅���ø>��Xrj����7�K��6��<�%��J^�p����߭����ާ6��ř����uy^��;ڷ������Ny�@�"*Wi:�����U�ճ�'�7ş��~�A7��P{��s:*ʙam-�NZ����������������]�5�8w��Ɗ��D��T�����4t�Q!2���p���@�%�\_GHJ�� \�ޚN�g�zf�eE�G�F4Y"����y3�Ͻ�b;y^3�.�溴zҩ��R��[�;�sES�\R,�Wq=��ثA#���o��\�����Ö���!$i@<Ƨb�cT�֍�t�z��yK)���8�������LInҦ^FB��攠S�=�ɿ��V}�S	�h�W�dAnҁ�W�d�@�K�u�oB}̜N�S����Q�4֤a��xW'[X�Z��ٯ�O��s��?��R��La-ӣ��9��?5�x���k��/���/�!P�LG�a�����j�ԏ{������V)�X�!kk���}��w:%�q=�R�F�a�{��t��7�>Q��B}U�`C 0a�����Yog�'��(��ϝl�y�O��_�e����J������3��V=�?+˷y���9I�%2�.�H���l:m�Ӕ���>j��$���0s������[��5���n���h�30�� 90���Q��?��{�Z�^�ʞ0-m��0�ʤ���^�TT���s�]F�%�3�s��^�� ��}�h� %]m�/��_�W�gr�w��\F��Љ�ms���<���*D��v-2-r�X�*��a$8T�x���7�qM�
u*W�&��-��&Y(,m\��R9v�VBjh�����i��UG���<䵚K@��/�o������Rz���?Lߗڼ:(�wƎ{��$[�@�y����7]=��JM�r��}�:CkxF����oO����m-��@K {
.QyI��y�+P1����D'�+�I���$+�@C첩p����R(�(���)��z�1X�-��a���@@����z�u��L����Q�B �,�a�{�7����Ԍ��ɩ"%�꼬�-C?�VI��������р�Z�Y��'iy���dz�dW�Ws?�6E`��t#8/�h���@�Ғ���M��x'&u2��Y$🀛#H��y�?�f�E�V��Tb���_��:��P;�Re��X���ao�j9պ7,p�8�:�S�3is�(s˪�2�A��ϸ�T��x�-0�j�G1�gv�x����0_F�3Րe@?*M�3���K!E*Z�����}��`pB���dwIBbD�-:�]���	C��b�4X�Ȏk�	�vc8�����r-���?����[��eq �vB�^%e��8���i	�AaM����Ӊf�#
��)2����b`){ZyG�3����-��� ��S�|Pݓ�2��x״IZ�����顂��4xD�.{8_�@�����TM��ݳ��`"l@�i�/c�q��l��gèdX�ņ��b��H�q��mPa�����3�U�Ԇc����n����w}7�I߯^+��˅4�'Fm�/^��l/&6fn�p�m���@�}�-��{'���+wT�qH|� ����z]l7+�L��Q3���"�/�C\QC������r6�e�~ƽp��ľ>
�|l!���0%��.��/�����r"�KZ�x��븡�����O����"�hZ�	�lmߐ��,�n