��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf��4Oᐢ��\����Ⱥ�UҚY]u��'%E���i�_s�v�؜�.A5�w]��o�8K��V\s��(cf�D#CA�h���^����ډwS�����o#���V�Ћ$�1 �2Yz��7t�K�������� [�+��%qm�0��C����S1 �ҭ�/�1lZ�`�'84��3u��U��"���>( ?��y�����8$�}�L��w���a:��5��ٞ�=Z��u�=M]�̎$�+������f�S��ȑ�\ipV��N��t���Ѩ����ī��(mNZ�l)S����h�����Z�ƙ�5ϼi�ˀ��|��|O�_2�G�Zh�d݊���&mvMP�3t���u�G��_%v�W��g�=[su��Y�+�DƦ�c^�o&+=����������n5zy����� ��ē<ad#�t�"lH���n�.*)

(��^��6�#������}4^��tWP�i�Ŗ���i��o'{�[��L9sz`}&
��(IG�F
b���Ud�쭣�j-���_�5D�������u�����ג��(�{��?E��E������Ei��H��E�~�Z���=
�crPk~V��,�՚��[X*守�N�� (�� r��Sb�vp�\�2�
�u�q�*R��g4{ G׼�_���Up���YÍv��2�/��9�� �Jq-��G�gu����q,Y��w囙^e����y��{D���0p� ߺ�He.��u:`��[�+��_����DDh�u�7}V��O���J԰�*s�%@Ρ|���(�Oh`���x�%��o&�8��A�� �������Ό�:c:I�]f�8�b��T��2
�-�,W��߹��D|�����y��!VV�j}�@��d����T��4	0����'������H�V��6���WD���D�@g��t��2�V]��N�p�����k�e�L���ηR�FQ(dROׂ���ȗZlf�)�+ ���� r�W�Ь=��`Q鸈I�����st�L���C���$�y���qh��NC�TMg���㕁c�PD[
�hc���;yn5
��:#`ƹ;���8St<�� ���d����(���:g����Bf��J�`N�?�_��bC��O��·Q7�x�ThJ!�"o�?.�R	f��2������GDe���� �Ӫ����+VI�~&q�c��:�?5i�!��^"TAF����n��`qm`Ul�UOY�C�L�%�g]k�k�Z�fMT ��o���%P��Q�[���L���ž�fXL$A}n�ː13����.�F��ƚ�7���'��q�F�O�$t Wm8��T�VXY:$�t��*�2��D͛�خitp�/^@ђM7��r�U�t��������#��,�0?���W��*r�Cދ8�:L�'�"���W�/��SjL3^��'9p���N@~�ҟ�+������I�X� ��)��>��å��V�춍hN�ǢƏ��S@a:3H[G�2��7���u����_r֛9r؇�l;���<��N16SU��v�����Xq����ξ�	�L��?D\��uDO;O�Q�!��;C��P��m���<�:�`">�Ƨ�a�Ͽa�8��1��J���c]ՙVZ[����3�7�F�4��]�P�e)ltY�3Y�q�2I4 Ɵ}�H�Cc#Xt^$oNY?w��|L�q�w#��8}��i��+�T֘x&��3E�%!��X|�{�L<���9'�+_��B��Zm>��J�/L�?��E��W� ��<H��I?Bͼ]�h%�Y�ʞ��_��꟩�L�OOٞ��q��;�梚�h�rj��I}�Џ��S��W�L9�B�>��L��2�!��r�漉�NC�_���)������� u��X�#�bR#/���Ї����FǑ�1���\�4�����.0��f�*���0⠝�Rz��4��Jl��&>�C�39-��O�4+�V|�_��Cؘ1�F�����!�$
hp_�?�#�e��CDp����'�����L�E-�Da�G�q����ۖ�(j��$C��o�5䇖�B`�h�u�Į��NB�5��Ÿ��-X����	½�s��fe��1m��D���DA+�'�_�)�
�%ߩJ�0�� ��2��BA���*�pS�l�zȇ�qv��NC��������x?����p�f��muM&D����6��$I����l�74K�o�Μp`L-��yY�7�2�Yb�a&V��U�J
���Mh�Y��?W�b0ǋ�;�f	m��=`(���^ߕ���v[q�����9�R�pYC�]ֳ���V��7�;�pdXB̺<�B�֧<��x�C總ݲ�ʚ}� Z��m2w+��I���v%�]�2C�1n[:e^%��t\RwV�3���`�l����Ǿ��!N�L�yM'�|ɽ�buf��ry��i3M|��o��w/�;���#��P fj���|r��s�.�ʤ̠��}	u�{���Y�Iy�v��"�;
����m�=�Ax�!/d:�q�%����Zy�!�Vr�t0٬&�[����.�J��scaKR�q��;z�h��Z$��1�:���tͿ*ċR���B��������W�Ds��S�d�%ױ�K��Y#�%�<2 �T��>K��<m���?�ޯs���¶A�+����*h�x�Nfʎ�'r��k���1��C�5�����L�KDl%hp�9C�*�#:��/�F	����2_%7i<--��&�x_�sqaj�@F���C�_�~փ�"o?��[��,5�7Ul}�1����Lik�,h��EZ�$�`Է��-#���;e����|��yE"\V����������$�H�0t��8�R}�L��w�QΧ<�jCJ7MVV�ӧ�А�#�GD@�^�MV��L/"DZ@�q�8z��z_��nݩr�/E���d޽�c2@H����)j�c:@ϯ>#x,�{B����z)��(;��/�U��/3�a�s�d���UⵗJQ`o���kͮ��o�c�-3�v$���s�>u�Jq��c��!���z��^3�:�;Ϟ��`���CB�K�u��{�)��RO�'���P'��"�}�˃�o��D�ؽd���aru�R�Z�$8�`���3�7�yjY�W<���UO�?g�G�0���Y���>п���� y��O`�p[���k�nɢ���4�Gn����W���+��K�iog�϶y�a�F_<�w���N�^�e�����9PN�5�B��I��r>B�H��+�|�Rܒ*pz���?o�z&�2z��3A���D�T���&_���F=��೚�\&Iy�lg2���#	s3��ܰ��v�ԙ@kjT�M�̊�N�ɐ���ט�+NRcz$���v� sJE���!>
��«dZ06��;x� ���S���^�W����g`K)��vrs;}pV��a�;� �c�u�����p\���9�g�tk�!ɡ@�ӫ�b<����:g���P	"��i�	0p~������'x��
sR��7[Fϭ$��A"�f� R6U\)b�ꥂ	GDXY|��s���Ή?����C��5F��D'ʟ\��'`:�(,�oښ�L���%K6���<�|x�!=�S�-:<�`�vM���-�=_��ؘ��	�[Ix���I�Mݶ�� ����� �6m~=Qaa$�<���i@�N��$7�~&�Z�H�V��h��AT�z\Zڮ��c$M<ɗm�_g	�G��wbCF��YQ���<�����Kzc��c�J��/b�Z9W���͟u�
y�U���ر�~`I�=V�%�l�UA��6��{9���-�����i����� 7�"9)D�e��x�e��Q�D���K�Y��Fa��>+P��P����v�,I�-�(���:gޝ��LS���@"p�x����'{!���R������~VI�@�m��O4��f�$*�^��7 �ܕC�6�~XB�:��I�Ldx�2:���ț��[�����^��=��	��9����~��l�+�{�7Eo�,(W�~����HDI[nX�=�R�kt�%2#H����~��饀�Ծ[7�uV�{�%kA�a-�l��;'�Lo�=���� [�l�thm�	?`H��d��n�N�B#Y�ֈ��JPnY�TW!�ѐ��K�@ʘ�|+j.}rt���n ����8�yi��fu��ޯ/~�Y�9����yc�1�����^�u��
mШ1b�����k����Q���S��eo�'v_>˥��G�x��S���o7H`�Ē4T<5D?Hoz6v�g���d������ѷʓ�̘�j_�ЕB~���A�L�-댉�T[j�%K��ٛ�9�8T�-4y���o%���kHn�<���+w\]@P�4y���T;ni��7�;�ݱA_�hg���k\ @[.$�W�~��$[ghyƁ姍jj֙�]���ZlGs�Q-�LNP��"�Xɺ� �4a�Q��)�lf"xT7%I�7�9T��C����s������@�g��}�C��!i�d�D��iA��
�ڥ�f�E���hv�~v���C�LS�s�����$�]DL|��0\wr����ia-��'�u�D����<���2k���G���J2;��T�f?Z~v�'�?R�G���P���eY���?0��68�h|]vv��,�d3��-D��R�4��s.xۺ ����@λMl>Qg�gˑU@��n-�(,��y
�72�ˆr�pl1����ڇz�l.�
A�)��ۀ�f��AԞ=z���u��]Lԥ��2�Cϝ���lc��%7�U;[W�V�}'���Ӌl��3���;�W��,��
�����<���U��c}$�.2glBC�1��ÁA�.t
�m���cx����ʤV���r�ݔI�I�6������x�����s��R�W@PX_C�XoGw7����1Xs�� ɕC�B�LcP�Oܼ����=�/VE�P�ۡ���1|�22@^fR�y��o�gA4��MJ�:nR�����W;H�οr��1T��C�n����V�r�?���3<Ɨa"D�h�+�v��kD��(�F'�@J�v�0��m�]�Z��f0�m~Z}��K��~%�w�J�R�G� LGDLX"
��4X�Y{B�y�V�Ju�/�^+ ˌ�s_��n�u������5�y�	���+6c���j�A-+�"ȵ��5�5�� (0� #sD���T^�k����u�0��h8ɪB�3��+=�n���p~�,�F7w�Z�|�,~Dӆf\�~©�K]Qg~l����c�k��q%��]-LTR�nL\���4�e�o4K�Sv�v��ۈ�5~x'�9�#����@Y}/�R՜�o�
��{s����t�"�_Kit�����a.ZZ���a8�9�Ԃ�^X\Eq�����%-/�����ߦPn6	R߶ƃqC�'��Ï\�$;y�K�����.N����a�7*Q%ث��d!�m?�|�ݾ�q�0X�W�>;-����	����L��x�>v��b�g���z[K+��xU
$�Go;Ģ,�(ۚ�0`��!
�v� ����97���:��T0�|���;ч��
�x����MD��N~�ٍ�� �#���}�z���Ê�r�D�ïվ1�9e^��a��jrL��Y��e�	�~��a�˼��1L[1eLQk���1Dvy��;lƞ�2ӊΫ������/O����ʦ�K�(	�pL̨�:��u�RT�e�����p� ժ2�]��z/�=�"(����z�L\�R��R���� ���-Z���	R��9��[9��/�=*�F��L빍�b#���l:�������+�z��]���\�a׎��Y��Q���h����|A{���s! �,q�X48��b�2����j]��~�q��D[������S��`���-<<�%Z,+���X�Y+%`��0@����c��-Q$ǂz��� k����+�WVzwBhR�Sb2��N#��g��&����[,>��+i��5wT�=u�d{�d<\�q��$&���;������Q3�*yT�sP�b��Gd���M����l�U	mjJx��=R�7�ݬG�r)`��A�ih��PVb;����Tr�Y�e�;g�w4oI������˻�N޲�$���i��A[�UcgW�@@�;ͱ��$n�\[���N���=o�c�jлuY�,��Z�'��\��A3M<�����kG�_�4"s{NO4&�S�Hx�P�j���`�FR1�Ky�7h�����ŏ^����G��vcJva��@4�(S>�O�r5����n��Ӟ=-tM�Q?�z�m�����#�Y$y��Ӽ!B5]����ԏ���f{M�fi��e�wf�����I�� m񏽅���;	SQ �0A �cT�zt�y�*�O�V.��+�:O���Huޫ�{W���-IKe�i�H���z����xI|^��rt4���^G���͇t���m��������R�����'��8�p�S��>�V�췉@�\g9gq���gb������(�hd���vD�Ȋ]�^�h:]8U��*�����M�R�)����p�yE5��Ҹ� p�[�:���U��]�˘�K/]F���-E9>|�	������Il$��\V���K"��G�~
|��zx�v#�ֱ�(�y�S
��}��q��b��.Ɍ�o� �sz��>�g;820[�s�83���H�}t��w>ڛ���j�>�����p=>���m����>&�ጕK��z�9���ϯ����;��H�n�v�!�������Ufih|�Y
�j����L�\tZ"��zAv��{/�6#�Һ��ǧL����b���/к0Ç9��_�#HG�����������a�F	���*]g'���n�v��U*'Bg�O���J��槶�����:�=H�*!�8�#) !eM�u~���Z�pm�0O*��n��yp
�"�<����;�I�㨹ȶ�H���i��羅�%He%͝g����ͷ*�;#7p�ު�[^.OhXhU��:�/�jE*�RF����[��_/H��e��o�y�{�t�V�A�`���2�9���������n�r����G�ԓ�no4� �L��m���jSe����<~$��:D�u���?��s}�'��_L*�d���}�{���>~��֋]�CD6J��-`O-֖S�>���(i���W�9a2���µn�u1�
s'b��Oo�ԭ
�Od��~�FR�&�<���'iU9��qr)#�V��zS��t
}(�rqa)2�&3�2�F�V�2Z��t�"�fg���i94�������Zd���V�N��T�9�Y"lp�i�vu�MK�*`i�l�E=�¾RuCZ��@��tA���u^R�Ӗ��{� �o�òp��'B�pu�K�������]p0�r�Ȏc��#�
D��X�.;gK�H]�nq7^u9p���EU��(:XbpZ>�	�"V;�?���u(Rc�<�S_*������fI�^0�Zdz^ NUY�Bs]�r�*c�p���u.�W',��'�����g9&Oް��5��;U#�P����mFB�dA6���#
Թ�p�`o�i���W�� ��1�.��Q��U=8g�������ʹ�aVIj`��65�P��=OAi\�=�B�����xq�l`v4�Vv�վy���\Jˈ���
]�RM�h��78&F�c����nC���l�9�RԀ�Rw�5t���=��49�p���0�2*ڶ8�4-ޕB;�A��H�(���E��	ڠ�˦�Ű��j]�A0[`��qI�h�D-��ggtP�	S��跧�M*�kn���ߧ���ߡ��R#I�7����l�jb��lf�[��RE���enP1��Ҡ5L��Y�ېD�v)@_�cv��}$J�e&����Q�vjn�x)xjӌ�o�����Q�u&�^Q^g>�9�s���H}�-A�*�"�H��P�'(j��H���V�+�k7�=�5�C�0]Q�<����S��;}I���%P�/z ^ ݨ�������J��B2��vVZR�%��e��P��\�ؐ�����Y��#�M���B&H�[���r1Qf�MT2MU�/��M��S[C�2�!	���XR_�?��{.r��nuqk�f*�MN[��"טd�)�+�}���@����i�q��%29] 
�����A[���c
�����N�D��h���x��8}�.�@'��7�.%+DT�o�@ZE���߲��q��Ȱ����<,"T�r;�+ƣ�EJ��Lt���B�g^�y��=l�~���{zy~/́��:�J�� /����]��k���S�DV�3m�	/ �;Di(/̤f����`7�Fh�_k�v�5ߛ�s�-�	�"&jﲞ����ֵ$~���?N�3W�"����_�vj�!#��c4�vX�e�J�(��z1���1�޿�����,Ї��npL}�o&��\��\R��}��\o�tw��F3s���2�5�����'{c,�cP��.$4`삃������Cs<���)�E�9w���Rn_�͗MC��Vl�jّ����z��H9�Uׁ����F��t�MO��`����h?��5V���q����)�oְw�7P��=_�����|��T{�P�\�顒l����w�(����ڄ4V,r�������	
���z �,3�W��]�p��̞wɖ�Ќ4������j~� �l������������?�r���"A
9 �6C��ԋwB��!�Ʀ�A���Ȩ�C�KkAo���`�t����Ӟ�Uh��HĲ��h_h�1->��@�P2!=&kِ�@��|�H[ҁ���|�!�"�A �ƻ"�{Z)���@"��r��X�8T���<Z��Y�Y[��ʏ�۟���1N4q�Ļ�f��c�w��p9���@qg^��h_T�Z��q�\�bG{�B@�纚̗U���ڹ��~����-/rۂ�BC��"RU�*}���a9��)&���T@�Yx�)����GyT~eBc�Լ�вz�x#�I�8�Zx�CR.]/`�/�Y�N�
�ΐG���h&�m�(ΙmH4�S��ƛB�si�k'����*�L�̅Q�"A<^5���9]�ը[�+	�)�������H*uTҞ�#�k�����n�p�KBٖ��@���D��q%�$�=���'~��.aL?9 ��~ᕣ������c��LYB����K%HhP$;���J�B�
���7} ]�;Dh����;_q�|A�k��g�T	lC�5�Bޞ��Je�B}���H����t+J�	�5�-#�R{ʋBX�;�},O�`�з���K]��'�n]X,^o-۱ў��gW��#��Sx���Ԛ�Cv[���J�\���C{�Kr�/Y���׬4���.�m��+�^�,3�`v��F���1E����Ź)(���o��!�.v�R����	&��Uy����U�ߒ�������0���Z2��:���_����0�i����4S�H�_1A�1V�u2z�m�Q�ŀ�ַ��~�4!��@)��/f#N�)��|�C�{�3r!P�ч��b��G'[��I��Z�s[��=ᘤ��nV��}*&sv9
b���Al!a�b�����;8�/1�A�=��]����HlT��E��>$��PPqA�#	Nx��TKP�[��8,߯�=��p��lO�l�\��k鸈�Z$0�*9��	CH�-��� �g��Z���< ��~�z�E2OB�%��W�J��{��dl�Z3-�i��3)v�-���	b�}/<UFY�]6^�(S���x�U��#@�Mu�?p��̀6����l��"���
��oH�~��0��,�ö~��3������pQ�R[�ol#��q1&#�=��+6ŨW?���M��ٵ��-I�O[8[�7�e��[��i�]L�&[�vmK�!�_�ܳ�.�d�wb�<���}K�<�|���O�W�t���e�c����<��5g�b	��������;�c���.�����IR-<��R��Y��BM���zX���p��j�wA���T�g�[��D�7�0��s��KJo'&�N-ge�f��cރ'ɔ��i�Q��c���ֱ�̅���6�X��kzx:���a�d���`��9>��3��������"�ʳ���Y��y��׎K��݌i1��e���c���fL��[>l��P ��/s��cJ��K�
I)!Df,4#ص��á�+x��z+f�����D�<%��#�{n�o� ��,��+	�a�my�VZ���3��i�s��'��5�̼�2>��v,�{k���{"=�y)�ǉ5��T��no�嶰3��Qo���t�2�ΐN�p���X��@��U%#�k�Dŵ[fl�3d3h�գ�MO=9z�_���~m�ltϓ��$L�}���Kq	��`���*��m�cU�1Q$k_�Qv����·�=�=Ԯ���S���n����C��"�7_�&q��TT��d����(y�+�E	��m'��_0G�7�o�ArJJ�pR�����ő{[_�m����4��j6/G��0^�!7<�
�� f��]`G�Ɣ�X"I��׺��ъ�����Z��٥���ɱ��2���P\o�\\��d��v�9-|Ќ�C������"�XBJ:?�%e ��d�}t��k��CF�0M��v[�M�����1F"} ��t6�|�_�������0�E�ֲ�,�ݩJ��jΘ�0j=q�X���7 XU���fN.�M�t�]B:��k�~s3��meO�Wc;4@VZ�����I�V�+�G;�R5|08�_���&���s|�/C5o��y�]F��?��H�c����%$9�xѳ�%��� ���:�}Iey�1C�M@9k����@�+v��cn���L
]VEr��x��_C@
��8l^���9;I!�jIװ�Y�.u4l�q�)Ⱦ�ۋ��Ĕ���̧��u���5�N�n��zD�K�D%��^vxPF 8N1i�q��z�P�T��ތ\�qt��9
E�Gh$�!]��2�7=������alh>���d�sSl�vr0�m
����p"N>��PS��{d���7����/{z�*�]ZhV+ȯ&�:��s�e:���]O��֌N�s���h�Ǧ�.|��gk8@��!�C���&�:��h�c��̻	�n�������G��Q1�"J:H0P�^BF�� 0(���3�{)����D�E[��h*�/�A��y�'�\c;H���@J����Ͱ^S<M��{Qpi=�BC�2��/OS��q5_J���)���8b�)�W�?���|�Y�����6]{)�@Z�A���Ғ-��wJ��!|�j�-�ה�(��M��Dۃ��$����&�2B��-jTl? �a#�Yy���P�h^�w{�	qĴ�R>j@63w[L8�@4�:e"?�MGH��	*C�=��}�x�`3(��܇A�
 <͕d����tn�^h����!h��Oڭ�F�[��YVW!�#�$�9��j�U:�����Z�o�����}�c6�ʐ�6���X��2H<����������V:�r�~C��m�7��=�Lۙ�7~p�P�nq�]�m�q�3M�R!��	��{���r�����N���
>$���Z���P�-�q5�|����N���$Vqpۮ����rT�^Up�B���K�e:3�� ��&��"�c��z�7(xk��T=�/�Gh-��������ޟ�2DD+ �+���'���� ��>Ќpb�md�'N,��;ss�?v�ʸ��=�E/�/U5�%�rF�v�a0���r������׆gvC�����ƅ?�EʏP�wl���H2Y������H{��: ��~w �aNFE��eiʸ[OrF�
<�~@4�i�)�4�}W�w��п�m�Z�.�_�,g�1]c���`2ǵ�D����&I���Q#ʱ���Sg�G^��!7��Oo�{�y��Y� �
n/� O�h���_��OH�X��x�>j2C�a�װ���z  �.�Lc�%F#��R�l����:8Ia[�%�k�M ��VW,,��d�y��N�>�a�#}��I��Uf���,E�ْ���x���RX����;z.���E���
�'��Aڴ�&0��r�#�(�V%~{z�x��� \��ͻ�%ƈ��2�_ǝ������ܝ;M��G;��AD�b�\�����9�ow&�fdJw�_j���Ij�aWR
ݰ�!�}�ݲ��Q�;�g�6Y&*��(���*@@4��5@O6��v��"t�A��(l��.ږ�zv����L�
��`�7�%^�q�z�w�S�a��aJ�J�PO�m"ʝш�� �_���巪��qV��kFv��le"6��%ۜ|F�������X䷄��֔�Q�la�����0x��}��D��e�_�bCƐ}LM�B�g~����G{�ޛ���hdk��3JO�)&˽2ה9����M(��R4�� S�<�m�`�8���%���s�JW� �Z:�͵���DX�a����~,�6F��"�h]�ׇ��5���h�{w�_���<֫�� ;K~O}������4s�px_7��d���#8�� Bp�������w��sc1�n5ٹ,@霺�(�xDFV�M�f]�qѡk������1���p�+(۹��1\�}`��_jV�����8)R2;t��S� ��\��q&1���FJ�5L��A��K2)��o�!5ֱ`���w^� �ᠿQ�ɩ��ek��@��=�Sn���uo��(�8~��R��62p�
Л�O�|Zl�m ��ܼ�ܷ���~���*��u�k4]P&���2b٠�8kYLR٧��0f��
uV��2�8aK�R�X<����#:R_ϏﰋKn��[9O�zš�4���U�`#��r���fH�F�+�.�>-�N���)��a�z$�i��?�<x�f�:�5�&�`@���D�X�S�y̐�4\I����Di���2Ӗ�5i����d'�dK'P����a�޲��5�rwv��]�O�2w��B̩g^r8aQp�1$���*�CeQ;��Y�a2��+|ey�?K�g���� ���Q31l���.��b����x��˯Ye��y����X�Ѥ���T cx��B�삏eX���I�>Hꢛ��"���v)����,������1�f����wz�3��k���E�1c���������-|��>��$Ԝל�:��951)g�yNo^*�L�.����n TI�8��Hdn��1����+r��ݱ~ZcG�vD@�2�#i��i�9G��-ꀭH���{�ɗ�}�W@�,?�!�!ώ��ñ��}�c���%��,�jYi�Q!g���0�Ƹ(��9	��xF��D�� }<����t?m�W] �ȕ-���v�ܬ����%�O2�5�+ݍ�3��sf�4`�vL߬��ƹ����)T�"a}�b��,�aI�-J`�� �9�f&���� �G�W���ѣ�w}���l؟�kTw�<(W����j���=8���V��:���U��_��5--�0B�۸}7�W��a��h����ƋF�>D��F�\\j^^m�xl;�e�������4Z��y��Y39��)0C�N�Vӷ�Un�[��n7��i#�[������4_h��V���5�g��V�LE���&�f�X���`f�k�v�D�j,�5�ѳ�,��xߤ�7B	,t?�/��_�[E�N	��%��b��yN��YI=���v�m�vEZe~%��\�8���޻�ZHݠW�wT\��ц��|VZ���'��P���I)Jz5��(��Bb��|�'��@�-l�;�^�	�Rh�S���N�2��Ƚ`�0m�v�m^a���8{K��$�xt.;"O��a8�ïc�� ��R��6�mϪn_��+�9�?E�&���➲U[��F�"U�\��W��m����G�s,�Cw
�I�R:ՠ?\zo��_K�,W�=�zI���߈�ۘ�\���r sVa��]Z��􈐆�`ݼ�=�0RI$������T�v�]9��l:J9-�N$�ꌬ�-�b6"5��5x{�h:�Q�;���d�Zd?1�2!m�<�I��U=�k���=����꽜���1�D��1�ag;\��dK_��#���v�*-�7k9s*U�}'��?���Fh����E�Bő��/+֨"C�,����ڪ�������9���2�v�R��a����;3������tr����px���qp�*���u�b_�Шt ����NG_ �N�3$?�j����g2;Fji�p�{yS��O
��<wO?�/�]���:�HEh���f���,,X�ژO�5�5/��(]u]���Ȱ���{b��-���"����  ��o)#y?���BO.��D�E'�?��gZa�qm���r��3�d{��k�*ޥ�}6�`x�/GRX2	<
����#l:_1(�KSA�Hx0��`9v��C.{<"@�7�n����V_�˗@�T��/�5��v�@�X�ջ�N�RK��::�����c�b�h�.�`\��r�h�]ᰞF��w�?�̷E��C6�f��WA���/�74�`�.���_�������k-ӽ�i��π�k�)J��p���軫��C��Cx.����&]jf�݄nH�`�� ɒ�.HTů q������M��ģ||z'j��=}N�Ű��2ۧ����N+n֕#��5����F�s_D��O���P�X�U�#L����1^p̢"�P,�����k�|r�������WeP��I^�@0n�6�y�\��,��X�.@���}�Qr {���1��7z�ʓC\�?����4o�ņ'\�.vSrN��U�?�D��F���h��QQ�>h]{�g�(�񫎋E��\҂�p���wt�▪�������,�P����Y}�F-{�=��E:.��������~�W��2@�/	�!��]��M,$�Q��
u�lLA`��GJ|�C����
��n��\Æ�ڎ L�=��ӑ��-���x0�/G��'�-��(*Kh�>�	Ҫ�VU�b������̡2D'����ذǦ�8��3c�3�$�ęG+6hF�+5�H!�6Ef��[�<��$��M��S�Һ$��:M��k���[	�'�f�	�� ,���`�Vf?�=v5��T�(�\����TR��k��w�!7��Pý��ꉑ�x������MO�A���P�A�_�NYI�����n�A����ۼ����F�G�Hv�>�T�[/����B�:��"-Iyg(>-2�������9�&}I� �&���4�.p�y���ǧ�~Τ(���p��l�x���us��N$%b{����?�B�$ͣW_VM+���"I������_.�W��Ah�?��B�۰�2LO�ڒ�jj���voʁ�VTݟ�6I��g��2֮J;�9p���@	7E'�VoS:v����9�,�z̡B􅕰�Ԍ��ɑ�V��3ڜ�"��A����Q����	��W�E����jm򗕻p�� 2����qՓ}�
�KPz��xu��K3���
*�ëo)��=�,ǲ�?��яj}��'�^?�}��e�&��SxF��B�`�~��G�ׂO�����o\��\�I`���C/e 4aK�-5"�6�H4]#v4�����c3�7�z)����r,<����iI@����� $�a�~�D���X�  �FD��P�C�6�����GCL�T��8��'�7��LG��n� ��\���>����^4�\�6���{�PI9Ӣť%W�A�%j:��/;B7c3�D�y� j
��u�\T��7����*�+���x�E�s!���j���q�桒1�C�Nu�1�u?$�m��Kۀ�ki:xF_ vD�_�fD'�N�_���� ��󱳜_a��Zҳo�i�>��ҡK����0V��b���8�����(<c�b�҃<2�����:��T_g���؅�z������L����$J��k2@�F��G�����l�����=�4�49hӋ��=�C&�9�pV����'�ŕ�0싶�́�C��לL�B���Ny?�)CD��ּ%>�ϗ��8��v��7g��;	�A�}���8�����XGO�jT 1s���P6�o��%�:Y��m���A_��a{���3�V���|p�>[믪����.��!NQQ�g}�3͡y�H��r��u	��|�\.�)��*!�ZƼD�o����E��ݟ�~�W�Gb��A�/�����{ӕX�ݲx�ue$|�_�ѣ�G� sf�Ȑh��'�ڔ��<o��5g���]�{W�YK#D��5�DV$�$30�98~dQ�Q�c��,.�_�|G�9nY|�&��&�KK�<2P��$�h�`�E��[�<)�_�)#��Z����Y��x�P�'��0�0e�X�#���*����sQ�^9�F_uf=�"Ҩ��z�"�fA�˨u���ʇ��`G^�$�#j�+h�M�X��x�fG�veRi��nt���-oz%6��;8��.�M}���j��~�Ǜ��rY�L�r�C�n��nZN�'�uj��Z$�Y*S�k�,wVӑ��'�j�*]��OV�m�|V����ぃH>g��e��
��4s�Lo�tHJ���%�U��p8���潲��P
0��0#�F71S�e�^���.�u�{�T>��\�k�U$���a��ﳕ�e��`���6=ą��|5�w�S����V[���̪ʑf]�A���y���=")ز���&��	��`u*r�������sS�V�u����{���C��w������Z5`DV����gI0���M=�
�j���D$_��z�A.v�L3
�RdǃZ���
�y%+b�@
0�P	|H�[(���.r&sO��'�5�c���*�=����b[X�A�핂��.	���on��%;̦sUe>v�/P��W��Ks�V{��t�P��ӊ���.�w����