��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*������j M����J����Cw&�u����Dg��>_�,��o��3�9=]�sn��5���A<�-��Y�,���AU�G���̻N�	�Ϩ�g�ϵ�w�Ω�k���R�9HO�o�u�(v�W�T�yVL �q^�Q�0/�����)1�cڵ�E
�W�D�t/�Ș���~x��R�X7�]0|��?ͭ�m׭��e��%\rN���H�i��8A(_�P��0];�ű
�0
�@�=�eH��j��闶�|���v��U�7��P�1(���?V�w�{�'�Uj�(�^/�Oc����\����+D�lDM�=
<k��y�t��8f&��I߯l�I�ZH�b��=h��<�e�nu���x��}h��|ǣ���`^�Xl��4���i� ����X��5�,���=?P2�Z��5��ɇZ�x�v^e���7� r8�(�������&�d>�WEp0�("����uD��nrȋ?��~�Fg �B\ػ�L
F��Ѓ���-�#H����0��^�T(�-~9K���>W�:������<	��i���ܲNy�숖��!�=H��Vt]��NDsӒy9��_�Hf���vF���-��I�*����3����pE������;G	�b�s����kKCy���=�9�i���VM>Sr�1cH����25*�_\��]esi;�>8�z�.X���R����iWU��d���	�Z��T���&++��paX.8����橮��<�flG� �M��J�e�(;�{�Aٓ���x6x.O�<�۸�gG�ޥ
��4��&�v��{J�UTq�!���'��`9%�Je�V)|D�'@f$:,�������?Mk{d+m\���4�+a9�Hq՟�C>�f�Sem���s���xI�a�j���;�6����>���
��y�|����CN�z��i��	���{�SIW(m��s�*�`0�i�]� 
�8����b!P?� �����)�6�z{�`9q�U^����c��Rg:�eYBN^g�o`/̀"M��V+�i�'���*�	�y`���[�a��'��6�!\c~V����M�*F��7B��Wg�Qp"��e@NJ�z�0��dt�^���u�4��5�$������3�����4@ʅ��m��_�^N�Ĺy�v+$�e��
��W����iG��a�����q:^�ų^bLu���!ѩ^����?����iJ�F�0Y�i��I�@���y�~ʽ�TV.9����bSu�,�ư�<�xz&�����a�x�m%#��A�|wӁ�����B��V��y<5B^�j.c���=iE����X��>�\�@���G�M�b�-B�w.�x��,+	��KZ9͵q,��S�-�=�2N�O�R��U�s�ORW�⥬r�����ԯ���.4M��M25��j&�bpZ�;����;.Y��<���?}�e�c-���#�iE������e��G�ǯ�F�4���\@W���{��7�#?.�W�R��Z���ܕ�� ��=�(��6����S�%���0=̲2� 59sG��4v[
%��u��/T9��p��{#j9��tٖ�b|�����ɢO��޴N�(ەEސ�{�X����g@%j6�����v�Έy�:�@&�ag�f6�/��FM�^et�r�$HF�����3ݺzw����	��<�[��xc��[�|%�T|���{���t���|}mji�5�@��")����� `��5�}N�CEX��7�z���@>To�DW�����D�?-�G�Y9�,�Cb�PԵ�7Y,��s�>����.�F��o[�P�@`�tx�&͛�GS��t���f�g�l��S.
���*����K��y��UG�'"
����˵$��B)�	頭�G=Z��\����|��]�h��),=�%�fp�]�6��dU�L�h�==Z��=Y!i�.'���	����Z��j~h��
�8C '�t�d�h�f�R=�55`NFeDSک�Ǩ����� �/�M�E�;��g��^�P���]"�]��@6�k#��?,'�˧ƹ�%0��g������i,?������7c��Ow^�T�ך^�j ʬ:h)��i�0�ӗ���EF�I��E۬�[�DʩĞ<���b�#E�wO���̉��e�2�p��5�H�+E���g~=�}���9n�*-��$w��?�xA� �١)󹓲BF2f��M*���U,��L<@������2�Y�.:5����r=FM��Jp|	4r���
���7y��(��'R�oU��J|���	ѧ�zއ� �*��))��7/�a��'-Q����ɞ5f{vx~:�]4�Q(��vC�p?h�i�U��R�j&U��]u��Mh
�r�I�3Y�����u(��G�[#X�g�W!��Ĥ�� !��%<wHo�	r���P2z�Q;%���!���y���*)G�`������c�ۨ}�A�% ��!���ÌA��oW�m�p�C�?=\(������<)�GK�2����������2z)ү��>>q�T��(���/׭l	��M��eu��
�ݾ��j�+~݃ ����r��ȡ/��ĕ�3�@it����
Mo.j�,���B�����j��6,`Nn��'M��U]��]�(C�x��a:�C#g���`����O�
�&���-� c���r�V}����ڙk�R?D���R^��踰}���U���u^�R��U
�1]X�3��1l��g��7K�3���G�-���Z�� A��Bэ?õ�"�؜�%��ׇ]�`��rM@ð�0��D�bX��-��3���W)@{uO*�!~��iC��ӂ֋���Dy�)��x�,�cQ%Зe��a����;'D����(F�� ���WEHC-M�7����b/{�0����Y�F����T��� ���� �F�^��P�v2�e�aE��#�j#�)�ؾS�~D'ʅzN��P�5����IP�k��%_]�B+8�OC5�[�ůM����Bջ�&T��B�Ǡ�GDxaHj:L�
V�鱐��������OH�dp $Q��,��D�%7��i�y#Qz����.A1�E�����B�z\a�s%+8p�X���	��{�js�����Xk���
D�8B���Ê��������=" #z�����NV�{�ϝpԍ�}�+g2����7��ٶ'��eo;O5���M@�GfG��?��D�����(��v�oi�Vƈ��Ks�-\s+�|�H���[z:���4��N���Oy�z��5��'L[���"Ve<��Ѿ�7���qN���K�v�B	�n�W�g��D�V�S���»��#��.L�!���e^2g]L촖�3�2R�A@�嵒$կH�������y�kg	��A���gu�ʹ�����;4��c�^0z��_	��ޥ@�L���SJh^���
�kpr�˄V��i�H�A;�}����|g
�@���+���)�S�	c G.�����[^�5A��:�4}\��)X�7ʵ[�Kq^WO�{?�$�t���&O:=��r���#�Z��仴2h��*���{X��+Lׄ�@�(l(�	�ha�^_�$�
��,Jq��>9��Pf�;)p*�M��]K����.�iz�?�ue�EPy����Eq�&�<���i�{mp2��8��������q$������	�^���� ��ս��I5���4������ߌ�	=)�B1l}��L��A*�S��8�3���*����Yy*��8���~��jS����^�傂�"��bQ+Q�+/��R�#����99Ӻ��~�l��ӱ]�f��'2�� ^g[C�����\< 6�w�wF�]e D�u��P�DI&��C�E�ݱ�T;
���.�W�)���'DUhwt7S�R�Y�镋��3�5
t��sbc��
`I+ҏ�XLwB�!
��a�����@ }N��;%�"!?�-�D��j�P3z�c���5!����b���^�D2+IX��e��u(�[�K����kF�'EF�5E�;�����
 m�~��y�L�����L������^Uڏ�r*�����^��c���׼��Ê�b);KZ��R�R �b]��&kU�����W�MX�*�����򽭐�U��'�x/�����\K�t<��A/�S��ͽ(�� ������	f=q�l�xh��xS�+ZP<`T� J��y?�s�ԥ۞�ֱ�$Z
`%I����/�o��!/b�T�o0�/?�E�=�Vk���d��Sk�T��C�Ks7&;�!K�rk���C���qi��j*��4�(@������������R������������:{��K��2W7jz�e
����#��F��o�V��Ka ��yLQ���{O��F�0��U�|�/��Z=KKP��Bp�������?E�bΑ8E�BV6�����Y����Gu5w�>�"|Lf��aH��w�̖ͪc����Ќ3�R������	�l�O=�ӏv<ډ6ku����m��|S�S�N	��ȝ�K�ț)�0��X����,���E�]r���IN$1���Gb0�?�>~��1y�Q�]�[
��*<onk��6Ak��PA�4����k�v���՜-�V��:��K���H�ʣ�W�[n}�]��Mͧ��o�×?_���S��N�bQ���<�h�*���Hj��}�e�ZX�!��%���]fÃ�@߱��$J��b�
���H��oqx|�9Hs�:���j�as�M�kIX[��DrN����$��a�]�T�!)�:�x�/�����_�T���S�ؙ��4Q@0Վ=�/%v��G��K����6�f�������\L�~n�LM���+�;�YY�0�_W�i̽I�{�i��ɛ���%+�ouzc>&v�xz��G� e��Z�1I��ˏ�u�dvb��+�p�y
��� ��%r�6��z��"l��}H;
�E�q�]�}�!\�w�μ���IB}���'"s�3xa��t�0��ӂz|��hl�}�,,��m\�W����%���������#��J�����q|3wX�N��<�/U��
8eF=*�Ր_^s�[[~��r��<��xT�6����4�%��<.? P�I<�P�$K���B�U���N:?�.�������?`���� z�KǦ�pU��#�q�Ԕ7Gbo/y��8�H� }��߽�
Vl~SP��5Û�t8�N�:GOU���T$�a��ۛ�q�d���J�kzB��_�;�	��R9��"q<0�.�
!5���.S���4l��ޟ�J��Q�5�v��oo�̗w4,��CݒJ. k�
���[WM�ߔe�(��6����� [�"���x`����u�h����B�N�����?�Y��˩��̮7�!��WזZ �\�j;��_�n1���W�HÒ�k�nO�y.�o�a���op<8U���g������խ8���S<�CP��Vb�����^	���OJ(��ra��YӘvZ�nm���~,��33h��JJ�v-��v���F4�<�'�ԖŲ!k}2����TKk�xPU>e�OG��\�T C���J��I�Y��߱L�)�)�[���i6��� Yr�W$E��t��ώ�l��w��R�7��z~rIod�����\?
&}�Z!4���v��	9�R�se>�X����Aek�;꧿<�HNZ}
&�m2��x������6!7�H�V�ō���o%��'���؎x�G,N�X�ۿ	��}�>_!듿�6NSD�o�����$Jj�5������2"��ͨ�����;��K�!�Bz$wD�>�.�I������l��%�IWf�R����d��x�g��I&pk��r
�y��wY���g��"#6H��H����r�,,�������	->����S6�`�@z�t(�Jy��W��{�\*>�.�KNef��{a��*���V�vR�N�"o����"����E�U�F����pWN|լw��QR�����xi�[��!֡�(aN�S���E������m �1�$]u0*wͣ5t�&�>��VS���9��y�3m�J�7v}<*4"� *p��҄z 43%�y�׺�;ת���O�3�f�����BK�D����n7;Y1v�㹂��c��D�O����)��;Z~�f�2C���{��p̡�j�W����]�CIbc�m�J5����e�����t����R�a��au��Ē�1��84��.
p;J�#2��Q%�e4f)O?o�Tsj[��`�ځz�;X�c �l�rh����D8��̟+WWn`��b�wi�#Va�ڴ.@'�[�	5��9���`헼f����!�����	g�,��p�dL|����(]�Q�����4bwtS��:�%o��ـ�y�C,�B�a�m	��B��z�^�F�����9Z.F���^��0���;ye��p�6%+{&T)���8{71�6
�^�������^@a&�5��-�Ë9�d��s�<�o�*f	����45_���બ2
�1�Q��������8� ��NxUk�g2E4�&����z�G�~i�Ql'�6��p���A+��q�}�д�f�Y��v����ʖ���x����Y��,��:����8���h
�C����by+�{�Zl�>Tl_�jv=R�ПCr&Տ�l��`�ir�� F������2�P�^W��9��]�2�ꋕ�	��De���P�8bu�x)h�~�������2 dTL�28���=�F�ҙ��^���ׅ#z�ʙ��?L�o���ǦC�s�H��K�4���P��m��;0�O��ס��[�T��L���8P����|�:��;B�ߔw�1�2�m��:)Q�
()��aHu����?c�o�����=�y�˦݇k�v?{l&�����H����,)�QX�2�����Q^����	���1���H<���3���D���N�weP���\��V��a��ԥ8�?\_�0�t%�Em��;}��ܶCT��XJ�Y��ƺ�������5.���oVՇ��GB����ud	�m����ģef�Ȧ5	�`�\�	H<�0Ѫ�z��S�F���AO`��N(��E�#dx��C�?�����2��Is�4N��c�0��f�p�	��'�(	b4
�����Wa�Mm��DtJ(�q�uBpf��¯�Zy�R@�7-�2�8%�K�W����C�
�08��bv���/��M-��̈́9Cc��z�v�b�e���.��K?.��xwa��&:���1�a�&���,_����~;�v��m��ů��d��;IFvD��a���f̎�c�&��yǢZ�M��痴ᣛ6��p�O�M���``p�J�n$Ną ����4����`Ɩ�V��Ϻ�{��3Zϥ��'�
=����n>�w�==d�@7Qi��G��{o�R���[U˿K�D��.a�i1ir|]@��Xq�˰��([^Uk��	�5�Hqv<��:���ݳ�!�D`�[��<=h�a�_�̃Ҹh�k�P�VT�*��P��`��[����񡫐.���7$��j:~��<�f�1�I��R"�3>C����]dQ��b��=���e��:"�Ky<	�e/����A8�,�Z�A��d�g^���!X�Y"ѳ�'�8����8k�*���߭J(�*]�z���W�m����+[�O��"_j��/��
e9u��[ra����7ǮR����������mz;g��5�kBL��
���V��v�NI���l�+�n������WnK��[/ǭ�~�.�ǲ+S�^
��e̛׺T<�5�/�����2�������]�MҘ6�������U�R����/�m��Ǯ�͠]�h>�ǺP8�p�!Dcdx�FY�/�c����ϐ8�aP���ɝ1�".�I��4��I;�?q�x �/�T��w�ތ�i�6|�	�U����e���z�)�|�ghvLl;+��r�$���n�N�R���3ù�������x�����c�H��*ō��H�,������F���{�,�7N��sC�$�+#��
"�.9H����?`����M3�si�j{zR��qmF~Qu�/:�z��a��a�>�͠N��jzvY0W�,���#slD���&�t7"g���Z5u��	��-�\s�hj��[��V���n ���RJ�=�3��E3�Jb�e�K7¥���TL�Y���"-(Z0��t�F�Åj�Q��q��xt��fܕszz�r}]o%��V���ʁa=�vEYv�M�\v��YZ(�b�����i��m�qe��/���#���s���5q��f�s�����v�m�V�_��%N*e��s�[�NE�Z�<�g*l1���m=څ����gY�|A�S�7�b��������<[�#{L�� ���$��C�'=� 
7��	�h��ܨL��z8��Q�	|�r�u�_O�+�Y���!�jE�Ia,U6���Md�&e�a��}�@T 
����G�vD���pƩ�����3��'/U״��S$I8�d�9�e�hm���
V�m����|%
P�;I^�O�t^�C���S�m�:t��$�	~L�WYQ��j��.��V����nGo���Q�L�Eacӹ�۲E��Z�(yW}�'p�Ǜ����JYi�����Vڗt1%�����ʾ���>S���˼w���%x��1d��1�I_�-���}[�L�x�S����/�F�<�ū��;�-������ ck�z~EG���:+g�VD�.�؍1�\88���l1�["".�)2�ٖ�%i���W����`��%M:d��k�\�q�z��-��x���d�XvVٶ\����L���&�?���&pa��ϽR���C����*>d_,%L�yL�nT�8����s����
"*���a�Va�?l'Y�T����䯸R�a��2�1�ْ�T��e\�~0���9GΓ	Ƽ���	�Q��J��oVUJ)�����^H�R��,KM|��x�C�{��װ:<%�U�/�W�v�r�P]@�Z�Ui�뱦������mNQ[aUT���1×������u"�]G������{|���!���q,�=�r�o2*��� #�,w\zp�o���^�f�5@o�mv��\�g]�j�q䣿,����s_յh�Y���pQ��u3��dS+ţ��&�3�j��}Z���5���P����2r?�7�����y�g�Ps����CQX�v��KP~
1�NcL�0H��T����4����5�<
�b���1��v���dؾ�����0�5E���0����DR&�!P�}v� ���/c�s��fZ츪G������p�Q7�i�aK����xxo��Do��ӝ�A,�ؿY��ə�6P ��ͱ�ԩ�����J��A�2<�UOO��D:�&#�e�-���v)�4����詠�8�������q~<W1�<5��5έ<�)���'zYZ ���<�^']�&i��܆bl=]:HHh|>�S�1���0~:�	Z�gJ-�F�|�]B�0u�_댳�ɘ���No�#BX�������T��<�oUآ�}&���{���q�Q~�.���x)�|lP����5	w���y,��I;��[��p���oUhr����dL���ݛv�X������1閭ŵ�eB�0�����Z�`�J�V�7�H�j���X�$`�A�C@|hA�	�%ЎC�m���/yP.G
���Цs�ԃ=g`�T�BU{���O9��P#��M)vŶ]�d4�tUU0�$	���Q�<�A�ʱ��#$�a)�J���etSL1;���<�i��'rA�^]�Qk�,��g7z�H?��ߨϙ_�~�(���}Sŝ�j�)�` #��^|�wYZ�}��9k����b�`M��XY�k������a��*ߐ��KW�ǒ�ّ�J��J9�� 1�n�
0������iM���^Vl��� �ޅͮ�HL&i�à��EW��{~8�O Q)5�&��|-�)�fiގٿg�xR"^�N��*������������O��v�	��ۣ��i&q��#;�э���i��T{$QM��1��`B��.��1��qȯ�}TW�}�?��確�߯�"��s2��J���6�^��f�[V��<�����V+DۃR(i}Tb;ZO�$iɯ6X�F3r,ql�T��ִ�L�8���t����n�%.�=m�x0�58����1>��}	�B�5�Pɹ'zJ���yv{�e8j�4�mu?��G~{�����-�P���0',Nk&�ANc�z�*�%4W�p`����)=�@����qAbsn�����d�k��-��_�yd��3 }�XP��w�S�JQ?���ؓb���0�4�
zHj�6�a:�4��>P�֓��r$A�J陏S�g9Ǎ6L��j�L;�컾|=0r�������r-x��Ր	R[���%jl�
��h~a1��?�X �r�m��]G��{ j+��9���r�u%㠄��y�urQ��WBN?���+�4��cѢ�T@��R���'�Z�?_Wޖ�,�)�j1�ܯ�E0mr ���PG�����T���y�ud��<�»�`��	9����.��He��?����-�|@����[x���Ě��_��m��|�js�;$hÛ^<c���ϱ�H�I�˝�_ޠ��jg��=
yt;�R�aI6�tfJjJ<�6D��1>k?sX��#r�N���S(�k��@l���jT���T��d�!UZ�໶d���>��(�Z�:���/d�wZӒ8� ��Bݘ̧^H��M��S1|�����r;���
׉�u޵��|��Fsa϶t�-���:t�8,0{o��K-�8��§&�Q߅�H�t� �����?���ɵ:�4uVm���
�*�e`���A����;����@��d�GΕ��U�����g���]#=�cyz�`���]D��;5٭T����9�oE��q�R�C�d�����yԿ8�]�>�J��C�ϕ��X�|5��C'Dw���l�O>(>�a�� ��L/�Zf{?6�b�1 �g���X�S{�]_V�G�����Ľ������$<��H� �
*^ ��aQ�o�sI{�̠\j�&�`f��K��O4�!^�z���]��l~0[�QR"����<�_r���_�B��v����,	��ix���� �6n�xjA�1M��!��l-�FyZ�j���[PA����⊎έzU2S�%Ú�&{*��c		���g}e.���{��u�2c���3��d��z�Hv��n��%(��UO�1���Kާ5��0�H>���X������:)��oj�רzd���V	2���<<�.Q��"�f��7R)@�`�����ԟP�-R'g�.1*�cIq�n3>�[<�ύㆌAQ�ME����EN�m)D�G����t��>�p��-��<�+��A�$�xܰ�ի@C?y�c3���Vo��\	e>�{[?S�r�K��1���
�D�K>����+���"h?������\����;��$��8���(`��=��+
+9�7p��\������O�,?��9ܧ0x$Sw��+�r�����q����hf�,A�D�W�0�>F܊��h���،]�߯���v��Ë�;�V3��<���
UH���'��Wl��/�b���j��v��4#'<ߡ���8�T��GΤ5Y����&��d{�X{��o�
�6V��'�RL�������4���|��<ݔ�R�T�g��_�����T�����(	���g�j�)�Õɑ�g{��K�^��(�q�\t�M@�15�Ij�� '��\�j��1_z��j08�>�u/+1>a#��5q(u�$�'��ٻxT�4����B�x}E�Ql�c�E��/�-���Ho��}&(]0�F��ǽ��;2:e㚰�\�����7�2���d�C�}�$j[r!�1RcFQt�j�T�!:���p$_�Xt1�)�a�����$�~^����VX�k��&h	��($)Xk�&�]C�[�O��bt1J��>8�W��>]U���k��������Q3�~��ۊ��M�K[�QF?B�Yl�=F~,]>�0��Lx����c����EkIX��F�8}���Q�|�������9jo��1��V Wjɺ(}�f��o f�<���
��Rh>��c���~-'�kbT�y6X�����}�3�����yH^J�^~]e�/o���D�1���gvo���KJ��G��D\H�-�	�O� Z2�g)��40�D˺�#L�V����l��i��x�Ƭ�_�o�o��ϣL����I4�DH����$3-�zU[˾�v6��R,99�s�+��^A����ɝո�?;j2�����ܫq��ޤvl+eA��U�$�\w.%d����T/:��8��@6�>=����Vx��iH����#p|���ģ=g����n+�:a,ƜIOSo���wcs9�+V�O�E��%���v圼�"��3yfq!���0�����8�K�z�N%�!��u
m����X���[���=�M]�鉶��`�enx���ur�i��"���<w�"|&�)�	�G� y��)��R���UB?�t��أ�3V́�"�祫�tt�*ĕ��!�6�{ۙمY�f�2&Vm0u|���@7控M��H�<D������I�%�u~Ǚ(*5�I@����ejt�^� � �w�(�Y~��v��vf���o�/�AC�/�^񩒥���s��-��`"*�B�� �����Bܐ2u�a�*A���Y������4,Q�<�>Eg�$s-ꆝ�#,����
�!��q��hμ�?ĽD���u����
���@��h�B#��Y��0</<��$��LJk}�wu���맏���� k�`�%��j���Մ��v��׿}A4���UW_�x(�ۑ�7Am&%�z0ny"c��Kt�3����CGv��۹�`D%�2롉�tHK�J�x!��"���yc�O+��&W�r(�\"��yK7��ӡ�w�xdoCc��	;�=�bGTf
�w��5��)�3�x����o�[G"9�f�:.���=sd�ހP���}����b	��d���z���t�1���p~�<� `��p��%�\㿉����#��~SN�{Sq ���Sd�$���6#G
�/ q3{�}p.���\��aE�%Y v���$��dOI��]����5J3�"��T[�n:��}��d��p���2�rA ��˩n���7������s�t��Ά,�os�|,�ʵ`9�.W�*�B�b���(�Uȉ�l�4xV2X zZcCջa�D���U�륣/Y4�JB濫6��p�߀�!������ ��Y�=�(�τ�u2*���������5

��w�������ۣ�sRқm�7ab-Y��`�\���gq-D��zYl�|�{
�s+���u��P��~g�	��J�,�O�H���}�BRw��Xgc�d*Z�R��hmޯ�����N��[2��q�f�s�@AY])r0����1�V�m��=@��E�����"׍V�2�y�~�m�!_���@�wC�r�\��s�[DBoFU9pU��T��Nw�4A�N=KZ#�s ,3��6h�6�~D��ދ.�K��r��>C��R�����5b�V���z�b�U�~s;
�]6&nr�'?�!V@���/�^ǹd�Gr}I�1JZ){=�����P��^}42`h���P�r���VÛ��2�>�}���KGº����_�R���^�VKms���_(�p��\�ؕ�H*@�Në��P�������O�~��[��&�(�Zn^�?��X�t�f���<ՓB����R�i�j�~�����^��wg_�+�C�o�m��`1�^Q9L����0�%�M9�v[��:�T�v���@���K�C�����S��@�}�X�ǍM{�Y�v��~��,�������=XC���R�n���az)�d���:0Zx�ٜ�q��$��\�-*���H9�ң�4U�j���5�!D�}s�gl=�NY�l����ޮ�jSʘ�:����!F�P^���U�~���瘔�uG83���I$�kQ�yK��Z����35b�5(�v��|�E�H�~"9Q�0�[w�y�8������QR(�"�4ً7��Uy΅]u�&_��`T��2};��{U*Dx�����pY���2�y%R��h�b����ܢ�n��V�ԣ�2�Qz<<_�x��.�x��-r��za�8(�KM���H���G�5��0ܩ�æ�F
���ɕ�lXd/���s�wacߣ�r�� 5�LM����w��{qfP�![�il�̥I��㽱��`�[��*�Ѩx]�<���_��X�T��ٴ@(��/l��3��@��Dn!�0|m1�/�����G�DPq�`p���kAޙV#=��ң_������qkSpo��-	�l�O�i�
G.��u�꬧��6x#�{G��L�%�Hc�Yr�]u������8{Nr��H�Ke5��'���pd�9 2Gnǝ�:v?�j��d�E[�V �����紞@��|���]�	��[��[�"���M"`)�������ܶ�J�>Ia�>Ր�&�fͮ����;����J�$�����,�L�%�Wk��kNN�so�~)h����(q:[�ɉ�Rv�0FL��L�E=���h��[)۔��0�t,�d�o�L�� ����T��̣�@
��]@�H�w2���&N�4B��{�� �!'S6?�^�0O����ʍ��[�)[�,X=��`��/� 0�W(6]�,Y�=�0'@ Y4"b��wgu� )�" <el̝Gީ�?!�S}����&H��<���퓟��`����Y2��IŝX�o�œ��Xо>Ş,�Qb�W=��P����s[�dy�[jǄ��F��}�DB�� k@���w�PO]��؅�lh`��W��[�J�zN���}F�j������-�Gy��h�ՑH����:�p�߀8
R&���c=x�%�E���#2��߆ "^�����X�4�4b�G���`8b��Y>�a���G��x�&Ұ;�Ulz�M�tÅ^�����bھ�˟�/������Z0|�mR�0*7L�5��im]��h�WL�����:7�fO9x���Ld�k�O���T�V�f�i6�8�ڕ��3�a�f�)]��[���t	{&BW����"�-��-2�7f!ݷ��+LF<�E��{ 55��&��D��P��s���������f�	����H�	}V�g�S�\�y&N�J�M�}��z_ȣ��{=غ���g��$�O�k�?�z���k�9*ar�H4�#�Hzp{W�|q%�+�nX�&���]v6��X�H��C��[�w���gT��t��
��$� ��%��ނ���|��&CC��y��l�!�w���X5�(F�M��� w����jod:� 52U�b�Zp��d,"�\s薥�uu��̕��!@�/��4�uN���0��;�T����:�ӖSd�v�H��n��ιH��Y,�+(�]k���H�1�π��%�`�1]?{ne�XKN�,L�hk:b1�<Z�8K��"x�=�<p����,OYn"x8�OP�!sʪHxz��l+��|�+ۇ�	��"�&����C�]�_�}�S��EX!T������jA��	Ͷ-T#�Ǿܓ*�X	s-��}H��o��#�G0�lu@P`����H"�}?���1nE[�@\*	���h�:�I�J�� A��h��(G�AZ��R>Qҷ��+���q�-��c>v�@��r�(��&I7���:s��Y$�x)�)Q����e�Wy�~����������	��C��07#��8��+������_���?[a60��ʱļrs3ow�[�Dŧ�V)��â*�{���lm�j�wz~�g��TPǘ��q�M^�L������ hh��J�;���ȁ�%
I� V2o��uE|�S�ބ	%r%���/̮h/�u���B]Ar ϧ�mX{R���+�k�����n��_-T6�̋*��(�!�3gql崃=E*S�y�����E�
?��
���!���f|h٢��^�jhl�É���=��� ����
0���a�^��\�&kpґ__�,,q�×U�/��%e�c%Y�V�?}����L	Ym9%3T��  ��x�^��M%ߦP�jH�|����'�J�����$ߤ����!@Ӥ[����gͥ�oڑ��Lg��J�OD��Xd����_/ܺ���0'�,��J��}�7�̅�O�����]g�d���f%+v��b��\�]�^��}܀"N��Q�����`pA���B�E�e��~���|)�]q���a�v�HJ�`��(��?H}!��/�]'��a�$�X�S%��}���ò'�.��P;?��3�z�����^d�e�"�S �'�O�o��s�m+!S�J���/Y2��M���<u"�f1*��MSYM���� 	}����p/b��
άC���<����^����c�`<��H���r̋w�Ē�q�Ec��Y�vv
=G$����<�dH�n��{�ߍ��β�M�T|�z*Xc�a4k�h��#�y�`A�nt"��O֖�}�a�~;��J���<�1w���jz�ed������Hy5�-��awg��(4{O�c��UFۮg&�莙��&��c��Pa�L�I��������"�ܜ2������;�[���+�F�� j:�w��H��GʠZ�5�ڹ��j(���oޖ*h�ү�R6���h��Oέ� Z��ɢQ{�'q����?� Mf�;�]��m���U�N��-�J@4z��3+�r�>�vҖA�X����!1
,�T#*Yw"���=�^\`��[��]�����H����8�2׼Mr�c̫��tG�A�YkY��y�V��M#� ��$�?�sgjm��1���3�F)��kT��WCPD�ݏ�)�؞'glo��ҧ?���f=�*JY��[0<tx����I8X�E�a��,��E���׶@�:�&�íPߊ�ͭ<�K���G��N1F
��}�F����+Y(p�L��?�����_9���+���:�[+n�2��5D3�dSe�ʉ���!�@KD�q�I�:�����%���P�P��Ji��_2��S�wWW��м"]����rZ���r�b�r+k�pq��N~Tq�l&��H9�a���������o�4w�=��x����*sS_X����q<�E�<8X�B'Ԙ}����������$�� =�js�l�;���ڣ�^=Y�z�8׋q:����I�\�~��XH^�_��f;E��@q8#�g�5�P�e����O&U�����Y��dd+�H���#K�i�)o���f��Fe����{�
��i���	q^�}U[�]]W#�u�6��~[<�
7�]k�@����9ֺvh
h�ى c̙f���7j�_�,��S���y���K~C�昵cX�o���4�<��ԜtY�}n���*R1=b��X4k�?[��p5��H��P�t��ݲb��p��&z�.�h�پ���r��귛�|�J!1�	f`��g#��at<���pC��0���^v`7�{6sI��]u6c����S�b�32��h��D1P������%���ǙP��%(�@�}v9��}��R�*]B��&16��*����/p�R��`��Ӈ�`R0q����V�X���0�K��Ή�#6�=8���D��N�Ԥ.u	>�O��B���Gc�Ŭ�Y�𾳔�" 
���H�l��;�m�TR�/Ou�JXp����(�'��t���l��m��k_ ��^/[T���]�i�a�B��8�p�XK�������m�j��T���`�7��4�$Q�i�l<����S���~R��z�H�&N��*?l1rx��w��b���P"U�T���r�鑵%��Sp�>�.e���q��ꭳ��_3�i/j��P{����m�k�W�����8�9���7z�~����D��qi��Q��������y�4Z�$Ӈ�Է	�ҖI�l�1L�آ�V���m���X,�Z}F����>m&r-���8'���$��k�o@�x�!�48z䩡�L�����
��9��.���L�����x���Ӥz��ۍG�t
����;S�!�_c�8���1�9E.�	�\S�	52�Z����Sa�q�]���m�2�̽+U���W��ɹ�͖"�&���z';�=ʓ�wv^Ƶ��5�@%���Qt�8Ko�<��õʳ3����$���l�k��N��QӘ+y��y,آn�s�i���qF��[�[�^C)�&�r���M�Q�,���B��7�w�i9���g%�m�I����50�+"�U鵂&���J�y�$�XkC�r��<�("aV�v�1��rX��b"W����0������	�/�����j�$�v��$D?��=eM��iF���#����	IvN�Ȣ:�5�;����+{���(�2//�P��5�[���]�z�L��N��m$8���)��6��JC�Н�^B�Ue�$z�5jC�S�����[�+
�(�Z80b��,�v)f(���)�, $,�����e� ܧ p��8L�ns@w����k��S��7U���28hh�Q��Ć�e�/��݈+��UA���X�^�.� ��~>��]I��LM}rv�ǡ٘)ӵ�E*���9�p#�Kd����Z�D���u��+��_=�SM	���=�zz}�Nf�W��"8k��,��!o	�����z�o �?L	�&Έ�B^g���E���D�(�w"�E)^�Xk�R��m�.��T����R���~����o; '�;�}x�
��?���:��JV\U��u~H=	�tI����$��D�]�rQ����[l�����C�%���c�o�m���T����l����ӆtMH�ߚxE�9!R/@%���:�$��hb?c��v�~|�u8�I�O^���t�-i���E��W�'4�'���U06�~v�ǳ��(mI������~����4%b��B%�}w�N</+��~�Ȟ�w%fo#�����n�Y �iM��a2���?6�F�Eԙ�c
��D4B�Ӻ�L�	�#t}���d	��X�C�9o�ފ�IOp�a�a_3o3ǒ� ���H�%���D�@��&N���?�(�M5CR[�x���%¿#GR嬁&��QU¹j6d���ͨL�ϟ'5 S�F���g���蛐��ֳ����ͯ�v#�z�w���� F����g>+��g���Cb���A!�T(�y��(i�HYV�k<�F�S��gC�͐�J�ϙș;�!��֍�i:.�)¶�1d�#��e�Z� ��L�f��,���	\^ik�([W|Zw{��OR�A�n����� 8�g�1Ē�;�fT�58$̝`�օ�@\L334�,��ZQ�V�7XD�V^�5����d� �&�g�Q��-�᫖�n�9��#Q�c�zm3lr'W�R,� DI��6�/��zU�x�&Ղ�P�L�9����zm���WCv&�u���
P����꒶��I .p�[+J ��(�i�f'�ᬶ�����lo���wH�)���)"ʦb��
�����Ŷ���|�zV�\�����ڱ��(��eƽ��
�l ֊ˌlC9�|i��֨B�iv�zI|,i��
��#"Jkօw�P��q}߉��>p�o�5�h�%P��DW ���W*��E�9����}ٝ�s����	b���.����S��PX��S4���2�����sU���X**�<�\Y��e�_��u&8�����O��#Qix����R�;���2�\v	g�֮<'m���TO�%�aòUg/2b���B��X]���#�1{ۮ���M�?q�/&�B�{����i��O�G!�G���=���A�!ٗ��~��(�oc-����xu��h칵��Js�އ��:of�i�G0��a�*�@)�˘n��!Y۠�!z���;���)�*�9DI���Q�W<�\�.�2-R�T��8���ԶM.�L�]�����lS��.����p���,D�em�s�Zq�����}+��P D'�E�M�ԝ�c�=��N�����3�A��T��V#��,�I@}M������ԒE�^��\�E;�B%�on_��rt�ǻq�NN��!5��\m��|�[�v�f�F�Fɇ6�;y�#�=���J+����� }W�"�� Y�-��U�����z埏σ�vg{���u�`=��ID�?��\J�+�]�a��6�2x�RG�z-mbMU}7 �z_7@=�8�
HaD.4��.�i�1IHt� ��2)OBW��Y5�������� ��&_2z�p`Q5����Z�+�Br�HȄc��=�3��쨝�*�Ǵ5�Ϊ�~�r�Ւ��c�Ѧnh��hn!u18sm5�B-�����t��L�+Ҫ��dD��M����	�OQ���N��ɒ6��3c���Cz� іǷ�7U��	1b �KN�\�B�� �����*�_v=#a"���N�5����<��Q�G�-��ݓ{���S�L�}�^vԤʽ-��RU���1"{�����=�]w��?Gֻ�����5��fDT%iG��37L�f fUJ�F�g��C��>6R�bh��4�@�j�T��2�c��L:���!vXb�B��q7%x~bס'�R� �~h����Ό�eϏ3f@Wמsr���7��-�\.�Ȋ�^�?��漣Y8{j�y�l�Tg
^��u���%��{'�&���e����B4+`�#��~K��������̱b���G�Y�	GQ�LA:��5$8����~��>�4M̤.s����!��[����O�Fpu-1Hj� uV�ZEk�:h_)ì��.0���۬k��7��?��^<�IDL��g";F�CI�H��T�j�q�".??�S1u���i��Xu��<IH���K���)��:��!�(5������5Sļ��[S�����}I`�IS?l�t��\���a`�8/k�mхA�/�W�:�t�Tς��]f�$bߓ塪��O<_�z-�=��Ti�V�`����X����_Aׁ�M��Qb��f2�b\s���yI�*�7��t��@sy1��s�^A<�\����;J��	9��09l�p�� �[-��o�
����X�v��ݥ<�j}^�aғ�)R�5)@1�קۃ��UR"��vQ(��7+����EY�T���|֘K̦v��4s�,��v�󋮭{��������{�C�u�M�ɭU3�ٯ���mъu$.7�����6��.����q� F�;�Gz�Z��0'�h��72���8ڃ�w��uٙ`9����o��^p�4Uj��k�.�xs*�"
a���Q���g.��y�>|��t�)�帔�C��J�DZǩ��;��K�!�m�#VmX���GA|�ENk�9���]�HÇ&ڦ��0���"D���pJ����*i�Q0����f�S=�p.RIM<an��w��dŵs����7��Ҏݘ�c�d��y(cd��5�Jս��KǯWP�a�|RyBlD�1�I�D�xvl�I����D�V�=��`���� vyª����o�<^'��ñ�Z��coZ�Ɠ�C�3�s����>׏{�Xo�N4TZo%I&��X���Oޢ�������)m�*�|�z��ުS�$i�1�H�(���~�>z�Wq�\vU+���lRs��K����ٸa�"鄸Y�a�۰�H�{z�[��Xb�
�S�>/;d��s޴Kv;z|��ڔU�����eŐR���='00�}�Yk�j>v�I����;�5ܴB-���O��YV ��(N���6��*3i5��RZ��v��捱=����+<�Ι��z���SD�R����*�-�Fj�	1��L�oA���ye��	�g��XM�\�8��}	J�Ì����ڦ�5y������K͋^���4#ed)K��}�x��uic/s����sb��x@�0\�[~�N�؃i����ŔvŏUC[,�m5�e�����Ģ��\=�o7�~J�Zᦼ>�m _W����e'G�V���z�>G�6���rg�T 3�\�!(�JH|�_HR�?E~����!a-5�U����T8�%=3\��2�M�J�	�6ȝ���֙c��s�힘s���m����>�9i������"�*I�b��]�i'b&���Z�!q�T2R�Z��%��V}�D�*բ�?Lg�g�?���{
_��������R3�1�u��{�@�h���ݶ��0ZFc낉,�<}�6�ƸRHm���e�ߨ����d�/��-W��j��ѝ=k7��dd���E��;����p�W����П[L��*`ʙ��Ҹ��^�^3��9�R����O���"�c��c��8D��w`�ε�'��ZK��>,^�����6Fu�Ӷ����2'l�����X���S�M�l��]q9���"������%/7�j�\+BA��P�k�@�
��0ti�&i�!�?RD�𮹿2��7�'۶#e$�:`���?�z�YzLD~��!M�_"~�&[G���b���GZK��7q*�nª�zY�oh���.���+6��p2��x���ó�����g-x�����b���{��A�4�Ƴ@���9�ⴋ^��S��(b�$�����$���
��s����1� �r�ۯ����zީ�'GEU��s髤�C���ٚ����O��_�Gh�3z�-��>��_a�+oF*!'l�sh�h��Ԧ� (�!��j�c@lL3P���#@��X�p�
�g�&&���yP�yg0N<3Sq���0\��(���x���M��A_�Y���mw9�?<3%���Q����G]i�l�ll�ݜWR�������Ӳ��lF{7��	��t�d+K��Ø�Qi�\�>�f�TgL"��\���?��ؗMlcR]��l�5 ����wה�1g��9���]����Y�0�C�H���2-ZI�N�d��)ьf=c~@G1���6"ZG�ܒP	=�ȢϢ���J���~-�cL�Ы
QRh��&3,��#��n���yU8ŋ����g,��)?x��lX��А���ٖ���Ё��~��	�������a�:y��H�Ydѷ�������(��2�w��g��Hnn3iH����b��gW��fN�q.g�U�/��"���M�Vi�Rn���ŒИߑtZ'�ݻ:����s��5w�,��&��_`�{������?�a����jYݼ�6cOo�_��+u둈�]��>q�e�U����N�-a�M߫�4���#_��t���_�T^%�<?p7� �btۛ�����aO�y�#�+�فƞ��H�2뿽�G�����>�&�A�%����Y�l:��C���磏��8A���nj���t��T�?�P��s��������se�Q��u���HqK���V%��;_����F؏�q�;��T��D��bk���7��})�JX:.q(ά�k�M�aK�� �)�°[�+� �͈`�C̿���;,�O���q����P�ī�IQ��C4��p��C��?H�L���@2��^D�"~�	3)#��~��)��w��_��8��s,ddS���N�EaU�p��[2$�"VF(��Sa�K�2����}��Vwv`������<���g*$�GO�bp��Ho�k��w�&\�O)e��;��Nj^MN�K�f�9��/�Oj��j�a�j��$�:PA�b��@k@7���[pSs���J�I���w�.�^$9����k�@m����ZG�M�*�y���\Q� ����z�J��\M:��.�4� ��b�ڜ�*ˁ�J0�Գ����СòėG�^�'W�xv0\�[_ޖ!�Úg[�})�C�vV�PQ�i���#-:�	NT�|�pvP[X.�%�o}�����_��l�@(�����3����C�*�a�N���IY7�d�"���Q1�����]n9�p�Tl�2Ur�츶����}��?���E�xM��sZvc��y7a<[}���7�4�/���c���>����YKYI��T'���i�$�!���p��8o����N��m���N8	��a}`�E��t�i��5�G6�p7���"�����A�P�fq��Y���E�����S�7��s��l4nH��ȰiW��\WQS�%��E���P>;�:���`.���(/q�m�����@H{]�Μ�Oe��eE�E&>zkg�D�4т��Ap[o��d�Vb�,�џ���	HѸo�aq+���$����aq�ؠ�`��w�/�(��J��.�o�v��������X:L��yT\�}��NF%p��;`,#�+����8��A�T�u�JY5�%낀�����O��tn$���hcfL��=ùʓ=�T��#\�y�/�ִQ�>A���e{-���sa��zo&	�@~�6�+����:JU��=lu�=���ᮄf}񘢔y(��l.ʥ�U���F?�2�+���lt� R���F�Z�|�sv���<O�%1DS'O�-z�=�77�A/��,g�YW	��Q=dPKUN�'���ݔ߷(��{�@!]tcԢ�Xvi��a���Rc�jk�����ؠ��qqc�قY	'�2i�~h)P�#�X�.g{���tF�k%�mcFC�k���-��V�nM�������rwN7~���h3\"H\�=ڟ�O�Ϟ>�
�vb%4p�ͷ1�H�^I�ޘPnک����e�f�jΤ��Y��X���)�'xg4 A��	�#S�{��K��.7qg� ����tn2�;u���N�:X͂�ů�,�!E�۞�G1��.���E��9�HH�Pm�w�U�,���֞�O�ĭ��+�ƹ)�#x{��CKN-�iT��Z7�&ܝd���|K����<D�Y�i�A����9T�#UT��
cx���4��s���\���F�B������TW�Rj�t��l� �t��LH_�ha�q:P��\�pQo���6�C�&�/���v�(�;���fw��_�M�:�A�!�P�u�>�뷸�/�d/u�t\�?�y@^8[:���FQV����� by���$���uB(�������	�Thy@�� 7幭/:�(��P�53J7���1{�@�NK���3TwGl�u�r�S�=�Z_����4po����g+bsz��#����Ī2�:_�n�
��<��D��]���ua<Q�w��*�Aƶ�v0�����j�f3Fe�ʑ^��� 	'��oT��rLC���P�Gܤ��T�9���՘"����Ҕ��j�G���+��X]�3>%*�@�0�481Q�s�|��,O�p����df"w��,�C%ǝ��<i����~,a2���L���`���ұ!+���H%y�v<�f�,|H�첗D�ۈ�ƀ��@�5q(���;s��"dd��]��V��F�wn$�1��e���Y��p��;���hIX��`f��;M>KL쌿�A}A*z|ٲr�� 5����H@M�OR=�D�l� g����9���#k��	�=uŠ6�����fE_�y�xC���v�u��c��{9i����K���x��\��
��*�p�̣��Ӓ2u-�;K���E���0������j�)ת�-+5�ES4�����H�䂚	(�6*s�߈�5@L�-���S'z�gr��R��`X��7�	FL�((p�i�� z����FK�	��1פ`פ^m�a�<GDX)8�N�!��t"U6, �,�I�7�����1�[-�X���Ὺ��|����[I���ܖ��͌���V�J���q��;�Աo�'B���L�sB�����eGyBX$MP��\`�#-oO�*���Z���_W���ޖ�������xs&���9�jņ�#`�?a��9���t�o��l����󢦖|���l)p"'j�킒�:$����ࡴ�/��W���t�yt�+J�5'#1���a����d��zg_��VZ�l>{22��*�~z}��^����-v&�����d��R�=��C`x����p�1e�N��ǃ�A���������BWŦ�9��gW���F�j����s3��:��H]m���B:p��ֱ�����*4E��o��2tp�����3�T.4�\��;�����X��	���H^e�Z	(�%�#��:i���	��xNVFw��;�I/Y��a4�?��-
D휿qO ��e��m�a8�V�čR<��~9-F	+E=���G�t��RF8W2eY$���8�e6OO�+l��A2��2E��%��W�Ϊ�4�l>�Qf�/��Cf���.C~H�ń�"���+@cj �G��ĭ�~u�"�1���0�ܘlqL�dJ�~�dզK���$��d )�B&0�]a�Ԥ�]���{!�2�w=��tfy�ߝz�0��&�l��7���@-�H��
�3c���\�Xc,З���D�g��2�A]x=�>����&��P�;�1��ê���Z��y�5m�r'��?�:�p�XH��-�����5�p�f�[�5�O�&_�3���K&�v���p�P�ՉS�Y�!�+υ��00��/����)����.����YoX3�U�MT��e�����s~JD�6���E�?�w�DRJ,�$_�u�HB7�WxG<gf�3�<\}�}�~�
�P�(�Jj���Uk�j�X5�� �^,)��W΋�P򑣞m]���E��=m5�(c�!KO_F�%�qC���t��t��/���jl��=�6�dǡ��2��#��$�,����
Z^��vM��턓4�/��i��W���Q�X��UcrW�&=@�'ػ����M2��z��(f�]�x7�`��G cX)��I{J��~��蛏S���Nͥ@��<��M�Ƣ-�x�5��&�.P�Dt����1Df���?b%)�Ks������Q}��VI <�JH�Kگ��<�Ta^�ʳ"�h���{��*�ᝀ� �OpX0��Q{��
K}�g��	%2�AӉw�7�׀�s9��0�M��$�L"M��"�<(Znk�~'}#g�vQQз�e����e�S4f�5�y��Tqz1*�u��Y�yj�]�L���5�gZB5P\iI�&=�������;��|!�w�(�y�\
1QH�u�zW�	
j����8���>/�h-y�lH4�_��_�:���nc�0^�º�[L&���T��}N饆u�~\��O��J��f2m�Bӽ=#��@�L�{IN^穩�4�՘�����{I��)@,�}�q�M�֍�b18���'-�ڼS?�s�m�I�#?�`��(���4N���}��mtI؀L��.���.����AߢB�9F��J�2Dz�H��=���C֋�~�y����C2�Apnp(-����x��o�uޔ�P���F~�P�z�����ʘ~�p�)��������,uH��r�I�K�>��^�ol]l-ck�F{C�?��䝐8��Ϋ���'������>�I���ۦ���\�56��;��I]C3t�i� �f+e����Ťs�0$��ͯ#u��嶨鲄PJ��¦l�j`V�el�3��@��C�����`�Qn�k3������>����8I���A�K��'� �0�`]���7Q�=�|ܢ?2�T��8���E��� 4���z;��<�*Ӥ1{���˚ �D0��[U��j�� 	���t���#�[�K���g�*Bt菤0�n���w�J�����c�X��B�B��G���B��:Pi��ݽ��?���^�d���T�ymD�l�A�y��2B6]��1��%��T�G�����גޤ���r�%��^`@
��k��ܳX1x�ڼn�D�Ӌ�M��/+ È�怗<��M�f9������M�$G��oU2Qr�OF	����	y�����|���QB�,�оd�F������5}�μW��5�PG��mޥ�te-��jg�p�����9���y��>�r`�#��{wͣݞ�`y�T �Ԑqua.v9&�y�-)�E��$��Ft�J����j��^Z�)-�[�#�
惴M��N�I��k��,1�nV�*߂�)�_���B�|�\�)�B��G_T(k�%]�;�~9-��[�?��+�b}Y�W5�&�^)�r�N��#�\">�L��|/���WE�����!HnwO��;*�@> �b;��8�ᾕ޾�巰cll�Vi��~����܅Gv:��Z�i�C�D�<m3R��?34-?˦AU��<'�z��6!V�o��q
��J�E��)�&g�>N�[�"��'2T��̅���^5X��[�a3b5�m��槔��4��4��R\�A�4��_����u����Y�tܗ��Q��AU�艭�n(���E͂_5�uq�Bm>��3�5�Z�sv���"T��]�1��r��:�B������nN6�=�4� glo�����#��P r:��i>����XX��f~�R���Z��(5�Dw<�f)!��a�������c�W(1jos�I�>jאq���No��4 ��e���?3�/a�E����g��ĥ�����g��\l����Dv��Fۤ0���56�{'�H�;.5�=(��N��۱���@���LQ�e�0b���e6��7d�Z)�Z �2��|�A�M��B4������1!���SG��V�A�gـ<�TRR1�����r��VAE��T�����!��l{�5��󍿩*�����K�D���?�W�y@�S_+�%j��X��3�����/k�~ABk��+~�o�`6���L0}TY�S~��l��z�5ϦoSpm����&q/�P�%�9�LU��n�����{k�������p^�;3a0��<@e�u�k�ߋ/����$�'���5������d���O�#�Ӣ+e�V0��x[�D9�7-ݚ�$�7��$\$����R�)���J�%���usG�bT�����h7��/oǄ{��Tc�	�8��J�\����q��z�%�mKð� ��-6|�q�hF��p�X�9�	t�m~�0��y�PO!�:az `U}BU�]�Y�N,��'�Wx�Y���@�2�U����u}<AC����.�y&t]J��L�Qo�� �37ãy���(㮭@?�8.n��E�KzK�|�Y)ȳ;�=���N��]��h�b�%�[�8rHav� RҘZu�m�3��4Zf�Ϫ�Fn���yˏ��Łq��ˉ�W��?1��֤�<�7Z-����6e7 o�j�ԭ�c���z�*�����)+�׀WR�YzE���FR#k���+��(���ڹ*��K.����a�ةz���i���jZ��ѐ]J
�g�b@��"������G`'1>���S�]��s��5�4���$<��W�#�ؙ��n_�t>�F��M�_	 ���>�./��(�g�B��Շl`�e��!}�d2����YM�\-��,9�>Yi_��h��P���[~G���6W8��T�% ��+^��;Ǚ����	v���L�p��ڎ��[�,��mL߲~�\������PV]�NU`!�P���J���:�����=��2�=�^�}'a�t�l�2�DD�(���ո�1��k@��=`���PT�m�7	 p��(��� y�I�j2��M^v��-� �(��[�����=��{Jv#Gj�x�2P�_�����&�У���XJ��ѻ�\�Ԣ O�i��	�ME��
H ��i��Z�0r��틅ȉ��"�_I6*fjWY��Bw:@�k�ɚ7X� �0b�ǝ�<i�9T^n#�U�/#H؏΂��p�g>�Q�\�	.�7g�qv�e~�ۦ�z�����V|Zv�qU �|E����Hߠlψr���r��-lu�Y�4�56��C����E����D�k��4�~���v�.�A���޻R��G1[�۝���2ۆn}2K��۽��ّ�<}����<�>����R��cnWo5�fb%�V��j��`���[���/3�b��%α=agaU�j���?�;q(�*�Ӷp�5��
����I�Wq�~�ކ�2�E���� ���ԍ�x������#I�q���3�n$�:(,�)��1Yk�+���5�ښ��2~�>��Y[Ӟ��J�~�VI��y�����*�L�$��^_�}���-�Ҿ~��v���1��5,��jBL	�|vlH:@i�� Ć��Wj���:8�#���-����2B�f�
�,P�<�Eꩻ��x���� >~r=,�Q�m�f�h�\
B<¤Edk8��`iS�9͓>�d����}�_f'���43��@�/J0����~��Έj��F�Lbk ��;�H��V�%=�&zO�)ڿ�-$�H6Z._G������,���r�۹�zb��'�$_c�����n�����T��]���v���sp {��%=����a�l,CJf���z���iԌ�9s�h�Fz42������L?�&u3�D{p��������A�����M6͒<�9�3W��*�Uo�x�foo(qx��f�&b�H��9sL�D��W������W &�=��^����6P�d�dA	�~�[J���Y�bąG��Oj*�[��h��.p ��W39�T�o[��n�Z�=M7A�ޜ��éyTgGk_�)�J`��Cg��o��X��]z��$<Ð�r�3Su���>D>����+�)q��U���m�6̗��Q���d�_�,I;����ky�8�H����&L�K-[3����t�?�+3}KL�kX,��{�$�X�[���s����ڜGH��
��ퟘ���B��A��Za2H`Л���3U���)�����zmH�71��m�01bN]�w�-)�0��ŏ�5�B���:�1D���񴁕zxu��e"z�5��e�e�Hk9�/��TВ�]�4Z7<��i3�.Lv2�ϨS2�2�cx��Ld��)N��R#p�`�w������I��1�z~`��}_�7EfT�D���ã� ^�b�x��J�)�qD	�C\�\N��!S��0q����.���%Ek.�'�t���s���o�V+�?�-E�#%�V�l A�j�/�Ć~θM���#c���G�Zt��ޤ��E"C>���	������N��CϘ,��؛��_3�Y�:��g|�<}~8+�H�"&園��s������!�e�!��2b#�f�rލ�TI�A�kj�������U���_7��N�b�N��g՞9�����ڪ�����xL�n��x#���5��O�5��xB�L�����S��1�&��j���Y���Q�?�z����Z+a���@����ƴ0N�� ��d0�|u�Ϥ&��l�g�})	{(�A`�q��-9�� (N�Y�n^��[ǟx-�-��\�=� ��h���%8 <�A�9LF��7JL�)�=�%���t�w5�7�QF��IOO�k@����>1Z����I_*Ma���:r���ZrZ�e��T�H��Ϸ�����{j������&֨
��۷��O�Ƹȏ��Ǽ��D�~��X �Ab�WBp�'{�2��C�����S��o�_Ӣ�WO��R���kK3�,z|�N>�@�B���eO؀��	EGY����}V��H��U��>oz����VU�o�U//�g��P�AӇ�D�6�HSF���������J?�u}�C6�fb��`i�.T.���N(�,Z:¦����g4T��E׃�,����|c f����5
��O��cc���`����ɠ�g��>�%8��N?\yM8���ɞ�4��B:��R�1�
��R�ИM�Iך��@fctsh�2bddr%^�'�la}�PRF%0�n'^8��$ʩ����厔7l r�'���o����E1�=V�~�s�@j�l2}Ol�`�T��s�\�@9�ͮ^���M��^Y���Z!@��`7G���u�]�HBr���_����>&2Z:~XD�D�@X���0�-���K�D�wv1�|�$�X���K��''�R��I8[�b��K:�}R��/��ߝ�:�-S����ơ�*@�rF���O�C�UBs�u�'���=>�)���2N"��߳�����n��S􃟭��*��-�vB���û1�gy�Жl�&�?�2k�bXQ�W�4�A���S{��K�n��y�չ�%��r����4����#�j֪U�\Y�,,;� ���(���/!)^��Y����Kz�*i�R��<w�t,p*�7�⟘n�=d��N�7�3!���r�7�;.���:�����#f�쎣�SƲ3ٟ KA�K��a뙍�w���w�u��p�kkL�H�O����t�kg����K�8&X��*F��}�]���8w�������4��*��ݥ ��^čH����~��|�mA{*��{ qԝ��*U�y�r-�a˃9���_��V8���g��
��%��a�۷^	�t�	<�>��$>�I
	)6��X�Ė��Qa�k�|��r�-߄S؜B�u�]��_�<(L���b�^����]3@����4�����. ��$���� ����W�����Ɉ�]
3 ���)���`(��V�'i�Wd�Ir��y��R�}�ZD�J,&�.yمv�&�wKD����D8�U����'2k���>J�XJԑ$�mT��~��:3h��a�QZ�[�a�j����v�[�!�V���d�X��JvX�� �S�U�Z�,�N'>`�C�[�H�����m���QH|�T��k�39.���h�������UB�x�����B<��B��m\���y�.�7�&��v@�К1��#h�ܩI��Q%~�cGHtG/Rw6)ť���C�u�@	�nz�B�Y��H</A�� f��@���R_6��b	2`n���V�;�L���U,�x;�9��zP_d�In{�R�O�m�lt�=eb�����=�.�Ѯ4~�D���k���-"�"#�%���7�5A�a[�>��ߜ��Z�mi�R��6~��{�z9H��6_tL���rϯlw�A�n��O��Mq��3��ˮ�}]׷?m�5��[G������ãcMV�WAL�9�B(�E���b�Fy���:OG����PQq�)���b����!R4ޙdӹN!7��N�+�:�y���x2��*��;�Y��K;�������`?�z��s%t���Qn��a{';��L:���ٕ�Q�ͪGuv~M�u���cc:	d����Z�C3�H����@R`e.	���g�s�%\6�֨���mg��?�Q+�Aa,;=�����i���
~���v�����vETƅ޽�q~A��e�y����*ڊ��_e�f4r�O+��Y���ͤ��B���uS��ہk����b�c�ſꅻ�|(�H�ib��t c׫r��k��wP-Z�`�4ͤ'	��x��o��1�ط�5.D�hSM ]H�.�*��*�6d?(����<����l�1����I*Q���3��äc��(4$� �Š�QT���/-�1�����z37Ѧ���.и�Zp]@����&D8F��6��a�n> �?/����l��+>�� �&g���ȕT�s������HM��	zq����]\�Raݭ�7��� ѕm���o	!���V��{�B�_�s��s�ќY}�[��Uw]���3LJS>���I����G�����x�p�w�.�ub��#˭���5�JS�PцL���('�Ht���;���܏0\��`
���;���Ӧ�]e��t����@pdr{�*n>%'+w@���<P��c�'?�Y!_��?�/��i��V�Kv����ܐ5�[���)��Q�2F8h�佪����ZC�F�85v��9�:���Ċ���Lhך<���4F+��j]��>PG1�������aQ�8p�,��WA ��ȉnV)�c�`N����W�jد�h�@U�J����������b��Z<�*Q����F]��Q�m#�O|6�η����/�K�~�^�:��Hq �����3�e���7=Fy�^�#-�V�>�h4Ec|�8I�z�]���8�Ҥ�v^�(�h&0�����NlVl�T� ��ߩ��;K��QP[�����K�eV��D��	z���
1O-T�7�6�1�J�ǫ���Ý�A�.�B�ݝN"3H�ݦDH�[$�+�Qe���� {����]� ��=H�Ŀ���/���ٺA��=�u��\K��0������h0��ǎ|'`F<���X�I#7������rA4Ζ��6�؝mLC;K���A�|��Wq��~�1pzZ{5��FD�t:�)�c�1�+��2 yڡ)��E����φ�l:������8�{O�KA�L�#�9�z�l�������)��U��`sH�Mx�Y4$����SP	`o �fW@E�`GHiD �Fbhi���F#�9w�\�>�,*�)�a�����<:��A	Gxנ�����m��ؑq���j��W�?�MU?ld�Ee$��Pk�T�b�����|CB嶗�uCu:�S71���T��e���C�9������{2�9Y�JL$��	�7�_D�J��4|�A�1=_�"q���Q�vP�8U��/M9-VC6�.��h^��?~��l������~vX#�F{�c�z���gE�X,�Y���ݡ�Ҿ-�*�.T]%0A��\�t[��kG/am�_,ryle6K��B�����Z�=D�!9�F�ԄM<��k��~����x��f�i��$��Mh��^��n7Q�]q<;�s���0����6��t��'�R�H�v'��9ur-�j7�3��p֜�#.UJM���>�Ο������*��mN���C����-�5d�¯�JʯO�d<�U�ƫ�`��˳Dv$��+��-|k�b$w9�ͨ�����R���Y������q���N��lߊ����L�)�/��	k@{���җ3�zq�t۽��"q��X�a��'��X\�C�!πN��H���x
���7ϴ����[�w E�rux;�y�%Ńg��1u��xS�v�>Ka�>�.�v�2XR/Nt�5�`pyh���}lɈk����w����<����+t��>ؚ�M�AC��яf��~^�*`���&��J�%|�gc2������6WK!@!�7�s9�A?o����kԒ	�}��E�gd�_Lͤ���h����s��J��2��&���h����SJr�#�-J��7�&5S���T�~�*��W�pi?��d��LD���L��h3ZM��*�s��O*�$q4�f�uΗ��DU���S��+�.;�Y6�8�|ͤ��6|�n����n�$�>� �N0]��c�R�=�7�p��V�t���_�K��@�	���� ��-���uA��D(E���Z�k����eU�m�E�̦�+���s���_^r=��$���a셫R߱�+U�ɕ���+��l�CQ�?�o�a�.\������m��
�K
fIz�b�p̪Y�ewy͠�� Ee�G���*Sg>lG���Q23��d��a�Lϣ�B����v�"�1x�tat0����>ڥ�ݵ��7��r��l�,MZ�|�Xr͠khL)�[��|�!�c]��1hnb�� Ѝ�X/nnl3^=������;�9�'����ȫ�<Ta�Q��=R���%�1��a��@;�ШE8��
+�/{z<�[�S�b�2⃋I��2���m�J?�<�rv�{]'h<��,���Һ��7Y�P���śp���ū����}j�#�au��aso23l�ـ����K��TH���,�����9�tj�/�Q'k��y�i��w�6Y�&����3������U�)�2Omܧ�f%�{�/�����ݫO��cZ�*ɓ6	]�L�ŉ@
u���>���N������#�x,���`J��i3U\ܬ�$if�f�*�Pg�	0R@at�#���oh7�'w��!�8�M8�A/���]�F�rpKjj��V7C�qQ��߈���60��!�� `8��W=�J3W���2)��I�d�O�/��CF�E�i�D����`�r?�"������!���ɻ�HuѠ?7�Wc���c��a�����}�v�7�A��X��ޅ�Xx���`^:]g���x��k�U��M�/9d�ͯh��P��9�����Y6/�����z�")��	g����`kx�se���-���Q\UT�X�J�s�y|�C'��Nk�+B�����f�$��B���v�~�?[ip�n,��(��-O7�f��/2MQ�=�� q���}�8�T��a`�F�(�<:�SlY|�;RH3..J\7A0f`3��������js������~�#$1G!�S e@q
��{������=��j�$��L�mVW=���|(?��[r���u%w%���N�/hd�&�$�'QTK��/o}���өA9�K�>���pSAv>Ā�	*�/j�0O�LH�+�W>^0�L@����#�>�������8B�2')�C�x���\lǒI�A��JC�.`W���+�;�~[[�����9K���>�ef���k�+�i�Ծ�^�^z�Q	��6[�q�	�Hι��ҟ���}3�ں3�Z`��t��eu)���[ش��gB�S�^����''�R�!
�	����x(Nc�u�N�j�U�ToA\�c�/�����"ٴXW
����w�� #fuB$)�[�yMKj��կ�A�cс�[sa1����;w��x�3�X��LN��೽��3eEZ��d;Ƃ��4�~[R31-J�Y���;9G�E"�����X�/p�o�.~l�O��G���s�1��V���[SɣU�=o�q�'�B���7P'�g&�j�rz�y�F-��-B�3�,ŖXc�"��v�7xm0���YX�M��A��t�3��}�eE�ā���D}��艵�{ ��'%��2��R�hY�"���E�J&6�*{Z"5IYm�̩�X�p�Z���!l5��5�4���"�3ĩm
O���{�3J�,��SD���buYAe`*��MKH.��o�!�)_����j&���g���s_(��:�6C#��Bw���T�fe�7[��r�8�]���Cގ_G��ht!;��x�G�%�d���E+^*�)<��(�F)�ǘ���즃�HL']_Q-������� .)�黤�:3�0�\
�@n�l�eS���Y2��W��X�O�o!�������s�7�wT�b.��`��
�r�|؄D��~<-�T�LZ���o[+,����&�5�G�Y@U�ztw��aP8EB����dF���8x�&S������q��!%�͇�2刿�)R#9�X�JOƀ»�����B��f�y���B�FH7��[�1�|@␕6��������>�6���i���#$�?�$d���g���c�߷�>6In?�����D䞽�Í�J�.����|�«�K�\Z� ks�T�Y&=j�u�I������?�#��u�@8n�4{���Ôt���v~K���ѕx�q1���U�5����ca�S�ם�)Cj����΢)IS ,��Ԯ\�6��>tH�=���_D7����vI�0<�R�2
xCu1¶�5w�]̎�J)���� t>�;���zC�-�͔�+�wBX��8��	��?F�dM��������X�H��Wd/�T���A������r5�s;�g��2��*^NxB��Z?"�� ��)��+�b�0�wa�%��f~zI3��	>�?��gl���
$�zsOk�vXh:{41���A�Qx�M���9t!q��_���z��������67�<D4W�a5�Pa�R!�8��x|�t�N�)A
�f���If�$+0J�� D��>��v���D�T��Q��w%MY����n�͋k�@��fLf�@��y/x+���h"�%m�
��J	0;�w5�j{�&Bh\��+	׺]�,r�d[@��	����~��z��*�uD
ˤS��跳��.P��	m�6�?D�lj�p;�DL�[w���ٺ�qޑQ�iW�AZ�pB�
��&�A�X�RG�����"I��?k�O+��}�4AVH���:"e���1��$�F��/}$Ap����[g�4��|�3�!�����7H�XdD�8��O�r k?D���u�}-�Z����n��"��̻'��j@�\Uz�ԙ_d�n��i��' Y��?�C2��.�֊B,�z����b��S�^i@����UI+"ҟ��j�%�$���e�Ś���j�05�4!��oo�W���+t���4;I<Lc^oa����{h?����p
Q2I���
L]��v���hv�[3w�Z|�K'���������em+l��	0����g����,���q���l�嫡?�Jboi�%g��M�a�=��{g���D�t���o;���u�m+��4��(KL����a��-d��}�Ϭ���"�;6�0Y��56��x-���(�0b��D�(♭���s��f�˂�
�t���������O��\�[�r� ��P��[}��L9e�tk����݅}C�E\}xŏW�;�?�9�K�¥�GL��>V�Q���H�&��?v�_���k�ܙѝ�PN�Տ�Uo��G�&
t��ٮ�<�$�Yw��)R	�	�IE�(m]U�ʱ�s1�6u>D��<T��04M�z������լ&Ͻ�	w0-~����Z!����+`��n�v7�b_��RLm�0Ѿp,Cd�-�s�������S�m�n�b�;�Xg֪��b���-�d�'K{w�^�����f�����d$6������H�] �Bڪ�o�~�;��UId��2X�\���T:����
��M.u��.�����"zV�I\�?��Ƥ�j�s8`��MԺ �$���� 8گ `M�EP�?�qь@-ث��S�j�{U������M+q+HI�Q��_k)J�w���3$�?\�����2��R��*�+���Z���H�uʃ����sK��[V��G���?�d�����u�M�F�xN E��ַ���nWݡ;�2E�t�Xޅ�ӾBI�j�X���Z�?�U�`�W�N����0�.̓I�|�9�ނa,:���%Y�U�<N1�;���V�� �W&B5�������Q�	�u�|>1��T�MyJ�U����C��6`˭�q��J�}@>����_E��/��g�����)C�ۢ���6؆_)��y���rJs0�e�R��YH͇�DL{��es�m8��L�˘����� s��� ��G�E=Q�����3vSD�?nf�����{0$��Q���U���G6&�� F�X�*�>�@ 3g��8]�7�7���U� %��{���#����"��&�� sx��Ҷ�`��u�trz�)��ΛaB��]<�T"r��e�^�V�9��*;�Z~�=����s����m��f͍sى�X�	Y�4�3�=�8���,嵞:3�cj/�i�Z��]"����Hmf�k��Ɖ�io����G��&��ׇG�2
��e��:�)�������1�vS�x7��D~g%�ᢎ��ox؀ex�!RR�9�6��lFz���B���|,�|�ߐ6�Z[�a`����d}�j��i\:3���*�ӵ�TW��[��G��g�����o��*.�⣐s
+�z��đ"'��*�g�N�\�+�S"�Q�\mm���:���+�~.�J>��ƁF9h����0
Ñۖ�𓣶S��T׈����9BnR�3�����e�#;/�e��6����l��o�c��g�=��ɖ99��4�Yi^o��R�[�p:a�ФE�=E#费(�`��_�Z#M9�,5F(e7����Y9�\dGc�
A�畧XYL���V���>:���.d��EXb�GP�S�p��[34؃�?�]���H�y5����O�_�>�elC���퐍���1]�1❨JQ��|T�lG��!Bq�S��۸�d�Z����$����*80��}}Y������d�x��ѩ'�/�:�?��,vF@fUG�����7�6S�Ş�b�oჹ�ә��|�*�$A����
�s�D�f�8��f�p�q:]V�D�~�&�� �U��`�!,��
b��=�A@�&�I�--��aX� ������� Q�4P0>��!�r�D%t �Z&P!3A����y�"��7*1ć*~�:��W�Z����vc�P��A�\����ʺ��*4	��ƟǠ�8�,pUa�K%y��`�?�C��&�\ݑ�sz2Ǔ���{,g��V�s'����\��ǚ��a�Ifݤ9�u�!�,ګ[�C��`a�$&l`�k�4)HS���J*%~>��ʴ&��u�b�m��m$�`ְ涆"PW+ty�({vR*�
����cr�ܒ���nC@1N��7�����P*@���2���ҫ>���,-�5IC�Tsg�,�Ȝ�^�K�͇	�
�h�
��Ǔ}x�u�(Mܼ:>�'S��AU
YC ��'R��d�$��T���n$M^���̀�|�o�<ĭrA�/��%��<k�i Z>Lں�U�V��E[��ӥ��n��,xb�����~� \���֖�|�����f�*��}���S�;Qv=��`ɕX�x?�7��?T��A)��
�������AKo4�#�#R�:��X*�=���i�i��f���qL�|"��������z_�����tH�͜��`����Z��F�7#�9o����5}��i�_��S�$ˋ)++���x��:��>@/4�q�11�h�O���I�7t�k�աQ��[e���jF�p�V�S�F�hC:�Q���*�۰��E��p�QP�j�A��Xz	���`C� �����B�I�I�Uz`�
��{�@�����<*�k�Oh
5Ҟ	�z����"����B 4PY���^�]��o����Lyv��I����6�3)��pw�GA���xNI�T��_�VI=�Ňo<��9@�4a�u� B^���Ԯ�5�"Fh�=-�F�%rմ��fS���amH1k���� |�d�W��?�Xmu���o�/|%Dv�Gm�?8��k�`��MI��I-��11��5���_:��A��.�F?���n��|?7 ����!�Dda���������9zE-����j��02o�W��ZGH��B�\�q��Y�9��&��ZX3_�.��t�3�M�2x6[��Δ���R���0�#E��-j��`�up��N�G�0 �	TP.�Iu^6C2���ncּ�����)��^���h�&��ۯ����W>@��.���̛;O�_Q	J�������%�m����r�_X3%Hr�0�r���p�k�ϛ)pn䢷)�z�PY=�p:���/�e1o�Hn}�Կ���q����j�|ʘ��r����O�����]+9/�k�5�NX���O����_��}*�1m���B�M ,��s�Q�mַ�L�>��g_��|���,[	J���d�B+��(W������T8V��de��|���#��0#5�0�}�3Q��Q+Y��O3Ji79�J[�g��y@:������F���K�b~ZF��Н���wH���&�Ȱ�x�L�U5E���\�v�������wT�}^D䓂�KMC�Y��Pr�F�:4�4���Վ�:��� JN�3�l�w|�s�^t�ŀf8:��[$h�4�k��D��
��Y�5��l��2���ש���Є �sX^=3{���z��'�����Pg��L��� ���2]�@�Y�h��L��F�����>�1�]Y�籦�CςJL�e������b���s�ۥ�t�j���*��mq���7-9�ן�-�}�6[
L��r��>���G�8��p�U�d	f���uǢ��F���<��pK,�z0��"��0*��#$$k�>7L^�����-`�7�Ѐ-��%�s~ћ��LK�6Wb�q?1U=��<] 9n�ҧ��[�u��	�/��ɽ���gu��:`�j�.6#����s�dǡ�LcY����(�EN CUD}�5\�t.���8��Lꩩ:�Փw[�X����8��5�p�G��a����u��@m �|���峛������~te���]��*&����
5����e�*�c7��p|`{�&�tת���"f�Ȯ��)(P�3�uReE��C]ά�qAQ&�@��r_�XiXf�bL���� ����"F���+��&��Qw�
O"A�ޜ.��/�Ŏ��9o����>b1"��r� ��H(�l�6EF�1[9��N|E��'�m���|}}�Dg���F��oMBH��[�vLmB�Y�>��/'�hd�1ood1��4G{�����)�Z�r��a7o�4��`?���B]�U�ݽ��q;Hp�{ �0-���|k��e��p�jjb�z>,%%��Bu���kI�����k�:l��toT�.�~�yPi|�%R��v�f�q$������U�K>��V��f���� �(�`����}�� �S�[.��n[���u���s�M�`Y)#�O����
 :b�pY�����p8���ӷ��>\�.��iɂq��~�i��9D���%c��Yi$��ܰ�]��ʃ<d�mgWeo��`= a�)���V�$�� �[���g�9�I���5]��蚺�	}Y �2����O�x����gG≣�<���н\�D]dL�#�c�*�h��Z�;�Z�S�А��X�5t�&O��c���Xmo4��SU��;Ч��
���{��&�	E��S�w�辦yZƓj�N�j�f~���!x��m`˰Y�qX����ڬc�\��]�{������hV�Y�1�j���1�n$(��5iYQܞ��t�i�*��+�MϘ����d�M�(�:ֱ��.�F�q�M�S6bߛt(���H4H��MJ�z-���	�6��u;Hfm�^��&�8cA�X[�����8�7W�z�0�ᯆC^d�t�-����f 3��=6������`.˂ө�s�|�[2���pis��}	���P�fm�m�����Id�7��N�0y~҅s�C�ډ�P-('֧�!������:!��di���Z�Ƙ��,Kk��6�Ŕ�6�
�?�yތ��mS��s��O���U]hO3?�`ل��Z��Yέ�e����dJ4*8��>��C���lM��� ����$��׹9���s轃�6:����f��Zk�M{b����뗚��:wa�(���@a{5�y ��T�RA��a2��|y�j�ɖ���+��=S����frMY�XNC���b�ߙޛ���')��iCr�`���Y��34���͒{�[Q�IuD�����^}O��S�XDy��hRzK�@3��J�^u�#ة�[ח��t�����6��(OzK*43���������1˚�S�^	�,I��:^(�]N��/��뿖�)H�������}��Ns�B_��.�9�n���':<�q?��&�]�%�>��'U)!Bq�s��\��T3!�d@2i����[o�-՛dÿ�hg�}�)"�Cm���)�Gk�7Q��� R�ݽ��!|�5dɱY�N=��;�Ԓ[3��0�c�rW7�[k����_�X{:���U �\W�Q&��x^<�08i ^��d���J�12�*�:r`�FX��r/��o<�	w��݂�°�v���d6��C^d���=y���ȌL���՗I1	�"W��1^���a>.wϣ�L�1C��w�<�� ,^�U@������J<C�ЕKAF*�p��ߞ�j�tI��Hݷ+3<��!{�A�c��-����_%������ߚ�V�am�[ Ғ�-�!-Co�0�N�Y�?����:,N�l�NaU*>��_e�����IB��O/������94 !��:��0�4b�$<� b�r֣>[����f��6�L�{Bb��>�2�f�gS7T��;��s�����@��J��"dV�w��>0Ͷe�����/�q�4�d����H��R��O4�j[p�c�jX�� :�]�B��<��w��aF��}K�tS��tl[иZ���Ǌ�J��Ea��w����8=l����E��?58E�� �!F�2����~G~����5vT�%_�>�GE3k鍂3�$��ifnZaV���=�/]s�?�~���XdƔV��^[�ھ �*w�dR�y�$Y��U|�+�dEu3�!��[�ŔQ�d�� �<bc���%xs	���*E!	��C����n�$�\_�|߮�����8Zl�k�l��a`�r� U���m�vY�aEp�E/�0��Nly�1U=k^��/,s��D}>r�r�_&=�!�ц?�5��N}u�3�:k� ��d�d�KF����sT`��E\�sH�S��2��<���]gu�9������oR6��wXG/���M]�c�l�AwDl�ɲ�v�*"��>�0)?�����خ�D����W��u\���h3�f,�G�z���D��a�vI�笌�Y�i�b}�,��	1\����i��;�Ţh+x��{��jű@##��6#]Eg��cU�7��{_�Qh��^�B�Xc�!�&�h�F��j;��a���1����2ўW?i���]�!��)M�����K!���9w_��ۨ'��X� ��.@.��aTɩ�E��G�L����]I���4E��~�b)x�?MXT\)�Ҕ���O�YPm����q(^c��ep;\���E���%j�9�����5� Su�F�iRTG򱂚jK��~L�H��@�z0�!	&XŐi�1�he��&Y���Жb@P�� �a���[��/	 p���|.�Ս���v�j� �!�MOĪ����+?�,74��NV,hIdo��ߋ���%�:8ӷ��z���¡a�*�Nw�:X���M���_�x�E���ψ��x���h^�|;�I�嗠�U7گ��R���
!���*�/�l����Q8��p�>�CL^T[�$��I�G�B�nH��v^�*u������7\3S�km>�K�x��;0�/5	�Q_�rb�\]��"��0��3�Z�+毷�ڻQf:�q�:�&���Tr�+R��s���<�G��w�Ȥ�Xe3��ؓ�R`��[YZ�	ɜi3hE��s风L�h ����y��kQn�yM���ک	Y,��;R��X�HC�~���+�A>V<lR��@pH�_�x����u�LG��hݚ�j�-�a�D"�-p��I���П'r"�!�WO!��nb�\�zp�!ȯ:�D����  �&�U�'�a��%���О��P�zx��]d���}�T���'���,��W��7���dŬ<i�*^Ń�#νcX��f#ak��C����%��<,_Rc;+��[�W�84|��%�;�^FM!�"6
��5"��Ou���N�[�E���T���X����j�-��0���1;��9���1`�~��ȇOb���)��L��`фf��I~p��݌�+�2	��l>%��,%�Lu;j�޴��0�kjq�T���w�x�D���S�~�R����ā�pm�:���0B�#�ɳJ��XH�D�6��#�����E5S��R�j٥�>�Xif����Vd[��w"忟�K]��(��6~���R�����aqR�����ԩfF$Y�J��%Jn���c��]i��yz
� ���`�"��$���#T�0�\C̀�/�Q��E܄��Xxۋ�x��������C�`i�O�, ;�tQ@.gf���y���<�+�-���i�ҜS��%��Dc�)������`����P���cۺ>ܣ�{��y�on��bMT:�c��Q����H�]�,}|���|��j:�X�m���Zı�0X�dҷu�L���<�F�I@S��z�Ά�[����c���6��x�ъ���xl�@���75O٤����"x!�x�;�M�����~;V�tנ��M��U��c;�>j�HE���j��kE9y������H.�����p­���хm��3���e�Q����Bp�ժG��!D�Ǡ�������w\$ 0��d=�����?jyJh�����v0F)-|���*{W;ENJ2t`&l� ^Og�,�����X8Ƞ�j��gߎEmiw��t���4�?f��!#E��V����5�F�	u��sPR_��F�9�GN@0��Wn�O׆f`c�Xz����A�/��눨&d�U����T�U	����IiE�f�3�)���>����^H�)DYm��rpu��/��)F�� ^8H&n�mJe���m֮�4��o�J�;��>2jw������n9�$��ul�dR���� C��������x�i��J8_%�sR��t����Fʁ�h@1���v�w��1��<@��ڸ����w%�����I����fz�2�.�b�?�=�w��_�u��_��Vp�������%�!W���^��"�+��F�
�e��������_�)�a1�� �b���g�lb�sNs�vn�2q�YF=�E�N�fr1G�p��ځ���~A��:�6i<�=�Oo��^X�u��(�E�+im��m$�.j������1�_�<��s�Ϻ�0U8ڟ&�ʉ&�J��������-:��I�X��P��p�Dd����w*�� �!#(�C%�Jw l��i�46�~R��<�oL�����ױl���͋��XK���Ѭj��/���ʲ�$%ʒ	w��>���nȄ�(�"e ��}<>Ԫ���?�O��Hq�9�t3��)����ċǡD��j���� {>�����G���9��*M�1�x!��.7�HcD��JE鹔C����5EȰ�FeQT��UPҺrx�\'�}˩Mh�K�w�N�|����c����l�O��7�X^ff���V� �?����m��y��*&�n3$ҹ.�|hlU��z��|���(�Hc|F�T?���c�8�t��W�*=t X{4A;��mp������:��]��tE�@�1hO��K�B�='f*IuV����UB��I�G�l��:I/s*6u�7���+]�ȧV�r�$=���eD���Ř�V�k�����&&P�Q���|��搰Jj�^��SS ����^r:��g�%�'\!���J�^�D�����������os����q��|�d�>خj�1��S3U���6��$<�n�}dJ��H��˩�'�����}i&�_0-";�p�`t$�f�.��Km��l��#2ujA�(�ȼa
,������E�pJ�UD��Hҭ�I��]�5)�_#vfMߓN$M}JQU4�G^eU��EIiz*��B�'�V�S��������9Kh�:���P�We_��2��E��l��}gߖ�u�j���TA#�7'F�}����ـ�װ�m��L�;^R�+&I�C5��_��� x!J��vY�L��x�+��λ�f1�*�M5VXy��<V��Om�?W�魧|(��j���r�~�n��oG����?V��d~
�I��.�H ����{�G�
�7̲@QT3ί�2r$`��c�y�@��.����V0ɑ��1ˌ���\��g�PdI���%Khn��p\]� �K�}S�Av.���
�n�e fPn���#O�s�W��π ��R��(��/-���nB ����	� 8w��~%�b)��;����۝�I�������b��FKu�
n���G�����@�
�/�dk�8�I��Ȃw��,��Յ��՗=Pv� !
�b?��*'|������M
�#� �\Xͱ�����d��`��MbrHx)�����-2��8�8 C�f��Kd9\� ��9n����p[���:]��p����rV���C0�jB)�����06��R�k¬�g�轮�F@|>!ie�Gg|��GjM\����B�t�ۺJ���a�,�]�;]�h���
ѪdI,��y'��BdeڧS��ۭA)ZlP���o��m�K�a\��q�-��k�<�5�&���
ۜ�`
�y�r�}��^	��!�u�/�� �D܊��oй�����@��A[7��t7����M��j��J5E��O0 �!yf��#N1{�:�zd�>���s��]AL3VY�BL+�i�������Zk�|��b��ئϝ}oSY� �j�
͢�Г�gYG�Q�`�L�/���2h�_�����B~����iEy�W��=�^��y�v�6�M�ǿ>m0�/�`Za۠W�p��m?��«a�"��S&��g�P.��'��狰 .����s�$�jhb��>;��M1r�nפR���v������>��4���a�-5��O�Z�tt�8s��P�z�n��Do9F��_=I��^i�:�h㒙꽵&v��[�VQ��Ķ��5����A�L;w0�8���5�$�<e�-h҆hM��親�Ez���j �Ù%NC��˞یT���$�}Ҕ��/�BR9T�^>�(�P�g(��3���ãũ|nx�I4�]<xdXui<N	�.7+g5
�X�aj��)Y����:�y��B�_�@����3<��k�L-u�mX
տm��������<(�99�>�C�(j�,E N��A�<8Ʒ׏@��Ė2mw�cʓE��Z�?<�|DA��?2V?>S8��yA�=�,e_`�3� ��Y.�_���!�g��,1!�#�wtq"��<�Ԍ�g� L3�l�/���$:���lPD7�ɹC*ޚu�M\��6S�,��TO��V~�K�)����_��e��>�
�,��F�;��߆*Y6a���b�G�n?'t�O��g�Pt��)&���1Eģ_�F���z��"���������|t����dI��wڟC���ܧ�(j�}B�:����i���gj �]+�m�6��-k�B�(>�p!<tˈ�#�Ω�[W�T!�AQ��(�	�3�rS�;�I$
|؏0���V��C'c8���kd8�M4����v^YKç��Z�vUjil��/�n�1V���?b$Fe�>�g �	��ܩ�WI�e�G�,Lh1�PC�l��~���ܺ8&V�S0����b�*E��NF���:1bP���v.��즠�١��t��������L���Ф�-f'��t�Ͻ�������c^K��� ��	�_�Nm� KJF�N�}�\[�L���}ډ4 ���<�*�P�����Y���I�ˋ���%rY՚��v��e�3%�%31H�i|m9��V�%�6�[e�\[�;��7��$����SiR���'��t��.&��Ά����oF;���J
�Ӌ�s�tNT�x7U�s�Υ���J��V��Zӟ�.�Ѯ��kH��1��k��,5�df�b^g6a8�ۯ��x*E����T�>57���Q�������ؗ|Y� -_��{5�}��
CwlL�]��F|�,c���R�\�T�����zS�#�����z��Èi����>�d���k,�~��ἳ��'a�[h�*ԍ�ٯ-=�sh\��d�F�bo1[}�w��}�)�����tE��lGV<��:�ӊ�R��R��68sU���k�־E�\Lt"�����-�F��İ�ǛХ�A]�`=?~>��w��P)�3��ǅHSψ�7��̶G���}����$vĪ;�����i� �v���'D���=(�:oZ��~ �}6�L���u��8�A{J)��`;�Ȩ q��8p����BfR ���!ƥ\J)s�AI%�Ȩ�K���ߋ�����Ʒ����
	�L	��b��A:��y�+ɸ�WX.����.˔�/�;�����H���-����[��`�R)�b!�P���l
��@�~7Y��_cnJ��qv"�Gc�E�)�5����^7���+���@�M���2�h�Q�>��8s��/j8�T�YUY�{r_�����z�Lv�{6�c� E��!�6{�3��6��yna�X��!��)�n��s{(|��O��4!��k������ͽ��i�1�qN#-�����=�*�
:���S�<G4���Y�JOvG��z�=8Ŏ۫v���#���ik������*�{���f���i~H��p��ʎ��ee�-��_������	0J�B����+7V6)
��V��Xg���L@�-���~�����?��}�\�l�F��~V.U�\��3�LVwi3N���L	E���..a����A���� ��dfHla^H`c�5�X�i)պ��\��'\~�ߣC�t���v�;���c�"��%�K�p�m