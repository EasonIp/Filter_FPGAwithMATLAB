��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�J��"4�=�7(�T�JѺ�ő��,\��s���ӣ�F�؏B�v1�fR�K�`gP�qʻ҉�aQXU@M�MՌ�ng[@˟&&ql_�8�eL����_�OL�&x;-�
����Q�F��J2O�I�_/a��Y�~�W�S�X�2��sGNaC���3β�����;{�x�8�w�_;Qu�m.�1'�i���;�an���
k,$VJ\�,���/�����B�oH���K�Z���䔊���e{�9&����T�,�R*� Stq�|Z�BH<�;�X�!���Dd�$�i��珡 �Pb�|~��^k�3�����AI��yd�yg�R����,�=�ڈ �/�<\�Q"���0(.��0V��O��1䩔��N�?��X+��(��u�>���-w���M�=��ؤh����f�|��YO��nnz���?-�O�}�lu�OU8n83b?��*�6L�� ��-TOb�Ȓ ��Ʊ!�����,Y����fm��!il�#�x�d�����#Y��x�yl-��dn��'����D,�k�������TX��
E��Kj��k<=�:S���&%��~�Z4N�t���Y�o(7�b�M���]�Y��,�����\f�'�
�B���l��I4yM|c:�;0N�r%����ѱ׎�|�d�#�k*Fv[��=���E��N����7 K?�r;O�A ��s1H^�9�HTWJq�;�c b	ml�7߻�3L"�kf����Z�!F�����(����y�AX��Ctp�GJZ(W��T�����K���K�a�Ё9�XvV6]��κ��EL��ܚ/�r��U����P�������o�V�ib|�� \�qaC�1<�U��ͦ�=Ԧ���� ���ѹh ӹ�Z����~]V�]��Z�Yg>w<���Wb/F%C�^���ߎ��q6I l�54b�Bΐ �����)�e*dʾ̠�vb�d|��{�ք���p>LF9�-������Ή�3���ؒ��1�I��:�W��/g!��O��+�"�Cd]�i����@�&�ʞ�qHN��8?��C'p���7S_SyL�������u �?[Au_��d-���t� ˅M��U�~��gJ����g��?�c\����g��xE�Fp�O������sfO��b����C��V_��SLw�~��$��6~��Ƭ�����|�$�=+�*vw��O��DHK����	���9�E�oP<�v]�wJ�q[�d3ܚ&�_}IhnC�=�țϣ5�-�Iz�
���?����Y	s,�5�����{�.�����1��|�[�S�?�I$��T�0�GK�J�nw���$��L���-��}�k�,����ß�W����G b|&�cI�l�6[0D\XTw�,!}.JH����%^�NB ����uR���@�҅S�7�ÿ�
�1m|�)�ҙ�6�:�[�[�J�#����,��8p.��ZDw��ZSqQ�&x���[�����c��¨02Y � �~�1,�t��#C3_�*Ґ�2{/�2iq��~a�����c�@n@�}��?���^X8�UY�Z"b4GK��d�pk?6n�K���`��{��W8����O!��QuxL�N���RJJ����kr��ɻ8Y�̥Iuf. ����j�uQ)�)������So�y����.���Tc�83Ky��! Z�~]��_��@��1�1T��������э�u77� x�`��}�lE�}��V���� {�X�G������<�:�	a���W��M��vL�1F�F����+��˒{�%�:w!���9 +�#����ԆFL�R��Snz����<�uXiu�q8'�c���@�������� %��)ހ���s��g(��f���6UJ<H�7\�_/�m�}c�=	 (��Vأ��Yޗ�d�s=�����#*���5�#���\��f�m���1'Š>7��<���@�I��:&v�4�}�i��vyX�
��V����u�+�~v ��D)smb�����.Q�d���������܅X8,��qb@�F��z!����&�N&r�D`�d��w,,��+m���p����Ga�]+ne{�ƐDC�Z���Z;s�.h8�Ǆ\�M'd �*���=�*֔�͖�G*�N؊�4<�qR�R7���X?������u��WT��/��&�o����'h�ӊb詵�P�A��d�i|�n�lg�d�_��$K8'N��#>����ͅ��^��NA�H���9=)_]�����ŊQ�b6D1�T��H�d��Jz&��O�ٞ%-��[�D��I�1I_�:]�E��"����R9Dy���� �m��c��˻������>�u��ο灸9������?R{wq`��:�,���^��br�~��B� �v�{T�?���p�s��g]�L�`>��"�z��	e�]�YA�AĈ�$�3CпP:!�ig�_�7=��������z1 P������q�L�FWt>ڲ�����6Ilzke�|�sB��c;0&�����y8+��n������c�6΂i+F�
f���4�=�q�i��56Q��8���M�YS�ΏVV>sK`L��#]��X5[WI��2��ӳ��C����J��3�F���-s�L{BZ���������0U�.V~x��3ӿ���8��B�PM�c��L��=�=��k�O�
7�#h�	 "'$b��������4�V�Ui0����
z��6���v��$�5ZU�Y�GĶ�o|�tҧ%���X����O��hX Jc��p,�)�l2w�O�������-���덉���ˌJl�f����Z�v�P�B]��^�t}��Y<�4��#S���el����\i�"=Ҡ�>�;��#z�ޯ�(����K��'�a��['ڣa���+���������q����97C����Q��T������"��{��G�s��<J&�䁴��z�
�_�۪L��,��=,�o[ -̆,�b��6�/Zѩ��ȴ�5S�5�۽���k&�@��?1�܄*�Ȓ�5Sz�a�[\�{�%R�(���QunA��t���R��D��0W����r+f��ϛ�:�1�l�5��pħ�l�d�Q�������񷟰Y�5SY6d��
c�6i�ܴ(������М\{d��s���05�6lf�S�dL@=٥�L��m�(��4�'�7�Rщz�ڲp��)�ּhzuoP ������^a)�6����}���7��K��	��$�HH쓅��_$l)�U����ɀ�����<�C����}Q�θdύn�����0$��h	�
�F���Z�'"��w�ȕ}�ڦ�g�؉�h���V�B�,��xJ?~WϢ���+�1j׽�;.~��!� 8e���[Uv�K����mT.g�V~[��+"x�d���c�>���
.e�;n��T�0��?���B�.b���b
%85铹B^�7$SP|���K���"��z�wT���}_ �{�I2h�3��Sp�/xuAYt�-Pjxѓi�=��]�d��b`��r�1!6u2�"�Խ�����hh���"3o��͞<�=8Q���s6���7��W�`>�qʚǉ�3���;��wt��Y$�!���R<<�1���˲�ĭ3�Ȟ���K��d��"�dx��z)�B�Kf���ބsqd+&�9-6V^1҆�h�T?���ڗRY�J���Ӿ ,X�"��|��W��Sp�kz�8�
=&3���"W��}���cE����y��~nI��C���)x��=��GFP�%�P"�1�/�f�D0��0�V����Lp�D`�G��}8n�n�?P����	�AzO�	ּ҅���w
�����=�Av"�c��5`���Jy�h�Z����aj*���8���D7Y�����^�س��~u�-9���Σ�N�O�ɉ	�@�u�|�֛��[�Q��D�=���Pl*�u$�%K
mX����&���"Ej�r�e<@%�L0�;���C	��ǌ5�:��%j$��|R�u������(K�qi�~	0��T�f��kb��1>m'����E��Q��sֳ����^:Bwt}oX����(���4���
M��Vk]��!li��!�fx�u���"����ӯ8�yب�SqR~���iQҡ������X�`9Kݥ�	�Nఙ'�Y+������Ye�5��y���ʋ� �֧��{��ѓT�і�
������1�V�3F��|�mG�7Y�e ^��|�i�l*y�D8R�h;�[EI��48~��ޔħ�2fPQ�Aj!n�$(�s�$�)yC��;6���[<�Iy�{�V��wu�lK,-��^�1��	7>��sd�B�П\-O�w��WY��{-eU�Z8��r�����V�%�[�8����:�ՠ���gK�ÿUŤC��5�ж5\��Nm�֕l#�A�I��LU�@��!er�I�7tMx��
c���*Z�.�����q \�s��J7��p�.��bE[w�@[���!L˥��aB�sT9^<$�9l�-�{� ?���/�D=�}� .~�f��+��77l�s��]�5�Ǽea����]�r��=i��`
�P��\P��蛑��ӆuA_�AW�b��;��b�!���E
�rڪ�=�{�C�/)�\�=ZA\�$?�\�Bt��#ne�@_(!�g�f:ݘ�i�|P�	Z�8ze	���~3����b�1Q�u( �]���_�ڷ�\ge'Ukʶq�&�ڌ�jEX���N>�H����Y�4b��T�(�j��b�vH�j=ae����d9��<N���9��+�?Eb4���vP>5`>��@�4Aq ��U��ӼN����q�37Ŧ�G���"��+�^C��%������ؕ��)�3baIR����8�h7~���+�*4S�@{���ꃥ�Ϗ/D���Z%�T�|�ss0����v�əģN��,8��$%��΃(6'.*�b���eEut���S�p�(����$�ڋ<&�*(�/��M�9�ۑ���ګ���s��<U��[���b�D��4Q�ֶŲz檹u"��N��4ҹ�L��Bmd�J��&�kvc������/mU�� �݈�G��i��}|X#�(��vJ�SFrf������X蔣�Kq�C��L�;�pp��̫l���ϵ/�<��k7��Y�|��5���9������J8����g��}�^�u�sqÅ���n�[�9��)����\�#������[��s�F�R���U���� 2r�1�9����XZ��@�`�o*@T5%ѿ�o��9�0��񛣖�W���?��8�~��%��9fi�X1�>&�v�S�m��p�q(�pdi�cX]4�e�Lٙn!����Z�\�p����)޿�K�Mk���L��%�"��̏'�~���t�;ł�5��j�.[S5�R�{/��'.�?�fZA��7���𾉠�ی#o�N*LLX�G5U>]L{_jXHtm�cT65�F6e�2M6�?��8����d���8S��k?)?/��V�5�
="��PY���KMK�ѫ!;p������e��r�9�y�4���k0/��߻����������5�о|��)r	��T���4�����h�PB���`�&��c��B5����_���h�S튺l��k��m4��`�8 �J2N�H5�f�<+����_?��*�%�}Z|N��{ഁ(��&O|���ᠺ���o�5-ތu�������.�O���,���\�Qx{4���0���"�,\_�&nDYSjT�Xu�����8VT���-����d��"���o?��{T(M�����N���ޛ.M-wr�|!�����ysG���A9�1%�1+��K����w=ߕff��@d�d�>��)]d�O�X�^���"��t/ �����ï�V����5Z�zG:�y	N�Z��$�l䮽�[=��Y+��N3��t�	�2`�}�m�8x���u;f��?�0C�A���X���4�7ž�R��A�PA9�1v'�-�y<-\d���Y�"��9\�����z+� >FVvK�l-T>������H�,$%�LWF���G�Q)D�]�%s?͞J9	!���%��00�{�%:ȓbk@�*Z��یtq��yb�'�(�*��g��ʬ7�w�Lw`jg&�ڨ�hA8 �`A�V�Nӧ��o��m��O�q�����[��x���I5��(����s-W�>�Δ�Z8�U7�ek�"�����at^���������8I�������,�\���I�g!ƥ�qDU#_���tv�u_=�+���jF_if��Q��2�#O������� ���W2��!���2����B�)*)Y�Jc�i������*kr�5{�/`Px~ �&�(��q��*��+'ˍd�����\9]���3��kG�N���[����������Q�Ɇ<n�{;��<��Z��`^{k�h��^�������͐K�m����
F�)BQ���&]��!�Ji�,6u��U����֒��<�_9l�J��Nc�"R�`{���W��^��C\�V<Sv�It�b-
^١�C�nr���t~.-�n`��΀�xQZ|��덫~���0�\w��g^��;�ֿ��o 류w]���� G��R����g�t-�<�V���в&��C�Ԅz�V�9Cq�� ��s=�"R���Aݷ&>�%���>L��ߓ�[��ρ��Z:����Iﯸt����M�6q�W�в�%-�e�9rN�?���Eg���H�g*��F����տ��(��`�:
"#w	ԩ"OH/���TX��Ć}��'.I%,f4�^PX�3"�T��w���BM��	�!/����I������� ,���;�2|����͈�]w�8(���q/�ƀ�ܿ�{׵����ty�e��c��ؓ�̴���!m�::�����4[�Lω�D��d�I����T��o�>"$�?��gЄ�b��;Ɇ/�{���_�AF{4�>�E�����o1�X��Ӕ�U��G��D�Fb��0B�7�/���EC^}nk� t��ܤ�M@�KfW����*b>ǸCy�a���I�3f!k�"<�c��~4R�tȹ�뭻����N�m/�S�
--�/�S������~j�5ʑ��K�h���x��4R��l����I��6he�\3����~g��#�B���è��
F��	'a�H�z�j���dAK��T�+�֢�tq�"m1���Y���r�6�ޞ�������t��5��s7ƺt5�	WC�W̾��]��";/�F��t��C'c��@8�L>N�gŧ�}U_B�,j�^�t��s�|�h�a_��F�c�zP`�w��\��"Q�Qv"e�_�T����� �o�*Z1��������{�%��*�o�&�\����wl��#i8`�\b�R%��c|1�QL���"���:��8������&���u3��	�	���]t5 C�b;ӳB��9�#��_�͌ۜfV��`F�+���6�|;��g`�v�S_��F��Cob+Z�urs¢����%������X�����f3������*�3�J�H?P-�@E�
 �^j�����f�g�|��p%�4�	�hq`|%�g��p�-q��_����Ȧ9^ݱ���79	/b�k����q]�$���-��ҵ�;���.ӟ6E��q��ѷ��Dwϱ���:��p:���W��FXɕ4�O�*G�0�d����r���h�Pf8P�2��v�WсFș�d� �-��9��L����k,����������m$֊�2���C�鴬�l*S���5/����j'<�0L��M�U� D�\���p��o��&����\�o�Z
��[*���;�u��H��f6G�;��M%�æ�X���j�sE��i�.�x���6��V
+$�u�F^xm�A����N/�^�3��a���R��������� �F!o�Z{A]X��k���E^���/��&T��~���M�8�tk�}�;#��t�� �&ؠ@�Vl���/�%�7���VU6Nі��/h�����X��ĵ�J+y~�-��ƃ���$g��D��B�N�1�a���U~)�9���<��"�?��q�����mKo-(�9�|�:lʲ��w���?fp��1.K}�v�?����ܕװ-�5b�r�������f�Q�w�����r�f�P�%�]��g[K�XJ��1GkC���^���b�̎��^9�h�~	�o����yjY�:��*�7�:S_�X��_S@�&}c���=�u��J�� �llOƒ��f�����:�J���|�9�6I7lq�G�x����~�_c�D\d��Y�;�N�������ۇ�s,g	=z�Z��0$ͅ4�f�	x��#jeG��ĩ�����i�mK8X�:�p���ņNw۷O_�&.:|��Q/�:�v���$��}����x�d��A���t#zt|�d���g3=�D&F<�0��`�B���pQ\���S��x�4/�66w�����@��ф�=��|��<��YZ�����˾)jZ������JD��{8n�FdX ��`����4�0��H�^;<YI1��d@1��h6��5[pd2͚����}�Y���-��o�h��b?�L��l����-�,������_8��G� ����G���Q5q����u����3޸�",A�R�WK��7)<���q��#�XPr; �B�l6�2z[4��8R��YU�Ƙۧ�kȒl<�4���aw>���p=�N�C��Or��2�Dk�.�Q
$���u��>��5��
E����8�W���E����H��wD����8ǂ�ޣ��
`	�is��f-���z�:}�����:�G҅#�	��L�ۖr�������\��D��t��S�dE�� FMS��E��杬�8�\֕���<XD�1뭮K�߷��ٷLso�A�9�o�Է=��y���X�SbsR؈���Fo5]+�����H��<v�Tn��f�T�?HτF��sS��$ae��u�`��[d��$-"�$x�BK��aQ,b�`�f��8\\��|=�كV����X���͋	lz[��;�s��*�nX����H��s�;�χbZ-��KY�_�V�;�
�����2�%��*ȹ"���k�>t$'�԰WS8zRP�pA=n��޷>�l�f��-b������~�հR2�h�P�n��θ���*�~��DQ���:���t:e��LB&�z��H��n0D���Q�rBL�0ͶآL˘%#��JL����@�+ĊJ�/��)f��uu(�۱��H�R%���+�I�j��~��Û,�eZʄ���X�qR�B]�|KD�u����4-~�~?�n�}(��ݸ����x�[_}+P�Z�`u��5�&�g���9�%�l��f7�=J�����p>KY3>�$C}ih���#�A�Mq���c���'���HX��^�q��8 ��×�$���BHϭ��R;2Q4tP���U�q�#Ҙ���0o�:W��vYC�[C��,�IP�i��u�� [!�A�
8N�_������},��(��A~my-������]��=���Ksy����OP �n�D�K5������y	�����-�7�d-�:�4f@�=�FF�)<=H��x@�>�n��v���;��͠�Hj]�ȧB4p6����|�����1R�p��߯��տ��?����X�`��t��^���M���Z:A����.�<zG��(�Fu	t�(;8w|��\��G��lS�-�1���o�kZ\K2<�̑����R[K���ڽ�XJxN�hZ��&��v7�]�_�*�=����hM����l<���?�i7��Q�Nj=��L\aE ;=�`�|5#�u�3�}E��!MR��Ɉ)��Tvy�џ(F����JW5�DJ�Rh��h�B)TU({��^�]�)�q�̕:O_���K��3Q����I�5���l����3�73_�IP���&��ﯭ���RJ̒���c��8B:|ᦲV��JL�f��^�G�4���zB��`&��a����	��V���s�T��
�t%:��$ݞ��EĒ���{�\ͮ4Z~7�<�L�U��_�k6�)�� m�]�d0�^8LI������q:�6��ZA&&g�^Ll�H:�b�%c�`��.��&7�0?�k|��6�d#nbߋQV ��k�Z-r�g��Md�.x�y�����݃���^^~/�m\��g�N,�U�p\_D!T�y m��zI��#_d�(����k�H.U�MU�yܧ<�cW�u[ا&��m�R���4/�giz��%�̍´G�Qڣ�o�Ma�l�h��M�!飂 ��4�����sC�e���������X��+5�	�v�t�}.��\�Z,�����|2&v�R}���a��#VJ�m�!w)�&O��S�1b:��6�ۼ%p�km��P�Gg�D��>�j]��:�)�Us�C愤WP|�'�@�,�o�Ϣ�ߋS��Zh�U��
����d#hz��&\	���F�Cݞ�4/�����
��D.�vfpJV"μ��x�Rd�� �=���W
w�c�l2ѸX�!P�w�<H��rq���q������/�-/�kQE~����'��䥱��t�(?Օt����/�����U��o�L�!�`��0m���*�"%HAF6��pL�nRe�e����<��8L�fI����q	�0��v��^����ٟ���+�='ٯ28�l�&{�i�w�%�+&��ҋ�f��K����s�8� ����2e�}��P�@8����e�˦��Q�)OX&�Aƌʏ���;e���6��RsO���M�v?\6���)�V�al���i"��]��kx��QW��y�Q7��U����-9̡��d
i������1O�W�����f�l�^�F������>��,|�p�hVbLK�� {��8��no�ѕ�2�|֌s�#��>�iLǶ�j9�L��u�?S�J��ɖ5W0>�ZV�ͽ_�*�攘���d��Z,2.�
���x�WZ��U�h�U�MږY��T\��Z_�i�4ɇ�L���נ��#�{�+M|�	����.S�"�d'����K[&��⊆�DheoӐtl�q1�ۻh;W���6U�F.c����k��q_Ҁ���l�u��V(X���T%�5B�0� �
�5P��oN�n���6z�Ƈ ������C��*�=´"iz��I��.}3����K�e���#��᳸��`�0ں���tB�������[d��,�P�Q�&�9��cPbEU���v�_�k�D��u���#��1��iR~])�C%���x�ɡ������١5�~7V��-7��T��[�,���q �}� ��
Z��dA'e��]�B/c�}����ɏ����8�Y�}�T�	�eD@O��@%�O�ZW ����d᚞�-z�\̖o���*����T�<��6x_Q��bq�u=���џ�Ȟ�K[K6vqW���T er=���LyTe��瓓M!��s�
�/���K��ϯg}~Rufǈ��D� )�4�����^�9إ�I��Nm��M͗�W�� ���@y%(�P/#�D��!ݘ�wkd���8Z���c�9,� ;mj����$���|�0�F�+Ǯ@�5D�÷�^ ����ä2ʁK�O.�aV�{6�H�)��(�J�[s���@t�� ���[��A�� �|���˱��AHSh���c������4�2�Lȹlt�"���z��?G{pB�-tl�$�mN�.X�g�e��G � �N.y"���r�pI�4�=�t����
�[��N�x��U��1�e�CN�@m�u*�L��}cn���A�ȭ�u{�U��Rؚc�$����ê<�)
H�T���Z��N9)�6����s� ߵ���3:4"�Ժe|��&�6���w�q�ИW�O�W6��P퇳�yTln�>B&�������h�Sn;ijЄ1��i ��xؽ��m9L��p;v��*,ĚUh���$�������0�~�g��uLD�GR���������Kl�oN�/����%��\IjT�	�1/�A�fo�DѴ�r��ZS�u�����=����z*U���i�`�)����v�]�g�6`u���D5����	�
�O���e�Z-?&��n��b|3�b[O������p@GQ�#�D��ͧ�AFS,�$`�y�+���`��0{��i^�<|mlLy�k��d�I�>�D����N�'��3�ჲ���|m4/;CI�#r�H$.@�%N�Ck�����
�Ak
ji�o�͝n�+b70kH?���&x����N:�T.���Gm�.��C]�~���ʏ��H�5��}���-��5��B��N���份�v�����qcɵ�=�+�;�Tn��G�PE�Y<�s%^{r^��q�������
��l�JM�٘����?n���l��Tt���.��@���5x���:���1��/"J�)��Qen����o�wa_�~�(�7����8��+;�l�g�QmD�<�@�G}9��@��K@J�z�Š}@�TY5�fAt�P���BR��k]{=���c�Ɔ�Ե�Ex)}��9�8�YF?�����t��%i����i��T�*����_���8a�QR����ŋ��%d��<��l��0xƛ�H�E��}*�G��#a�?����B�' ��ge�4RE SS��v��2�v/Ե��k[2�P�18�+FL��@�Ⴤ*��lc?'H�-msY�D����L튗��EE�Zb�_�?8�v�f=yc/��u�I�O�E� [REn��|}�T�4�/a�W��JX�a��
���^?���~���=���3qE#C���߸X`���РU=F��@ǵ㉡�$?#��nū?��b_��(�!��S�D- ����c��̱�����䶦:�;��w�1�����
�^
S-S~�޳C 8m�xU��?S5Ri'Z1{U�����[H�g{S��B��`"�ދ���[�'�p��ρ��^�a"�g�ݠ�WR~�qqt��y6���qV�~��V��H��_�~e��aV{UeS(��F%��N����)@ѱ2: H�o��w��go��:�j�v��@y1����z�;�?��e|��5��"A-��l�{ڳؐC�3~��o�{B
PC2�Jr�hm��F���v2F�*\M��y�����6�4a5C���IS�<�ʾ�'E���nT(�)��95	 4���X�[ A'����S!cef��mʙ-�pd-��*�Xlb������?�K��7k��z�m<n�l���bO�X@/�e��Y.�@��#> m�K|KXN�E�g�d0k_�e�^b�|�����f>�9�.f��ː�h�9��X���H�2��s3�ӄ��s��R��p��(���o�8LtB�;������9�B�e�U��>���w��- &-{7<�Q�d��"o�L��������O�v���Rq��<~9m�]��՟�i`6��#|�I��|ڟi\�J(�ފ��=T��u/�rH Z6R���?�j�����6�\� \��\�GgN:���ꉗe`~%-�[���y�Ե�Yh�Vd�a�A�S�S�� ���'	>���wA��վ�2Z�%�"NڇvH�ߢ
~�B�A���;|�yo�O>Eg<�����a�[���Y��!"��:}9N��H��]��Djn�<YWO�l�-�HBdĎ�-v����k9H�V�a�����.�+''G��O��$�j]��ڦ/���w�괞�ۗ	�oY�
0=u��'�����K �ҙ;��lg��2������F�~�.bQ��s��K�i�j�	�p���~w�z
����i/�5�F��z"��=d9>l��	�.m�	�D��W�$��[�����õ���m�6iFe�*�_{Y�޶s4!�y\�� ��ķ'�6.>�v��G�`!��u.�03U6��~�ͫ���5�ҏ{�}l�q��\b�x�%\ܯ�7�{�I�X��I:�3=�S\|R�R+n�̙i�p%T02�8�6Ϥ���5���g�otEheh�����>~_k��c`�x��|U@;�z�W�����r�T���zB8��<!�D��xx4��gg8���O�e�C������Ft�tS�wą(f�TS;�,�@*6�Bßc_v*�؀H���J�I��q�?�ާ_,�Z�F]Ѯj�kxǕ�Cl�dxuj�4�6C�F����1��	2v����g�ͪ�J4�vq��e����Ŵi1Ow�h��K>�㼄�Zc���,=f�DN�!�bi�ŏأ�;$��3�C.����GM^�{dy�e�wl��p�Ө�q�A�ڮ�X'�6�o8�SI$� ҫ�ĀuA�/��$փ�r��{TX20l��N�uثc+F�����Ƨ���Q(��U�TAwW]j��p�M��w�*Ttۦ�z�r�9+�v��쒝jA,d�ˑ<���RT����H��t�K|�'y�SD����35��
�W����������
����Ǥ1Ĳo����9T����j�º��#�rr��R�� ��S��?��Y��_��Q����yk7�d�'�;G�&�� �?�]�Ezx�><mj������d[�֯�yX"6����X/߫]���n8��݌�����+X!%�OE�5*c��^��5��o������q�I�sg_(���x���k:����r�E%E��E�f����suݧ&��G�`#�:��-e_B�*�}�]?�>F��7���0�	[;Y)��n�J�� KWY
%8o���e �� �d�hf�(���"�	�Byh�0��E8��ڣj��7��Ԁe�T�e�~)�*�vB�l9�Z6O�	���O�"��P"�aS���)x��� ��c���^ ��>H�ƕ0=C�A)�|�qQ�4?a�1H>���������Zm�	p�J��6T�%1Cv�Lp�}@d��d햜�;�#ڤe7 �q2l"I��>!-}e�-���ޏ��Q~7I�zM!����F!��Q��v9y�/�p��2���S�j�������Ԓ��C�79G�5]ڭ��)'`C���#�_�)IˎI��~8�߫�W�q ��`X����x�u�}h67�z��C,����uQ��xQ���0,��!�O�2z��~Ơ�Z�,��"{��g�u��4��Uøso	�}(V痊�>�o�?��-��b�.���j;K�P�".dVy�4M��W1
Rśμk�9�&�gm���P@v��rR��JpSܙ��էz�D<�l��U�����9O{������O�J)Ě�������{G?�R8;w���bVv�j�Υ��̤�8�A6�D��^�	!H�� ^Raû_����+y�6�x��ђ�Sv5�'I�S���`j��������f��i�����:�7S�W?�@�%[����d��ԇ�k�8D��[��UN ����"d�=@JuV��A"n�{�j/u��L:F|�
i���NW����:��Pv�[�J��H|��8@��H�)������[�� �s�&�������0���F�?�&��,�r�N���-��仉���B����J�E+�2	��#���I�Àa��o=�>*^
�D�~�����zd��4q#�a.�B��[a� T�G�)JH���E�_�����䂬n#�	�9j�x�4��'��컐��$gqltE�E��=8
z��sA������P8�v��Y�ņ6"N��nco�!-Ls��a"����c��>6Z&h�?'q7�1���AB���b���8��X~jD��9���T6�+�6ٍ/K��'H�O���NA��u��L�{$G��@����QD?��>���@����a׉���O#���t�ⓥm�Z�8
����s�RqM��>���a}�B�׀���.�g|��	�٥Y�C<x�ߏPWkbi�n�%�����X�L�&��N�w���_�!H��cN�-�t�lٶ�m&�es��wem��?Q��yD��m�\`��(��
g>
	LŰB�.`��
w0mƯ����n��*>�V��`�R�5��T�@��Yi�%.귢{�V�?mC����U\�^"����WbR��$� ]�QM�L͂oKY�%_����дë~ځ�u��E��s�q�d�߰������q"�[L�֌�l�y࢟hF�*�n���G~l�$�V7�͉�8��H1��<����� �� z�J�\�8o^nR\[�����*�P���)����� ���T�r�e��w+w���"����<��ΞV2�X۳�-��-I�ª�|�.\�^�䠉�[l���k���� 8�t�Rѓ���A��r֨�G��Y��K��S�o�|�wў^��*l6��#��|�B,�U`�H�鿖��!�u��k��cI�bdO�{��p���Z[�ʠ�4UAic\=P�D��'7���* YM�P��^�duS�߸�Z� �=��<�n̈́���l�[ ��p:����y{���Iz�_X �uH1k5*c�
�ni�}�ي�j�\לu���`]c��1�Fn��;-��y���̘�Z�Åw;�S'���ﴄ�C��2j�Ɇ��3D��F�9!��uS��<�4�C���C�|BA���V�l�Oq�ʃЌ�>G)i��ef |9�kn�t%pEd�6�?GY�.� �o�Q�jW�xR8_��'k���'��ae2n�H;Loś�bJfoP��ԼVS��m�  c|9�3���C�r�B�H�I�=�$a2�������C�P�$��*c�k���Q"�.|~c*����M�)%ɔ�;�K�ý�myK�����6p�#��F��qb?2!b����jdp$U<
��i����j\A�O�L��=��g��p�h�`l:����3�_u�$>���)�u"5�s�(C�IC��=E�"be���@����&�kq�w�W7���Q�?����Ӄߺ�n[�7�{9�y]ǀ�&��T�9&A��8�:Ä9l��q�)�-ȃx@�W*�G��5�Dy��k��pժ����4�z+��O6�5Зp�AQ�����!�⊡�?� �jql��r���Dip�ꤧ�}��C��N-E��9�i�; ~���-H����[x�JzO��
����t�TH����X�e�-��J�Z) �1Tʼo���_L��z h���)C>{���E�H]��TW�ܿ��e6�3m��֖�=�p����<2��s����
�>9��=C���!ٔt�M�v=D0�4x���/o��#v� �	�h���2�h�VG�6�ϫ)Sc�a�2�C�t�r����W�yPo �{��R΂j��/D�U���?��[�J��9��52n�����&��T�N���2LD;�'�ylrw�l��13�`}��,����e��%���i�t���n�սJ�d�MEhrԏ��z+�t	]��mG��M�K��`�0��Q����Cx<����&��_�5���ACq���)e���Ӊ{Pw�p!��\�p;�&�AK7�]c�����2U}Nz�wI�(A�Xw1���<%��=�p_���!�9٨H��6u���#��f�
��R0p#�ˇǇ��]|����͢
>(��hm��AuNz��"y�3�j�8�]�����ڋd�� �r�����3G�u�d�\J���~<��F�P��$����j�fr��s��q�	���]w�敿р
�
��b��BfW��4W+�I���8��5Z��;�4�/��'K��)Q
���_}����~}�0{�z����)�{��2�lX����|�d�+�qS������s�v��Ȑ�����F�A��=��!Qe�AO��C��Kl�)}��Q�;g�4�Y��#d�ct��SN�����2B�iJ�|�'�a�eO��vViU��n���$b�6���:�:��lb�I<`z�'�t�i��|3[r��<��	L�n�b�)sI��W�I�ūn�/~.�ݍ� Ɉ�Te�#��6�3�	��N�GdD�l�?E���yZ���
�wb$��W����uřw��Nk ��^r�8�SxE.�s�]�C\��*Q���獍|kAS�{��e�@����C/ی��/�?�`��>��A��&߽�-kI�K�����{�QP��p����ƙ�`�Lۏxb��M"Ո/agL~�B�O�mv}��q^<��m7N���|I�{���p�B�<���y�S&�c�Q���q�	��za���E�v/�ȩ�Q�1!��*��3P�'�7^�m�	C?�@0z���S���Z$��
�
Wp�+�JH�Ӆ�ٟh����c�[�����K�V�0CLy+�[��5w.��5�'�t��1�,�|�.Y�:ZbA0�m�mqwNUƵ�p�U��4ᛍx��rOq��N�bKZ��?�M���IE#N|~.�wX�Q�QZH�aP��u�nǍg���k�&�/X��o Ҍc9�V�l��S/��41��v|��(U��2Y�Л ��]��=53�]�r:o�c�������Z��֥�4����{ƍD7Ϛ��#`$�;�8�6~��e-u^��	�^���L�ǻ'�ً ���� �3�F����ŖeݹV���t4�0x�b@�N�oн��H��<����J&��p�)|�1����:�M$ys}\�aYag�h鸲כ6׮vĞ	��x(�v>~1�W�ڊŊ���D�b���3*	R��	�W8W�!1��A��G�Ϟޏ  �-�9i���:"JY�����9[g��5c�?2���6�I������L��(O���7�'��lz�g@{���^�f58]q&17Q�~�q��E�Og��$藽?�Xg�D�<P��[��ED��h~4��([��{d��6:&��d��]217��'���V[��1r}lA!���(r�5�.��䑻�Â��+TW�~?���eb.=x������`ʣ4��)Pj����֭�����j�px�8m>/!�ͺ��M���:Tߚ����*���3��X���5�;�5Ʉ�����:�K���̦/D����Y%�r��U��׏P\��)&qaU�[�,�/0� e��4\n@�x$߳� ���Ea2�4�Q�.p�6^ְ��,��Y'0*�i�T�a-�wșΔ�':V�e} o��dkE'Osf�-=���B�۝����Z���!����>�;���7�3��:��]���Yg�������캊�܀iH#���e�	}ƶ�j�^�,�9`�S��w(�`�U|���'26��2D����f��e���~���f6�Z�@����W��ȳ��,T-6��jo��9�ߘ��L�y��=��4ރ`�_h�8����篛����=I�_�ۻ�C%OO�R��S�tdԊAY�O��	���I��b+�ƻ��j�3�!�k�#��|HluΓs�l�}����lLՌ,��Ϗ!�
ᰄD�^&=%}M�����}�M��&����nx5pS�OD�m�⟽��<1zW沃,ޮ,!�y�a,��T�{Z�� *bi�YnU�LB |bQ�:P��o#���ü%p5\���F��rg�&Y��ٸ�W�8�wD?h�O���oX�M�#zq`h��}�}��P(��a�
J��E��EjJ��Ӕ����T���W���"�%�����we#c��j9�����L_��4d�}G���)y��cA�΄|�^̇ǳK�Օ|����W��PhC�|�YTbQ*����
�

��n�eda�V~֬�E�;����'`|�'p����0��1a]n����O�2�u�]��L��U�!��}��S�;��Lr��{s����$�,U�(����:�}LF�,��B����#j_�ty�|N/
G�P	��|�q��U/�!�R���^���>�5<�� yO�(\��a�2��럊mu �7�-3Y!9i��ő�,��I}�*��O�⮷�����O��fS�����
����$Z����,"��8U�!���S�����/�C��i����(q��iT@%��6��-�=,yi-�v�*�HZl�5\k��ӑ���UťUT����M;���gAlE�lv%��f���H����- �kD=�^l��ѹ�;l/A-�.�pW�����*F���uW=�D�^�P~C�!�b�u�"� >l��)��ǜ���߿Ɇ�#~�V�̦(l\{���JD�E�b58��JK�o�l�p{-� ��z	���l����N�ƽW������"쌇&f�9H��$~��c���F,<
�º�[W��|Sr��6#`�j_�{G�N�B��2�ֽ�a����!��'�(��1���VI�D ��)9����qE^����QC�*�̺t�y�珅��| �J����q��籍H�@����IY�dӎme�ʣ
�T�B���벵�`~~=5/�K�\g�:Y�GLYui�����A�<� �4TLL2��f�_�φ<�&Nj5���m+1�	��Z(�5�@V���}������t�G�*"�o�kf��k�W2�r�Y�G� `ƪ3N�8��?tJ��1�"W�tQG�u��m�l��z�9:�⢎�� ��j�'@��P	�N=i�K��VoG��8+ƌ��a���*�,TID�'n�����X�t2 ��v��[՗p�"������VT�m� K�e�w�����V���t|M�q�ԋ1�v�cD��1��L{4��V��{��]`ov�eF5��s������-k-o����*��N���T���?�k��.O��/q�gi��Q��BRG�@�j����T�]	f�G��O�nޜ��KX\�3ee�������7�@�P���[:�{WC~:,(#G} qNRq����\=fpگQ�W�m��Nh`����K�rϓ��B��:dE�D�o��^d����vTc=�Ɂ̠X�OmQ&�p1R����d��%��f��  m'Y���H�����l�׆�x�s��=tsNf���n&)�(�{e}����_�6\0���{��ro������Xy�ri��z����-s����zB�^Х�ﺹ?����7���5?���A%I�Yi�2l8��õ�˸'$M�d�k@2sed�Rc�5o[�q���%'�'r/�MK' �u�>����)�\
���B�����R���s�>��c�7N^�bA�-��8�Gh�UV�|f�����"B]�>����r�� `���u���SSb��E���⢈k��򷤳���h�s.���K�R����k�t���ĀZ�1ڡ�i���H8E#8�G����o����ۖ,�w�K��ԑgl|�5���+����ܤ\�I�zM��CJ��Ӳ6u�.�KS��	��xF�@���h�Q�#S�U��i���qɾ1<=���E���봽�u�U89�����5e�u�|���V������L_-<΍5�4R&r@���TK�"=F����H��b��[��/�ƉN���=��
�?]Bm�r������i��q�|��ۭ)�X��_%{�M���{�E��l��'J8T����PT»������(�t�xk��mC&�������NN�h�������ճ<j�\�2G�s+���UsK��LA�W��p͍�,�9�S/�0!(�Q �8�8B@�uq�%E����d��@�i�M��]1��-b�f��x3��NbMZ��{7�=��f�ʀ��췈�WN�~MSA�3�?��vzh=X��A`1�	�d�{��8�,䁆�*e�̆�+��HF�I��u��*�����W���3 Õ�Q�)t�IzP���OO�by�5�������?T7F/����>>9���b��bgU¶�Pbm��L�S;���b<�C��K�hR���o�O-5Q���B�#	V�/`�/E���ݓ}����ʜp�YO��n	�	E#�2�E4��E]�jli�exb+��9�y�!�"���JE�!f���Y�ya}�H�j� ����޾�b!����ﱅL�z_W�d��c�;hE{����D�z���N�u������9�(upԲ�0����?��:+Cw�}�01��5�Uǅ��]����y,Pp�t0/A�oQ".&$Һz��1���>^60 �n˻�� _C"ا��w@�g��O+�����f
~\$�,lM�X޽Q��f�@��Vl�e{���Vnc��K�����d�5E/�&P[F��a(FO��E:'|�ud�>���m�����1 �%�C������?ڨM�{��V��@����8k��Kg��@�@�ZK��.�_��7�ό�4�tL�N�����(^�3��1���y�µ�B��3��f�ɑu�1�$.�Һ
B�0� ��g�]�l'h1���N�P3:#�2�ݭ�<eɒ��$=�G=$�耪��(*����f�ΓJ�6C�qnFΜ�g�}0�22�A@7�6:�[T�:^2Z���m��*CƩ=� u���de�]��JX+�	����N:�%X�*���d��z���Օi��i�y��"tw�x���y�T:�vM#/��C��9��g8q4��Q���|X۽E�A�o�>��rڛ7��'1�U��@������v�/����= �o7��y�y�	�Q�)���2}��HN(�I_�.��X]m���]9 XjI#[�8W�v���1�ŭp�r���f����s}Yz�+�1I���s��`�v/��%���	_�8�@��;�h�P)�;��~M�3�r��( �����L$벖�C-��PkD�����)A�ӷ+UA� fI�֊�zX�P%	�8�KD�î8GP��w?E ���<}Ť"��9�P���v���$��6��#>�P̵�>��P'�e׍=o���
�쟜�� 0h;{W1��(u�#�b9��,P�o 1v<݀{��aĠ��U�
V䳺+�݈��@ϣ��$� 1��Ǘ�:���?5�*�>��<��G��X�����	i��"J�ф$٢*�F0��;��^���4E�$Adv]�T�=�7�������7�B9����%JrMH,�T+	م�f�`��sƺ��7 �n��ѫ���j+�x��r^ّ��<*�.�@;�Z�J%�D?��`�ӮJ��'�IB�-q�VV����Y*�a7$t͙cɢ����4�#(��[��:T
�����g����j;YdJ�.6����#M>�8�ö�*S�V6c}�������//{��N�<Y��a ��=Y����6C۲����Gw�(��29C"��a�x���,a���T��K��:����Z�m�����i9�>�P<	����pդ�fVY�^H�'MMc�{X\tG;(K0����j f	V%�x-���⫂�mu�~�üG8*�Yz3��t�cj_z�I?�qߤ���_'H�u����sPA$��)�: (�o���P�h�N;�{M�f���o
�Zuw���aY�"ъ�M8v��G.S�{��t���`L�-㦩���,�+�
��%�El��b����R��c&���U0��� �IG��\�/� �T
�4��u��f�.�f>�×��yH����c�w��!Scح�g�;H5x��r�����~�L�xÁ-�tq�A��C(��JL�>��\��vҨ�L7;���[k5�#�61�V�� �q@¤����o��q0�b7"o�����9�}������K����0�#3L�ScV����z'ܘ?�Η8�T@�b�Lēt�4�
���w��� �̲�'X׹7;$�`+F*����W�� ���hrl#��V�y�}������t�ʲ���B��_w]�����\M��J�ґ��HU*-��~�f�ω��y���.Bh҄S�l&}L`HdQ]q�p���!6{�q	eD�ZQ^Μ�Փ�i��]�	��	$+u��F�<�ި�C�4%�~�'#�ob������nL&�Z�nn�oKk��u�0.V�r�1!��s��!-VH��C��n[�(��B���2pnІ���1b��SL��6�+k�gi���dDr<>�j��=��$QL�9��� ���8+&��cI�NC�q#�n���Q�Nd��f,ڒ��*�bJ�g&ƾ]]z?*\�v�e �c
)�`��{3d
����V:|P膂O=�˿ؘʝO�ͦ�����#5��а���S�$nsw�`�k����~�m�w�	?��ܡm����$[��c��"{-0f���r�?$dk��O*_7�i���F�b~�?�b%�@)���*�T��m�pϴ���$c���t|o�fe)��ܴ��DD�RT��Ȳ4l�ʠ�&���1��E����
4�,�7(�4RkG��t�����_/O�`X��uW�E�Q�����qC��� 4��G��N���J3�%V���`�mX{+G����;Wƈa���J�07)oё_YcN�&c`�/����/-���7>=��
���9aTf��� M��я�!JZFul��0* �q �Gu�[ͳ�ċ��:�*$��ؙT-;�".u� P��3"v`UEd[e�
JӶMҽ������oiy�'ґ�e��E�*ԍ^�����=_Fs���Q缑M�<�����6�yq�	e�@Lhr�rj��@���G(����A����i�E	T19/;� 㟗�]��}
侜N�@���ܳ�qf0R�F�\����Eb��[� ��<f�w��W�M>�sJ:��c�������a�
�v�F������yJ�Ir.�D�!$�Z�2-�y,���k(�F�ʢ)F9�M�M猠Y��"�I�0O?��-�O�N�A6��pן��-RSS�G�@��G����?��,F����-����<#?�D�4^�П����)�ӌ>�s�Qd��Q2�7Ծ��P9O�f�:y+?/"�հ��y����������#D�!�bh~�|�L=)K�C��}�+)�Ήp���#@MP�$˺~�#b�y�����@�ZAV���[˿���q^�F��W���}"p+�������sE*l��6f��	�X��i�U!�¯�u{%��� 0����C�-)"A��(� �+��E�.�N���o~������PL1�=Rn��k�F��B��ݱj������r�����sG���}M�lӸ�����RL�I�/8d=�.j���fٹ���g������.Ӹ��(�������E�F�r{�k���ӈ"s� %%��8P ��k`�R�AiTh=�x�v��A��<��_�*]�t�����79y�+��8��B����w*vx��Ë�n�E���>� =f��3�u��_��ϥVf�sY~.iE�,�W���&�
TL��j���.~2�yҪ��AZU�t��!0��z���4��u�Uޭ����� ��.���v�z���c��G):�^�N/�k��Y'4���^��ebF�G_��9Yi�k�`�h�H[} �'�~�b�������Т`S�sʂ5��>$Y'�>g��NEڎ~��ws��U�I'Gp�[��?��0����]�hV��&�uyɜ�g�[
9F�Y�eݯ�����؎U��E�zc��S~.yl܌h�ee��E]��>�
�X5#ʃ�˱L%�1��
���Qq���*���]���D��u��
�0H�;[�g�a��~�цi�jW�Q����m�/+���z,���h܉t���2��N�������Y=�"�ݴ����n�0ή�
v��i�Έy�����.NmJj��I!�����	��|m9>�,���5#9X���n1cq���Q���ـ4�k�(t��d��9d�d��"�����ERZmEdqnc���%D�oǾ�܃s����6�E�咚��	����꒚ � �>M�(�����D'�k ��1�xg1$���A��gc��%�aס<�Q�]4�
^%�qN;����_n偿;�!?7��g�2�{�֙?l�f�Dk�#+iU���%���̝	�'�-"�(̏^*�Yt��{�b�&�Ÿ��¿�I�]?~j��< ��ͷ�ޜ!�:8�����<H�,�SF��> �k-�������?>�G2����`u(�W� �u�|�b4�jP���:�y�R�9�.B��ї����c��ad\:g2�B���LYVL���VX�(4ɇ�C��Ԇ�Ï���<��w����D���+WF������"�ЈM���f�!{/��}&Vʕ·�[ڵmB�bz?��ݶ��ӡ��0��6��d`j�1��I����jl9Q�A����,��폖/J�������������vCt��.t����¹4�N��)��XV�F��e�j~Kh�Ru`8mF���ѴI��u���T��*8���'���.d�~Y�m9����
�Z���Y��WQ�2�TE�v�GA�$��U��@�Y��G�Y�ؕ��ۊ��L��ޮ���I�of�)�����be�8/5v��}\O�9���&����!�A�B��=뙯�L���p�^<�f¸5�M��z�/�rR/犼(� ��R��L�7J��ZJiI��g$�?j��Po=nY�^���9H������X�[�, �^����a�;N�qK��_�2&��{x5�.��G[,�G��D�$���G��2��iX��(�ӱuwGb�;�:MD2?�����pS�Q0g�Ws( �I�V�Hm���u�x�/pf������.�J_�Q�-L]���U��ߚ��K�Xs�c��T��7�a���/Hv��\l��1�/M�cgǓ9uR#��e0����zQ��a}Je)�#Pf%-��WP��A@8 Q�_�*��Ի�n�W�HBQ��)��?Hћ�J/��ך��7�����v���;�����K����#B4���ruޒ��̎ۊ�6SR��'l#H��A˵;�+�q�=��ɰ��j'Ķ�+!,:�]��cq��7�` ��;�^�,	S�"0f0��_b�^Lz<����?6��g��u]���/��W>�ѝ�l���K���Z�+ˊD�3�LV��zj�BmP���B��q�+�>��º�Kzz}G(��T�1���ض�	��]Ʈ$��&7�8���6/���6
3��ز�����������W�%�V+���UFrߍD�럴dW!`H1ւ�C�B�������邭�RS��?�vy�J��G�eپ���lV�� ��*��!����&]���Y	) �eI���]����5A%6�����ҕ��iZn蘿
�����z�{1�񕘯^�D���(5���V+!�;�yBX��#�sh���+�D�4������j��}�3ܗ�%�x�wu�� }`U���Z�(QI�#y��K��>�1*�U�JR�n�
����g`���d-�?�$��y�4�z�A^T{=�U�<�،@�֋���97��!H�Cě�lti��u���lx��D<ؿ!M)(�&z&a(�~IYqA[]��hm&^M����������Z�cb^pBR\��e���
AZX{_S�G`i���CR�z� �7��ްÆb�)BB���9��p3n�$�+��m ��2�#�T=RJ1ѕ�!�y�R"Ǥ 5?���	�c<M����c���e��Qn��g�@+2)]�2���+�u>��jl\;z�7i��Vq$nQjȞ�> V̄�c���.�sS��_��˩t'�ȯ�+�������q���F�2ߌiH �����G���V��u��T�)��/
'�r}W����� 'K���;����{F_�1ɕ!k �)VUK���rb��qj3���t���ʧz��ޮ�J����ߤ����ކeD&����2�}�Zk�Z����δ����T4����"���ק�:j��
bT�]C�7W���E������A�ЮzcԶ�����63l����|�ύ�D�Vv�+�����)�����cA/8���8�(�6L%B�s2��-�7k�7�'<�$ܸ��(��6R[������:�Z�	+�ė�F�J���¼J׬{�\��&��
�\b�Ә%���kH�q���.�a�B:��Fg����&�ќt|��8�"�o�Ak�\�-}�I�����Ql�6ud ��RǑ��]�PC�c��/���/D�k/f֥��r���N��-+��*L:JJ(��b��Oj�<�	x�L;L����ʿ�l�AʃhZ�;.�bƽ�u�_��X<�]}�E��R�P�Iv/g�W%_�T�H���	��(�Q�ዐ���J���h�F��7�a��2�Z]쎟��M�ݶz���y+wG��ɞ2�H*)��H미z]4�o�� q����G[�#�A��ʓqǥ穑�/����E�G�a�U��P��J@��B�d� n����G��T���k�sG�]C(3�0f�c�T#�"����<���7\o�*[��;/�e<^�b�L5[�4�%���-��VLc�]Q8�LP���/Q�z�����Qw���Q�ʘ��u���82b�;.ґ�5l�}$�j3���t��}�֋���p�b�Q����˙ej�%��D� I�"?�8�JOJ]vB��d0��)����}��ߠ9�b��]:��8-�Ý��љ�B@��D+|�K�rkz98���,�r��[5�sp�B��  n$�.6���6<�l8I�52���cײ�[�&�^�+���Z�1�΂yN�FT��:����[B>��b�0oo|$���ṫ��wo6��0��Ď�,�%A��s��@�i�P{�A�H�&�H�]�c�rU�Լ���&=?�$b��j��"=<{6�D;�u�5�D~�����e �ߺ�P�0�U�wWr�ntI��\J�?P�$�<;�+����E�?P6?�v�p��h>أESK������V��[�ek�����~��S>X/X]��&R_\�G�F ո`\��t��'���K�k���C�P%&�S@ϕ��D�� 8�'�:
+�H/聇/(/BkE�(`��p���V���(|E;�%�VOg*ǲl��fO-�m?1���Vz���T̀�o��!��>�;q��N�{�%�$
�����+ :3cٰ�Q�^-�XK����9<���v����`�z \�:o��2����*˲pQ�Dc��z�l��%3o�#��!-����j=��纃�i$鱢�`���c{��ޖS�p:%���8K����i��*�Q�r<
qr}����o�G�>�/�?��o�[$�F��Z`������u�^�߷���ʔ!`�4X�$
九t;H��rl��Tm88PS4��aj�����~՝�[��	;��sey[����q�*ѳ=D�$i�o��L��K쁦��|� !���AAZ;J��i�StT�柃��釭��*{�3��g=+:=q?��������#R�ox�����i/$*P�1���|��x��.�;�5 ������|M���hv,�P��Õ����LWb����+�}����o/O:��Am��8�H��y��%⤣��,��.]�-��Xҳ���p
E��f�]��7a� �ps���cI��s)�5�|/��[�%��%>����J�l8@N��0���w6�C�
Z�]]��˼���'ūV 2���hB�$(���9]c�p�V��g�x��2I3���P�b�sn�:-`�P�K����U�Q"p�Nۜ���U�,�q>��5�+F�%vh�����U��`R�x�ׁU!{�ƨ
ߍ'�CQ��+ U6R�sQ7�~O�~z��*��\0�	LO���=k"�X_�*���R��v�?��w�4'N����.Qx,tn��C���X�������K3159��g�	7��jb�_�=�*,9$�pvDM\�.��X���R��Z��^��f�b����ѯY:�7`�ں԰+@5W����A�yU�nڄ�AB��� X��v�#��[��%̥�^�'R�َ,�]i2����l��+r
�M�*�Q+69��mO��|���*�e��u�Vo��*Q?�;ҧ��Yٗ�.=��s__;�JE��K��YBq4�S7�7߅Dk�]�/����csݥ�}W������n������U+�!�#HwQXqY3��"���I?)	;�p��H0y���.!�E��v\������<:F1���_�����Z�b �V.��Կ��g��F��3���p=	Bk���h�%o^-<v#�h�l�U�Wb���f�qM����ꏞ�V�[���N�����d�wR�oM䃃9�a��V�w �b������.�QgX��L�d.��æ`�PмM���t)��[e�a(��?!~��j
\,:�dZ�Q����1n;s�b ��P�]>~�dfYW���Por����?�(��'�?7>�/��m�B���d��
�c�/|?W]U��g��?.��Ħ����ebΒ%�Kk?"5�T/��a�&Ή|��)�s�*�Q����%�ɴ/��
>�����no
:����OM:�����,P@C��<��Y��;�+���{�k_�����i�&��8�׊���Dv[�����	��y��Ȍ�FK\�Dta��Rt���"�AP��2$%ɸ > �ۂ�%��\(�} V�]�}�ր�_ӂ�����S�.�����o���p��W���\�g 9�<:lhjn�Ț|����h����$�#��u�=�C5����uǦE�>�qX�:��lcN�ԝ�g�l��t��P�Mљ��R�Ҡe�*v��b�K�GR׃��<B�tiw��qJ��Z�x��S,��K�*7M�n��n�_.@k�=c�+�	i7����+� ^O|���s.7��>Jܻ)FR'@�1ۚ�"v�괡�GI�v�NҠ�R����l#x�I���!��8�U�EC�e��E>���~`���1�L��~��S�Us֭�~�v�����DM �_̈�
����D̂��6���;/t��rf.H�	gM��{D{�*R�??�m��;�����[D��W;��Tz�����3/���,U/�ѱ�������ό�}��70_��kr���1Q0�a�˚��S���E��m��	�0���M�/��h�䞤��o�{�V)yt%���kI����� �p/9��$�͸v��I�������@��'t���`Oa;2>��<\�A���)��l�9҂�Î.�ì�v�a^��V0��[l���h)��!i}��A^������X^wKp����[TG�m^��#�����a��Y���;�æT���������/؞+��2���~�.�;fM��=�V� הJ�m��)� �Ksr��p��5H&#���'k���P,����YE�{g�~�ڰ����j�{=�Q�T�p�|-ܑ���ϝ�OXd�M�~ܘk*4� a���٦�m���k��~0k#�G��;�%��AN����a��
��2�ln?M6_��U^}$���#P�:>[Qk����vRC�u���_�޾nw�j4�6�
d<=�;<��73��cy�p�V��Ǉ���/C(��df�ni���aW�g�w0����W��.���W������m�'���]-�`>g�y3<�O�D�n��U2h�T^~�rCXzl�ݚs7�����Ct��x�%eJ+�%O%�WmKa��Ī"fs�A�_�����y���9��R}�k"�TƐ���Au޿)��跻_��񡦾<�<�0�n�'�w�ֵ���:�a��ж�~U:w�.V'o_F!<�������'ʉ{�ȫ���C^s�+ s�\�� {�X�i�b!��9��?p��"���i_	G@�Qc�[���7~}2���(~}\�߀rm��t��e�w���􊅂��-�e0ݾŜ8�6Zn)!��U�e~A��_ڌ����Q7f�󹛠w���.
?��9�i,8|-*
܉����c0����Oʭ��v���ݏQ��O�8�y�?�Ϙ�UwS�D���J��4�����UYlˈ������z�D���G��s�qi��#��5�������
@�T5iGB1��z/%�,���*��[5��8v��fV���W��ª��0Z����t�d��"�PE��02����'KB��K�V��Li�#[��g+bf3*B�o��ƙ�V\��k�Z��7�ݧ�?Iċ`��tm��n�F��=�6,�Lv��{�Z��"�Z_�����˪�:�6����|$x���@D�V>���`�0��S�oK�n�L�� �9�S�GH�n �W��؇6'I�j�b#�)rծw�;�!��c�ݞ��y����
5�q�L?M�>_�H��l�z����	~�)uFi�T���8��!�jG������`��ԗ�����/}a������aǎ�u�a�PE��d@����ޯ�9{ۺ{9>O��`	���ZN���4����R&t�f�H��3�#�"
��*ۭG��P���m�6��%cQV��Λ<A��T$�-)�(��t��(�d��NF-�%S;Ӣ�d����.��l�/�U�=�/XA���@�j�����q��;o���鄒\0]�	⓽`0WQSP�tͿ��#��%�������'YW�L��V��q�P�-��!7�H%���C�ʢc]NK���_�w��ب,���oA���>(ܤ����#�{��Z��l����M�By�7��|~�v�v�~���ȡT���Pl�O�o���F�a�w[��{>.��e���U0`��=+��tmq�)��#-��(�,:�N��Ԅ�q)��jD����Z�xo�����M^�tD̖�m� 9}<��Ҭ�����8A	2�T�]��)��Z�W<���;X�6QP@���8Ӛ��R.M�M����T�e�j�}���dO�
Tt�Ua�@���B��� +���_�����ٮ���EOߢ���+~����tƓ�)�F�z&<�"�È5�GkĐ���h��n��� (�E@��5t"Θ��}Yl����s8s�Ԉ��i6�N���Ɵ��sX��qI�7�GX�I��5�Ҕ�NJ0�y&˨�t�5[]����s�f���Z�5�S/��LS�T�9.�KHA�K1�1=�]��@�^���_@�F�g�7o��_�����0�jRJ5?ȁ�n4��}�P��p�)>V��$��|������,�V0G� P_Ls�n�;���P��*'#ݘ���nm7O)I��0�>� K4p�I�Ёk^��˭Z���Ũ\����Q�C�����.9 $F��#�I�����!xP5j��Q�Y���E�t!/CӇ�O�$���6��׾���W�˰I�#Wy�3� W�d+��&*k)��1Mf�J��1\"���]���*6>��O�2�jTu2���@�s�ʬ�c�Mư�WyjCMT�� K ��^��c�����T'��}o��}8Gq2�ZS��d�e���}�͡"ހ�ߝ�}+�w�OJuG���س�3Z�)q_(�ӘƯc	��]�>��^��ش�9�^��\�"A��|��Y
 ���ܱG�C^&�rږ�-]�;JQSM��!R�{m�8^� �xgc��:`��9��B��?|di�s^Yjzy�R� �	�?��0�]�+�{P�� ��9�.4���zB�>p�����*a�ҹ<�60��h�dH1kt���S���P�� '��KpI��t�~&bh���H���u����'��Mt��ix�a��SWH ���j؞��&>�.g�:�#����F�����G�����q���=�)����b��k��y�V)y1�=�+�ʭ/p#��M�b���p����E+�=� Y/����6�{�q{��eve��Q��-��6���m3�����R�l)�\�=��0����,ф�ɳH�� ��Чt:R����^��"�
����22~����B�=>q��A>���nee�b ���6Xm�~.�x2G��ݱ+��p��vw,���_�<�G�0���ց������_�[|<~-��{�?w-eY��hk�W0�I���!�O������QN�����֦�W~FI��&�r�6m(z`Ut�9њ��h ��7�ˡG�vo ���L|��k��26��z��C���բt����RPӬb=����c(\MFA�Q�g�s�v瀳nB����
nƶ�.�PgC`~H[��$���}�lr��a���f��QM�d&-������J LRW �$}���A�U��t��-� �m�X�u�$.�b(���?1a�W��T�1��mM&S�����j���:Ǹ5]�5�N� .��2�i�w����!� �؟㵎!�y��[�0������c���'��Y���'���}����%MB`!a[�`8���`*bo��>\Oqœ�č0��O?�Òյf��u���(`�g'�:U�&�n��'���7����p:����R��WB��o�I�|@��~8V��IO+C�NBnBǿ���}���r���zc�I��V{0	8j�(�J�����F��5kc��l
�ԣ)���Cӯ+z����m�Pgw㻆�S	=)_��[v��ξ���8��RH0�� k.=��%����D�u�	P�7mD��M��o+���bbV�4��iK�[�� ��VǮ�	�+���N(D1�W�
Y�6^�r��_W�9Y�v��)a(�;�B.F �2m�ؒ�� ��I$xu/Za/}�;�0v���Լ���),�Ĩ�����+�{q����>gj/$�R��I&W �3~�
F���S�{EZS|�>ژc�H�'ګ��5�����?�ɆT���3�}<�K<'{��o�D�d�� h�`E��!�D�LiS��4�Fr�IEc���2�4W��y��A9� �?��n��Z�u�wg��ֺ)GV���'�X�y�ڢ��L��
F��%��1A�u0X9��'�b{B�s�J�Pʚ.��I)m\�6��Xd[���P���q����D�Δ]x:]��^�&Gs���x��C�P�Y���4=�2sh[-"���CA+k��)�+U���R��2�.`�uCN �t<�w2*04(�ӡ�-��1��"L�R����J�Җ"����v��x��?@�,��.��jD�Ȥ�7���_����x_+Қo#G;��+>-�uj�g�T���况�m'
^.�6cӺ�)3/�rIo/)fa]��ZZ��0<��gQ6�w���w���	>�F�r|�G��a\<K=E�}[�{;����QK%�-A}9a�g����Sۥlqf���@]�B[����R-�F(4��ު:,G3��E��ZQUU�i�?��Ws�֮���D��OF�-ľB����ς�S"��^�B�.Kr�C�#(���}���w�1�*���!�!�5�M�N� ���k+G�7��%ܮ�����uHT�w�T)_� �n�m��@�[c~;�H�yJ�:�x㫈	IH�~d�k��D���p��H��B�:zX��gbw����c�<�����#m@i�����ߗ��w�@��On7���۔��NDn �$V{9���V;L�a�g�N �`��F4��5�������C��n�F�Ϸ�-'ƛ����m��9��'/"5v��	��"�A)�Lę�W�t������ErU�˔H�N����_���-�]��K��р�G��M�ć�����c��v�������I'�o��M�2�8�c 7���8+;DE�y��ꇯ��Q��Kki�%p�+y٩����Y�J}E����6�N����x3L�b@���8�H�I���$�Mџ�Z��g}���Z,���ˋ���ewx®�����$���6�{����/�j�����Qr�k��{�L�X�X�g��"Ccod;qO�ez��*?�#�X�g����Guh8=�[Uµ,�X�]�76簷��;ʐ��*l^O�S�3?�5�'1_X��Q�^�[7쏣@�;�3'¾%�/��?���r#j 6˱��8eU��@�)Wz�hW_v�"O����c�eWC5�rˢ(�G(��1v:�3�u�޵�J�ߝ	[�[��&Mƥ� i� �E�)���x�����1M:��=¢��r����#"?�A.`B;e��q��>��� �w�`�]}E"*�7�*	Ģ!���=�N@:঍�M	2y-��"�n!I3�Ar[�c��Ȓ��XNkI�@^@6@�5���QSj$�s�	!_�t����:/���έK>�R�2���+����qy"s�
���?����Y�L*�B�`��_Ř�}1b�É\�h�rx|o��3/6�YE�&ny�J��oD�2`�����Z��(��,fX_A]-�tr��8_�D�l���w+۝��9��d�}A��� f<`���[5~��S�g���	�ЄԤHR�^�3��:�4�Y"���2�i{i����{M����i t�akp��*�t^�0B!��յm᳄�U\q���A(��������N��S���e�w#����l�:%��8�-''�E���ҝok��:{��|/RW��������{F?�	�	qi].�|��OZڍ��ز��Ü����]��
�Ł�^B����玧�n�-T�͑��!c����Sܶ�,�ʦ� �ʙ�M���*�p�8Dwl�k/nA�Η�%�ih��μ%����)�ʬX�U�¶��4�bpEJm���^�p���cE��l/�WӤ4����/�g5	)�Y���ing0�LP��Z9��:b����Da�~�in� ����rD޺Pg�H�-�����L��	�dw�����醦��@&x;jo�
h������^�	���xӭ���z]�Y�t��y*�8`��t�!/[%�@�/�@�����H��ȹ�r@mE�r���%dս������A�ɹ��3�idF�P�p����g[7,�]� �͌ޮ{�_qwE~#��hw���W^�D�Fz��(��ܣ0"��Ib�f����qJs ������F�zzeZ{�OxD�ݶ�H�	��mEuak��v��L���9v�2��u�J)�?An��S �n-ϔ�z_9�{���T�� �k��p��e��[�Te�_hM����]�cJ��k�S�r�����v���`�s������O>�#�$�lZ�	�
�@�����!T*wb�`6��A�Y�ؔ*��&p(��C�!i?��$��|_?��0�Pz���;0h�Y���n���Г��wY�)VZ�?�Oو<Ď�G�
���}xM>J� x2�.�~��M1����S
BM�h�������g�w�:����(�SY�]bH�\o���w w�Ds�"��^�ڒ���vQj���s�����E����3����jp�d$ ]]b=0>c�S�C���m�9b?r�qlf�����'R&��c!�	^8�{��s��P��gX�^lgn�K�[�����S[��J���?po7%@��?b}�~=3��g["�Z�~�g�AhD����Y��-ݦ�<�P<3{���"aY�@U�+;�����W�*�7������E�ǥܣ���}���8��}����O</��d����Iy�(�&c���j��,ȱH3�=�ޚ����kX֑�!���^/��sl��1��ɫ���B�k����[s ˏK*��.@�X_x���l�NSR�I ���pn5���N1����1�JH�uIʾJ2 B��	��)6ރ�rE(L���GVgeZ��I��:�"'z�0-^������~��Rp�S�Ka��<�Zre���4��njis���X�^E��=��f5���	�����^��1�e��{��3��� :�-c���݅n}-�{cV�zth3����,￝y�� -�D+�����p��^�`<1�ƌ��VC�9������ (��#�d�_դ���b{̭7 !�5�^ݼ���Z�h���=��8w�`WJ���Y�lѐ�ZJ���V�Q
�x�������3�P�׸��5h����һ�ve7�u��d�[x(M6�:�"���
��xŴk�-���EE��{jA�p��V˞��w@�w�z�Nۨ���8����D�3!�N0n̚ ���*�sc���� �wO����ލ}���}���zn�7|okS�)zC�͢ݞ��t�-
F�׿;QG�HO�RB%w������8l$���̢��� 1{�9�W�	�[��
C7z�!��6�v��Z�ұGQE������`�Ȇ�F�I�BJ�;�I��M ��j��\S�-:������@u������a_��h\/��fvv��q�B���`i�eL�Vޣu�s��
�P^��gy���F*�z�yOj�J�i�v��$�c��?ʌ�V��O���_��X:�k����d@7d����R(H�8��څ��d/�%�YeĬT��a:�Rjh�&6������2�է�[��v��������ۥǉ��:˻̓���>���{C1����:�vV�������<)���=�TjR��+������gb�
b�����.��Z��5�H�}��mq"v�$��LBXG~��oԍ^���t#�(�Ӿ��eо��S���ģ��j�|0d�!�P���m��vHsQ���.2T#O��M���V2�
�c��t��e�:�y88�,�������>*� u'�m:��'O��u%7٠�+�OnN5KT��'�4���h,���?�G� TX��8�r���q��+�1~�<���^M���<xl(%D�*�lt:�܃JD#f8>�:��g̰�i��'k�㞖��c�İBs�(���kZ���$���'
�j� ��$���R��}L$_`6�yr�O�A���ͧ��uC��n%BTe*t4�p%3����K�7IF>=�����#��Tjo{�tLf��A����$Q�5'�'�O}�M��rP��|��L�ԅ��y�}�u���e�E$A�f����#7"��y&��k+!,�X��h�`�<O�����Չ!)��/:����(^ơD���rc�H[��HE}�"�����Q2V9�M���<�j�*��mZ�q��԰!�,Fۖ{�y�k�y��LsLu��f�t'���Y�\����7QZF�N(���T��ȕ?P���ԉB�����8�}��?�Q�V�@([�\�������Z��'�k(la�H�ٲ�g���Q���Oj�RK�Zmw4�B��4�S)�te�Ǭ��(@�B���01�������H ZY��냛��-���(��.D�ډ+N�F'���9:��|]��G6�u�1��zwY��F�h�fC�:�����ʾ��+��E�L��S���>�Y��&���17ߔSn�	�{�*�����������Z{�����g�l<Y	���	�d�q䝙�M;�����>^.~ß��+���O���¤��@�ݚ�7���6Q��V%��=B�*�NS���	�O,� �@bO��yi�[[U /m.<1�qP�p�z�3H�<pSD`<OWa7���[�Gk8��,2�K|����'Ð5��J��;�}�Bۄ�w�Ӳ1�6�L����Q5LQ	&!�:S��GY:���=�v�����r
�}TBm�||LD'�~z��`�N�*���Fʝ��B/���s�ͶX��
��p�Xe�΁��H����ij��Y!�i�&�u	��w�8�_ey�.Rڞ1�S�;����������~Z0s0\��� Ñ9n�c[�}��2� ���s�{���_��/���Y�b�a2#��<<f��^�8�3k?YG���v�d��:����I'�݌x`�
�ɤ'aOO��p�t�[��.�RXܱ>�{��itZ*��Xz�\^L��)��c�&�©�8�s�+y=��@����[�f��F��*7i�(�/&M�Ĺ2�Lq�}��U�\Ky�=�R|��@jr�F��ʩկ9�o��ލźA1x~�-�<y�?�aN�F�(){�.�K�%A��/��	Զ�*�l쁞����n���_Q�ɂ~�z�������&�g:��O@��$�W���o�d��G�Z^�[�	E�9�ChTV�P°b�q�A�8���*/��Hɱ7Rp���Hx����p��PR��:n�� qeH4VMђ�8]S8��Y���L��[/{P�h�£�~�v�
e��#7I�nx�J=�<F��Y��A�Z6�J���@L՚F�5�{��x �����!�O7&�[����A��~OV����Kp����Pm2��ޛ�R&4S�u� �:kY�� �ݚ�!8���N9���@s�-�����Ζݩ0��T��(t�=�<�����ߧ�9�Ng�����z~���#����}"�/8k'�4�M���E�p����Kٵ��/Z�8�I\�0�e��F�!�Q�|�	9 [�)�l:�=>c���s����uқy���k��H5��Z4��HL`�Q���7cl�S���?��"��,����免؆����-��).hmB���Y�r?�]��h�?�+�P�B�Zc���uN���ȓaL)��w�|Z�����!Z�ĸ%웝e��������������OG*�I3͂��Η�x������Nٓ&"�b���vcDG��F1�����U*b�0�a68u32ف�_�*{�N����jaE��h����z�5��ar/�N����}z`���}5�:T�1	h���x��m5� ��;F�A�)��m�+��9z�<�/q��p3�%�4O6����^�����}t7�i���r)ǂ���IqN��	��S��.R}>�)\�At̾Ve��(N&b臩F�'�Cl?�>�]�C�oU@��»�!A���.A癯,s���z�[�;�Ax:w��T�tMm׃�����$����Ք��}�<)@��H!��ߏ�͝昲�3�ׁ=���ϕ!U`�*<D�C��2íI�Cfo5�x�%���N�撃��F�+�I�����:	��OU�WB�������\� -,5&-Ll4ll��Z�B� '�����o�H{�fģu�߀��]�?u���`�<RҜ'�:���'K��&��M�����kqe����+�8��IL��8r�����*|����ߴiؙ>jE�
z]+JA����Ah?���j{�u�Vv��v �?�&΋�"b<��*���J��R$��#Nkv!���?�&f���ؙ-� �ג�`����b���%J�'=�bBB�Am�
��+�!�)�,�5��H�S���Q��$�1)�O֜ �FJ�(�{��_�CeS&����PT�����kw<�Q�|Q2~�7%>���9��-#�=Qy�	�s[u8������oc>
��S���� ^�RT��D�<�E�v���5g��I f��ٖ��ҼЭpw�Y����'����N��_��(=���$�z.�c�i)FD�E@���];���Y���Y�%)�Y�ʍv{�Y�,oE����>K��i����=��!�9^:�Ƙ���;p�v9�;Rey�E�|P�>��$.9��^	��Ȧ��U�н�3�_$ݴ�8TbZ���%��ͯ�:aAA?KffOj���2!�G]%�u���*]X�*PoP��B�p:� �s��ŏF�qrK5�m�j�������ɄЭr��v��(�6��!Ȏ��4��jf��Pe���ĔSe�������h�O�K� ���n��S��3���1�Q�Mc��R�(}�|��v�/H� 	P(_����$�&��j��H(�7!��羟��l�{N
�M��sM�.F��GB�2�ԇj�긦�i��c�լ�+�"/��<_`���~��%tn�Vk���ɷ�EffY�g��<: #�c��Xr���h���;�v���y��?I?Q�+	t����T2k��K���yC!T��l�`��o������MkvP����zJ�5H*^C<��P���X��w>kg�2i,��)�.�DZ=�v���^�&u�@~g�L:�oJ�A���$��`[ω�GO�Nw�|�9��h��`�X�K�I,�D#'S�ч��������άbc.���(��WU�Q�ف��;`�rb��MͲ7�U)����Hz��H|���r�!�"��D�(C_%�PV�b�7kd정�^a� ���Tm;�i5>�qV�d(r`=C,+ӷ�y���e,[7	А�]L�!WXjdL�����!%�jh��q�g�09�ng���2������� op��=��~�R>�B5v�:xS�ގ�@�='X,��0�p�wC�^��a&�^�;��]ؚK�0�6���4�ʛ���`���'�o��F �eB�w�U��qA,z���oΪ*{T�@Y���3�,�|_k�t/kUR.̀ˡ���Y4��gA�P�:��H��Vn`����mf���!r%[�C����:Ӧ{I-#�	��>!z�bn��K��rA��R����:�.��n���gWS��(E���DC'+�.�A0�ת�Q8$�#r�LF>�� X��j���Q�I�⺘�ւ;Gf4z�� _����E"�!�a^�sE.% ��[�����W;�k
��|��q��Pa�@�Ќ{�&a�Z,���I��<��M�d�bl�;,'F1�Wl����o�qˬ��n6p�����)��~�w4-=�k꯱�\��q�G���tɤm����E����q0�C�3`4���~㌥��c�jpx3� �w���>�,@D�:�bΙǖ����'�U
y�Eŏk��p,_ɑ�p��������B�ņm<r=��iR�@b7�o^��6K�:�4c���ڒ��g�ع�	)7hp��%��sDW61v��`C����ZX���kw(-����_��*G�����k	�/H�U-^�	�6�J���NƏ��"��NqU� 1g1��v��&r�RѧuA�U�Z5�4��Д6��˽Oh,�/��_���la�'*��MB��Ҧ�I�	QE��P4a��U��p ��������<˻W���ޅ��c>�A.j6�2�y�6��Z0ޙ� ����ң ���u���H��ƿ��ͻF�'�, ��sn7/Q�ѱ,I3ud���1��x&3�,R�ߪ�c�ܙ `{��:nUȒE��kU��2pl>�^�U��L.�O&d��Ʃ�Q�	�q�3Ǭz(��b�Bt�����0
�])*��ix�����&a��k��H#�f2�գ���!٪"�ˆ�`���A#;rz:��&� M����;[�)�|E�ы�· p��pmy��yK��u\�
�}�hH��D�G������ �"�8R�r6>ً�懖�B�+�O"-xk�@�V��Ѩ��²�B!�� �1SV4�}F���X_�^�[�:��@�'t�V�!�U��;�>��eX�w�!�!\�v�%����=!Y���l�����V^|rf5����"��ii��Y=���O�52��YcǄ �+��L������(�ͷ������������$���h�v�ˍ���U��S'a�󨖡�)0"���	�r�ί'��j�.�o��Y��~<WQK�#i$��9(����@�Ό����Qy�� F��;�vP���t!Զ��T�3��m~�x�^��8��Ģ��ĝ�_���T�Ó!S�J�:�H}\�oO�`�p��]�H��W� ��,���0�.��uy!P5'���_�gΌP�*��l����-
����Q����J�G�A �;��Uw�=ٛ�ڭ�1����"��d���
{~�Au˩$�iju�	u�R��v����W�'�����&���/�t���-���|�3�3dW��B��P_}�a�]�|z��*&�)Ji��1X�K+�����1��*�׎��<<Eq��W2KO������S	�:��v9C�yb�mf=�]��� �V4�b��k��}��
0���~N� _"��8,p�@$j�y��6��Q�&T⺏�-�A��n�ߐ��dTF��b���	ʕYZ��%����3+���cHG�(�<�;�?��P�;-�V�6��c��=6L ���>�[
@���a`��'�NF����n�9�rJim^����������"���T�]W�u�=�M"u��{h�;�p�v�����l-���aߐ�;s� ��g�6��Cw=+�P;��7B%�8�|(��H�#�6
mlh0���~r���= �L1]=�0��J�I �+Pv ���.�;�Q�����?�m���0DY����Ȧؖ����Gw�uQ���|t���|���M3�;L�t�	����|���"Q�����p$�44c��;k���ML`��*�)���`#=�J�`ѳB�Ul�����e�~���m;�C:����Bc��=��D!ܱ������K���]�������ٝ�$�_@Oo@�G���U�uS�k��:7����Ƃ����5��K�j�$�&z���H9VR���(=��W�Js\�� p�3eMp����]�*�5%��>��3�J�Q��<wKX>��q	���V1���ɤ������#|�;���] ��W��7f�ߛw�Y��!t�P�{V�S��s��+����U�!����]e�P>;��-�S�� ����vg:B҄!��2�WUj�  5O�?8뻏�=Ǔ�uس��R�}�*Q%1,���'��TZ6o�A�T���~�������y��5��ΦT~f���R��Ź�̽/JO0C��7m��f2T��{�k���P��V������F��\��F
*�ykg�2��],#�������vR3Ж��4}�e��I��kmN������l�3�	�%�6W�����h�Xs�I��J��kʓ�,7���h�O�@y����V饅Ps�A�5�T�)�YC�U�=59�D�=&题�"_�~ ����O�K�	����7cg��I��R]�W�~�ش}��tq،�N�愖�ӯ\��"��yQ��V/�C[�)i�qq�(�n��=eı7Qɑ����쿊k�(�XC!�/���\S-D]_�H�G0�u~ӗhh|�N�n�9e@�"��9rm�T懠�,����Y��a���������D�iym��V �Kj�_�e]��E�(`��I�2�/�����A���F4��
~�l+t;	�^e�~{\;r&���|B�o�*�M�!����_����T辞R?�ZHWN7ݙ#�D���֫���T��vD"����7K�S����b��͝�����b'1�D (K>?��
ܮ�e����`&��;�d�SA~ͪS�3���x4lm~�{Q.�V�n	<aŋ��i�,�!���/�Pa\�q���z����C7f���s$��tLM�g�l�}�ll�L1s�/�`�6�t'x)�����Wdtq�q�a~�U���<)ᶥ]�}&�bJs$�F�8s��'-T�=�D��l8ƒn��C7���ݢ䗮��Ql����!�]�%+�&���H�Nn�V)\d�(�R/��9��(�z��������|�������T��������)�.��5����SU��z_n�J�1��q9�{�sQ��޸�Ղ���ic�.�vx��Œ�̼��\�/�WId�~i"��r�z��{�!e������TD�en�ea�{�.�D�|ߋM�h���y�at��!u�d�������f��S��S�h�@���>���H+�<�Ƌ��vC�&�TH��5����z{�?�E}�Q���%P�Bǚ��]K��0�w��]�5��A�(zW�^�������&ҳ��*�W�ԞpMJ��D�75"�5�4a7>����I��gI�s ��O�NA7x�"��.��|��B]w�
�#�G깆��~T��Q,��m͚����ئ��W����r��>�n�� b�Il*�0c?j`ڃd�vCTދ�9Q�VPٗt΂�{��Kι��"��%Q=�cOp
��a�	��~��Us�H�����h�8k:���B���)-�z������E{/$�H��,HO��"�v��d�-�J1#�T���;s�n���g�,���Y��,l��q�c�t�mM�䰻0D��G$M8�f���UE��ؕ^��@��N��
�V_�)��K3柬��/ǗCDox��S�����1�޺�HDi�����Ζڨ0@w"�r�`?;';�^P<�7s��(��I�%f�C?%�N;25̂i�B3�44>	<Bc�O��FL�� -�)n�M�� �I�.����������5"�]��p��3X�-(��<V�����:옓P�귞��/l���ټ,S���,�	k�$(6{�f�*.��g�G��p�i�dG����"iCr�ȸvlP�����q�qP���ڎ�WT���T5kbX���6�W�s#� �;)d�;a���l�[{����Gg�-���`oݽ��u�������7��Wx\?�&�\@J՘_�r?���R"�,�G�-����K�O�57�Y��z$WC�b�z�v�3��,����=������Fp��HCIK�8��E�0��F#���J@Ӭ��V�FY�Z� ���f���e�w����[+���]����ֺ{	J��}��6/G�~��9���w��A�|���wpR��Uv�癥f��܊u�2\r�Q r9�%��P�s��q�XJ,L���G��Hm:��"��. 	3�F� 3��r���v�khI��r��V��Ԋ'జ����Fo{Q1��!c�`�g�I�;Yd�O�&����Q�5lD��m��no�!�?$��É���xZ��?TVa��&˿M�[��R���#5g�3qyN���1������;�k�<�*�]���lƖΖ�S��Q`
�f���I��"Q^nΈ��%�g�e������P�Z��e��E�#d�L��4��ĢA
�^��yC=ghG��(��CQC���-�6kY���/o,�� :��&>8�G�e�#7V'��m�~�p2P���]>&�������B�|�/�|���x4���x�r:�/��k��"F�m��d.P�*x�@	$I&��E�Լs]m�ߓ�XϤ�"�R��������iV�>٫�C|����B-d�A�~*��c�[e��Vg�%t�þf}��V�i@Ǧ��K�q���M�k�m�c�9���L$�l���F�JF�1-�I��,dFs�/p��^X/�PA�^;6h��"�	d�˚����z�G�N5}~3%�{��'�C\�F8��y�E����8�wZ!Ӭ�j-yIGU�2.��YG#�E�b]օ�ؤ¦q���`�#���>׽�s�i�uw�&Td,��t?S��"l���(V�����f�Ҍ�9u�2~1{�����F�"�"��y�|/B���nl�n�!<�nnwm����|Q�$�7AD���ilt�m�Fj8=�Zˍ����^=��oc���n���*2�y �P��o�Ĝ���-���3�L�h�?���h�^K ��+@�?����3�b��
/;��O.7�y81��Ȯ�����/�����P|�ۅaSS�sU���D�:�E�U�J�jt�+AT�y�c�8�Ɇcx��ç�n��/�c~{�ǈ����P�¨����n�ڸbrLw*$�c�n�6 ��Z<� ���7<��|����*���(r��f�V���% ��e��P3!�:TQE.�pou�b�E��`������\rx���)Y��Xԫň�]��c]�<?����5/zn/��������R9vy�}\gg���Q)QՉ�kՈ*�ׁ�K5�[Ck�;%N�FLv5�	�����>M���_��i�α�:��m��R�d��(���gn���$
��D��b������kKsc5�D��X���p%�$�9�

�s���h��˴��$������>��<����L�b�,�­Q��K����?mK^����%��M%�"��4=
�4�>�]s�wP;9��R,.Ӯ�}.�z���<&j
c�s���I�dz|/ܼ=�(h{*��ۈS՞g�����`���l<��Hoc�� (5V'��)7���~�]g��ʘ���a�P�z3z�ﲚ��<RZ	B�D��wNR���߳~HYj���Γp�/\�����~�9��ґ�i���^{�Z�i}7���>#��t,!�f�p���k��I���Ӟ��+��p#��J��Oe\WD�R`��)���MZV��s�An��^�]D�r�ŋ�;	��Į3ݱ;�7z�c�5���WF@%�M�p;?��wv)����@��2/LZ�)eG�!�2�ӟsr_�����T���� <D\��	>�9?�-m�0����,��{N��:�	�y�k)p�F ���^^#���A9�YH�a5���˨y��5.��F��Tu�X�G��4���]y��#r~�MB��3�;����b�qkf,y[���R�X2d���W�L�/w��m]Z�Js4�����9��`�ƞ&���sT��U����`���++�VK��Ȭ�e�����n3�s�F��I���ƊM��$F�8�G�����F]���K����j��jZ}t�iv`�vfp��[��<�1:T)?��J)w��p`-��8XAZ��a��n,5�a�ˮ��!��5���j��7���z�\y'�Բ��/��� 0�-�c8NrN^��D@-�)d�������+Z��S�i��3m�7`w�j��>�E����2��ݞN1aO�86&"ƥ���J��?���5׾�Ky)���W~u�m��B�����?0�Nf悄���D&��\B	����7�y�C��i�%��?l�R��C�VdT4(9Eƾu,n�E���T�� ���ocПJC�+d:1={�ɵ�W?��~Vn���<��[�Y����9�%���Q�wXm:�D��4f Ӯ�Ə��0����3�;��N��
?W�]����G�z�bJ��Hoާ�툃�-|q�p%$�ZB.��GoV���Q���L~4EG!��*)p��W��&�� `�]�� :7Ϭ�^��b���Vү>E����S �qz�J�r�up���Ǩ{�oP�Z4̹�1�������� �\�7b�6�ߊ{v�?�:��{+0�L��!�c(P�yz�+VK��dn���٩����G�r�.�)l6�G3�~�ڻ�G~�v�(M)/:��$՝�9��'U�L ��}I�%�2��g�3�{F���}�{�{�����W��UB ?�s9�<���F5�U�n�eݝ"��h-�B6��}(Z9�[�z>	�����N/�O��;�ؐ�@�ۈƩ���u@Tv��M��iַ!0S|�b��Lҧ��d����.oob��7Ĩ��+o����Ss(�(���/�_fX\DN�����{�����s;y�Km`>�9�B;5�&E��p}8�_��9�&�`��T�=A����y���s�e��)9�9�J��/m]z��>�������B�o5V�Q��7p��K�Ԕ%l:�^���I��)4Z�ȃ!���X(��?W���{��eZX�L����#�E�	|�nƓ�9���Xːct^��c�p�? ':�a'���ôCL�-"j?8}\�-�2��R6����f�R/!��"j��x�$Z�;�L�#+&H�m�ē^vw�pR��.��>I@ݾ���J���Wm)m�Ð$a��	��WA��������(i���l���>��_�j�������(w�7��)D�~��F%����w�kmwR����#Io#��X�\ n��Sc����(�=0���B�{8<�,��hijr�S`��W.��E3������]�H�u�H��_x�,�-��;e����XH��J���M0�d�^�4;��LN���m����?i>w�}1�c��:�#o���'9�URG���������D��bn���-�4xM�I�W�B�O~;���Se]�n��4��u������_MaՔ�м1��&�2��@�q�P�U{;�(�๶�؀el�Gs�(���"������䍫�+g�1-	���������!��{g5��qDpb ��7
�
Q��$�F�&x��9k�ȝCی���Z�q������V�9����,5�$J�<Q���G��p�L�j�pQI�q�ha��nL���7��{�6)~xNxQ�3�B��w�p�*�f(�n�w"�=��+�(f�{���1��GS�U/Bh��a��G"|G`����m�2�;S"Jϰi� �!
��߈p�ih�6�����\��&f�*�M����ɌFM��\��	�h7 �����,V��W���R�dlU���:�eE@�pb顖���`�>�ݽ����s&g5��d��rE��#a<��R�œ��b����:و���rK�p1��0`i�)��i�ћ.�a'wG?�6� �ܡ�wŵ�zm�$E6-c�	 D,W��Zڙ�p+8��P*��,2 ~�2�wZ�D�>
�Uve,X�]��8����)��Ƈ2G���T�p�c I�,��./EŧRPj&��8�4̉�r�Ԕ���P�:s�T��Z8|�y��H:�r����yi���
�WA��[#�É||8%�I ��2�ܦ���n���n0�W����]�"Җ~D�����k��%��%����ͻr�9K�
��4*�E�LB����^+����6�E�;* q>tsm������JP�a(���z���ER�Q�R-�$���_Ԧukwe�w��{���eˏ��x--�W�^�kQBJ�`���5 �#��� "��'���{���D�t-Sc��U�����)�'4s��]��H�7N�v��?E1�Ȅ�Z_kU��i�I�M�����J&r�m�&��B]�� d<Xmga�����t��ƑE�� >��k�W&�+X��4��zkN?!_z&_��}����
�hW%���2��4 �]�C��Q�ҵ��̶_ne�z�o&x4)�L4�ud�������-M�|��/�ˍ��������vA���r7���{��RpXL��ç���@�
�	�cy�|��5܎��B�`�1�ͳ3�Y�7�pg����wDe��`]�W��!�{z�a�f��H��$���t$��%.A1C�����h��XʷS̴�GO�A���b��v�B��N��\�� ����1��C��#��j*�D���k �&���m�./���(|���_�� ��,b�������;�q<���/,�<�ѿӄ�A�ٝCA�-^<���F��U�c�b��KWhs'���]�� u#ҧ�U��p�ז�� ��6~yz�A�t��D{g���9���DG�ƃ'�[����)R���f���h��ìX�˥.�.
�e}���V��:�)С���(%���t �Y\٢�[UI"�����=�F�p1����5NZ���e�ٶ��V�E�?�ow_L3]PlH/&q}7�"����6��t!D[���`z��No�4��r�.�o�����l��#��<�{�$bT�Yf�"�g�7�n�Aؤ5,>~Ǣ�w	��sa�"s��06&��l(&x�"���@<Ứ�[m�����/2�aVb���[ �>{��'�_Z(��8���\�R�F���M�դᴢ>�f��<��{�����J4��b�I�YA�U�-d�
"2V�젪D7��H��pY�~*>u��qy�������K��`ʭD�~�"Q~�@C���ҫ@߻��\���-{�5���hZ�RhB6�0z�x����Q³j�X7A���U}����QT�`������<H�x�1��5a�c�<���lQ� �n ���WN��͋q�LN�ܷp��:�ȳC����v���͛��Y����)�h���.z��?�8��L�Շ����c�p�@^x�v���r���L�)�{Z��Hw�� ����������۔�����W���r�oO7T�k��`�v\���4�6Zg��|:�8
�����r��T�:��&o,p[�E|2��F�<�x�c!<�Gy��K�Դ��K�Q��Y�S	 �:i�ݤ�&�Ƙ�ٕ����&����Y��~@�W���㲘��j��N�!�Zz���q�c��,�"�*2��]	���L(M�e�Gu��M^�p��zb�����Z̒��Lx����,;���_�E��8#HD����R�V�1��g#9�Qj���Ș6�V�nB�t��T�o��W!?f/3���V���]f9�V�5@��h�׆g2�^��&j�4�aJ�r� s�Abt�wJ���l,�����N�ʿ��.Lt%y��0�������[I\�6��\��ct	H,��==b�p�R*�0	������V:s?�ܗ��8�{s�͋���y��jg{y�3���v���:�_��(c�]ż��u��� �▇�$nꓶ���{£p�*c�ѿ������7�����+������� �4^���Z9��$�P�����N�/9����S$������Qx9�aźO"�(�bx$�!����q5ڔ�)z��g�q����~����U�5S�ZHw�t6cc�Va0P����v�� �H-ְɒ:��]O��y_�Zΐ���E0q�G��\_w�z�lW�(�?�b��˅�}����0�6�k���9���D1 Ջ`�]��*�ǂb�岐[*�	�-�z�ҁ�P��z�ߗX	����RM��K������,�|���l��Mg=4AK4�r/�&�	s��˚/39ohcV��Wh��d2�r� �@���D}�� �ɇ���8����1��ΐ�Q���r�>���\��#�YA��rɃ\�31�U����"��������,�272�}�N����C4��� n.q�u�UPDdF~�\��E�&=W�ny+4hNĺ�V�~=*<.��ZŐ��K��E�G/F�=�oUw�6��{86d���4Jv�t�r��`��γ�e8B�k��1�J�3��>\=��To�o�>k�@iTMJ��I�����|}uXZ[w;;(�ʿ�+�YZeԥ���ܓ��:�=��� ���x��t�#��y��XD������ڪ�h�O8��Yg�"�,��N��b<��������h���j�u���+��*�2v���KZZ\�/�Y�
��q�?�Y�`V�T�����h:7���AN��ѓ��� ����=��5���Ɲ���F��5�C���+�F2W>w��f���2H���5U�)*���3Du�`2l���H$���#[E�����|����V����_��w+��bf*(ee:�i��W��cB�K:�,�c�����i;Qe�ڰsF����4���8Qo��U�����ѭq=�X�쉋"��8�ޗ�F���kg��B5��:x��z)�&���5;٭�8߀��2��*E:C:/ydq��w�i� Jl߆̸�t����C��i�~�l����|%�PJF
�����#�|��~\�l��ZL:�H����� �ga�^�?RLT�靱-˔\�6�����+��0�5v(L�+��<��t��� �x?m��GO<-�U/L��إ\!�%h"+�op�5fA�F�ϔ����� �/tz��|,�<K�4?{��������� ����j�w�:ʌ�/�QY���)8�B�U�M�[3"v:Y�����9�K8X�ԭ�0i.� M���d�UN�fm�p���a��[�1�wI� �6��M[�x��:��-U��lIM�mX��q����t��r!�lA�5�Ѥ}?�Tׁ�I�����$b��[ϕCw|�惒V]Lf5s���m�g=Q�?k�C%6,y������j\��$)GQn:��e����nG�i0JEb��Y��b��4_G��d�E��Oqt��K��� Q��h[�*�ع�����;Z=�<�uV�)�^f�9���čWrCk��̋�M�W����e�
%�lt�2���S��:���l02��m%��&ܹ��C'���Za��d�_�a4�W=�ް�Ѽ�	��#?�����8#az�_�*'����SD�����"��r׉�NX��%Z��-�I�l��-:wUlt�����V�u̒Mb2!X�S����2:�)p4�_�i�q�i�e���Eu$#� ��aC��%�c��	|�W녊�6\r� ���d�5Q�0��fK�A��(x�� f��h�S�O�v$�d70k��M�6���X�Z����b9LU1.�Pm�x��4����eR�c:�}������pϞ��q�����a��ʜB�������T��^���nM�����	�g�q(�9b![D���*ٌ����Z�0+^a2s���KlMר��F�6�Iҥ6��he}C[z��!FE����=�Y��CZc�?�"��d<���=���������\�A|̞~�6�� n��ߠ��e��Aڂ�)����V����lJ?H��UL0�״�y�X�?ՠ>
(y(\O����ѕ/�X�&�,ų+�3�z*�ܭ\����[���q�#�b��=��-�u6move{���';��k
ʋS�� �'��_l�M$�9.X�%D?i�`�Hz��:|5� XE��\HW0���,1;���:+��`c����(Њ�띅���P�Ay+��#�(ȣ1|���e]�򄂡\�YWB�RH���d'�\���F#zن����wf��=��͓{�F�JU:P���)���%U�k%F�͒�1x���k0�}f��-�5�p����N���U,�e����{�����--COc�y~��5;���)� �C����!���^��j�u_v_��j�Z��g���ˆh�w\�a�� �l4���+��"���b��^�,궫Nw�U���{m+����E9���]�$��J���9�kbF�&�,_Z�pׁ�h-���O~]S��8I���Js��7~Ea���6>���ɑ$�c/�� ��`�3��+���:�����Skg���d2����qy���m斅�pRĢDQ��u���Ѻ�;��:9e̪g;��pС�v�Et�g�1�q(�w:�qI!�-!�a�YT�Z?'�JJz0c��%mlMXf����|FZ|��i���M5��/4�&��8e�D�|+Z�{͜Ov`y�d��$;/�*����ئ��3.&�H��K��� .�fp���mCܻKB�9��V��o�l�B�I#���هz��B�v�ㅢ�Q��{�s����S��B�R�0ӽ�p kv�"~�����
���V�z��;*�[���L�D��4��~\_5:_�K��G�Vc|�Egd�bԳ�Xa�]| ��&��F�c��jP�_�d�j�Clv0t��ۮ�ʑ٩@����+	+"+����� _��9ӪQr��1S\zIS��rH�\&]�Z�llo�O��1�*Y�?܍����Eh�b�o�^�y}����GT�R�>N$�d�K�jT�NM�L��|6�ur6��S�	�(�̀R�vJ�cǵ���|{#g�t@�j\�!��J�H9bτ>� �K:��:H|	����5Ҧ�t�4�kͨh��e��V9UN�۲����*���)�˚�A��o[h�� F��7����#:.r!������[� �C�<5���{F|ۙ�c�ʩ�����鑁�s9���O�?)��P���Uj�lL�qB����F4;�3/u�s�nvh��3;F&���u��o��ѳ*͖Ӵ]�M�3`vd�JRg19�sV��Aq5��*�ÝT[��兇'��	��4k��	�O�f
U�W�6���XzZ����Jɾ�@Ι:Q���%r1�o��E��2��L��*�iO�<ڔkW<�m�(��Jؿ�������}�(��G企gZO�Sc/�[C��!+�g�eZ&A��6u<�)ߎ-l����X��Ѧ&�(�'��4�H^5D�K��@i�Er:�J��aWy��R`�l��N}u�������GTǽ�a�]��BP0���
]u���F�dPLϝ�5���ӑ�_J�^)�A� x�:��X4Q� �xI�@��H��D����Q1�/���ӊ����~�p���q'�W,�r_-[!��~��`R��1�H�v'��W<�J�,���:D��TC��%?詞�5V�%~��%� tֱ8��������:ĩvG-'�k�y�p���	AT��@|H~��;Z�è���5�ɚ|y��dB�@*�k�BR5k���|�lD�	�y{5y�
��z$X��v��]��y��]=��^�?��7�p�,@A7����U����]#��>��W�KG�Σ�Ct����Jy�4jګ��u��ݕ6]�x����r��
v�+�vː
`9�XyN�b��3��))�B��.{��IO)M���x+�K$���s҉we+ZkW~Z��� k��WM����	n�n���p7@=[��/ /��1e��M7�d7���{q�X�.ឥNbk~BcرH��( ��y�+�#����O� ��2�����*���se�<l��U?�f���f�����k�0��j�}�5��"cK�M�}Qד��*��0U���퍤� .pd�Ɋ�(�p����nr�F�ҝG���I�nl���(`dט��i�����ig�z%wN�k� S�J��|ܙ�@#%�eƆ646�YNk��q�f�0��s�N'Os���L؜X��~�1& 
��R(�/pFFK�ݜ��t$?1��vK�2�?:MT/�(�}g~̯��ƕ�� D�ct΀�'�so��NW��,~�f��+@N-�< 3)K���>�ߌ�r��f^�9��]ε�n�E+8�E�X��:���ҵp!��I�1�A�4��ՠ�ɹ��pL�����N���Na�(=�T�����srt�i�kC��g��/ޜrO��</oH�.֦Ek�w 	ģܝ�;����x!��;�ő>�8Z��� ��Е$a���-�j�>gEF.�\�V��O|���T"�5!�ު�<{��7�6x<�����WI�U�a =h��$p�w�-�~��ɿ��4��u���C�Z/_w�wm��)���k��'��pt|���d��W��m��m����Yj-C���Y&����j�Op⴫�^$.�ɍ�y�Q)�I��W�X�Ma7o[��]��}^2��0������v���͊���
s]v�(���&١)Pv�(�׀3�}[�����0=��}� �ܓ�R�bWa@S߶��\�xS�]�#�<��D�/}2AW߄��֘PJ	#����Ȕ���m5�_!���L>����=�޳�D2��WO�#��WH�չ!�S�3'�*p�S��*��/�c/�K]�,�� V�����F�#��0������K.ۤ��aGg�5��F��İG����aP���� ��)=͗����$Z:���=����ο�c�s��J��J�2�Q���։|���&��W�����A�����`ԨMn�0�-!�����n F���AjK:�X���K/��1-m�=Y��+�|��b�^�7��)�=x�9J#F �ѯiaO&�D�ᇴea�ؾF��<�ڝ�`�ێ���ty?sG� nS��������|<񤃛�F�X)��jВ诂�Bw��X$k�:�zJ�]23�]M"y8Ѯ=� ۋqB�ٰT����l�W=���6԰7Ǳ��f�8ܖ��g�t��[@3�	�!8����x:���Qʗ}a�%���RH�eלA9�XgL��ײ�[�����d�9���C�?�\2�I��V����e�l}����6t�^J��6�P�xW�'m'��` �������{�Pa��;��?R�$g�vҰ2ۍ�牼&���c��x?�_}��C""̔�>���N���� ��̘�n@IG��� �D-�a)6���%��5�?Aӑ��uo���ʼP��
�s�[��x��9^�-�<���6����M�.DW���٨�Z�?%�}|�8b�	������1�׸���1 L#|�M�k�d.�$��*A&��¯���O�J�H=�EG��s�R�Ki�R@�G0.�5ϖ,A��t���F�ָP��z3v�V�+�4��Ed�ْ�~�T-���n�S��5`�����n�O������f�� ���(�Ý����c/33@�f$�]yaTI��p�~ʯ�P,}N��$3��^���>O���\�|����ǳW�rKJ\|�˓R߉NLە~C���z�z�s��>g������ƹ�����TV��w��dN5��:��s�J(-7A����Y�_9�>{ -aI\�VG ػt3�	�m�M+��t�0��M �b>t��Wenr��ٯ���su���1�/��)K�D����e�b���މb��5�8U����X����v�f��jdg���ߚ�B�<�&e�RHu{��,J!G,p�sQ�̖����#
b�܁x�:��.a��!���tn�S���qj��d�m,T����}��3��e���'���m��,�D��ϡJv}bLu�8�
xO�P���� �O���=���2(f14���;)#Kh��go�����S�Kج�UWw�`fj�^� G���[75�Ŀ���זzK�Dȏ6ޠ�2"�(�������ɼ�`�s���>�P@|*�q����UW���Ġx���j��%b��R�r��N����TZ���@m�� � ���V=T�mVfy7�F��"�P��A�S
EǁZx!7���ti�/UK4��t��r|pX�q�@���l��Y5d{�?ϸ�����Re�>�]M�CV�l�V!�L
QQH����=�?bW�����n�%1ݳ2� g ~�b����HKmA�}��TقUT
"�ڑ��-�Z�!��"��J���3�&��L
%g4FPZ����������&�ǘo��6FT�5Q8��Fa	��t��H괥����[ -�Qd�`��1ڕ6p������n�,@#�+
	�V
-����]�KAM���&�X����=��Ԧ�QA7s����Y�(��_���s<肼��X��X3Fd����!���e/>�ܲ�G�H� ��Q:��dN}��ٙ��3M�w�	�L�o̾{���QI:���iϧ�I�ZFhuc����IW/Ѭh�P��M��7�o��̸��7����'cgz������\�8�o56��V2n�c��`�')���.!̝�q�}1r�j��u�	��B�Qȅ�/�i��>�
V`��Ca�[���sͬ�}hC��G%w΢���B���=v�U_Y�x]5pԢ�M�F+�i͈N���_h/�"�,�������m1�lyJ�;.9B9�3���ŊsN���9��.	(^a-��p6�$Y�8���+�h~5�7��U����!炜!%�栂��^	i��_�W0�fX�M��HD�IҾWòx��.�̖$���Ū���J���s[Ҡ�����h�	-��U����p�؂�:�'����`��DMmPF�yU@
g;�yM�_�r�ĭ@H^�.	!��jnJ��sn,�(D��^���>�1����Zv�$�G�������;HY^�p됩��Ut�_���\�$��'��R�7:�{���DP��cE��l�vaT<���4�,�{G|��L�}:�d��H._���"�����Y��-j�`2�����W��Hƥ��Q:��@�zg�/ ���n4�>���k��w��yn�z���B^��{bE����-�A*���� Ҁ�&>˙��(�e�BOH�4{�����CԹ����<�ŝ���?��v�}�0y�	�N�KL]���!�VKf���Z��e��\P�4aM�؅U8�=�4p.ɾf�ea�PK�%��D.ڬ�a2�1����B�3������k$�wF�J�Y�����_�|m���kj�}׹F\�T/�2t7<Y)Q�6f�r�/q���$@���ͰD�"l噓�d�֘�NR_u�K��^�y�Ɇ��)����aޢH�9	�v%F���u�����E�S~�%7�
ic���`�K�A`�o\$����oHϴ��0�k|":���Q���GQS&��c�j_|U�UA��uq�ϓ���tjl�"V�	^����^�T/$���'���*���xs���L�u�	̫�4����Ģ:�?<��w�)�떾+��r��m3�[ۤ���Ia�#q*Nj��7J�8���v����1���r�L�x��~aeG}�������؍�@�?��V�~�Ē�9���:����\K� k�5�Qо�{MOO;�E���&�]E�,��W+��2�2�!Is2s�'��Z�˚�,0�ARYA?��=��ak�����2��'����tz%�Ko2ʄ�^zݲR�0#���7��G��Z�H�-B P�q�M:�H�����W���j�՘p���F�JG��OV�,U�t(h����2���Qc�٠Ҁ�j�U6�B�Ȑ~�p/�V@�9��Kd�B�.�D�X���`����'��A,$*�p�d�S��<�^ �^�Z�O�z,�?~�qz�ܱ�k���^C���X���ex�[��P���F�6����ˎuM[TQ�9D�K��:������y�\��<��C�>(�eT�;U�f�J��������J��8�뢹c�݂�oq�H�ȡQ5~�L��n��ի�)�C�>W��(t�����i�{�ua�tΒP��dȔL�F)�����!�z�ԛ������fv���i�#V?�*K(��7ʳG�*r �D���u#+n�3e:5�HF�����d�_ݟ��]_�����ߑ�h*��� 
�>l�4z�����A�.�cU��K3�gѪ��q/��:�����^�Ц�q�ʷ�_׏�׺��ɫ��v��uӚ$&��]5?ωpy3t�]�.�~8.�H��q�����h���u�a{�N��6�7(������?����).��("6�����?�6������˚���LN3-�}m�D&A�6�t�D1
Ɔ��qI�Q ��8St9����;\I��1&ǒ:�gr���	�n�z��\���+�#�G0ײ��1��uC��LL	l�(�����y6���x٫ ��[رܣ8mn�
��{OX���Y��J{�A�*p\�O��{m�W90�<����02��f{���˘ػ���z2(k�O��&H"̐!�f���G1�%����d�?/ !FO��QPL�)��rU�g�0 )�!��C"_�1z1�+x�bT��P��-迻�,��k�մ<��<���J���E���#���������)ې�	~d��b2RK��O�IO��ڋ���C=`�R9���i��M��k�	<��l��x_���t@��3uCT��1X�켙p�t֨�!d�M�䟤6��9:�Xl�0����Xճ�eF�6���]���M)&j<�c4�W����L��ƒp��NQ��r�C�	&T� �+����X-�C� g��E�rÿ6�����#1�x7qtG���w�Sъ����#���7/�)Ʒs�=4��49�������q0���}���T��BHOo�qW���Q��q�K�H���4gm�Ӵ{�;�h���;n����E�9QJ}��8���㬤��A1j�ζդO��c�Sv�!iX�W����y���\�ok��ӏ2
!��?�;u%n���5��r7�*���$��Zݲ�+wҙ0s���U�xq��z�/��0˞ 4(.��|z;Z���N��
9����8��ؗa�������ኸ$���'U�:��m�|����]��{ }Rg�cڴf�ҒDM��n�}����\�ĭ>�Y�{��t{�D'�x�H��{T�3�`�v�[ν��vj0T�k�ZO�GA�i4%5S��Y ?�Q�RbV�=�D%�����0�w��-y�Vx\��䒴��|šay�	����p��O�e���W���{�����djVٹ%@,�5���;�+R��߹f�ۥ�0�pt� �X6�먌��B����J��:��:�d+��tf���9�eH��l���JO�x{��x��ܚ,p����d��wu��(��k˓)�� �'�[���ɖM�0���oܬ7�]�=D����U_�����n9dZH�`:�����f[=z r4g�F�TF�ͽ�&-"!PoÒ
o�E�J&Lsc;6Jn�dyy�5��O$��� �TL����?��.�­�\!�4�� �^&�w�"�A"����7ɜe*4i@�L��J��hm0�Me�U0�h�R�cШ��ڐd/��d%���\���SDR�\�0Sd9z��x��1#^�Y�SjS�L`�8T_f��3q��6��0� �h�1�zI&/�Ocf]pt �>�\���Ydwr���.�G7���ac��<׼�I�5�T�"�FdX�C���.�)mR�g�?x�eu[be38M7�8��nw�w�,�P�`��S�hg�ݒ6�,�ȩv[, ����n�k�&'Q�U�t�?�d �=iy^��6j�N՛X����R�n\p�T���(�2�X��ST�^}U%�Nd��I�.G�/�2���M��_�樣^��⨞��X�vq�Jx��je*�}�f�8��$R�.m6�ߌ�b�Z\^�=\�ᔣtկ�3��}���C���I>�m�Sd^�·���1�}�y[����o�`P�+z��<�����Q�I1ٚ%iɯ0m�w3V)��A�fjm�o3v8�c��L�nڍh�k��c^���:�Ȅj���p�)��`��4�*u~X�%�$y���C����_�뺛ܜ����^N���V����9Ѻ��`�x;��5�
 �^��DEHa�ޗ�ui9	��a�I�T�,rf��I�nv���G����yۍ1,�jy�b+�~EN�5���
ds$�l��B{���5]#�����9���й��;j[�5�Kc}X����"��@6��ڏ�vhVAu�O�O��?YMՉ�b{�Z����	���e��ԚM CI��;��C.�B-�+ˮq�8p�N���� �N
��6H뚍?ߪ�Fx����bT��WmZ�f����x����O�Ʌ��t�,Ó�j�$tt�-�$��E��BN(�?=����G�7��c��yk��qIo��+��v`ϑGu\J���%��v��A�����^Ѫ��fCr�_�*y�$ʹ�T�R?�)�d�2��ʳ�
V1J9�S�TZ���Ǖ�9�2c!��n#��^���\��bXcL57ܝ��w��g�ϳ�M��W]�W��� ���U�,��e�X��FbЫ���}4�!�`T�0�;F� u�3�Wx�i���|͔���[�:B�!��������r�������	��S�#d6+�X4��6��^.u��<�0)W�gaB5� �Z/����Q�A�֗n(٫�/����`C8g�Y1��&R��>�vB�<L��:�-��*���Ř�ҡ8��R�-ם-�*L��>�zĶ�Ѽ;�.z���6�ܩy2�9��Q���|zS�a��������[-�t���#�o��:�"�c���؞��*�c˕�֖h�'��A��W.�t�f_���p�m#���M0:!%�K�!���G�lj��O	��7�ظ��Z�a+Ƅ��xx��/��s/�\�� jL"F�oX�*ݭ4!u���=cز�\5$ɳF��5�c%�z� �K�q�t
��~JE�3�K���l�}BP�����U%x�[�#`�M�FV�Ũ�����C���H�p鬫�5*-2�w�F،f�Lf
zB�A��X�:}c�"�1]�[6���A$]ل��#˧j�1&YY^S-\�6˽g,쓛P}@r��p�Q�%O?�����r:���7(����R�q�B�}X-�v{��}}0��F����R�ײ�@�_]L����R�mG�_��d�;�)��#�-[^��'����5�d�7j5�i���)~[�)ya�Ć���r$:�'-B^T�"<|�D��pɑxT���*�ɡJ�����b�="K��ԟ�����2�[ZM����8�p�e4��Vc�Hb��D.��V�J��W�j���z�7��������c�\A(L�S����k}F�hvTp����o�Z����#Q�*U���A��Y�/�6vs���},��І_$bG�䙔��d\�ވ�$���UW;��X/�"
�Z�jL��:��Tq�H+�WXQ;L>K}Aל�X��}s�z��P�xCK���wL���9)�*��_��э�.���m�m�!_n�%�uO��C�
io��m��MGǊ( �HfPCi��Yy�{5k�"��L�ƛ4�m&�XN��MCԹI� ��X�����Jv&#�U�<,���h[K�]��� %�iGo�h:����3��������ҏ/t�_�nMb�hȣ �:��t����=(�Wߠ�;� �����S�]� w@ �)ް�I6�7>���.����]��0����q�yGE�4~���!��h������5	����<��Ϗ*��drc��F��F]�u����2�}4.��j���c�� ��X���g5���������/z���a��ԉ6Е��|���\����"�kȟ�%��^�l�����r��i���T�2
�[�� ߳~�쿥�y�N'��JQ����r.R"�
�3�����X������ד���2��)�.Gs�:��\�3�s֑����M!eӺ����.�o��ǜo� �1%p��(�� ��V��>�G��,�f�9��� ��:E�aB��l�~ץQ}��Hx~��~���|�?^~�M�(��,�k��	����t�`�h��"�W���O[/d�t@��L�9� ���X@7���A�gOi�:�%l+ �Ja��~��^�G8,�'����Wy�y�����\w�l�� ��|�tg���O^���'��0�^i�&N���^z�I��sυ��D�B)L.}Ő�����ݪ�0|�<2֔ʍ�Nۨvx{��$��0c#��dh]�ԃ	��)@C@�.��H �����k�t
�3Q-xhǷ/�jn*���6��n��L�~��M?���ZFR�Pjk���^�ZD�N��A۔1�tt��2S��T��F;.sH=k/0K�Kb�i�J�X��7��mH|��<.ӹ-jh����*�Y���/'��R�ig�I�����.rl�T�0l��_�p�"�%��L�:�-�����r������Fd�sca!��?J��y�������\z\��R�/���@�4�x ^@��+�����-�U{2�B���Ý���P�[�)�`�`1Wܵ�XJ��w�!�H_����U��y����Ǟ+kM?92uV]���Hnؙ8D���G7�.�YD��4*e��HF%+�٪>)��B�m�Xq��2u��_nb_���Y�K-��_l��)�o��L˂��B-r��K���u��"@�N�k�W�Hy���J��C�.�~hT{a�J�@�R�*��q��w���tv.���qq9���vMG�����T�X��:t,�^ee�%��x}p�⛝x���O��\k���H$yV��;��MZ�ж��=�� 2uW��v�/Ie�$"���Q˶	�������m곑��"�]�`J�Wu�ĺd8�i�*W=s����dh{㑠<6�K���.�R"�i2��)��E���C�������#0��[ �����}�)dx9<t7v����Q ��!&�T�}~���?j_�����5�H�m�`�kB��.YzH��T�e����*-���L��x���&�Gc�_����ʱm��;�k��I�[+J�I�����9%9�c]  K�Ryna���C.C~��l�o���f��ִ��8M�+b#M.4��E�'(�ur�hE�H�P���-u,�J^�5��X�ɋ&�B�M�}�U��^�K�4̓WT�AH�tL��N�^
?�2�=�弨����ߟ򀜠��g׊�fDw��ݠ��
UV�X���~A��/����()Ĵ�7qZ���n���^����\W3�P�<�3�JE�פ�^���q 񹵿�jR=桚}��z�P�ց�Bֿ��i���m�O^�0t�^�)������s��p� �@?�9��`��0F��fMu$O�N��QN��s���Af�Y|����SX&���j?�c���|�*��\֢0d�"6���zC���_�yY΂���l����U��<�c)�"K�]�jSW��;b�O�EX�R��V�>��q�B~�~tI���6�WV8��f��w˴�LS�
1��J6�p3��<�_C�
��VP�1�ɒ�����Üv��vv�՟�I��5^I���� _��sN����>M�lkH-���|jAF�FWc�1��<md3>+�Cِ0�p]�vΒ�\�kw�O!Uj����xrR�f��w���re�ʦY�B��玸Y��&{(��>nuG��6iA�s@x����.�Nк��q��yG~��7D%=��%��B=�<Ky��K\Z�w��-�S���/�]ǨW<�"��<bz�0�~
*�n���0���$ �&�
?`C����k�A �%h�RH����S���y7���v��w�Z<O(Ϙ~�;��a���� ����6�e�H��>h�^������a{#%�)3H��1���&8�yޓ��s�,�G<�[���r���Io�����<?w/�ݚ���v�M�^���)�P�V�H���|��c���n'��D`�������,��!���u:d�~�?-崷|�(�x��k�����'4{���aR�v(��W���	KD��ÝAÞ�;D�Ͱt���������L���q��.�ak���$�m0#𤳲��О\B��9QV�VX�~��"�����\��mv܎t�����H�x��� �K2��m��i���ؒ�a�|4���yKCr��sX-Ρ�c�� ~3�Z���a������i5`�j�)�e��%M�V�-$����i�d�t�����0�&�Z�!��fp<8R���	U�4)F!m�	:j�w�qG�C���?+[�T�:��	�;N�^MC��NTb_�x
�����qJ��/��{<�iv�n���U6\�_XJ�x4"�˓6��4j\�1��YV�y+���O����Տ��$Xn��DoM��<�=��<�qnw���Φ�8�i���a^�y��\0;�Tԏ
�+p/8���zw�oK�;E�9��H��ڊ�y�`���xpG�g�d�p������)�:��9,�qF?=1�Z��M�E�:���=مу�|�Ux�w���#��U�x��n��	E=���{�8�Zh�ב��}p@��(q�$f��0��?_�3|X�
��N��z�>k�������|j<�#�����-T��{�
��MH�A\[@��3Ý�I�V;u
���W��� ���aLj)�����V���a���W�K�d�����Ű��֐-U+���ܴ�~@_�g!��7�8$[Io|(��"��K�H$F&�}e�Rc�zF���O�.X�q ��sߩQO��K�H l̥]����᠇1t\m���I���٦��AT�2������J�g�r��QhjF�T���D���&/Iׁ_P�;Z����������U�� =��k��>�����7( N��P�2n�V��+#���q_JBA	-K/�����p�	�BQ陋�Ob��Y��hNѶ�a�-'׿*è�VF�.�O=�~��C��f����g�-3���7ƌn,=�޾�El�Qs�Q��p�ô�Fp_�&��Y|._��u��N�L�(�<@�9�5�m~�Q�;��TU,�.�T��)�!��)�ǬVJ�-<������0����X�WH__ܴ�Ҋ�0o��8v���2��(�,�*�y�%湯iql�Jӱ5T5���؜����0��OL���ƪ؝l�3g��#p���Ձ�O�d��������m�̳:��X�p#��%�K�m�89M����/�d�a/�g����X���~t�ٳ'�5�����*f&\����t����{mU�����/�X�����[H6�+h']	���	�m��އ5�� D�?�Ƙ�_��E�o�qփ�'��S�*�$wu��rK%�^�\�Y�rߒ��@�p��)�|��?��L7⏂I#;���>x^v��ئ�-����=2�1�JE��������XP(r�K������,z�x��T�b[��!�m7���q���+%���AK���Di1ꛨ/(�mhLR��Q��G��<�WY��[�G_ "��#_a(G3�o7����!�"��{�AI�A�^��cvum(0�S����ɂ.�|��z>0V;���M;>9�4
Q������M��??B��+/����o��"i��µ<qGa۲���.�Dt<��iI�W��f��� �t�H;K��R�Lz�쁉$M\����{F�����r�������_���P�cwh4�m˩z��z==���:��٧�%F�-[��ū��E}º���u�N��g%��i����eh�K�dD����Y|��RW �������̄�p_�E��q	�w��z�����T���@?�亊M��|h��sP9�cD�D�}�z�����3�94��nI,�9��B�F�?�Tw�N��xl���C��C�@�,rW��a��_�G����(	��N����o^d,a6��)����A��H�^��<��and/�?U�K+�V*Tq_N�vÂ�F�NM��G�[���f^� V(�X���������柭����Xݰ~4.�HV�q�K�?�:��g��1�	�p���k�7A���p���s����@i�(��t4@ȫ���?~W��?kY����>�-rܕcd�k9;�	���W����<IͿ��O�'"�E}v�5W��r���.�4���B v�8�G�T5��W�U���rmJ�$9FE9�Y�>��׮��q�v#��k�}��vv!a�L炀�R��,:NF
����;�6�|��5�ב��P_pH�m�֤<���,�n�����{+�q��F�#�({
OZM;�/R�㎃������n���EPE�g;
ЃdGr��v����Ye��؊��8��W�6��3��N!���&�_'I@�"	��F4\#�@u��ka�C]q��&b�g�>a��+7�!Zf��t����CsL~Zo)B^xa4	Re�?=pYUpّ�?�����9&(6�Т��Fc�|�I}Љ,�y=9���<-���50P.�L_<���F	�+�!6?x,(P9��"Cg��(��֨j���JW3�o3�ٟߊZU���:��Z-������	f���}��ԧ�x�t�X5�s�'Oa���{�� �#Bﮔw`��u�x�,��!�ĉȝ�h��>o���(����r����Z)�m��m������s�Y!1�gДr�9���Ą�c�>nՁ>��Ol�\�EK) ?2R����`���H��������"��A�AxM�a]��ļ��Iiӱ���=3ŋ���ͽȀX���X���7U�ۚb�R�Í���g0L'F_��$�#9�ދ���ӯ+pʫ.���5H9r���@��o��X��F'	����q���H�,@�
mm��ٹ�='�����d�yA���$�4_d������f��ȿ�v�����|s�$��9Du���D�Z�;pQ_x̼cO��Y�7��?r㞗"�1�����mw+DMd��$������x��kX�w�<���G�#ɧ1˗ߤwu��S���u� ���j��W��j��W�tO�J�O9K]������N�@�� ���V�VgtP�&e�Ye��|S:��4r0?n�3��ۘ���Ʊ�=�N�p� R���.�S�#̡}���/*!�D)��j��a
I��1%S�08�9��[�in���X��r��x���3��k����pU#
X8�J&�C��]oK���E
4���u��2M�]ą�%�@MՈA��,.��$�������q�X��`�yK ]bu�@O�b|�:�Bo��5��%�s��� C(���c��|�7��Y9���A������y4F��F��z����7Ъ`*�����_Lb��$����\�y�fGAP��O�\�*�	�Q ��--��;^u{�*���:�4�Q����,��\�'Z)&�y� �r( �WU���yF�xk��ٿ� ��%��&�(���N���X��}�p-���rj-&�s�L���Ē� @���q�|G���Xؔ^.\��M��h$]��]Qۻ�I>"\֔_e9W����1",��I�S5�t�u¥���M>z�a��ކ�]m۩���L��m�v�DB\�t&��N:��q��7HÆ�wd��٫���!$`:���a40���,MARnj�	0��Ԩҳ?|��ex��8�^df�$�۴����(^/|�d��?`�V����E�d�3-�.7-�E���ދ�v����756��:k!�ݓć��'ȟƣ�[^5�DBl���lZ�����[�4�G	f	��=�ʂ-��7A;�yx'�}DL!���x_N�A�a`3��k���i���`�?{n�u-1|��q����c��y�O��)6H�d����>�EL���� N��!
�1J)��F?�Ntk� >"A\&�$3E��f�,�  �+�)׎�w������o����[g��,��F��3
��*^V�qz92y���]#(�?v��ml�W��j��:(ɔ޾3n��[ʢ��W��D�V��vD��/��!O����l�c�cx��hT���� �M
A��(�P�S�'kV!	w�G�f����-�ME'y�W����F5�b�2��gū09�*�
��<eĉ������	h���A6��>�t<����[YPS�W<^2bu���Pk��s�k�lY��C��5��֐l4�����~͈ 3�%< �����L��}<�2t-��s�@�/��t�+)\&z�ʶ�?���zg�3�I��d`VQp��nA��[��n�	>K7FA#2CvS���뺱8�o�uQ�x6 *%���皠�E^a���v����"���?5�*f�%�k���q�	W�߂���O�&���d���J��6�W0%c ���-,vkL˙  :�zv��Yu%Ǵ��q� ,����67�A
w�����9p��V��άF"������ʢ�`�ng+�L>\���)��>��2�p]�Io�
��ֿU ��$]R�]�pw.Ft��]
W4��$8�k�!�������Y��𐍄��jT �?@yܚ5B{E�gf��5�N~�n�����^p�&c��0H����ª�V\6�n��K�e�D���]!��(}k�u��j������$-�ВX0�E��R�X �A���;�}�d�=b�(c�jJ�vÂх�ـS�!�W��C3r�!���X�"0���O<����<�j ]��w��T^��w��>�%��x���\��H��a#ls�&s+�ioMĤƹ�FM��N�?���w4'X�M�ٗ�'2��-��\��Y���z����[��2�=�~3��N��>g�D����#�m�X}v3����)=��r�jk��\��;����ęQa��rv��G4XӉ�Ƒ�(�h�#jo����`g�a1�R����]}�[��:#Ʀ�m{Rΐ�I���\�����e�z��o��b�V3��`�.�Y)�x诩@�9c��b�I���5�������3���5���T��`<�/�fd�/�-.IdT#99|~�H�f����MeT��f�@���������[�:֕^(>��5�D�m�{4X2%�^V�-<T[V���6B��:����f�]���ƛI�����vƶY�G�@(�vcQ�0o
��D��E%+dލi�Q���xHz)F{;�M��y�C^�U�2XN"'�T��N��쪡���1�}[B/c�M��^����k�P�h9-��'�f9%?�U�����)�_����Bw��7"�F�sg7�?"R=(���9Ʉbg���R�&s�L�/y�ݘCX�&��	=�ƴn^��I%pW�[f�.�3�]�DxP
3�a>���H��#���\����U��6I#�������/T'Pc�X�f������.]��] \��Vr r(�# t"�ې�+Di.��ˋD�'�M���0��Д�9 �����`��u�A$����0���ZA	�:-Y1�I��𛦳ѐ�n�`�:�Ѭw*�}+G�f�54بjOP��d�N���D����Zj�ϲLc�t�~�P�!F '.�N�Vh'��g���g&$��(:��2�':�	(XńQ�f�&�X��c�8�M�ȀkL�KO�e���S�>fJ"h9��(�d�ƫ����^b�k�g]y�y��Y���羷�w	D��/o�U�	�|�=0P�ј/��B���r����N�{�<�ↁqPK��;�H���p�S�H��F//���W�řb2��ؓ^G�+��m��eʑ:ʙQ����7upEp��ol�M潈H��/^��5����9\��S��qr�	���H��8��-;;KT��;��{s��(=ܜ��р/Z����#��Q�.l_F�ɨ�� ʉ�d�k�ind��c� ��=Ϙ7>�.�	m��:�Y=�n�*����'�H�,r�LN�Vazh�%����|�����UWȥ.���涊)̜B.�T�nպ���4A:$����d��&G��F�P�L��qǁ��%�A��ӝ��}�;4�f��;�YB�O&�@b��,�3� ֜��k �7�a���g�XN~k��	���=)�O�hq�����T�˓p悚%М!��%���v�v(�4�i)<M`�=c�Κ@��n\Gf��\L��w����'h���e���YSUݙ�M�h�Hn<#9"�"51&H�H��w��<�^�@��pb�9*U`A�_��/G{&^��P��L�1�-U\*�˛ 7 ݌�k�[4�����y��>��rr�+R<W!qM^�z�E�G�s1�:�yQ���P����y�Jߌ��-⎇+<�T��V*����FPCs��y"�!��W��-��u:�����F.�Ԓ9��F��<`wnt	i���"�fƅ����)B���W$7v#��DI�a6�����	n �DD�~djn%ޫ��n��^?��IK��X��C����QZy�B'Ӝp�>t^��H�ŀ��0P���UɌ���o~Ye�g�h����Y�E�(��,`��h/�6�Q�>0��I��ѸP���m� �k�x^-j&]S�@�p0O�&u��X���3#�	e�3t�
��#������~r��P]એ%YӺ�����,��=l���]��h�I=�|�����n�Z�uE ��.�nO��f�f1�� ��dl��Sk�/X�N�[O�4$M� ��c��H���4m7�v�<�@+�RY|�>�Q��}�����&_�Uh/����;��=f8��"<�SQ��a����+�UW��Ԕ2֒*[h��!��͸�G�qi��d Ȓ2� �_��Gr�;��*���� S����Mw����`gט�@�m���Ha�=����&��5�k����9Y�b������ݔ`�L0הA坃�r�}��:��x��o=a�?D>�����ң�,�&]|s�ع)�������㪢w1�+�I^e(B��Τr�b|��hÈ�^�Y���1b������T�ZN�h����5�y��
G2�.H�g�%���j�V��kta!)�qOw[.N��BA�?���#�Yߖ�E�b��6�x��F�O��;���-��'�T����]:>9�'*.j���	l>t�\���{�*�i�����g7ՖZ�^�~)����qO)��ͬ��eX���4��瓴�\��&�#J��8�_� {��ہ�>6�ز�����C*y�y���9j����n�[������L�LT�`�\J�0�O��|�n8���O�؎GĲ��$
�����I&	�6M�Q��%�R����AM��mX�1�&ڙ��5!e��ʜ}��)���A��De��u�84f^�<s�������()��?���C1�9�_G#d �p��b�"�x���iԗfr�6�b�
 �O��6��tEЕ�����ug O��&7�1ʗ�Ȇ����J���޲#_��t��IGf?"�Ḿ��'R�����j����D����=P�H������)&5���f�
x��5@�G�l�ی��J���T��b��7��(������u�[|GF�(�W3��f���j����<y���0��+[��:�p��O��"�l[�`��˻�3�̦3�M����Lj~�g��*4�!�݉DG��|��}��¥�Eg!i�=z��� c1U��3���^	tV�核G$��v�`�q�(��1(i��B�ﺫ*B���J���O7��OOb��M�B,)\)Z�B�`-�o߲����&�����P6#�t���m�]��|YP���1�������Z!N���Ix��)̘Џ����J'��^�)m��S�}�A?��ds���.�?�
ϢD����"�
��)%�l�*z������3tƈ��(�z)�Z����Ǒe���Q�;���E�K�3TE���c�U��q��mX7JӜ�GNI@xJ@�,7q�[��󎣬ШP�b\�2�h�?�աՉ ����)��v��-}��A���V�Ѷ����1��$�o��p�W�}�R��v4N���P���sU}���e����t�g������|B��C'����8����|����`}�iE}Mr��� Edÿ�l$urn�V��aВ�ߎ�uM�n�i����} VP��Q *B)��ܼ^O��?���;t�q����A���AϪ�2U'�0��K��4��2Ϫ�t��.���P2P�Y�Gj�as38�b���ĮG�`u�nh�C�0�nV�I��f��KE��C-o�>Ģ���i���]O�A�.~���C3OVOI�SZ;Q�_�
.�Tl K���&��'(�x�%O��^��ǧ���L�ź߬-�6��y>�ML���c7退���'����c�G7]�x�+��z����H���[H��?X�c������n��ꓗЁ��Y���=�����ޏ'�2��,��l���7K|�1�T��y���)�q�P����K�l���e��}؞�r�'۾r�Twq1���������̄���r�����/[��:3��fh!*���X8�;�cP��� ̶U��~������=늣�#͏����C�r^�^;�W7j;��b�$5��5�������Wd�:>M�1΢;����+�yk@��N,���|Gy��h�JJ.����,����pX}� %0�"�m����	|gr�h����+���М��Ǝ�Z�=-�������V�k��c�6rl.��)���a���9�`7dDU�����5M�+�5-�I����tM�`�դjە	Cz\g��j5�{���p�bGn%�}���"<�!ӣ���[��nJ�Jh![��P�@u��+���/>>�4o�PP-4U���wsk�̚S��s��_��2	�k��!�G�@3�υ��M�A�ڻ�$Zn����춠n�woڤ�[_]��Dd�VE�[Q|��dQ=�Ub���0�'&�X�-�
gr��J��v���������fU��l�����v�O�w4y&q�����'Tcc�$I%>��	g�;�U ��j�'M�������]1�>.B(L�gm������A|��Ҿ^���	����������!	��oVJ�b���!�Z ZF�co��^���s�������X�0��Nr�h�S6�4n 	^)�R��R��fK�?�/��T�81��m �,y���ƒ�^��w��T�T�Z�2��a�q��
���]CJ�d�_�raځ�N���?Eד*��>�$��\nN�}��z o1���N�Y��E&m���hP�s|(4����ww���V]��h���Obox;�F�����.żtk=�\㘍�֟��1\}�aLe���1��s]J��/���s��_�<D2��w��BB�M�2B�_mͲ�C(�ޅ8L|S�K��0_���K�ᐤmu�jf?i�1�H�Y��Y/�p����`zy�Gg{�=�21�:=w�J(	��u(�I�[�����$cT�ePКVryUV�S9)m�B>����91����ҙ�,�g~R'�c}���9�$��Y�c����l��cu�ݺ�i�C��o1�o]�|���L5����X��Q��q�0�xMW��H�e��
��`#��dȘ9rT:�-o�SH�*��A;W��0��+�� ���	��@|��.!�@��T�z)|�F��ww�)���5'�/�L�\*TE������k"=+"n��s� eQS 7)8@e�׍���BEa)0�t?���y��K\��ɿ��N�nONV�;.��U9�_G�e̒��!XD+�6���Ġ;�U�����?�K�6�\�p+Z-x"Z��w��q1����m1��1@�x싆�V[��B�k�J9p	��k�<�$��E0���i�=�cYc�ic�M@W\���~�q�WĖ��p�kXW2�	=$\�^��t���iPf�p�j}���� �C��)F?ꖴ���Z�kK�ȏ�k�Z� �aeR��g�&>�=�J��?�=E���<�H��rx3�0��~������[%��rW����M��P�a�o�o�J��>f�-+߉���=k�f��"��abP�=��$�ט�$F]����P���CS��W��nĉ��k����$U��o �A�)�>�]�1��Mi�;�B��<9���m�׈�7(<��(i]���I��9k /�7zjFŵ���zy��;|�hN��Ī@6~��u��j2�Ŷ۴�a�/}<��*�G1{fm_��W�ި'��7���Uk픠~����O���4����$�=�"�ݔy����NF�Md% 0\ ��:�S�bE���sg�Z����I���U�C{j����i�@��fyɸM	-�[-��u��0[��"
C�y)T ]T/�EE6�1Ls� �fɒːߊ�Q�Z;kԯE����&�]��.�`h*��A�&� �ƳZ������4�à�"�Ff;�/n=ca���V�H��V0�q�������-�^9�a)�6<�!E�5@�Ʋ�z���]����2#1�� h�}�Q��_v����*��GѲ��B��X�g�l�&��L؟1u�U�C��3><�W���f��V��h��r��$@''��zU�V��<�%e*C����8�!�i#ӝ�b�D�]�5r��v�G�|��O^��\��q��S#+20;��)���.��iB��0v�!ܴb1����z���FL��f۹fHV�6�%�Ҏq�$>h��Os�Peg_?TpKl&2~�4| Y���[6���v�U�&[R�ߥ<�_�W7� ç~�3��Q����rq�U���LS"�ڋ|e7�R�&��s:
�<o�\����`AO���/���x@g���D/�f�[	$<� x�Gd��ʬ��y���&�lixxHU�P�u�Vx]m����.��Rxa@��$T�T����˜�P����mc�����i�L�(_UݶE��e��4���,�^WJ�-�:wC��<eȀ����h�q0�M����B�[�l�X8�m�x޶�v��o��I�ن�w�aHkJ��v3A����l!�n�0:?�u\��[�z��|ŝ��ԑLN�7�[����r�}}t��;���>>B�	��z�|+������O�	���=	��n���}iWJ�	*�'b���AZ&W�)ɟ���P��w��W�O�������$��?��w��;.K�2@����e�!r���.������#b�H��%����\?�B�T.�V�Uc�_���
SV�ɴB㎱><`�;Q�2� ���k7+��܄D1�]\��KH��5�L�Si��δ����F�tϗx�v�;s��\������5�}�c���0?�i�VE̯nLS(/���\���ἤ�|�t��_�w�0r�H7 U�a��'��w� ����:�޻s���9\��5�^;��.�kWV�W㏴
��n9PD�=_�4k�� lD�'�������y�^2/�j��͜;.
������X�/�eGy�Sp�Su�)&�
�
RT��gY,�H@7����k����4�CTX�F%-�1�.UZ�?�� ��p�_�����N��\�do��ZĎ��c��c#K0���*V�x[�n��iR�gb��,����P�n�A�i���7��P�ݪ��~�S�����������3q$M�n��CT�WM>��@��).����w�PO��d����S�g}�]9e��mv�K&4B.g1��;���G�|���/y)�!��ݰJ�=/�L�N{!�O:�/J�����8?*�k�ֽ��U_��U ��-D�~�m[��V��<!�&(����>�hC��2��q�/l�;�^Qt��MI�J�jj�23=��y1�=^�����v�S����si����O �����R����e [�+���U��u�M�S���h�+9��ڗ/�}z��f�b���H�Y��s���H���v�(C���C,�����.�#Gh�P�3jlt��A)o���C���� �2���~�ͦÀ���A)�CN�W����a����r͋��A�*�M������Up���y�I���u�g���ոy�	 ob�@L�d�m�`FR2�AG,q�/��=�P�'�9�D,�����G������=�H���5��"Q>ju�hoo\��ⳋ�翐8���;�Q���އ�HPK�)E�#���D�d�8���fk��R}�S�[�ȡ���z��F���k!��"�Ú�|桟��Ɩua3Ș����2�܈�v���*�����X���W{�	��E�2�Z���S��@���Q*<�������?�?��P���1/D̟tE� G���E�O	Zsܽ%�A�E�q�rf�[e�y݃\����V �U5;6V�?��5��s!:ӝJu���,'U��7���<�q�e�8;PuɊ!n+�1���=A�Fu<']�R���9\�²=���p�~^���1�TD"Y(߫�B� �� ;��Y�1�E�MU�}>��y�p?�^U��)��/S�������R�-��)A�����	�􍰧�qkFiQk{�u��n��61��#�c�?U�9ņ���H�UC&����,��G��rc��1E"?K�YEs:�*莬��P�ss��@�_�����E�c���m`q	�.�uO�*� \����vHG�E���G��F[_��Q.7%Ђ��o�K�KYZ�8g��o,��r��f���������6"P|�e���ټ��fJ�����=�ڧw�g]=`P铳�?~��̠�dS��7�H_����%O��R����G���Z�L�u�N�W�ߴ��>��(F�@��-�����	��g_����g��=�q�diۍ��k�Z#���H6|.GbU�Cyl#Wv@���g�k�P{���zpDft����ڒo�$�&�v���c�Bn�J�����wP1F��	QL�x	D_e��/���&��Zs����nf曋�¼�ݶ�t:��{������:�0Ʒ���[���4������Vɣ[[T. ����D������93]e�	�͒7���J,�=f��M�a
���m�O��t)hn�'[�U@���00�RU����g�5�W�b�����]ګ��N8t,�OEfD $�����k��9��K9���dR����Lh����BP����^���-�}��/E�큨f�Ew���`�x�ހ|j��7�K���~r����Ɠ�W�����A��o/ܻ��ݥ����b�\��SWF'�@���H�������𓳋j�.��\�}+�2��e]�ji�
1v�,�m�E>�����6�
r#�,7^Q0/�����$;j
J�NO���1��gh�q����h�����<Y�!���Q�s�S� �䋲o:E��1�YZ-��%W���l֫�e|�SV�*��-)�8S+��^�8�ႺQ��Z񅧣�l:�9keb˿2�AX��^3R(X}�ǈ�&'սc�9�.�L������^C Ǧ
���2QI#A�����^��42�a9o�f�Lg�F	�2!��`۠�PH�����eՋ��=��v�N'�,i/�=���ri��M������R���`$��fO�� H�>y&�(]�}��rPboB�^h�WSmH`���zmC�Nc�DO^���@��<[������αyX�hUhX�3��ߵkr6b
B�M�.�ٖ~�)3�:&-s1"+}��j�m;������ kT��k<uj �_�vW�=
�����zf��ݗQrp���L�K����ć_�q�-U��-��`ٵ�Vv8�V�;�NM�'�wV�IT�3;��
�(a�K2z���հ�{��*!���QcB��I�g��VL��8)�ˋ�Z�R��D4�65��m��8D��݁�Ü��}m ��������A^�e#���JI��i	y����?(�ō.�ݽ�q�%����j&s�(�k��޼J�Xv��6�
F�t9�$`�`���n#��[�f��+~�����e/��O��S �br��͖��:/:+H'5�r���M\r�N���R9������s7⎒�n���<x�����q�X�K|{��<^��o#����CU��#2�3u6oN���ٹ*��	��ac��F>Bf�mX�< [Eo"U�#�lBǓ݌e�e���&�q�@�bu�*;��
c�4.g�0B����cz��U_��	�s�
��<��~�(������l�Uv����_d��(l�����~����k��
Q��I�O}�'h:�"(��H�[�\/}����UeP�wFŋKJR�������FP�hO�
�9=5�!�m���!]�d�
`W�t�e��li�$��L�6x���#j�5C��y�JL���aԆ!���Ú���2<`�DGng�a �ܳ �l����0/t/I��F?���*xq����X����4�K�+}���J;�"0p\�^*�?���% ��7ebh6E�*j�� �(��4�;�Toz|�� �n��%����"�:�^�`Xf�K>B�c���YLl�\fR�|÷x١��Yd�E$�R���D�~��Sc3x��02/��y6��vW{x.��7����;鋲!��\�w��d&�R?�����W'L��I���^����av0ѓWz��q�Dx���<ڛ�fT��i0�x���=�ʑ�D\��"�@&ǙU��s���YEٓj����eV���>H�������-?�	�4�%Yͯ��L7�(0]��*A���覔�L1҇Xd��.TV3�5eƒi<d���"���(/=U�o��/D�E%D �<��5+�+���Rz��¼�߸����������