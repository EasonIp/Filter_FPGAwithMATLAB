��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�P	����6��<����`V:�Ufv#�խ����!��O���$�opB����n����\5��<`dQ!1O�VK3.u��q�Fy��g|l�RQ̒�jv�
3�-U����X�A���G@�B΄6������{$:@�>��*(E��¶�����u(�,&�P9��3DH�c߈�sAzx�k����� ����/�kp��;ɪ�}n�LrU�ZH���g��0��X�Xe��^j�����Mٱ��j7E	�V�tzK`pB�i#�u���V^�р^K3��AM�d`�����g�)�Y�����[IЋF;D�X�%8�y	:���#Ѳ���Q0K[>#���+]�nԳxD��J�CsjK��3=����@j�=B�"Hl"M��|)bf��j3�"g�}� t�E#����47��Q�ߴ�RI�Q�.ԛ�.-h�����8q�|�T�6s۰�R�$a!���oͩ�%�qb� �掊�����}��6
���H�}٬��
�XJ�I0QoQ�LL�4$m%,f�ȹ�O>��{��k�Ɍ��Մ�g��>U�o(�3���2��L?ZF������H@_}�G;�2 �-Y(��������k�\���x��kկw3Sl͑M�G�~'D�!�-곓0Ki�V �d��x�>o�EW���BW��j�7�h8�E�鄐-��L[:�R1���G���(\s���_};��P�'�>�^��(�IW�$\,"�{��5A�z{B�n�}���� �nh���؅8W�Mln����ʛp-�N=g�7�r�7W��n!\���n�b�6;�n�G�H��I�7�X3'�;�Y� ��b��)�.k�������(�2�/Z1�lO�<7'6H�Py@v���R������!�cGB悸׎`X��pb�����S�+VJi����e��`C0�d4|ܺ�| ��6��rT�&T�K4�}�'�����~�ӈ��H����4ժ���@m#��	���c°#�z��R��_��[��яև�T�� r=� AGo�O��rLs�u��?鮥�$�c�V�S���j�H,����i/ۚ�ϰ���7�i��8U�Z�5����,R��w1�0�xG��W��n��
iu���!��˓k8X���^�<�v8`���.�]qA���SLk1�8�S?)�K��ųz6^�ED'VI	��Du�Z��q,X�cpkG���b"�s�돽��u��n]��U>��!�;|���(�n�ؖ��P^o_oJf�X�+�<Wl�ѷj�6�"Q������6����v��Q�&LnVPW����ͮZEs9�y ���ͮXG �X��_x;%�T���Ǣ���ÿ����#��b*��t�F�9��| ��sR���U�w�M	bd��y���>���`��hB1�TH�� B�@�S{ۈmI&�\�&+.��9�=l�QD�Y���V����t��	L���Ey_�m¨[lv�[���C])�6����V���WV�#M<�u��Bl��2�Y���[����s�?��U#�q�pRW����a�� fF]������
�֛zw�Χy�s�wt@^tWP�p�C�C�׻�;qL�l�Rs���x4���жe u��r��}�[�n�!�(Ɓ���=[S��ϔ�[����^���c���`uY3�^y͠���QH���+?d!M���.�<����v����p��$�A�D`%%@z5Ā�G��a�T��R�EF��#Q�Ta+�����6#e"|��H��W;����o���ti�{�@���ě�dBg�'�X�
)��'d�\gF�<	�olA��{Bb�T �"���>xoK4Z~�=���YB�|p��6|�Y�Vk@�l�m6�`����o� O��H�� áC�Y�X_a}$�5��<d-Á��X븵mS�m=����|w kYx�3�m^��"0�~��.�?zl����?2�,D?���κ�g�6;Z��z���.�6"�v�I���-��Ԋ_�;�T�̶�:rؒk���^P�6!y�u1O���t��k[���k�FS�#Aި4�T����^��+�������>O��1,�'p�]W���F�}�V\�� Y��D�`6��8�O�gR#��9j'f/R~�̋L��ͧ�v��o!�&��.'�e�����e)|'��ǐuH����ϔm�)��J���Jv��";ܔIK ��}-ʹD���;}s&��X#o8�B�&`!�k�����pH�ͤ����7ў6o�� H�*��8��N�5�n�9�̓�/]v�0F:v�B�G�\�D�$5wD�>��ݾ�VBז��ͨ�T�'�珋/��?����/ڔ��*�+��o���ᜈ�#%��N�V�'3Ċ�3���t#�4؞�p$���A��2��
Ps����W]�n���P�r�H�t�t�qҥ�X����k�2���1�*t���� &>^�	6W��ɔ�Q���vj�W��Bb�eua�ȭ��h��!��xu��a�?��1����'���+-�R)�F�����|s�2����n��f��c�{��8��,!p�G���8����|���������t{c�Go<L�S/�`qٻ��7�o�/$TR܇B@��I<:������.C�	e�)��'B@���P�6J��D�6��o�+5���?+�_f�>s��j5�]!؄Ѕ������.�����)�J?Q��-e�R<��o��*s�Nv!����#��+{�念�5H������X�]�!8��~ߕ���?R�_�p��J�*r�� %��E7���~��$1b��>8��\O4x�?>0vO3,��<D@%��aum�'[I9&���{��S�}f��C�RJ�}��k0sS��N\<(C���e|��xg}��,Ao�d�E�>P�2�Qu���Ni>F�m"�qg��ּf��Ԙ2eg)�אi[M��$���X������էx������9��C*7	c0��6��,�z��˽`uA�@5��5�Y��d�N��2�����:����0��T4%�3A���!�xz�������C�7	����{cz$�[�S')��!_P[󀜹|q%���s]�6nӁ�"�!��A�:��=��tBD=@L�H�E=�Z-�p�om"勆��XN��o	|5Z�azHE�n�H%�c��9M��s3�l���W�8kR�Җ���f@�;�_J�?�/��,i1��@�h,w�᧽�7���8��U�w�@<O�ok<�\��z��hӓ� �8BԲ�F����X"�V���E�\3[�B�@����ol��<�K�6ѤA�)�ѧ~�����a����3�����֟>�J�ދT<��)��=P
����Dj�H:�����CqS�T��n����S|����P3t����Y|�5�6�ˆ�M^�/k��!���˱h�R���b0s:_�҈��x)?M:q�|6s���gƳ�B��Ɯ4^Mب~xT'%6'N�0�o�=[ ��˄#r���Y��]�"�c:�~��Y�_I�H�Qp,�����~���<P���HU�9:<[���X�O����&?��U:N��"��^+�:�|����e�;=	۲��mI��	�&�L-^�9��GP�r�{Z?p�HQv���vJ�[�ri�_�[��>˂H��*���q�O]2�D���ߟB%[f橳"�O��[�-��PoN�+��=����uJ��j��?�눗L���f��2Ԍƅ��7�{�[d��#�ŷ�RDx���Q���c92/���xW�\��&��?<(
�"�P��,1����kTHiL#�~ !R���;�0�OFB�p&���`��kT�Ȋ?WB����j>�&4�Q���K��%I��y�|�����`,]��y �!r3���{
Ԅ[���v�_��˼��؋�^�q����G���`����OK�e��H#j,����5���ܓʽ2M]֫n�ҫU�N_�����u�-�����r�@5��$����؂-]ҥ��+S�?X8՜�Z�̕߷^�Vo:��Ku�8'$�h:�HŢ���S���uv���{��Y�if��ř�Ė�)�=�r#���M�S���b����|�
F�dT �x���$	 L��Õ�&��W��S�����TA�QQ��-��OI%��9�_�;�\��`�v��oS�ߢ}��q�E��4b��X�Wڄ¤���a&�n}�˳������p�Ψ߄{�Җ|�WI���Ќ�\�R�� ȴ�'�pL�[X��:�͝q�xK��-��G�W�M��U$2?f�16h��0ܢ���Gr��<n�Ϲ3��Z�ې"��|2߶j��Pr1s�tVlh�Ky����W�"�p�$�r�
��9d\�<rل۳�	��Re��2R�>q��4��K/M,�>�m#�c!�mCf��E��W�F5�2�W���,�&Y����`����`ꘉ��CQk?��d�n�8m�j+?{�>�A�JF�b���M<�6����J9�FD�Pࡱ�]�X�Ï��ut��N�q��ӤZ�w^@3;Z]���P|]v��������UG�\~��4��7���}������F�A�6Vw��2(�H{�<���=�Zγ����1���L{��hE"������Fcp3������ID38�|?��Ֆehuʣ"��J̼���z|�>zxI�;7������	cY�?JwA)RD3�b�N7vr��S�~������jP���;���vӨlҤ@�I�*+煖%ncXb&ޏj�4�%=t3�r���cPr��H��Q�7&��k�f/�)ҕ��h��l��'�b�}0]�L��l.E�W�e�2���䢤Р�zo6��9{�J��:�b�=�s������iI�Ջ�1Z]���5��^�I����?������67��^ҌPO�P
�k�	?0��x@���VgQ�����vz��c*�\4���n�;e��EŐ!"��Y(N�xa
W�ӕ}d��T����~��9�nh��[F6�N/|�W�m},���ܙ"�ȳ�w�#�Q^'T�C�Ԯ�T������_O�P���
�!ꯈ�"�Kh�N���2����t��6Kޕhg�Z�t������w3q������Ʀ �5L= &	��S&����{~�!R��<��K�����,/Kj�Tn���O�d�b��y���fRS�G���*v�����3��ω?���J Ue���?�9ߺ?�p��]7�������$����;X)m@�S��w.���15O�"�A����Y�b	b����q�6�o�"yk9�1���\�rRW�1�߃���O�h��7{�臱��r�f���|L��X`f
�Bdd�������� O��<�o��6�Pk��}��������yLv��K�ۃQ��1,���n'#034��8c��R+�p��!�:
D,"&r?�������(�@���m8��'a����/*!��0X�l	��	��EF���Q{�An.<��"�Fg�6J% 4�2�9�:�Őq���.Gy �FG�����6P�h��9�ڀ�,{��DI� �0\��r/�vQ̇�p{���R����*��&���\�Q'	O��)2�Eugi���u�� �@ �6˙�;�����G�-���߀��`�i *,&.
/�[�[%u�E��ދ	���Z�Ԓ��*,ނ h�����x��Ħ�����1C>|@Z>_�=*����590m����^,J��I�|�2{s>�I��S�S����ӖM&��ŝf�6��/�9�Ё}LS�$P�ª���rgf��XW~"��
n���:V�щ�I�]ި�wpI�cխ ��X�����~O����\��]Q��k���-�g�ʓ*i����s�.��_ˮ\��B򢅠ܴZ�TA/3e����O}`�����SσJ���r]� ��8�K��2�.\HM���(q������H<�?�x�uAPw�z�!7np��s������_j�w\���1�r�3�g?b��m��C0�S
��D�� �8�b?J��~%���s�n'�]��޶�(���4cL1R�6GI��o��I�.��c%;�P���Ӽ�-q�5t^Z�BT$f�Jk���f���� ��y.�Q#�& Tj���u�o��$�c��Ie�cr�҃r!$��Sv����졤�x�B�u����{<A��Į.�{�i�R�?����«�|c�5��8�,�yM`8#+I3���M6&�"\M�J/�b��c	w���I,4�l��O�V��
�V2�	�cW�w�}3<HF��|VĬ\~�4B��{%�D��]����)=$y�v�EL�_!թ�=[5w��ȱO�/A��(�>[����FSt��58��%�ʷy��`��og��F�O|mF��D��Ƴ