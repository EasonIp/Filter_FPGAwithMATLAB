��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$�ʆ�YVc؆y��2��/3�pĮ;ߴ�6g�6����a�QD5��ub�^a�q1�o���gB�MF2�'��)�59==�N��MOڸy� � �j�|���Zq4Fy�)�fˣ4���%���L��^b�@���6��of"?��"k��7�!rs�5�=�B�z��d��,C�Y�1KA��v��I�5�ޓ���w%�I������)�Ģ��&t���b?3rp�2Q����2�ǧ�U�f��7tҲ�][��Y�����Ě�OC�̙���)�4G�3U���4V*���S�G��yl��}���bq��D"XTW�W�����w��#5)��Q�m�^7,�t})�[��@�����|�&� �aPɾ�r��w~/�e�n9�a4'J|ߡ��,=�so��@3��K�$c��>�a�*Q��b�<Ft�
-V�=/����:g��UW<ȩyQ�`�����g����$B^?׮�o�9�#���&�M2g +��J>�*��Ҿ&�*�Q��t���~��Ģ	E�����������K�/�ͧk
C����ß�ީLd�)!T��n=@��M�"�W�i��Ϯ�:����i�6�v���T��%���&�r�}%�-��g���@B����7�¸6�ʽ+(�;�a������+6 C����ꕯ�`Ct�����O\up��{"�;���soY�\�eoV�����y�yzTŜ�W"��o&Y�z�߱t�KOA��� �5{&d�6m��?�q󖪂G�{Pi#i���	�鄨�?���l�j2���T�T�/����@1i$��w� ��g7�P�*�p:�6W	)S��.G�b����e�x���'���P㡚e��K��6��⻘��w1�0QeK.2���P�T��8;�n\KlUV#�j���;qX�L�~EK-I6��6�dW��ź���5��k$����-*��rX��A�[�9���}p�9�X��wz6�r����`�z�t�b�,5]�uaa�e�Œ�R�r��|�<�mJ`��R���r�V9k�G��B
��lQ��'��^O^Yd���u"R�o/���k��U]���| �����u�L1�gcS����(c|'�<F�.e�"���_|�/m
��;��׈F�P_t;l-�� �A��?��y�`���|��՜�L<L�W&���Fu����@% ����XN�ڇ���������W:�<I��w��|��\�.&�ёXL>��k�zK�=�����F�8��N�~�;�n�Ln�C�����\b����?x-R.����No�vx��]���X��y��q��0@�G>��:�ë���O~�����
e�*T�a�F¼�z�QZ,�+FR���O����]]�C���G��E��;��TWey��H\�����_N5[i���˩c��(.60��A,���`����.����\+IuWR\��~TGV��_,���>�"�NQ��%�1�x�qz��q���C�i@%���n�0���q�9�팣��T;l%�:'�L!�yw��RV5�_ֆ~�upYl4�Q��8����}�����71rl�Y�ۦx��k��l0ɁdqaM/��zD%��p5ʻC�_ڸט���/�]ɐz��RlHIq�<`�s��E�'���Ց@��\��������+�����|��p�0�+ �o��{�c-ܖvY�2��g�[ٲ���x���T�$�?��ѓé� �Oi��$��QԌ���#�9�l�9 ����V��&1�?�����dM�v�^�R�3]&�%���CǁF�W��5��ɬ��lɥ�u�(��S����ّ�%'v���.C+I�԰V�A�qè^ѯq*XYa�iPy��^��������>�g>լJ@���~�����������=L���J�r᠄�.(t��Ϩ��h�/�-�����-s�7vL����EMLl���T���i�"Cp7�����<�ym�6F����a�s�v����k��9g]��{�#u$:���2���V^{=��!D�#3:�>���S�N^M�t
�ډZ����Tm�b�kZ��7SR|�OVa�HZtf9��Ǵ�om2���z3ek����^X�<�-��}ju�!7!a`l�`��\��� ����f}w�L��6�-o>\0@3w�g�*h�� R�e��t���_���D�%�����?d��wzJ��O��1�D �����LSwN��8�~�B^3�:�͹�g���c�<���`��F��K/� '����K�[.�Ѕ/Eo�МD\z��2�vc: 9i(d�p�ڀ\��wؖ?�1H��4o_�v};���2����]����H��q���>k����Kq�H�>�]�o,�z�!�H$��4%��zn�f����cJ�|���K�a�jqZ����#���P�
T�m=�j�`�� �gHo���,���fǔ�]��J�2@	;��ϬSd޵�9%��~�;�%9��DD�T��'bu���d|�-���Ҋ�QD>��=mm�vl��1�r������.����e���(Cg.3{~�ݔ\�r�}���]�k�AuS�x|��=���}�&��~ʷ��|!��!0���|W��wrjʮ虊��IԸ��T��M9��(P�Z8'7�Uh(sf�S����c���I�3{{�koӻ,�$w����:W��4� ��9#�B�墕�۷5�l߇�\����}��%�`�2�9@�WO�V�׽�����40�DiehYH8����@?���13T�qS�V(z �%i����/���/��qG)���M&��q�[=9����f:.���;��-�v�L�{ǚ�l_�̈�fS�xoO���P��Z�%M���8;���S� ��	���e��Q�v�/n�fHef��~�k���5�3U��!�G�2d��"^��ŷ�L����,�$Q_K&^�[����	�d�m�p���H�"D-ܮ��5i
;��>���wH8�Ov_]���p���z��v2 2��[��a��w�E�r��У������
>N�Qj�b���^?ȶ/S^@�Y���U��@�wR^!��_��*)�d�ܪ��?�a���;���-ٟN����i���{�B�Ӌ �֪�$���8�#�@����Sg��K:ܹ�5d0�����4ԀT�g3:T���\�^���T�z���B!�;D�`hh���ydE؇r��mK��ɏ���V���ٽx"�U�N���g[��Vh%�V!	�$o��.t��GM����#ҵl8�f����c
E��\�cu��x�mY��t1�Ug�����.��1�m�n^�x�6��V�ݠ�xPD�C��b��D��V�w��T�{���BG��W����T��'��<���Lc+���� =Fd����R���Y:x��"�ވ2u���P��$�����u��R�,��c��̞[_e%?�β��*�X�]�;
�;{0)��V�b�����@����	���M�vo-16π��Ѯ��aӵ�q����_�M�i��β�9Uy�w9�=��!K�F �6F�?C~�pI\��?���Q)��l?o�!��p�L�'y8y;���C�f�+k^k��_rH�a�NT+���F�}�;�J>n��	��3K#-�˪*gX�$���)�$-�\6P��aԼ��ab�a�Xo?C,�:���(�W������Yf��0TT��9`�ö�M�L���hvP>JP0��Dw�\��R�+��F����Z�� ,��:J�MF!S5�DY��m#ò�W)4���k0<�:u��P,���}��Fx0�$���9G�����H�A*���(1WZQ��<�dZj6䮂p��N����8�ʤ̣�	i ����ov�"
���}�[��]m�l�I�h63j���dO����c �?�zt���:�ܴ�R%�8˅_���h��*�Uf|3*�g�عFf@W�L�j��ʸ0nE��_8½�-�/XMx��^4[�<CqE��?���U���[��N�xj }R�.��7��"�6���AT%��hjȫ6R��!_3�&�+���.�HUb��t:���Q�;fm�N�j
�>`��MB֓7�0B^kؿRѵ�8���i�&"�q1h@{�Ҷ��-n9�X�ƴ��8��I�]'喏�JH+I��b,���SK��lcA�cv�PH.���\�+�N��M���/[��	j��4�?���
|1^zEx�Kģ��q]�0�h
i:뇪��9�q4\����Z���ziL�vg[���#�ʥ�f�@�󒃏?/c�gBHD>\jW�괴�j���1MM��ų���5a�*r}���'�PdJ��O8j�O�eh1m�L�x���[2HS�VTj�m��b��7Dvٳ!��E� �y�I�tP�$.ʊ���[P\j}�
��Ϧ+ t�v�;5����s4��޴��J��e�4�Nm��c`ʝv#��}�@x��$tC(�x�Y`V�ʅo�kXv,l����<,��\�#��OY:�]��t��.��'==�;�s�?� �+7�ܵS%����e�'��͸4��\�e��!���������,��1Mcn��ݔq��Q�Hv�GYg�E�0��[�K�;��6elY�����3x�M��7l^��'��@����ia�1���%�����̕/4�'��,�.�_1��z	e��L8K�|��+�eɸ�4��U�N����[g�D�M�U��=aӾ���4�֭���H�*�M0�n��<�:����a�OAӦ&\�X}1�4!(�4������­����+�6�~Z�c_�Vf��z/��C �qL�e/�Qo�M�}���4�b��뙓�����ܪ�E�[�c��
3!w��V9�45�+�dv�-謓F��v�>�!.|�Jt���:�l}9�����'����q�F;+:׮��hI��V|1_�V�r)�'��?�5H��<�f��ɦ� ��~5C�Y@�!��4r��Q�K^,�o��n�;h?�0�5�Y35��}Ϣ�Yܪ8n��ɹc?�V� N��rie��@�2���uIL�^LE��͗��A��Z�#Ȅ�GH�S�Fi��2��2z->���.>�g!}	��7����e%w�)9Xn�<J��A�FB��Ԧ��g�Z�疚l�'h�=��Ew��vd(���ɲ�� ���H~a�iL��J�(�2�!�)o��ٵ��Ӱ!c�����[�6"Ԧ�fiSulB%�y��� 6.�Z-��i�s������O���{��/|�ެ��VyTQ�wp�G���;�4.�>:0B���_T0�k�Vgݛ�$�:�1�����+>���bH��}�c;��T7����4��E�~VD�O���gõ�3��&�V���lO����:�p�\�Q�G���g��IhjTn���挌?�A��9:�y�m��S6��n=��n�xa)8�[rRL{e���_[������J�E�<pQ5�z�ҵ�����k�p���y��Ϻ��m�2��3�,��W!O(����Ԣ��8�BnJ�Gu�	Ri�: 'Ć�_�#����M�����D�.#֢��h�?X���}B��~h'��F#g%'Tmhd�7ˋڞYP&�<�0�'���Ow�S�
��]�v$5�"������i]r`������~JӖ"7!ݿ�8&;��"��Ήt���5�+y�p�aGdN�([��~�TvV�6|�j�8�{V���++�����j
�ѡ���<����+H�癙��W���4�	��<�Q�ugǧ^ON���1+���kT�c�/�ῠ�aݷ�N�����W�	kM��������(�nQv��1��Ug] ?/��r:�����c�ɿ�7���~��u��[a�~��AO�K�E�Z��^5�7����\q�b��#�������zi	�9�����N)�\��X�7�˗;��p���є�Πt��̑I#����[�%�_du4��V�ܘ(�k�H�+�H����:�v{��Q�>��Q�؏|�������%�5
�[��6�a�:F�Mv����_�+�*�L'���֎�@:q��m�m��TzJ:OEE�)9w�b�Pٌ�_���������N���]�Wgm�(�\ތ3��C�Ϊ���?��(��ɖj@�FX�h�!p(0NځB�9Q̪��\��`�Ra��"׃ӳ��	�g���g���c�h�c�m��ʿȯX�$��%�-j�g�W&��\N�mD��j��hBqPl��o��/�d�&�Bn5����Ӫ��*Pj
tӞ�����V�:}�v�����4٨c~�j-27���%:�l��mYl�\�˗ޓD�~�s�0�D���%��l�M��s�$ȪJ3=�dt W6�*�i]�mx"��U���}C]�XVz%��=�M��gy?t���T���z��N�c� �e�vd��7����=<=�d�s�l{^�o��>�3�=c YJ:g��{�`R�"��ԕ�->C T"������;��<1[���s��w��"܁w����r���Q�-<�
��E�3�^�^,�ȳ2ܲ��~	�l�@C ��{�L�k�R��Х�nʫ�[d�K�z0�Y�NE�nej���E���1��������/��ϴ�V	���08Q�����[ki�RQLY�>�������#��9�#�G���������g@��~!O�@��q�DE3h����Y����Ǜ�vZdf�0z��&94"Р���7��)�F)De��ʔ�w(>[�[�fU/��']��}�>�җ����o�(���!/���N���4I�!�!���@jNLQ>���f�Ja^����PA�$q�,zW%C�AHI�&>bT�[v��֤IYg�����=��=Md���*�j�>�" �(�.^��ͧ4D��z\;�ZV��o�.��w*J�9�쭞���h�,�,3'�{�U��WN�v�D��.(��7F�m½�:����v�<] ����Ww�o8ه�38�Fw�Q�f`k�}�h�aO ��W���Z4?�����pS+~D�b�w%*0����C�`g�+�㸘]��ɑ�Z����D���������}�5��f��E�-�S9��K+����Z��?���\��M���&f�I0`&#y�7V��8��&���S�W��:;T��"��#L��Y����>nҕ�}i�ε՚J �A�2V}*�q5<�&��b�-����nA�j|P\.��,� �*�*�M�k"���ks�fN��A�\�. 䟻�tHN�Z0�EK��1�#e�Ria0⿎�����_�WpP�퍲�� ڇ�X��m�?��Eg���ͣ��� ʁ���X2���m�H���x��lFGZ=�O#��91C��vk�^
B����Ꜿ0A*�7�-E�� hA�{d�i��7��ܼ>���)���5А��(l�P��oU�(>���e�kF������=��HP�i���[}C~�{q���X���Yi%�s�xG�u
�����>o<Z�I"�v�w-C�CSՍL4���T_�E�uٰ�U��$K�偃�v%��G7/3I�ct	�!��7�c�!"5�a�G��Ϛ{t��zR�b�d�����$S�q�jt��"<;�!�ق�|��� �j�fs��M�	X�קf#1��3yС$�]�'Ә+��RC�'v˝0����i�Ҫ>�����������&4kb���u[]�7-��T��p�C��N]����B{|�>w#X"7X�\�������"����m�����m��b���������8�����n�>�mx�*��
��ݰ��A@�.�F0�i�c�'�@�u�U�o"zm�^�M9G����]~*���b���t�+]?��;FG�����z�)�	m������#S��Ür���y��)#o�s��/�޲w���w���������ֳ#��°4l=��^7$��6lw��2PN?�p+�8�ܿI$1u����_�7��o���ؒ�P`7�r��=t� +��u���#�;��I/�ꗻ���q��w8�\8�{)M\4��0a��v$r ��ݿ�XFW�i�#ECA�!W������QG�/3�"�fnU�r�<D�r)��b�j/�����
茶�g5`D(�����jd;�	���2#����
	#��)Iy!��,<5>�$��׶_��O�E۾�+!f��b������ֈ<�����Y4�F�b~���x�'П�eN��@�ۄ��7�1��D��(�θ����+���Ϛ���g�g#0��C�Vw/�]Ղ}<�٥Y+�s��}���FE�h�r��,+�4��2<ښ�Mn0�|���[���#Z	5��Y���ב2�DdQn"����_"1D�Pq�[��5bf��@���7?p�}p�Ƽ$�e;:��	-J�;���h|�(ц#���z��.j���bm�G�>�S]�mtk�s[��bf:o��u��[�+yA�*�zH݄��nmg��)9"v��\�0[�%*��	�j��Y��/AH�a���M����jm?!��{�iJ膷���M�v �0)E���8�V*Us��iZ�����u� ���޹\Ӏ�)�G&��9���,��˕�δ٬|8#��~�Yʿ>�9����)���tn���B��_/I:ss���Yo�������uX�` ���˼	^�	�]��EȬ���C�SD��c78��[(��4��r����;\7��0Ṭ���ܹ(c�ۚ&v�I�K���$�nٲ:]�5TD9��LSF�����gDF��V6���	�
����~�c@;磄|�H����<��$��'8vCy�������Y
ڢ�S��S�QNt�,5RA��06p(�(i�N������Y'�$,������tԚy��;�z����\smp�, bV��(����/����%�8-ar�C?��zN21���#6��g�n�%s�3�u.�b��jjQA]ob��C� �4�.�nW+:��h��Y���x͔И�-�5Z�Yr?<�ec�[�Zʾ9� B*�Q�k!^P�B)�D`����˧�nÒ���E��~�ޫ��jl+�I5-噡t1�F�2�nZs��>JV{k�K밫�j��g�"��at�+u���Z3S���؃�x��Q^����9�*㑇p�>>o��nw��
4η�[A����M��}��"�G�v��`^;�t�e�M�[�:�Y7�sp�&��$�qBF����7l��B�x�	�T̿Ce��`�4�?��;�4hI�M����ʤ��S�:HE��t���:�x�O�4n�7�����-��i P�g��u�ֽiL���ʹ��G~0^��&Y��pZ�O���,�!�'����V%����f�;�M8P���/-�0��#;������dm��̩���� ��m��
;p�q�#��ɢ��)2(R-�46},y���R��Y�G��"��/ۓ���`���!��P�h.[�y)�>4%��X�L&�W�%`�gX����-�Vc�pR�0�'C��C?r���4��;T��ҏ"�n�ꯤ��ۢ��.��?Y��X�v.�ZD.�:�8�M	`�o ^����n�Θ58�b㇩�ً�P�Z���� �x�ce���]�Ԝ�J�
`J^:��uy��ј/�4W̨U�q�|)���x�'�S%K�/�������K�ߩ(�p�Y�L�(�j�[�P��Q��,~����R�7)4[;pp��W��٫a�0��|X��~��V��3��Q��?�m�׺��8q;��C�����_�Ns��[�*��PY�9hSK�xv���i[�&	ãޭ0&8>�j�[����Ʉ��]&<�5���IQ��HtV����|���R��a�
I��z�gy
�!�ڪ���Һ0�U��Y
��ζ�fWq�}���y��.��Q��t�'��Fb�O�<R�8G&�W����&X|���J;ON�y^���>4��دDɨ`֊_.���4��Ed�mD��9�r0�Z�����_\���%(����z�_P	N���{��EZ�!��s�lmVl�|e(�Җ�¡3��>|7(8k��� JB�b~�]�I�z��~����MZ�F">��U�ٚ�<��Νi�ٍN�]7OX/��oYVt�j��̰k��%��8��{e��������*��o�)�u� �&�g��e�lks�Ig>�R�X�� %a5���w�<X��b$b�k=/�ѳ#n �����b���P�R��sř��r�R�M<���ZOY+�z��Q���/G�,�[��j �:`�`f��9d�
^�k>��(�� n�E����x9U��
V�|."F)W�����;H�>�(��!V�,��OH�7�&� �K��w/�i4B}�A�W�s2ݥ�v��/ˑN��u7�&~���YW�o�1�Ӥ(�#�S� ���GX��`��������ՙ:�-<�w�`�d���Hҕ�,�61�ē:� l��ْTb1��DT�7e�ǁ�e޽�ddΑc�:5N7t��W̃�@�,�nz"���s�����c΅�_H�	*\3Ӽ����&�_=��a:�_��u�k`z�ǟ�N"R�4�� �c"�e��T�F�F(�M�Z78���d2�:��+�rGڹ`���&y*��9V�h�mG*�)=�K�Y>�ڤa<��V[���e@a����C���M\��f������B���Ͷi���I�/[&���S~!%?0��m����9{=��ļ@�,��ͿZ�5��i*VԛPW�~׻z���<o+ ��>�����.�����5v��)V0�y1Gr��~�a)˔Y݂7�^�˪�,���u���4���)�M��@&Ɩ����:���8�@h�B�ϻ����|����Uq"T���嘼\���Ҕ	��m�/���~8 ��� @�������0lP>u@q	�+�����?l�[�s)��v�AtC��Yu�1�b��ARw�9�!s~�AM]&��O��B�#Z6���bj��e��u��������P���;˼m��(Q�߬"���n�ēP]>��!��)F3S��5�c#���2����I�,~��=ъ؟�'{�8%�6H=�׌=sU�P,�!�:᛽��X��W����R6��K�oP�/oω��Fk�A�miQ ���u�9V�o�������t�n��q�2�YG紜��G{�/M�/k��o���9���* 6�������f���Wv��7t��`���2���pl��Y�1v�Mz����]?5*��?�D�Yf��
�n���0�a1�b!'?�?��Pl��M�� �5�<=�����<A��M�2���1��i�����.g��-z�9��������2֦<�����`�(g8�����+�4�a��A�X�d:�����E�-Ǽ���fl�[�S^K�2=���sθ����ȋ� ��r/��ZOW?x�����2���{3��4�F��)ua��~αI�aoj!K~R+����h��+Ī ���W0�PsU����r�.�(��Ʒ�gH���Vl���k��A��,�H'_'���猰R+�U(��!�D�l)�R=�����.��� �G�
%8uҥr��V�@��B
l����a	�()��
�F#�>y���	W(��V'+Ew�FW
r��Ha6NE{�lECe]a�Fw9��FX�bu�RI�����h(��V��Z��j$�n����#��{�)��]�v�~�5$��]ɹ��f�`5:��S��DD��=�����~�po��-���|��]���,���u�4�@�w��޽<S�\�W�m���p�;�����9� 	�L�]̫,�w�e̸͝�qC��-�Λ2P	�du��P���:�YZ~<��SXr��W�`�&-��~�ۀ���_*j���O4Ϧ�>���������1������>�N��_u$�������VqRv���䆬T�M��]��K�?C_�n$<.!ԇ�@DU�xZu����d��,�c,`��O�@a�ֹ�x<�UxD��LO�o��_�-9���[��7��ukB)ju���Ϙ3Z�%#촞�ֶ�p.G�!�� ���&��y�4f2��KOJ5.���$�#NC�	I��Q�wװ�l'i�ʺ�q�����F�|��<ˊ4{z�m���5��6�y�{�����[�j���=޽����؈<e&=��I,�)��~���P�M]�6�^�6�D�&�tkkS��)���XªVt��]]���ǎ�P��[AE��F���؂��P�v�l���7mi%�RB��CN&�����/iѣ�	@��O�3?����&��$�.Ћ#ڞ�)(1 �}��w��"� ���́��r5��*^^��%��/y�;�d�w�*��}#m�'Jw\lQ;@��̺��2�~�6p��m{��K�$�BE+oCD�s�Um�-=K�)�������j�=�ETUq
�����C�E�[h��� U�N E,�M6C�3����q�h! �0Q�H��v���Ĵ1)*
�� ,��x��A�Af���w���x��BYW�`AQ�H��q?���K}��Rr3�MsU�%c�ﰈn��E�����H/D/���$�T#�KO;;N�����kX���U�Zwh�ٿ �`�Z�O���ț�N�J,��r`��|Ʃ��"�8^;ɟ��ӗ�T#��d�Sx�	��!,'d��	��ф`��o�6�)�%1�j���w�{��Gb;��E-U��� ֲI/�@�78��o1�6G����?�A�s6�$#�� �=G�e�Vj�==��@,4��9�??_�Y�?0"�KN��_!O�T.��51\�k"<�A�����2��_(��ڌ'�"H��$�2�U��j�l�C��㖡���iT[��|�y�B�,�HQH��QG����A
��-_#~�`��'j�)��^��2���y��W�ޚ�a�*\�Y�O r��U{}g���]�8� ��<B8���2���(��օ�ʮ�f�L��1Xf����a��hJ���zM���0�UZoiL����O�,�F��79�K�Eg�/�t-�F@u�N=��B^B�4A���)��
�3�ȑ�$�:��+MI\��a�L��ѓ��ԃr�~��HK���_�B��ZdX��@,K������e����L��a3�*� 
1�J���G1�/�L��l�:��'�g(���f��g��b/�Ȏ����� �Dث9m:�ݐ�{k�M����*>L&�|�^g��;�XT�%f�o\7��v�@��E~��5!�u���u.�2�uC\+eZ � !�xt�޺����(�GvY@�}�a�u�p�i��L�P�ևZ<��c�W6�2Q5r)���_A���u'��a'3~��g�6։T{k[�/A��ڊFy��C��L� |mP*�H�{߹��Ι����!K� Ϭ�?c��IPO�ecH�=�U0�	�\����1�b+��4Xk�A9�I�ڼp8���k�`IǙp�i��n�r?����7��tHx��me�Id=�}�����B �S�ZR�?I{r)3������C��~�&�1��������F01�� !kw�k�؇���18эϥ/�c�01��C�f�����M$r����@�T۬E!}lK�M	F��hb�Z��p�Pǆ1�`�I���)��]V�����CY�h�M��Ԭ�P��dd�/�]��hĦI�A�A��4��V�%�,g<�C��  �s�~Flk��k��6�#��ɳ,����Y�1��i�7�n�$�xEV���FǸ�h)����d�{�Z4�w	\
Lz7Rۥ@-z�;�^���{w�8���̰V؁y�jϱ�����������f�.9m�8�r�͠G=���^di,�CW�0��=�D��/���� gC6�ِ$Pd���A'Z�vYW@D�@pZ�{[�~�_|�c�����cWW�B�9��G	�P�y5R����?��j�����B�|���'�h��H�˄/  ��	�1���:p ��ݳQAх
_�C\	��c�	N��@�fP�rz�xf�N�W�v�ExĤ䅊����m�t(N@۪v�!�����1B���w��e'���^ 8��t��(��S(����� ������X)<����� �]#���y��W��wjFÝN�9𙨵���qx&WN���*[^��Go/����:�ptA�>/Z��2N��K��p�h���(����p����w�7�o���X��c�v.e�;d�J&�&�g�!r겝<o3��x6�߂�̝������6�Y��DWRY��n���4t�-��V
��4q�yK�!)�p���K�7�p֞�w-	d���^��.Ɉ؃l��2J�f��$m��41Q
�|-�q̰@���I���X����q�#�[=����dS�+�&D�߫�G=��@n��^y�����dՂ��j�*�lL���ֿvQ!7����g	 cn`g�u4bO�=�0�F$6�� ���4�is�6PӲ7�a G�h���p5$��X�z�Apvx�cX�}q�m��D���C���������a���`���P�7{�æp�S1#������ �)túp�j]G���a�e�z�eV�!��Z_Cy;|�����ɏ�����' u�iO�]���8|��j���\'�\�8�!0�:a���l �U���Ti�F�6f���a�-C9SL��4����ل�A�d�c�k"a���P�̩<�Mp�kL�����N��.w������kk8y[Uz;�.�����{sQC���7��0S{V��1���u\�SŰ�g��Dz�_G�
g<�1@:�z���v^�p�U����>C�K��}��r<K������@��F� �1��A�? �6,����\Vh���f莟)>t�}Ow5`j%"K��@%�6�v� ������5�R1r�b��U$Vۜ��<z��b�I��2��xGV +4�Z�ׄT����2&���y�C�{�f�ƫ����LR�x�y�ґԈ�]��%��@Wbd��@�,��e����dʏ$/5-����/?	YD 8ّ�nM�mh jw�V9�0HL>e���"9(��c����t�j�GiQ終.Fvb�b 7z���p�~�0vZ��i��u(m[�����@⇆w3�Y���г>���+����T��^�c�~[�CطmvnY��F�X�������t�V���[����/����������KPce1�dD�s�Z��(���ɍSi,��9� �6����������I��Me�M�tKKw��R�V�JC���c1�n�����+�l�5�|jXϠxE���+"�*���Ц3ي��ie���_60��C������s��_&x��u�1�<����Q�l���-97�Υ��&˭�����U�FvB�����
?z�!+��K���ˋ�t��:���	�2{�aN(���%�ӌv����������~ ����p�ng|�
FAO�N+1�r��D7W5��˜ͼO�X����5 ���+]s�٨Gqt/q.JM_8:�y�R3�>��"jϧ���ﳻ��r���H`��v��IQZ�v�Z���u�B���-�)��`#pH
t��ţ���N�f~��-��MZ �H��Xӭ'4��q��AL�(>Lמ���M�����#��K[�^r��;7ӻ޼}BbH�Q 9B���d�gd���o�3���X����|Tc���0�3�]/�"1gxC�c������g??&�wX�C�_�u������*0J ���>0�*9N��39kŨ\1�݌�����Mm�KY���8�kk��$(W�*5��7Yg:���~������G�2�/HKu�8q�#��J묤C���/�R���� ��Ue��b��Re��o�G�]v�@�߼(�eԜ��7 r�@���{��q!�J��<�u�Y�q�Bѡ�x��?Cs��#�!$1����Uf�C�h%r֏J\�q.��o���: �I3g^��W"W(�4ȉ���>���陎1��D X#�U�>�*r�n� ���.5��g����0�J��_�c7�\����b����W�-7F������r��7�Y�S"l�9~�Ʒ���R���rZ��!��2J�w���g�;[����4П?6�[`yC����P�J�=���i��^%�B����Rĸ�.b�'�^��|�6�&�����a�!������*]�%uHc=�@����`p�HC�"ĚFΔ�$�V
<�A��'
)�P���]Q�.)�u�����Ο^��~,{�ؓA�	��153tr`�y��|��o��$tLl@�ҡ�Ch��/!��Rn<މ���}@+��BtsA�7F]�X�	=�T -Q7�0�&4s��
x�k &�B���P3A�'\M]��v�nm�-���(i6������fUM���N���l�|�����Ǉ�	�q��6^A��/v�d����0O�����!�ў~�Md�E�~�=�؃�ǳ�`S�B�k)�n�d�׿�{ 펺/�e�a� �o��.V0��S�P\2h<�׀|<b��YJW��A��6Ɫ|�c���"�t~�T�`e��V������6�5�e�N�}�-X"�Me6K�̗�M��������3>�I��s�a�=�\��g�C�m���ARQyu�m"��kQ��`��La@ik��*Ki�+V���<�U|Q���eW|F���
�{����4h�ڰ�C�9Zk�����
�W��g#�)R��_;�D�xw�>�j:)�;�	Ŝn���[u���n����O�{�X![ηev.�}��c*�_�Ѭ�� ��E�%�/L'J�py���(8���Y㙈�ӌSc��>;��m���>��u����77��X)���!1(^�=π���8>Iރ�מ��5�n�Y��b-0�� ��^��GW���&��9q&$�A(&��Lȯ�PS��α���3r<���<���Y��B�E���l���uv��C�q0����I.�(�a5� �U��} ��K����8������
T���g�����y/+]�(}��/p�<�z�% �_� �=,��Eq��[%G>p��s�2��`_��� �Zd�VH�~*�W�<�7!mP}ƙ�G�:羉�M�p�K�T�20�=��@IE�/��<^vt�>���
�"�Ή��С;< �؉�W["�d���S|�^
Ef�8ٷ�SͲ� ��(��K����y!�2�����$�R�H��t�@o�����#�=�z� W�ۋ'SY?��ԩR���>(�_���(\?1)6��F���!?� �`�B� ��̀�$�6^�v�#<���-[d�$|��7H��VЕ|"��7� 
\��X)h�R��uş�0��&>�L��2�IJ�NP�6���+�'shF���8�y}�.�yD���t�#ͮ:����#'��]��iU���e$�,k9 �A �ب���"S�K)�Q�j�}4m��-����e�����X��Ӧ�hsct�là%�",�Ɣ���k�.�ܵ�����&�l�V"9_�>�|@�̷㪷�}�pRn�����R�����)�n�8m#�1)Z��nOVp��LM�w^��O�O�?�Vθ�o2%��9+ D(� ��w�y�ĚV�j"7E�Qf-RV_6@��H�W�5�������x��5EN������D�T�"�t
�t�C@�'$+��*�i�r�� �d��ѥӠl	�p�X�z@�����tn�P�X��=�K��H�E�n�vҵ�n���W�Zz�ǯ��Mv}X�s���uw���]`�R��Pcݮ;8�oB�L��W�Ii��������^Xɰ5������:��G`�Z[i1���>��y�Φ��'puj����^Y�#	������_CAo�=�r�GP����.�#�I���4�|V.�-ۂ6F.2��щ�bCk�*���j�/��9�ȳ���}U�Lx��T��cC1�atFw�r�*晿9�p�q/�Џ��JVQ$��2L=�X̓��(O��Ygomx��R`+h	~�u�us���D��ڣ�/�@|I>4g{�9ޅ�a'�y>�P,}�\P �5�POH9�c�sӦ��$^2@��V�`��ϑ��]����A���[���wU��ȅ�0�
*?��IJЙ�[�����LM�d���}��[�Ea��A\�*z��,�B#��yP��������he�\���Oh�4뚼�8u����9��ɷ�pL��\L�_��nB\��_ޒ��9pAN8�kQ�m&WG�����nX���"1��j*�e�*s���Qn��H��ӑ�L1 ���V0�{T�TS+��L�~
#����1��ƙo5�$�;�:�`�����얓T=X�yf�H��pտ��c��x%��J6�𼏇q6���o������r ק�Hb�؁�h�7�7B���Go�E�ʉ|H-��"�7K~����w9&#��
=x�\���#_:{��/7�q�"uؑA���,w97O�e�޷��D�g���Ӷ�eX/��[��"�3ٿ�;m�;�n�N�4�
�^����_̘���cfs��2��N�*Pn�.�">�߉���ў^�ї(�B�G�W���q�y�|X-�ȁ�!�2��yC���m�Q�Vd�8��%44
��۪�m"�,��L�P�;@��"�Ixō\���IqdSE����m�PVˍ��޿��������}�K:��f8��%m����H?B�#9���veV��9����5x��@���� c�y)����7ďc���:l4�mF]�~� �p퍒�Qb膒U�{aR��_�q�Ȝl���?G��Q	�˸��(�T0@�}�t���+�,T�	��>�&�V/�����82�ې}��������j�t�� ��P<t{���<xd�Q=}㇟��^W�K�I�<U�0%�E�fy�0�<�?l
O{h�.gh�78)��|ˊ��>q�s'��t:!}Zߐ��&���o:J��(�w�!�3_�uü�3Ɛ@��@[�����(U%��}$���j���۠F�ze1t���t�/�o-��\1��C>�N�<���}��������_������ ��%�}b�ú�V��O��T�E��2�����t�d;.��A�0"Y�]K��ꖌKd2��\�fvgݘ�:��ߛ��g7oX���7�h�i8-�J��S�K�;��v,�֏�uNЍ`΋߹�XW0(2��.�e����o~a�A�5ɪ��p��n�=����/����b�M+�����	"=������^!@�4|=�hU��"ǆ�$!A�Ss>?	�˽�BCP7t��V+7�2���F��>��t�z����!(+�hs��D^}`GK�=p�m{��jƖV�u*ғ�*�Ta��P ��¤em�_�=�IR��ߺ,	]V���U��W$u�Zn��2�;?�_h���kj7��s��k�g�k�WJ����@Q��G�;Ǆ��CP��d=�(����r����BF�k����(M�R����@ASx�l�]fR�|7�x@���*��i|���ˉ��S99\�l��	�zp���6��kM�Xf�3GÖ�����D�'o�3w���C���8 '�d[�Z��b8:�%{�,��C\�(�*�\l�0�7�m&���m]����a��^&$mG�$H�Ŝ9�%P��C�@Ηn��[���{2y���M�q�����=Pӂ�/��J����ʝ�s8p9ZX^��ex��g���X��G���ܗS&���7#����d��b�ʶ}����B�!�y�{@�ފA2_�e^���C����#a�1U,]�L��C�E*�]���i�D�L?�2�v�Dn�*A�J̯+�LJ~��	EG،�3x�s�ݎ��q�\�d���ǞV�)m�t9���f�9���VFM���I4r؀(��%爭�R��N�|N�LK��7k�����qT��]�廧�@��_Mx�F��� �4IW�T8���NK;J1�2����`w��~��"��k��.O�E�!+y����Jh��}@\���J�.�?6����<ծl����G��:¨"<;�旡��й��ώ%8 ���ʛ��d>:�_1r՘�M���CFIr��ޛ�?�����C���l/*H��%�0J[rLYa� �7��u�t���k�����E;S$ɒ��̢������1|���@3��`*���Qxf��OS(	iAi�錢pwEh���v���wm��j_*�xQ�^$��^k28�����#n��S��]�b&�Ѩ� ��Wc������������иD���R�^Ӳ��R�q4)�֏E�y�t0m��Q	��tX�3�s��.�������vm}�a)���v����c�h~$��`z���7d�����,���ۿ��Mj:��!�g)j�G�Zb}%�A�Nr�j�$�Ox4ś����8,yٙfˢbHV���;{(�_e�[CwR'�����:+Y.@UL*���r���6v�!g8cZd��|Dg?��]���\��"���nk�y�,Zx3mH�O%�zL�m	J��ۇ��~�o��L\D{�Q�3�5fq
N,ۗ ��
ۑ�=�l�ĭ��]��ZrX6x�KjE�m�.��(^b���Ծ:�mC�vBU&�(�r�8:��ip?����P�b����Ճ. ��Ѝ.s�7j
������|[m=�6y��,s�QgG�h�rgHɄ�3O��s5aeɼ��h�P��l.�,L��U	��g�)��
fm.�D��߫�&�e��7�������'�z�g!x<�zӓX	T�E��E��ۀ��oG���2a.;�6h�!"%S���R�d$�ǆvWW<b<�/MZ�C@�Cƕ�нSG��
o2{�۪*6U�R�1��B1o�*^TЇ��I3�o������N�J �	�Z�ĥw �A�5v�.��>����~"�����+��` lB�,�"N��Eq�����ٹN�i��A��_S�~7A0�|�\�+mv&�w�!	e�u<�~ۓ��Lz	ǹ�j9W�{��gO�j����OL�F�X��B�Ǆ@��p�fkmc3|�]!Cڇ/�@sX��E���͖t(�P�jf�N�/�����y�y*�\�{���?�ڍ]�˔�c)���hO��B��{F��&�%Zr��m��n���	B�r~�>�գ��f�����P/��5�{�4�#��'l�^D��oH��	8V5��8�O3#���i��(��J�ˣ�HS�a,�����Sn#(Y	���>T^i\]�{0t�~��xv+ёu�M��j��SO
1�坚Q�JM��}���s�UI�	`�ZF�[�#v:@X��ɼP���5$�D���?� ����z�Ν���%�����OX�#_	,&a�MP�#߰&��m�i�kB�ˮx�6E+����=�ʎ���y����ȗ�=d�&]��\���B�w��K�H�eQ�^��צ���^7K3O�[ZZ� �>�>Y���q#�y�H�|�iM;�*��%q��;��l�N�?��=`�@C�L|T����yj{�%�|��
��CrX�ҙ�m[CG��
!��4I�sJ�Zo	�g�n�	Ft�@�H$�$��1���JCƲ+����S���+�y�ꦶ�����gU%n��	�n�~���4�6`����6}�bN�暌B����fM�#ۼ���5`�2�[��b���rKN`�Xͥ��f��:TN����(̷^�}f�4H)ޤ5O�B���m�q^ag6�k(ڊ!PI�}�춌B<�����NG`��-Λl�j���V]�Z� @~��ߐW�Q��SH֦���ρ�)��M�MǹS��lCF�?��5|hK�A!xYB�������	�[C߮��F�(�ph����t�t�բ�IQt��~�VwZ���@��=����.�CqS�+;���5b~Q��E��k�:��k8�^KY��"�0E1��^��F�W����?��í �+)yj?_u@Y-b����g`��g�.��b�)2lۯ</�Z>V�Ŵ)�m\3�&>����S�	��A��(���W+<S����v�u'�5�+Y�^�w�7��9���ӡ8͖,~�Ծ��d&��5&��ժ�l^'өy�?\�9�?"�*G�Ѯ��}���j]C�W��bqEH��7ڿ���<�u�8H�!(����P\�厾�x�z����h�]�ۧΔ@�#_�j7A,i���~.�8�ɇ#�V1^��ձ#��f*,���%�`Czn����ס�¤`�^V����uQ]�g\����M�v-��
	LZ |"�ce��O�	�ɸ�i(���x��n�)DaD�[�J�&i�A�.#���[�&u4w|Φ*���u�F�WJ����ʡ%�?y�� x�_��=���<���*Y���fy� ��A���i�
	T\�E��_�e���-�D6�x�}b���Q������?�=��.�M0Rh����(���|����6�@�z�F;��ͮ�"?�uȾ�@��c{N���Z�S�Tk�'vW�o���_k��E9]�*h<��G��,��)wN1-�T<oZ޾)G՚')���
�2�ӧn���
�;F��h<��]�1��C5��U���Tͣ�+%��a����� �zѽ��5����x]����϶��0)�yޗܿ�ZJP�,b��,޻1_�p�&��@��*AOVՄ$I�y-�)g����ˀ�&<㈣���wQKb�a��>���4~��E4P,������~,W�^��.�ġ�qf�|)����$�Y�]�
K����\���]�ҡ��Ԥi�!f�>����1ūNou����f�Cö��V�QC_z�d��|��^R�1˱0N0z�	P���Z}�,���M��($u���%
i����ñ��K��
�i��2�����jPOs8�:S	J��%|�B�����A�2n���/y:���O!(z��C������YRM���fF=�����s��:*�k¤H�
|�w!ү������S��	A㺇�
�k���Zp;�
������%�<m��'0�8*���1	ƫӈ`h��%������EU��j�љ켓22[]#���>��_Mnf�E���gtU(3�c1,J�wul��0����ۜ,�O0PҞ��L��N1Ԡ.�*�(`9J�^cٕVaO�ʨI��TF�,���4-���={hi��սڢ���i�{ב�tS�/qv���0�����q������5���r)Sh�[˥�Q�
�m��g:��	����T��-�S��kd�֖�&�*K�9��"遘��o�8e��f7]��9B����H�Ŭ%����Kb�,�y�qx*�ʻ+3��4ں ��cA�~��YV�2��}��j!���X�"'T�ZK~_���U��;rC�Z0_�(��Up���[yZ#m�l	���u�`���`�c����~�l\Qs"���� D�C՘c�������sS\hP�N���񠐩��������0���\����`����GV=XK������w�h�ـ�[�~���;n�cX�Á~� k�U�Fz��	i|����j�m��7�)8/(��^1���fC��X�),��\��޷�|4�N�4�ČP`��] -�ΣI�Mr��Ðf�t���qgzn��c��6�]��qb���8��.���%c(�ƷaQK�ḥ�t�p3��0����V�[�tI5�[��T�6��ꁛ&A\�뛚��K>qѤ��ƀ��D��-��Z�"��ބ�t���zJ	�l��_/�*4�(���5����5"Y��������wѯEp+���#I�~!�.��Hj:Ъ�N��W�F��+��[}��̥mN ����=�v�t2����&*h���Z�KO�������#@�%�5��uƈ��jj%�M�2���~����kf=Ru�'B�T�T m�YP�bj* ���	���0�.�^y�ti������ڟAR똹�S&�B
"=Ʊ�vK��E
���u�%K�g���j�F�T\K�X-�}�4��
ө��ԗb��
>eN�q��?r֘����:�2���c��5��02�n��7xյLڨ\4P�t�0�����Zc�8��o�EU)�5������W�?��!]�=�%�o�D����s�jjԉ=�y���4M�̕�w��O��c����u?�M�(Rǘ�)���M?�-���R��*��?B���(��m%�Tt�ÉЫ�X� ��5ϙ�b�ϛLF\]��������� ����Q �M��;'�F�#�ޕ?�����
H���YTf�B���A?��\�ؽ�w��x�������f#��$�_@��<Ϡ��ż��{֒38'��C���39�)$V�y��7"�~[����c�O��M� ��s�K3q�4�V����s2Rǈ�j��L���>d�2(�#r*(�("={�a� ��J��'�j� i4��XP����4f�#�p���\��ם*����������F��T\7&���,��Sų��[����/����2�k��J��}r�X-�鉫�I=G	������n��ڈ����]]�⻬���r}�&�Ik�7K�m="��	H( n�Z�ۣq�wEo'�-�d���`%�i.~�i�^��j�#���J$^9�?4��m�;�����U8Z��cd_̲FeRJ�@�\���C^� ��mi�!�G�/R��1ͻ�\b��.)y����vӯB��~�+;Z��o���
��X�>�ES	�E�rKu@�z4����[H�ԗA���rV���,>��wĩ�d_��n�>�9��O�Q����[3=�9l��t�&������?���4��wx��7�>1-���N%��r%��nd	��믄I���Qǀ&n�4��r�Y�!Q@
��������Ո�.n��pt�z���X���1VL�kl��l��td��N��v�v�RT��I��U�:ᵴCqU����F�~7O�Tޡ]e��U������Œ�_��:35����ohf��vi!R�m�K*�y�La��B���r�9��jБa����F=��~�2�x%,d����9g+Ӏ� ś1����o��=��q�J$g���`�8�H�n�Q0S}��V6)>���!
�A� �T��v޲9&�h�~�>}!��fh ���;��Gױ�bQ�S�2.�<w֣����diu��_���`/{I�Y�5�3�8���J�!c�{�C��
J��}�b̤�K��+#QC�Y�����@�]A2E:�r��0���`�+�D ���s\[x�C� ��p!���~W�z�iE�q����8p�W8R�� =��:���6
��V�z�J{n�3HǱ��-&%���iX�F1��A��XM�F#.xa2T2|>�z��	Z7¥у�j?�~�h�"�5,���?��sLϷ_D�u�b��&���N-V���k��������|�K�v>�W��g�Ʉ ���1�H�ҷYҤ���e��Vѥ����[�ZS�4�ϣ�<� Ҕ�E����z����M�3},��Yƚ��QH��[s��� ��o}���U�)���]�٘��GS��ō��43���F������ǯ�[��O-�������gQ`�C�m��c����ѣ���)�{��Aa�jt�V�2�
:���c+��W(�����x.[(�s��y��\���=g1ޡ7�e�EK��&�SJD�g����A'#M�Ƅ�����A׀�AB��yf�,m��>�p��چ@�rTFK��K�)���⭸�j�����D�U�yf������IJ�WCѳ��3T[*.�KQ������O2���(vjk1�1���7��AlGL�?��=
���T�I�vx�&č	�l��C_�	 nŨ7�4?w������!���1-�Դ��A�Th�b�"��������JL{��:V<��������7��c�Vp����9�k�?��H��-3�-�ehEn�4��y�dM~?,H*_"��T��煖;��VuwU龦�7w(�\�Q���w�ۺ���1�kg;��������'�/7?;l~�{�7�� �!��=���`�-���H���?S���u�Z�e�t��`a�o������շ֑J�2���|=~Ȋ7�&R3�O�S\�%pT��{1$�.��]"B%%�:%Kv���)b	C p:O�#7�BU�_�#g��������u`��q2x��ۑ���r��;����/������E �
~hN��-{�,��6��R^��UN�t)����u�%[9�������@����ATH۽إɁs�+xi��֘�g�S��%�����ի.FW��,!D)�;����t3��� s�3JjN�Ҧ��2GS;���{��jp�ʥu�zP�v�e@�-��4�7;À�0Q��оv���Ao=�['9L��1=�����T��n�s&�I����5��;�*�B=� ��L�u��YÔiի��y�FB�i�,`dg�(�Ռm.���Òk�BW#��R�vJ��YIOl�^�'@A01D����>����Hd�ɹ ֒���S\���?k�!s1\|���\rQl��z��\��5���7��S��9H��|�J^x�bq�{�g��(������	�b��.����(4"�ln�%A#�N�ZLo��@^9Wt�I [�3z}}��Gj�e@�݋�
Xe�g��<=��"�86�s2���m�3@.G�ō��t@X�n�i���`�]��q���o̢!��f�"�\9$W�n`��������t��E��`��\��_�0�5�rF�gз�Ln��8*1�|��+G�:uZҒd�е
�1��X�s�;���q�b�z�8zi�&#O�AW��ۈ�%6zcg'-G?V���}�55
�]i�VZ|��C9�1{�������b{Gx��#+#�>���^��	��qˣ_:&[�'?�����{J�4 �!8�,�Z̐<�'�=!F�r���q���T_�G%X^���TCɛr��7������?��(�JC�,�W��My⓯H2f�&�¹���$CZ裞��3ۦ���8ݖy-�O2�U�kD�+�����X���wԝ����~eq������<���@`&$��4qlKS��k:/`�)-#;hS̒�m��J���?8q��AhT4��ń0�+���Z	Ǜ�](����\St�F��vެN%G�u<^IIJT>{<h��"g�M��Ԋl<@K�g��@;3���R^��IYn��sk�U>|��-��JK��������]� �f^�����Rq@�i�^�4ι�u�`l]>4oL���þ�jZ<$�8~ ��1��l�z�[ڭ�fȘ����G��e�x[�<�I�U��}���x�_ባfv�u�(m :�.-��KH�b������5#=�&��e��p���p.Ş���Q a�Ҝ�<�`�s�0�6j�)��|��tp?w� Ѭ���ƂͰt�T�Y�ܔh�e�pp�f��_�S�/+r��^a��;/����J��a�V�����D9��d!���K S�m����jC3�@h�rO���.��e�T��0@��[��~b��%��:[aղA�Yy�)ӷ�+��0��l�0Q��)�� 6�ِ4(�ȕ +;Ȭv�%�)����WTxqj}����G�l�I�|��Ví��G �
@_�βiE��Vqp�[t�t�T���G��N��I�$�Tc�mr[���s�<DW!�S�۵?<z���<y���}�duiTO���b���L�Q�(��e�e搮1�����P2�p���a��Ju�]�w�϶[�����{���!/HɰS�؄x��f�f�^UfH���a�����{|'�*��Hų1�I���M;9:��LhY��
k�m�x�m1�x�����s|~���#��_����4���>�b\�{�����Q�q����ɡu����*��jn�nަ�����.�R�W�1g�V����W��/o=��1�G�+�\���2Z�"dM��SZ�_0�p.Χk1 9g�on��6g�Xg.����n�+\��]"��Xؐ�߸̒v��(u'�@���!��g��G��e*Sl�������i��YE9*ܻ�Q�����4��ە7R�Dve+1r�{�X��-�M��Q�Ko˔��pU�s�e��'�i�Eƪ���2��1��ۅ[�dK� N%�$�\eޒ�;F}iJǗd?%x�k��Q����ox���Z� Ĩ��k2��c]O_�)�#�UE2+l�WG�T�Lbs8����[�k4-A�V+�n���Ou`i�`
^f�b|���<W�p��Y��Z%��qot���hp0�(��@y�'2��?v��0�_}R���3��\@�j���*Z!� !@�:�K��ND�7`F�"3NH7½�q&�h��Km�T��Ei��; $L\�_������O%�3�ۨW���/��&�[\m�3Z��g���7V�0"O��r/��SFBS�K�Icit!T�y�z��@ =�����c[�v:l��dP6@js1bq�@aG��["�)�d)þ�E�=Tֿ����{#:3�S�7K<W��s�ڴJ�2A
Y�/U O���S�%���N�_����&�~�y~Y��/��.��;/�˗SyS=d�J���g�b�`Ǒ��	�KzprB���Qj���e��ǟJ�]0��<�JZ@ԡ�Հ�:�P�;}ud���wF��������%f�~�h�-�:c/��" �)�^�)����,�!�4����0�~�4�1�H��J��I?��xphX������n�Fi{ъ��}�!g('��e��*D��s��?��y�*Ï@F"*~��⡮{�$�q�\J�5	�}�f]���FW��+�S `ˋ��G�����
Ta��Zy�a��{zÇ�d"��g���4�p�����1/��I��15����r�kŒ*[k�D�h�uã�d~0��=V| ��q�7���r5�0A����j��]�*#ϩ��NIbL�#���<	Pn8S�����z��M銡Z|���i�1烓��F����S�Iʗ�y���`�m.�W���M�;wCh�ZwO�$�bw�]=��B��R�3��}��oi��������)���:������MQӳ{G\�v�������ͷ��M?R���K�nf�{����](��Դ<�^��ș��k�P�]><���hr^]K�ZEռ��u�����CO��'�m)e���,����<r)�u�5���D���v8�dM�x�v��H�;'z۪��^��{�C����/q7��M��1I����-�y���x.�L��neP��f�������9���ǟF[����;��)1�9/��ǣ:]��{9kU���q'�yO���7ɾ�=��Η�0�6�o��.������ʮ�g&�y^r�_�ì9��fBp�C">�iZ�\���j�+h]S5E_%h�bBdU�>�XS��J�y�=�D����ǵ�8y���Ǜ�1�IN��&Y�:9��W�#�-���\��F��
w�!��ϊH�"C�@�.8�p�٣*�
Yi1�R�%�6��|GT��-�����,�i�B*�9�Tw!5F�s��AХF6�{B�1��|GB�$��W���g��#�FOI�jX </�t�i#f]Т���G�c��xq	4�Pu��C��M�y��8����w,��U��
��W����������YY
πS��@gG�?KŊ�gBQ@�����mvA�ai�����,�f�^�]"P�=�Q�5xi�ڙ�ڲ̼O �[�^��i!]l�|r_.�]�x���xt�CluB?���@��z��vt�YkWM���Di����Q�l� g8� _V��K�1�K����L��i�NGB�J�l�΢�A.�Tu y���ݪ�"�t&��n,ߊ��ُ3�/4�Or����G��vs�4e�춎��o��o��~	*j 4>�{u���?����Ãj��q��Ϯ.�n�2�4�%1;G��8n��H��r_�s�)&��c��c� j��-�#b�۝x�ϻ�H8�C��WZ��T?����k����Zrp�ِX�-L$���U��c��UN�=S&�Z]T;��ٺ:ts3(�Z�(��_uO�~�=]����ɻ�Nr^��Z|]��=@�}^r����]GL�w���I�)���d�N.>#;��q����k}j�����tL8�j�k�#]�����B�U<����̷��Ԝ����T\+���v���I��;��,�i�#���b����]r+}�^BWX���(�����)q'h�@�F�NWG�܈���ID`�)(N���{�! #r^������=
w�W\~�����v�~���[���ƖΈ3�Y*��Ҏ7��IL��k�K6$�%C���(8����<[���'�O�Sܢp?3�Y4\Y}:�,"]��=��>�u ^(�y��Y�\��C�g�$�f��#�mҊ��E��t�1_4��\^<H��2p�	�U���|�Kvdrk��Y�����=��	�BXv��1��="x`�ye\=�sj��t"�+��9��-��boN��X�:�~�vQ%o��Ϡ�g$e�A-R*�%���8�J�z�^�N���4���Z�Ԥ	��ʒ+�N6A�9}XE�2[���D	�C� V��|Wg�/���C_C���M'@��.����>�vχ���8��;�s�v[$Dؑ
Y��J'W����8�ׁ}� W�A6�5�2�ݷ�����iE܆�Zp*	Hw���)���i�)��wm��!kZ�9��d�{=�.��{���
7��c��T�Tc�����?���n�h�M�p�Y9wOI�5@@��g(�E�����_���~RW���<�sMu��c]��;!nJ���=>�v��AO��&]�t��\��#�V�Y�/�rtf}WcD�&y��{��E����Z��+�OY�ˬ���Җ�PP��_�dߠ�߂���%�g����T]�I�	������7?�~�MUTѺv��
�DA�⛜�9E�Y��Z��}8�Eiģ>�������*8��0?����b��B�ht'p��
(f��E8ae����hH"(��c� 4��:uRtw��c�Ɦ����Ht����;�y  ��ǭ�X0�Jz�س�W��gE1H�p��.�j�o� ��m��N�r��Uc"�j�L@�q;�?������l�:�'�k\*�g�3�1���ʫ��,��V�#1t��1��Q������b�1�Χӟ$���j��)�fڿ�	p�� &s�F����q�1ww5/%!U��)U&����������cP�ߩ�ӫ]wvK%1�P�:���y6��Y���/D#��:��x�&�.֩�CD���h#t,$�b=F�����$�U��uK�!���@s.%�K��� �fI�����VU]�w* �^�zl�c� C$*��	 B��gh��JP_�\�~�z7����5�=a����P"iz$������wT�3&��.1TOқ����ǂvD��+�?�/�ǘQ1;9n8�-�� �2@5ާL�������?viЮX�&i֏��R�욯��Fo�@x��A8�H�R���yf�:��8S�m�d4���$��Jc�Ƌk��A���%cz��"e����J��KR��uB��ו�ijdلF���4��J��1rid�	N��v<_LH(x>Zu�\Y/�j�~d��Ԑp��k��1��E�]6<(/�vYl)7�8�	[7I���u�jO [@�ڎ��K�ʸMҵq# =L���;�����N��ƺ�i�9##d�Qɬ�G:��ۤQ����1���\Ža��͔��s�J'e��xR�L��H��W����"���Ok�ȝ����a��l7���j��>! �W�J:�-�Y�����"�dQ5uM�����>G9�X��v��G +m�-��68ݺJPU0w��BA|�z��c����U�a��Y�����e%}y"���C��8�rn��v���� "���5s0B�v�N�凵�x��|���5s^ ɢ9;�y���e�~L��;�&����H3.�����{�ȸ>��6=7}����FRz���i� #So�꜃BE!QPv-�ٷЂ�^dof��za�P8'^[�տ�h3��=X�g���-�9�MaG\�K�s�����c��{���]|��*���:��.s]�� j֠0 ���`�XV����4E7�#Q^�7��X=��<����\�c{Д�T�l�`��I
�Ѷ�;�g*}ۋ8Q��?�
�G��A�m3&��M���^>G����a��#&�$B7��W.	�C���L��,���nO��oQ�@?�Z���}��=����H����C�{;�;�1�|H�y��=�i�_:,W!Sq��"ڌ���"������.�W1暰xDn<���a{̖��-Q%R�
���lԾz��z��tI�F�O�y3��$�%D' #N�Ѳ�3��H�kbI�<э���=�|m��٘�����eA��6KhT�?���=��ۇ��|��bdp*��l�*P	{{6 {��-�[ƌ�H!:*�uJ$�?%�y���� �
9i1�)�ݶj�5�-�'��bg��P2w���� %���ˉeU��8�5Ԁ3�(d�c	��y�F��26�✈�Axn�w�H�a\*��`p�<1�1�����dbPi�=���ãh��։�0�-v�����Y��E1q�>��{����S	0k�4Z���U�A���x���mZ���T3�'��+��5���7J>�|wc���5z�\���#~3�6=�i��2E�~�^��P̩��.hoИ�Fŗ+:.��ˊ�IN�G�ݓ�M	mU�ƏH�0��a!��FX���Y�4�[��Z@����aH⶝�FLO-���Y���5>�kR��|�ЄH!�;Z5������0�)�����;`s.�	���~��տ��f�� >Ӣ��9'��5
P���,���2������qH;�bt'c>B��wQ�4�>�eҩRs�v��wL[٪ �k�Ol"��"���\���������t�Ug���.�Q�T��i�|�;��<���$�iE��'����S��zCYҫ$,1��t��mFF �ы�(�qy�i�4Q	�Ohk��fPj;�Z����)����AϖpD��bBM7��@ީx�!~i:���ӄw�
w6�T�K�(�$�h69*�4���]����V(:���/gXn�B��q^֚?�R/���X����s��m&�>�"ԃśқ��XdB�� x���r���AT}K���3|T�r����]��-�F}B��U`Ң�@aM_yN}��,�A�
K�� Ϣ!�9|N_R�6�:Rd�g�a�����	��娒�~G+�B���E�1�_�aY��y�#�����r��#���Fku(��[P�# �p���*^B}u�ڵ76��!������m�i�U`���8�G�.�r���U!"��K�	���ȁlܮd�(����`���1�oeբ_����ق��C��L�*�O����z�} ��/;��H��g�8kt	�zI�次�Ɲ���I���/��V�]��Y�&�L�������?{A���֑�82`�aeco8'��s"��6vaG��o���T.$B�b[rZ�M�b�<s.b}?��������Ow�r���6sYi����"�}���`S;4��>��[ �mb��bހ�~hđ@�<^��,D�1��-�
�}B�"�O��Y2���E2'�A�/m��+�ܭ��7�E2-ݘ�RC6��?�k�rۍ�H��A�cY��Ud��:�K+�ٵW4m�r4����b�8����G�x$���c��}���KY��-)��-�4��_�*%2;�ʷ_?�Jf�GR�8#�=�-���W�	�Mz-�`�F@bCH�9]�8c�*`�ޖz`r7]~]c���^m"�S.ɍpI;�~5��
#�6�V��I�	��������g��b �}���c��=jGl�F�7��?�ޛ'��r�cw����f4N�"}X���Q�0�mU?`մ��zV����uo��Ӣ#6�g����0��E<CD�?���`�z�G��n�yC=~o
�5�5��ה�����rx�lԚ���_��b�H1&�v���J<�������;h��;��ɮBa�LY�lCK:/y"h���p�i �H�i��_���Mjș�07����@��إ�	��l��M4�q��	�ZȇZצ�w�#���3��_���F�V(Gm8��e�?,�����,b!É��ƬWⒹT��Ī�Ǩ�u�����wۤ?���A%U�#�r���:[�k�X^� �ڎ�wU��5A+Pk�,���w��D��E���A��/�і�	�(�N����Ȭ���Q������.�+���{z0m�9ڏ�|�p�q���ct��,H��x"c@d�T+Jo�3���ʮ7|�J�����sO���y���C}���m%zf5���g=t�8	P��F�:1�o��	:��4~Z0�;�m�t�k�50�Y ?*���������!n����_m�:!�#	g_�S�G�۪�_�<���^~��/?n\�i���a8	�-��lU��ź8��o3ݖ*,���?��-@`O��̘o�;���ͺK>i��Ӧ+�Y����܃R��J_Ѻ4G>�t� �'��%M; <�Miv���ɧі�S���3�{����cܖ
�\�i�,�J~����1�NI����Lc��vAhSE�5�{w��Q���.ˏ8�<�*u����	[J��g�E�tp�ʞ�0�y����?bSa�Y�0`��T�+��f�y�o��5�!��L(3ң���s��L/����ٗ�?���O�IZ|_�-��,�ڡ��Ę�.�3e��o��� U@�����8�!x�?~����"����3��\o��,y9)�&VTv�".��Ċ֎��]U7��{KD*�u� ��l��G<��()-�@.�j+��`��c,�tq�ٶ�Rx�������C��;�0�K��欖
XQ��������N���Y5BF�F���R]�Zm�s �����!�b0ېU� !�*�ђL��	�\L�^o�7uW¯��fZA�<�V�Y�*�Sf����� �r��T�k䥯�W-���b�u1�#�����/)�|�l�u��=�_?9C4?�^W�S�x�F0�g.W[Mr���<$ �w�1��B�@�߮�QXkU͐���3' 5=�IVe3UF,�D����� qt-���~+~�ڤh�=4�GiSu�u �:�7�/˛ �{��᪏��H��W,�����y�Bd�f�t�oq��û��US6Ia��ߝ*�H~�i���ݸ"1�E=<u����6��q��!��"si��BX�j3p�yXq�1
���!sWC姴�Q|��.�k;R-8��"xFX=)��4�ċ���Qf=z�k��T�������]������Dڽ�F� �΄H�8ٝ���n)7:]d5�s 9߮JX��~c��������ԔFRhRc.c�	D��\͏n�L����aZ}5���N *J�A�{I���6��u��x��M�-��<�=�DS�8v�x>�n�����%��M	����06�\.�"���}9#:˷ �N%����&��M1�H������Zf֭ޡ����?�ݼm��d���NL^a��pŠ���J��9@k���=�A�y����	2���P�9x�Un/O�7�PȌ��{�r������)ӴO�>������R)Y-��ϫ�E^��R�4���N���jhh��<��݊���w%&)�K�ڱ��{��#�u�o羰֦A���!����]R�[�B1"�r��mld@�s�1c�܂�G�O��F�ST��z��]�����u�&�����;�BN��c�j� cn�L�9��m���ޢ���W�u���b��Ø$�G��%�q���'6u݀��Zo���0�d%�pS��qV��R��{_�D�ٮ	AJ���!]��=�ƨ�lP�ma�i��JkզB�堩�T�ȭ����{u�����j�y���7E�(!���n[��A����$��g�~9f��� %��
�oqM���ڠ=l6LWV/��ͼ)^�Gmrq�@C�c`\;�+dɛw|���o����wT�2��JxK��q���|~���Xl��~��=��mR��F��~/PK�N9!E���N�7q^$c��@H�W*�~�o�� *̌����Vc�((:s^˛:`���f��W�'1K�I�\�"u17@ݯ:�3�{0�Hw̽`�ʃ
�y!��� ��/���Ld�C@��S��j��IqB)�����?l�X���t ��E����x�8ɂ��m/moX�C�{�����C#k�v-_7*�!�B��Q&6���|QϨU�|}��%/�
�yf{�[dA_\�%�Oђ �j�X���#�6@s0�$����4�
�����uW�>9��ʙY[�u=��[,hQ�2/���!�#=�{��ȡ�^�����[��0�� HDJ#N�&��_QT���v.˯������������8'v����_)�
�%�y�v�2)xٰ�ci�6o��ד0�W5<�k�ƴy�tK���Ke�f��!l����g:�%ڸxi]������{��c�~�ŵ%�4��_�䲈��=�ީ����#�4��XXR^`c�MU�]r�[�g���ExjL�Px�6��R�5=���f��y���P��Kn�Q�h���WF�JVmL�!��6?�s`�'�&|Lt�LI=�Q���=��˘O�*�9��8IX�����4�� ��.�}�*�6A�A�pf���ЀT��J�#\8P��խ�I9��Sz��] �K�.�;,�c8U�>�����N��%N�.8$�� e4��������JS��N��-�����-+����z�{��gMc���B�S!��e�[$��t:>�/N0��RDͩ(i6���0m�%�����[u����>p� ;A_�������=YBށ�
}��H`�#��}��C��h�<a�jbM/��z���|T�O��C&&�g������[��J0tNV�$X&I�eWz��t�ni�?H�\Z�}9u��,�{I�ƿ�V�tx��&jHc���� k�֎W�7`i�-� ����~�f�l�`��Ѵ�BrWp�*���顇:b�o�4�!v��x�sB
����k��Gz>shʺ�dF��ȭ�"��.�B��ǹ]6C�鸛ۻ�2"���*t���U��b.��N�3��4>���=�$:��m�q��L�or�gbY���i1��~tҁ�����]Ps�G��C��6:A��E�=D�"�V�� V_4�Vt�v�Z0A�e��8-9���_4��*;�~����5�"�1ײ�r�)�@BVr��6�V��/7}�� WF��F�Cimiَ�v2h�
�0>G'�
�����,�BC��i5�V��1I���k����	 ڏT��V�t�2����ø�\�r֪+��;څ�|U���YV$Ɩ�[M1<L�v��r�4s��. ��.'�]�=���9�҇>���Sg1}�+&ݺ=�Y��xE�#*��53��5����3�0�4�%�E5������"���̙�7������3I� �%�H0C�\����е!��@�݇���j{��������O�jQtM9[v�Y)g�^тu<k���8疀�S�Eh��e��08�w�Y��4h3��#Nl���u��P�Gn+!=�P1���@���f�'���@��B�49s�M]���*������v���0�ks���x���� o�ǾO���pf>��Q����*B�Q\������~�z�U��%�D����h^�"��؜�G9�f
��䓎@K�ђex��!��5Xg|ͭ(�l�.�,���gH"]RTm9dr�u�SQ5̄(�7iq߸��Ǣ xل[.��1e!�dB�1����)���c�/�.a܎�I,��$6�M���F�ͩ[����{q�D`��µ�v������]+O����U��l��-�:IW��wn	��#��""M��6���?�͵���P�,e��̾���m1 $P���P�S@���i����d�Ѽg��`_��E����;���������RN���}���2�,����J��
����g�ȯ���3�j�C��K�VCQ��ͯ�'�|��>�;<��
Υ��1+����e�yt�^�D%]��?@��JdX�r�mv��-��Ȓ0,VQj�7$=��!�:�h��E�C�N�Rn�Y��y���ݐ}	�.H�Kz�C5n��80���!Z���.׼(}��Jhw__/|��*�)�^��*N ���YJ����a��yj�$�pL�0� "�Ҡ�%��e�:��a�d��*�W�w��\�:�w�n�o^��h���?�o�u2j�P��BN�4��O���n������- 8���Tw�.���s�\�Jvt�s}�T��uD<"��Kw+�'1d�מ����>4�8�����Z���.��8��%��Pe�[o ?��z
-�<�;y����L���&�A���Ҍؙ��r���F	��m"Z�K�[�pR�l�T%ׁ2&"Hs/����'CpˉʕK����z��m�[M��{��Pԉ�gś<���p����si�c}l�$�2���LM������m��C6���7��c�
~ #��J�@���OOf�FF��R�'�"=cl�8�|}P�Ѓ �NZ��Ƭ!wr\���"\e����4H3�UOjZ���i��)�E�N��à��!����U������,��\��J��Jo����1��H!�^��*��=�����m77[=�v��y��ԢIY�J�O�ȗS$��X�.o�ˍ-�'g+������\�?
5�N1�c�8�R��։q�⠆�pt3��}��A���Q{?�!H���]�2QEu��?�ˮR%wS�o��t�@d���EmN�ֲ J21ѝ��'�W�ddݟ,ϧihOuf��jI,u;$1 q���r���m�P��h�}�2\=��[��+��ۧqN��N�وObǅ�΢��v��0�d�,�T':b�ﴰ7�L`Y7Z�.0�J�ސ7���I�΢fm�E0瞘�ˀ��b8)�h}I%����L�d�(Hّ�Fڼ��pձ�˅�\0�M�(�&�E����c:%��X�g㕭�]_���3+ޘp�<��g�;�ze�C|gq�s��Kt�lBv������lW5��u�/~n�ۘJ�Gl���q�i'��۞��w�Z�Nh�8�c7�۟G��7����D>����ȗW�K���3Z2�𡩬�����8�Ѡ;/�f{0J��"޼(%��t�8C��p}G�Ӄ���}����=0��yB!�j}z���z��ǁH��PF.���;�� ���?,-2�M)T53�'	e|?�#�Ɇ3V�5ŭ��a}m<���{*r#����I�a����М�E��gf�	��]QK�� #���=��,֚������s"�{�^�?]�5!f��5���o�1f��w�o�aFkH�;����q*nޜ���R8�i�V`<yȕ��+��S��\»��ҒY�7���|�.Le�?C�[��2�?��yݨ�Fb] ��"P̕f��s+�v	��2������W(��ܱg�-5b��4��uA�M�gQ�hx��:��D)���w�m�Q���J��×�O�3�B_�7Ɲ5�|ѽ��>�¨��dޘ��{e�K�4y��6]�6���.)$ 	�#f.4����t4^�%$ی���	�!)�I뵜��PF�Y����j\EQ��\�U��°HJCQY��:!t��!��+pf,��3�4��b(����Jdg>��3S�iB+mb}�T��h�9	��MZ�Y3�3b)9�P�A�Cix�8����v.��sNI]L���z�
���#��"#�3غl�� �rخ��oA��D*�P��-��T�Q�-�E�uS+�?+�y�[@ŋ]��}gch���`\ �s�Hn�� �����~�Ď�9���6�?�#�O�nЊ*K�����2:�y
vk�\<�;)� �Y5�#z�8��K�ı�-� ��* �����>o><�����_=�"7��������s�b����|�Ex��_PQ��ǜ�}:��1@:��,���象a���<��3�p{dH���W�Y�	�������T�)���%h�wY7�c���J��k�}�P!2qǽ�EF��L�� �c��
^��)r�'H�2��¬F˿�����`�Q.�]�#v#�!;Z�/�
 )���]DJ�)�սa���B�֮uhZ���|��V�x��ǐ��+`C���*!���5�5'�q-��7.��|��l�����oa�~�;-� �ڎ�H�M�(���;n�H�@�m4�2�fɷ�˘VhO��N{���6&�f�� �i��`:tw�|x�
4�	H�-mj#h�!179%G��y9B)fֿ%	Ƣ�3ؗ�����a���[��/e�N6]5��áa��6q��Q�핾�`�*Vw��A�WqS��;aϧ�8�Uͨ���*�����9�=����Ss���1�k��_0r�DZ��%�Ca����L],�8��I��.�X�"MN���>���y�Tu�u�C�(��J�ڟr���R��#����U]l�����z}'�v�E���8�f����y�q�������Hc�>)�XH�n?�O�L4ȷ���*OXW�/�K4yK9E�ëuL�Ǎ��1�=�C�q�TP �w���B`�{�DROt* �n]#������\���Rk��5U2~p�����yZq_�Uj��'Fy<n�Ў��/t�w�[�ў�k5�R\qzPv��:��9�_B�3�O�^�<�^��Z"U�� �vf~�O��t�����X�%[���c��~{� |����7�?��|̒����Ӟ%D��?�Z�i��-=2vF�6���1�]M��͵�!:h��>����z	���H�Q�f; O�jbCc.\s�o�ȯ��)�P�*��]6��V?���s��6�����xp��`&�P�y�7����'�@'U88)��t�x/]�)�_���w��5d,��2��-�Y,IJ���39���A|��`��.����X��.Yu7�Xg�B�b۲D�mfե�W��f�> K��\�Wö���9-���AE޼i��Z�_�!��۔7�-��Z�&�I��D*H��4T��x��~�V!���!S�Rmf���U.���gP�p���(:5D�
�ۨ��@�P�����n݊r��S�[���$�5P� o���5�Z������.H�n}�*�T*Yp�V��f]$�(�<w{�AO`fC�ֵ����1��E�L@�C
h�f��{z��;#N�#hՊ����Y���|�Gx����А����7����oȔ�����[|n���>�.�$�7�BN�� �|i�X��b
`���t��&a�\��~��1��.#�R!$�oк}SRѲ:�y��ZiT7�cǋ��v��w��+�8�M���Z�u]t�����Z��q�(X��DYT����5�3 ��ۤd�[��ܟ��挭,=�2N���Y`�7C+E@�7�������p��|ǲ\I��\&�S}����,������a���%���p�����(��A�W+���� ���������6��5�Be�{"�c�>��va|!�w-j�����V�˪�v�l�7vP*^߭�����
�Af�ʢn,3��HB�	�ְ��$��p{b���	�qT��(y�'��h��φl+�4�y�U� �ryMw�E c�/�I�������~�1HK%y�.�_49����@�[��X�	/�9%�}��R9��lS"��XN��=P���#m���=�=���Ab��'��LfV�y��̡o�%'q��4���);�E�QwIR����%�ڕ�R��)Ga���N/&KD�J���ff�e�z�2,P97S�����u�{w�Q<�oFv�b���s�{A��@4	P8
�(kCQ�)� �H<u���:ũ�Ȉ�#q33��'ZsB����ޑF�_��j$b�|-�׌t�f~�+F���m�Y��g/=�����^�2҈&�7���/��Ov�z_)�4��O��r�5��@,��Y��)�Va[Q���5�W#W&S?>�3���\��1Ǘ��q�Y��4�U�9&�����Zc��ۣrk7���N�Pa�b~m�V�M�w�
EO���]��H�P�wQ[1���&kd�[��F����Λ&��p4�P�&�[&�Ga֤R���Li�َ�2�Hxv9�t���V�KitNn52">*Z��e�C_HS�D@�n4�5�۵��S�:;����Pv|Z�[Sk�߀��޳!�篡TGl�M�."����(c�������0�xB�T�Wv3vԢ�+�}���43B�A'�%�z�e9����b����#o�N�51���{k�KS(�*���#U;�8��ֆ�Yj�A�aB6qxFC��S�U.Ἣ��O�1������,J4�x0����hdH�-��Ь;.<k�sE�d�RV'a%gk.`Xwޯ@��)i�):���,λ$���&H� ��:�����b��s�nʯ�8��c��0� ��8���'��o��2���RG����\�~�
(�W9B�
�l�]M!�A�u�9����w�c�q᷀j����^`\ K�b�j�*�W-�v�?A`-W,&�30/!�� "�F;D:O��FbdE���q�.��3�_ ��W�&���U����3����n~q�q�@�30��}����y��o�:�M#����Я$���v���S��驶���|�����Ms�����[ ����^�J�N��mɼK�)[l͵��R�~K���&��<ҝ���jr�w^�sD���pJ�/�GVJ���ǳ�pA���BL�vڻ@`̈�N�.q�wQZ�=t��{:��˓�Z���j��:�h#�U<����E\����CL���bO�{��:�?����Rs%��{z�_�.�����Pkޔ9�.v�?�."�_!��u�Dh�X]�G�����y��I�<ЫU�0+�8Ă�L#���'d��z�`���-d?�����1JJ}�q]�:0k�u��*��U@�h�cȖ�1�U�p�T�f���4i���Mz�zYϟ�慄ͦ?�ͣ�v]H�]���tJ��Q�5�Ԥ<�P�!�:�\�}�[rk"��L�e�l�> 7� P���n'��q��p B�F����r�O��Iau�6���x��
�T�AB_g�7��`i�gNӞ�-�ai��xO�G�����76u3c�VXp�
:�[�GT��t7���Cٽ�ܻ�Zr��J/+ݘ���K�*�Dj�_\:���h�x�Δ�6�0�9��z@���ʜ�o����"
��6��GW�S�"5�;R���B ׯ,O��fsҶ���n
���c^��9�� ���]�����d^���3��Ͳ%D���¿����z�_03#A��.�G�v��&�}Y&"v�:V�!xx��F��<��F/@���ՎTx�8�<4���8��_�ƷTp)h'������_@+	��w�/�(��\����+	�*����fCY��A���^��F.9�^ꋽ�.�7�F�D]B�uD�<*ko2� �ү��Ni݌V��B��KΚ�>)M��v��<�֔��o��t�pDh�����v�Z���{XH(FE��oD�0��SX����ۗB����=3��~����N����I	M�kg ��Mt�J�SYoQ�l5�Á{DI�� pA�Sym��ܕ��m2���,��3�XT��0aG��G�]K9�ez���Y��g�uǆy�eE-�(ʊW|�(�1��_��dd��tZ_���Xϟ\,�4�BD�o��
�za��������P���[l�#?x�n�9X!�n�B�Y�9��C�����8��g��Eʷ98ō�2߿�f�o�@:�`b-��s42���y@�P��7m�2�֢ͽ%���ܨ��&��#�cT���Kb��ȿ[_�0Zd�p0�>;����o{1,�2 �r::�g�xҬ��b�T�0j*d��9��vIW�OV�;���S��B􀔰������dPH@k��'5���(51�s�ߏi{d��L 
��kc~}8��_�z�f���Q��ӷ�#�=lhW �$a��FE���xQ@^H���3����s�'xib��2R���H�QFs�H�އ�b��yh�z��89�Z{�W�����X�ٮ
���p�Ci�6kN���ӧ�+S�7�z�҄u!PӀK7�W�m~��}6�/�{�6��t���ut��͒��h2~\���h7Z<��nu���� �D's$����,�;���w �UO�j(
�O���Z,��H�m�IU�Q�h��"��D�?
N�2��%c�f�*�4�5�R��JB�-�t�/�6>�7u��]�l��d.0q�H����[��6/�mnW��:c�G�0c����+ؤ��J~$�Vk�j=���� I�H�.a[f:��g�l�������i�� �t��C7;	h8�Tȹ�s�I�������L�����9��<?S��v=�x�x����'?k�x�%�7*q���\.@�~��NL��T���^%=�M��CP��&��b9�%%��1�C���jH���Z��g�,�>���k��d[4��B�n�ţ��(%�+>�n%�7ׯQi
ԑ���}��@�gm2{���Sr�U�΋��6P���&qH�ۈ�VU����E��c��Ҷ� 6�����s�~Ȧ-.͒���	�eS���l՜��J��I�ڌ��ߠ
���m ?��n�δ�0���R9�����`!�42lHB����_��f�7�0D0�iQ֨���}��?8��c	��j=�5v��nc�e(T�w<({ ��9�kcbL�ix�r���"������M�8��q�5a@W]P�-��D�F��#kFR�m�("V~�^c.�T�[�>i'혓�B�'�:�_�������݁�#�1�9X�����E���A!μ��,Y����"�h����E �e���>,�4��5<d�}�BrL�~ΙV2��v�`Ô �9�B����c���$W�
�1��$J�V���G�]B�j}GqP�\D)v%���
j��Y�2�I|rs�M�a�����BJ�Q���Wb��ﳺL%��[�d�8�e4���vlDhb��{{�uL�$��D_�>�� !(A��I�\���PR��	��?x�g ��Z�u�z�'�.$D/�
��oER��j7&�ej(����]�;W�(On�"�Md��2�����I�%;�"��dG���*q���z��	�g���Kަ�\��@�3�K �u���2r�R�`Ol��L��u�9�4=*Lм���	�9lH_d�)'�ɽ��3��#�E������f�ˡ�u���!�F�|��U+�.8�t�W��H��A���N�_I��3�f
�D��I�+�J_R<"��V���*Fx�&��.��������q4;�����J����aX��,�g���ޤ�ρ�@0�<p�W�d��Mz�hGk�3����'���� a�|�{$c�rf �e��g[�����Ó�/5�>���+֗ ��R��������.�\�y��;N�J��`�S��cN��;@Z�^U�	0�`�ˊ�W���EBy�l"VO_J��e��ޞn�p.��L�ئ������n&�Xq:�	�_��f[������N��+Qō$�U��|����S�ѧ�Uf�Z� T��G�[H��"�r^��E^��#l���CqK���"�e@[YtO�'ҵh� ����,nB���:��_�mО
��gh�c���o8Z ��9u'�����dtV�C^p�W���zē���y]1�+^�9"uAQX{�dokx>k�~k��i1C�!�.�#�l�c	]��\),�f����Եߞ�_����"`�$����3n����Л24Or��Z�J�d%J���y�D�V�~�kxS�YՀb�����ؕb#ucp'�N�C4�m�����:0˃�ٽ�����n�^� A�zk�H�Y�J/�8`=S<C�UW[��(�|#j�Xk6������TVQ�zI5�%���������>x��ƃvh�E�����@�Q+C�pc���Լc\%��5���m�ң�6�&8?;�1Qo����td6�d�!}�V�o�@����Z��T�G4#UX,!�GJ���'��к�E'I��&t�_��C�+�!��}����!Z
{���) zl�m����%Ͳ8m��$m����b��\S�Y�'[;����@�:|p$�ة�q�(�Ϳ�й���[(�:~�F�Lg��O���.O�8�?�"�y��"e�3��{�ꢟ)��'����#Ƃ��ܥ�72�y���r[*��A����#@d�f'��g�m�O�	��5�$n�s����X歰ħ\}���׀�s�
�v�U�cK֢(X�lȐݍc�h�0�M���lgK��N�;�(��D�A�Đ�+�q�ܭ-���b)靖`�n�1ܻ;3դ�������d��<ܷb�����w�j��%'HJ��͸T� �A�uE[�����1��*��ڞ����SÇ��[��8���rH�>�V\7��68�6#�k.2L����"����-��(�j�oJ���~k��1�>����Rс��2��=��z>���l!S6�J��Ъ�kV~�kM+���
���J�c�;
y����D�z{Į��=���(���N�`	S{fU��~6s��U:�� Ǉ�7����K>���&��X��p�E��N�7�p=B~����D{&���qe�������V��[W�`Sp��yο�|�j���l�O0{�����?�� ��6����(�D{9\�%[�����뼻{m�=���l�h�}6������D����	l*~�:���I�@��H��jC������Fxg�b4� 4[	_�ϣ�X���4������:�^~MW��$��?X����������_�_�2����'B��
%E�`f�ũ�
A�C�5L�4Ǩ�S\ڒ1������'�������I���y%�濆̼��Dc�.�`��f=�]tx�"l�уirQ-/��.��e#6cS5��E�����`*�0���fAN!�⟵V�c��œ��{��D� ����X;�k/j*T���f#G5�s��C1��n�
�%�i>Jx6������wU�u1ϻ�i��E���]�$T��� wW�$����G����0'u���Yg�u���5��`��/I�G��UHЛ]��;9�K���8�m�gI 3���&Yu��� �6\������{�=duڶ��1��%�:̗��7S��f��H��4/k��'0p�;��v�n[�V��'xg~@/C�)seg{B����`Ⱦ��#���6�}�P	��ߙ<�o�&Cm���Q��lV�d6<��%��.�6�_@�j9E_��4�!y��7]
������|���� �C�V�&���R���r���!:�l��9�{(�W��L?iW�L�x�흲��o��8��ߵ8L&�Rt�s(�R�y
ϫ���VqH�udDiJmr���ʱcr����a���e\?_A.��e�9�ݐ��9�M�ؓN�ÅрAfE����ԣ�'����P@&�2�f���(��K�͏h�%��?�v���$7\:�H�n�^��!e4�=����($�֮�-왬�4�_$�D��#3��z� Q%F�a��5���$]����R/BCe����k7m0m�v��|��|��^��9j��/;eV�E��7�+�CHVD������[�����5�.��/� �l^�$Gذ�j:�%)����ҍ�#|R�E�[T�s������i��\u�c��ᤨA��x#�l
*e������_�Ӫ��	���.�:�'��c[.Tp�f���%d�0��آ�n�+�ף�"R��rQ�3D�hL��� ǅE�ߪ=(��J ��n|��\֝,^�����v������1����͗$x�� M�ݮ�!<�%6׌���� �5���aP븕ǌ��j���&�/��p�.������p�@�� 0�qa/uѼY�K��ejUJ<}
�"�oۼ�n�*��$wu�l����>����<HT�ojj�M�b�8$Y��3�����A$��_y]�J���w=��{�~`�ѷe��\/φl�֓\�?O�q����7��
��ʉ-��q_1��m8�|��ܖ��Q�)���m�F3н�U��I���Km"��a@&:K-�*����w�(V����뿓NS�!�B��I�/��u��I��L��Vc8�
�qe�P��>a�
�Y"�lLf;Z�UwFGSfCB���9K���{|�D#�.�r�C~zg#��i6M�wRm�L�}썐�����vl�����e�B�U4�>)ʆ4�Mu��p�d�V�Yo�� ��(��$W��q㈎�L�l���
��FX��>Ǎ�|\j��uK��p���̼,=�G� K'���X}Hn����=;E�u�z��Ә�:��J�4�G���uh��\��sCA�qs.423��=����r�ɇ��*�����'��BͧNE���2�4^�r�:�߉�^�94r�A���ǘ�JD0��n񁀎!�v_��/�����(���3K
�SK�e��כ�d�!�ߖ��֚?TP���\cq2�-��w����(��	�_G�R}�T�aF��#��`N�s��˧ћ<B�����g��J�εtf-Z������ɫW�����@`��(Y � l�l���}�pb!d�_+y�N�zu(alJ^O�xPq\����|m��e�����|�)�$��MuN��BDP�������e�������zm9Ν���3���1�L2�����ڶ'p����f`�>
�A��C�"@sA�Ukw����b��$qL��]�<�_���ŁVٙvl��k��(�Ϊ��M�2ɾ���.��&}̥�m�Zj����l�Zjᤵ�M�b�C��!n[�4B���dC�jN�)s��#�e�Zm7��d���0Q�����Q3^�� K�u]���w�����I���9���3.&�'��h
7�>:L�FT�*�� `z�JI˽]�8� o��1����#��d�&����� 	�)��b���V07��`�z5b�)��%]�$L������Y��Ǚa�qDf�H �l�W��Ӭۓ������/a[�8��Cb������f3=ލ��c-�6ph=�K���,�T�z�v68w�
�Y����	#�:�k�bn��z��t�>2w�nj���Ӄ �jN����f��q������t��B���S�i�-�s�辄R�ֈU�$�=���7�F.�]uV�FD���n�Q\b:+���"����,)�=����{g�^(�s�L���x�ʹ�v���%��L�-�ʇs�������,L�I�4BM�
4Y��S38�0��0��I�0���x;����'ڐϯ�2E���0��B[���*{qO�eW�t��P��?�_����H�Wp
��:��L]�O�Tϥ�<�M>�������I{y�ae�R�b:vB�4�N�'�qQ�PU�@�����mt$N�5,�A����q��+M�׳o4�.�	��+3>^�h(`�������7���+�5��'���'д���6�����m�'N���o�@����D�8.���p(�Ԅv)�P���H�Ҕ20	vz$h������qw_Dg����iӥ	�ެT:�_���X��v��s�3�x���*O8T�3�$x�)G����9RE��.	�d�j�˪��KB�O �#P�I�{�̪mB<
���ֱF�̈P���s���$n��K�0�u�����ʺD\̅h9�l�WN�)U�cE�BW�Xm��~���+�Zf[�G�i���&93�/	�Ih��Y>Ҏx���jn�{ܘh�i���~z(Y	���}j���6��޳���T�VO.&�)F��\�����[֭���^��}��P�7�����U��}����~���E�#Ĕ��STz�����m��5��h7øs>(l?u'�l=y:���؄h3C����vPɴ�N���͊{�4����ъ@�S�g�ƪ�ZWO��	����ј�����Ժ������O�
�/�V�bS�I�;���>���g�����F�.Qe�r�q>ip)V���Y��.���~�}6e:�u�]�l�����zQ#u<������<�� ��@�}�Y T8�Ҩu�%-~�"�EG7Ry(|5F��6� �~�w�j*��(����{�/��P��HW��B|k�>,�iDя��st/�� #����s�|ҚB.�&���硳��;:�@�H��wg�o���4|��6���L����%�78vs6�+HcQZGB\��O{����!R��b_�}�_6FB!Mے��x�BK���߄N"�a�0:����z<�3�}�eن�s\����?�Ev��}���:�j��oړ�fTb�U뿺@�� ���^}4�@���.��Ïc!���<EeÎ���|�,!�l��v���k�.��̅^��Fٻ�D3��`��	�	��x����R�`�LK�G�O�2}u�3������=Ujʔ-��c9�����3#d�Y�1���ͮk%/��g���A7 {Q{�{��3��EM��� �<��	tM��qd{=�.=�A�tf�\o��.������v�iF��)&�����}/��8L5�b[f˲��+¿9�����7d�6N]<�*�v�XZ��/YmJ�d7J����z�t�@-�l6%Q�2G�H�uؽp���hKxS���k|er6�<�qr� tqu;S��P5o7l''���h���XB�G�7`�����x�F#8|]�W�g���o��g[�[�nP�'.�8h ��M�Ȗ�����2	c@�6Fǃm*$KG�M�x�x�;�l0](�+IQ�;����M׌h_8���x��$�E`��)'���ѵ� }9\�ͷ�����piCXPg��t�|qӗޙkL�;�Lg3%ͼ,&�^��hy��5�ЫQ�ѹRe�Z��q�p�M��+=�b�5��P�.�&l�>�E5�1�Q�D��0�;�H��	]���Yx�N�����gf�9$�E��%� ��D��U�{q���3FXm'�M1�"�P�Oåzh��g�!7beWI�TO]�BY�2����oN���Y{Bso	��O],��KFB�s���fA��Ѯ�b��VѠ��	G�_�Y�����bY>��m�D�>�P�_�p���t��d���Ii�ֺ�{���Q��mP2SL�ArNjl(�C�&� ���	2�26��z{ v�m3�+��@�}�/�O\�*�˭�򵬦?gG�y,F�s��y,��T̆ϓn��،���䨵{z��А1��t�rD�)c{����b"�unp��\�0
o�!+��'�������o�N*��%���� ��~oھ9�o�qض��X��H�#��T�C�w+p[�yA�W��|W��E��;��*��#Y�cHwk���f|/���^<��%͕�Z�$?��)�H!���QP�f\d2��KGr��:���R[�#�-}���B�7�O���Tx�!-m��_�����0�u;���A�8e�Y�����&�n����L1��Tdq��/^��&�m�C�-,��m֘���٢H��/��
"
F(h��%~��b,�l�s�Q>�k'���SGj��߯�����jh"�͘�J�!c����8�T��-�Җ�4�
���"ȧ�^`.ŉy��1��.DnW ��z���J7˕���W��6�ٯ]H�I�(oLeZ�&~��Q��)�!�o{�����Zk�$�!��J�q�We�vqԏ%���>=�z8�+�}�IE�TG���yh�3���O�����N������07)���\���,���N���1�|���I�7��Ņ|���L�?����+	*�g$_���N=�c�6��۷e�`�,�|��5���zЖ'�;r��Rvڱ� ��1WM�e���+t�J����0@~](�J��Fi�Sž��7����jE�J>1rܦ���#�� @���C��j�����V8��45���8Կ�:A�W��E��.��6!��>�ސ��Ɒ#�����y��>�����3�9�Ưy�HQ�F㊳mAy����z��{��{��L���F�]��hav+R�aܒ��������B�?��ه��spa(��N��O����v��nM��^�����S~����~}��1��X��[q�u�a��7��?��+��ك�aM@Q��k�֎I̮$�T�#��ҝ��^Á�h�d�f�u��t2+'C��j(d[eN�+jXv۰o�P�)x�+ܶ\�����&�d!�G�u;CtG�N�<<����[ RB�7�G]�M�Y�?/<Xry�Vn\Z��w�;I��A-�ql{il�	'աB��P�
���F��YOɼ1޺����]�r-5bEn��,f>i_�H�2{Ls��:��L���Ҝ��N(r��H0K�(�FƵ����������p���W�LE�E��ӏw&v����-b6��σ�Vq�직�/TZ,��Ǩ�Hc�����KOep�A��ӵ�ԇSog�X^|����
�+؅�u���V��;��iQ�kKN�φ��V?��3a����ǇsT���{IE���[�������m��@�)� R嬵}�S�I��&��胪���2k�-���t���Y
X9��͆E�a��Ə��.�D�Hd�Y7��Iވ��7���l��7��&�$I(snQ}z��Ǳ'���jj�	*z�k�gm�VD�u��^/�[���U�d�Z�ۤZ1SҦ�%/�
���;Z�q����z�in�!$�,n�ˈ5B�tZ����������ʈ$j��������\b�`�_� f��+��
%4�֧\�ɘ����9���^)�HιΞ�H����(�< kx:�־M�e	-�8�~̝��b2��m���g�_g��@���W�/�/N����{��`9YR��r�Jᤋy�x���ƙo�<C��Wσ� ~�'�!2߯A��`F �&p/	�4k�nJY�}��βm�B�p��G��jAtG���A8���_��8&�F���-��{��m���-EVΟ��YU��k0� ���Zy��-oO"��*¯�,�埯��Nw&�2���L��%+s�v�><���0{  h9|�#���\B6<Dy/gmO�QL��,���o;���N�W�Y����|� �4�eKb:}��7��]�^d�U�f�1ӪO*w�,����;Z�(��`Ht�4 ��wt�GJj��a07Қ��"�׵�k@4���%����u0#��;Q�y��L�����P��v���kP^�-%z8A���sdIS��6
��ڻ�"�	�,�|�JK�FL'���3�+��x̦_f�VǷ�**����&����3��2����"�_~^Sˌ��\Pu�F*��
�ʑZs=rLL(�y��9�\���D#�D��Lt��dT�V���>�Ӄ�'|���^m8LWA�f:�V�J�f�k,����%i�	%����L��{������&�#�|-@��iJ|�3�?�-��h��o��1EH�ɊR�|M"G�ɶ�Ʃ!B�s�O����|�p{
���S� >��mʿ�B�x��D����vp譆D�uٞ�P�b~C�L�HpD�����&�4��%���S ��g1gK���ѩ0�S�/���ٕm������C�	Y�W:kl�?>!� '�릶� o�5��GP��J�٣��SZ��Gφ�Yf����,n[F����o�nF^��3���|	ԣ��U��6�Y�Y��6,~����j�ċ��rKH^�2nЌn���!�}���?,�%�Eޓ�b'`)�:���(��Rm!�B8�vm��|eЊ�f��R�hG�?��J9�?���4ӽ���tu?:�l��G�eL����r��P��"壃R��;{�6�!ڝΜ���*zĢ�E%>(��>"2�Q׫�!���9#Ŋg�$����^��m���ckc�Q�!���@�z�⾐�-��&;��a�Aqk�r7�'Q�It�;��l��vT?��A���`ϑ�2���x�F�!Đ=a��[[i<of��	rD�sZqK�ȿ<��~#���\�5T�
!�C�4R1���e�]�U&wI��s���t\%�<�-/I���V�;\+b�n�gZ�?���U�����یed&����+�^mE~���%e���X��|�{��1�1���Īm�Tc_f}����6W$xŝ��>D�&��V����v�-��{33A�`�M-���&rӘwN(zr�{�QdZ a�+�!��|%�@� w��n68V��FF�ϱ�J �Xht�8ĞZ�o�`G��|�v��{w>r̋p����:� ��'U��l2\!ZD6x1]9�X4exww�u�
">��c��r��c{��0ԙ�6��'����C�"��ee{�o�-�\El&�ji����6R�#�Ԑv�R;��A?���u)H��fk�[L�S�sC�Yy�=� n*�tۡ�b��ECF����������@�[�r:��}���d�8�����Xt0�ؒ�>�y��� I
��fQl�L�r}y��-�x}��C��13�L�8y
����U6w��ӌn�]�K�Q���{l�/L ��A�+踠�c~����i
$��f?�VU�qO��G��e��U�,����3(�PF��h�����;�R'`�Z��� E��"7r�+����}N��W�=��м��=e�}�a�;�H�+n��jp=�a)��P�GG�]�����"�Ͱ(�[G;�������̀iU�=io:B�b�=�{���]�g��^��9�p����ti���7��m�QT�[�[�����H�/Ȋ�|�_����#�&�2H`�w:H�`�Tr�,����H (�Oa�b���j֊��{����,��C��Y���}3����4�w��<��?�;��[�^�L�n�Q��.�-0T��G��h d������
?���M�q-��$���!���ߠ�E������~-
�CH<�t�f��N�^�; Z�:G��=tK��S$��>���M�����Q*�^-�
���Ǵp���I�eU�:��U�OS|�ć2T���j�22��-W	1��R�ؖ�'1��N��n���q� "��i���!������a`G[#�Ҕ�8ar�X���j/ri��ޗ�>�ť�&ĸ�8vu�n�b?�_��Յd�eQ+�-��b�M����T���`�؉���p�9kK�DN]��f�Y��s�B{�IS�N��p.:�B�y�����Y���������W��)��Q�^��#�gf���l��BS`��gb	�OՅ[��l���YV�a#�#���Wm�Bz���.dwy=�Went�a�F���h��"�_�4�#v��F�����#K����^���PМJ\T���_o �Z��3��v�*l׍�M퓚�������ۇW-z����G��^L���Y~�v	�I�G�-.T^.��2��6�a<B����w��&���� ���^��@����բ.� �P���*ƐGxX	�a3���W��%��8�q�� G.(&60*a��K�Gh��Fe5�)1I�2'�CGN)c���h�"���j.���0`y��� \�j�z��W �˧c:��{r%.�F<���x��4Щތm4z�X'K��Vd�Q-����#"��od�!<��ͭ�0�sO#����]���ca�����)���6J�:�Dܗɓ`w�/X�2�.&Ǭ���D��s�'�L�z��L#|IBwH�D�?�O�Bܛ�b����c,tA�D���,Jp������	u���;4�?>	��x�8� $����d�c~�qR�[�
/����CY� -�h����]b�>i.�2�2]\�0= Q��2̅����d?���`���>@�w��ZPH�-}��ԑb>P G��N�k�h(�K��^���d�a�Y�2|�ۢ|�t:'�W��.q�i��h{� ���J8�j��{��+�u��++��4��E�N+s;��˂' �6��]_v�-,�/9�g�Q�����;�&O��ȋ?=��W������s.av��� 3�e� i��k��Z�F�mFņ8�Z������4W(�Ë�R�H�L�q�P��1�`X�J��;a�ʊ��8�I���eU}�?N��mɧ����:���sn!����e�y�~bTV�$���q�&!��(�����Fti�)�k�����8!w�itŴ9���;I��r8�������>a�FEӯgaD@8�q���L�>p�Ś�i<�ѻ�>rS�|%�ī�#���n���f�,S��Iܐe�؅��r
��%ud�l%�� �m�^ 	����]�5�VF�KhE��w�.d�.��yY�NS(rs��Í�k������,�g�φ�lЇ|��ZLքѼ5>�t�!� M��߮�HO0QTOѭ��v�vmp�Ch��D3ɛ��P�I	KB��z��K��ХV����g3qTX����].�쐊���%�΁}`ZoD�&oF��{GO>u����r��Լ	z�:�/;��\�E�N%� {��JC��٦4�{~�����4�{1�էnS�??���T�$3�����o7$*Cg�2�@Ƌu�/����r$�hs����@��]So'���U2Z⯒x�m��̸��;��pc����@�썢)�(\~0��V��✰�X��o5vS#F1�����<��T�k��Ԝ�Z
��uj�G��L��ZU3�}v��]�hH��x�7�P�� ���ǟ�k�f8���2b��?�׹�:t�ݡ)e���u�A-Hp+8��H�-�X<='?��'�/o��i��;l���@a��Y�!�Dwo@�Q��u�|��`�yU���f�4B���l8L���W:�M��-��������`RP'�S�k�P�^m]Xۘh��M� <������$���Y�_��0V��^'�3�}I=��ؿZ��Yq���IJp0�m��;۞8r�ۈ�,0͓���p��P).h(���^�aN�	`���gll�g�X��'kѻD�%��_{��3cXv�t��Q`�XVkh��+����4�>��h'J�����JiuJنk�'��i��M���k[�c���^XC*��Az��D�(Y�|w�d!Wu�Kq�]�����ߟ� �r��g:H��y�f�#=�#��c
iݫ~���qx��w�P�P���q�kd�FkW�`\nyO|P�|�{��U;�)%��}��Ɉ�(����m_�T�U �v���J�&3��>o�t�~.��~�	z���N��)���޶�|ʢ�
ZC2��� E��o'���#�KHt�شy-��5�2
��˔K���=�8?�C��Z��8&�|��Z�����������QP��7JQ���g���xn.�2��q1�>�\ ���2Wn�5ԏ3M�	Κh��DeQ����	�*��~��w'iPB��ety ]Cd*��I�c �7	[�o.�׵n_/�VvoXa�^1��e2�x����9Q�$1hbrւE`��^�!��?�)1����@]��LO������z_�e�oR��[�~Z�m�7O�1�Wr @Q?7�D � �Zo8��eΓ���B��
�	��3	#Đ%����C����^[ �ş�G��5yg�:�`������/�B�3��uT�	8�d>D�p�I����Τ߷o�i���d���T����,i��u������=���j�Ad���嬌l_�捱vٞ\�Y���?�϶m�/㮯���K����۾���Ki�#��@%?�a�6���i�?[���x;�������@�Y���4xx�Z)M�!��솀�
�����1��	+�m��7|V`U���z�%is�r�j��I�1�V�� ��$�>��>s���8s D�m#��}����#?��5�˫��l��O�Ͻ����[���Q�b�}+��s]kΛ$���O�5 �oz�+|?�.�(���h��::YXu�&�T���w���Ϡj��[�ܷ6� �����}���؛}�!y�hW
br������ͷ�K�29��>.Y�v�/aT����5�ܒ�:��W����6�cBq��T�q�-����V���U��-~�0��$����V=[O�#ytW�M�m;`C����R�R��`�)�I2��oH��mB�	�m+CǒaME��A�a��$����㓖�cD�����^���`��}{yM�iQ�cCj%�M��������zOL�≇�d��U��ҩb�cƵ~� ʟ ?�����\����(Q�M��l5���v�[�:���ͭ� ƣ��i^8���v�<���XҘnX(x`����0��R���{p��GQ�L�{T��֋���i\t�N<�8��Bɥl�j��F-��1Mf�n'.	��S�di� 1�H���b��!��zUd�J� x�ٻJ
� 4�'*��teCI����l����Ֆ7h��,�!n��g� ���2hCs��EhGR �l�L�"�����x<����F�����at��o�D�<����!�j���>1�3���H^��B����sc+��DD�"�8^��|��.eT�p���1���Q3�h���NM�p�����`��q_Vd��W"�L�&e��8ϝ�a\\��M�Xե��x�l!x4���8�[�#�2^����x�l�dv�h��g�Y���������T�J��2�"�<�K�C��722g�}�����n����#��qב�9}8�����,�eZ.� �l!ˢ2`�1����H4��ߥqS�_9C��S��+���K0��񏵼'���jqI�;�Ib+.󵢬þ��i�!
�/��9&��f�n���ne@����_��ц������U��Nɼf���� �����K�[����;�:���)������r��Q�<s^©V/v[~qO��:e�e��ܴJ�k������u�������Â$�d�S� `�P+i��?����G��0��g~t��!�)�&����ḅ��.��j��V#�\�\�UBu��	�6%}
!��J�"�r�f��Vdw��vU�����Eu��m�p��D�V՜?��} 0�=A���̣���h�����7����+rq��A^�b��i#c�U��E��_Ԙ?ѻ�s6��͈���j��h�v��/��q0Ú���Y�T4�&�E��Z�΀<sL�^F����5��(4��cO���-��2c� �/��Y_��D�Ho�UJ��� �'(�hi`�)$���A<LJ�������c׺��b,ex���fZ%��?���$��l�V8f�Ҽ	R)T�aS������ʀ�AgC����^��+"y�o���ߙ�Ub�6F �v�]���A�B8h�:s�O$\2�8�n�3+�Μ<c
����h�Mn�A�Ϥ��D`}q??TV�/~�wk�W�+�G0��&�@��$|���z��B�]�P�K�������H'f������%��x̌��ҋ��Ą8�b�{F���z���K�M�����!�'�j����e��[�o�M�dqU�*A7��μ��F��2i+��TMB '��m���=����n��%(鋒~�/���uO����P���.�ǻ�~۴0�����X}��a�[sX7���yK]k:˓ہK%-e4�ޖ���G�MrC�?�\̴I��k�Y/��~1a�{��s��hL2��<SBB�罝�o:8���M�&��Ĳ��] ġ���w0�]�6A��j�*��gH��*��>��o5&������f�Ԯ��G��v}��j����/�9]{S�s�6�b��9����V�����)�s��=�_��S���Bjbװ�Mw2�^!� ��E#�F�'��I&u���ip��3��8nw��#��Ǎb�EK�D�[�M�xq�[S�S]T�4�z߻�[:�>y������ຶ�j9k ��3��|#��'x���0�2ş���9�4��p����nh�I�:�u�pqh���������<�S�Z�]�e��Jv����B��c�n߉OAe�y.�K��\�8���oȐ3���浺�'
�ٱ��V<�Y�`T�L�"��bK�+`J>�#
vK�����6�\R��&��=$b�����mH��ƫ�w��=�k�͟|�N�%���ۆ�*��yi��_Σ���Y�O����nZ�o�����d�o��AT�B�rju�ǀ�?f�A�g�JX�����s*{9v�BO>�5XO˫gf:	G���f���3C��i���������cDK��`���ތ{���=�J���]& �P�ە�����/��`9+^��A�T�Z�-<������v�ج��:�:7�2�[)ʊ�qv���i@�G��P���$�u�S2m������0�֪ђ7uI�Ԉd�[�F;�#U�E�%c;�8���]�u���~�/�������r�$�H��H��{\ v�\D�����O�W�MNi1�o�DiM�VHp;EW'JRv���1	~��;��u`U Y)U�*����{�Ŗ9�j]�?�����Y悕��,||��+e���[��,*�~֛'
$�o��|����j�(iZKB�az}M�!<W:ϘL��@���h�Z�h��سcBMdt�2~٣��;����p�z?�a�t����.��j�j���]�-�PR��0��+͐��I�d��9W�h� �>�m�a�FY�Sa�wgX����0��7m7���;Cb��G�w�mg�����Tg��νO58l�V�ռ#�1�`W�߰AHk��0]�Q9F��=��^T�:k%ؔjb���ތ&�+Ig�����,#LR�i��93j��2�U�Pj`hM�&r:đ�Nn|AjN��*��,̓�9H�tL=�k<��m�a�8r���R6�3l���Qh�}M�P����]�����䶋W)�iIXU��4�gZ��i���u�C�&������:]Í�_	���ߛ- �����췑�'�����Mk��E*�xq�u� ���Y�E�f���}�e�8k�"����4���PK��R
C�R���f����/Y���k���W@�J�	H�9�^��(RnхҬ�!9^��k�_�	�t��{�׏�2p�:�4Lo�f�}��>�����:0J���P7�!��A{�D�����&�刉5	�L��M�[ΏU�s��3��l�Ŵ/wo�ۼ����ȑ�cA�-�o.�A��)n������uRlŻ���������������5*W
�5���$��G��ǆ�Mo�Ev�r��I�0�p"��z9�}$.`P� �7m
P ���d
~U��ik��|8�Z�gs�����$9��/��v9���i�����W�4X�3����赍=9rB��r9eBN���sH�R�jtf�4�!�P0�D)�:_���F�0dG���g:n&�ɟY���.�v�dw?@C��a=4��Ak��C�x����c"��b���P�_A�t�<>BSRc�v5��b�~
�Q��ohr�T���U�Ɇ�m��|g��*#架��%�Eؖ�Sk�Џ�wc%��v�|�y»N8/��'6�P�<���Z�s�],�ӏ����d��g�L[�R&�eφ'�ri%�&���m,�=Z�3[8��Z/��wZ!BIF3�k��B��,�Z�"9_�@g���{^���~)��ף5�,��v`p�h.�	��!���0RU��v4��~��th�)�@�i��������6d�0A�3����Ǻċ/lrv���"�#Zlij���4
�ư~|�:�>��	p_�a���c�"��(~ҏ�V��$���z���K(z��}�ʼ���OO�f.�4't� :Z�8�0�ՙ�9�׿s�u��ZC;��a 6bÞ7ͤJ=��,��<�5�{Q��@��ꈓ��`��Nj�/f�Z������c+�����ͭ��P�ʞ>�̇�er<!RT��o�/�!S�·Bߥ�Pxe�����Jdϐ�Į,(�>�`�ø�c���8*�!;{��2�NL�?Q��Gg�(�Q
32�ynڞ��q��Yn���Q�2r�3�\����5�0�⯘Q��g���`�N��nh#F�y��^�p-
kE&-��wxʸ�o�q;:�:�B\�j:���8�XH�Y/��;V>���Fn8��T߷�f�x+��WT�_��F��]��+�����y�U��M��Op`�7���ż�}�+o���y:I��>�3��E�ߛ���43ZA~�����������.���)T0���3��]�� ��}����e�u�mGSL�+��,�L�<�j�&�;�@Ff��N��v�PS�;U�H��#�Z�
��r��z'Ly�
/��Xa�c���39=�,��+��-��"��]���~�Y�5��)
*ԏ�^c��� �8��cQ
X��Wy��`T#����)e��'�<UIE�-}��m���>|�q �~"��CW���A1�.��w�b��"���/0�b�!wf��	�d{�����1�ק�f��t�P�0L����y�)���.Ҫw�H]�y�
eQ�c�)͌	�ᫀ%���Z<�^�;���M�gX��ؓ��$ǽ���_�%gǪ�g�4|C&�N����)��^�Z.̌u�F�3ɉ,�+�L�+t�� SA��6Ȼ3	tĂY=D�a:Γ�������<��.�RG�']p���e�|�c	�	�h�@�|A����b4-J�����/��,�&P����ɟM�����mj�QW>�5H��|���"��M@ȵ�=�#��= ��������B�'�e�R��N$:C��ƃ��Ǆ�z�A�ΐ6s���Y�٘\�k4%YW�N�x���rROW5��q��Q�� �+|U�^Q�3���֌6��L�o��ƚ�u:'durt8���S"`������7�z�]	�4��l�?>�Hk�͝���#x=��~ܮ0m�5G������N�v��h��;y�;���G�}J��:���'t�Rϱ��B$�����#��9�VJ��x6%(''��t�a��l��#�>�^}*Q ��A��H�ʵ����9�0�}��ZK?d��.��������æm�s/T����T
7uM$��F9R�U#ȵ�f0�4�Q(f�q�C0c�`�u���j9L�re(�R�¬�ma3�OZ�ھ���=�0`����!{��׃��t����TU?v"�z��6��� ��m�����,i�x89�S4�M��tPu��\+�aZ�1����"V��]�v��֞k��/�s�]zY��?�;�"�i�w�>�	!���_ʣm;��W��rnGs0?�9f�۷#��*����m����Yf\e�o)��hL�T�\��F��/6D (����g���V^��;��o4�:��<�"�fǦ�.A{e�}$/�����������?�C��NKx�"�ԝ����m\����q�oMk�����-!ac4����pp�K���@W���[o��BtJ$�Dw9��7w7|�����1A{�Ԩ5������ώ�%�Ď$�źi��#����vKi��D�A�`�D��I�J
}:�N�ڴ���i�YT'@�����2r�U�E�\J� �Ӫ}�O��˖h�g��zHJ�%� cgO���6<��=3�����Y܂��-$����3� .��x4A�GaUG�G����o�~�/�b���	��^3<d�!��n}�s�y{w۷�*�"�ZKc��?軙QjKD��J�"�M"˸;�VpKأtb*yg�F�{�j�I��S3� -jlRР<٫}��sfso�&EO�]4��JK۞�4"R�Q�dϑ�[B�vYF��>
�=��.�6���#8�E����i:�hpt�H5���3=sB��2f�nz6`��$W��'�>��%������`/��KyCL�uSn���^`�j�����I����c�;��3Ժ���ӈ��{V�	�H��L�o�`eL�?a���9�u\Ė'�ٻ	�Ë����A(�ۨl��ѡ۝���(;��\�K�4���
����t_����H��qg��g*DC<! A��Y��'0�2>�����%W�i�D�Ͼ�~8T~>>V�~�ID���t3��N@���غ�'-	4��1`�1;��f��T���խh���/�W�)g���e�ڏ�}�x��9�\zXY���ɒ`��W��sZ�[XSW��gi��d�U97�e'�&c
)��*�@�h�݉X�7��Su�w%��R_"����$��w�@FQ�8�!LHW>��\Rk��$��@�nI
M���(%bޭ��[�u�F�ʇ����?�� �h]�n�M*`�.�g\yW㽤��\s /�ƪ�7<g�������E#w���ʈ||��{�ñ�Ҷ�{��MO�`%W��'�i�����@�ݠNa��(
Ti����I���:��´��/�`��oVn.���A�\(4��0�
����\x��O�*�I��]>������^������]��n2:� df�Z%x!�U d��=׵�m�[��|[��]Kw������CN����px�"��@o���}ku�9*��$Z_^ej��:�����۲[�"�q�J��}���^��[0�u���(Uo7����Hi�D�{�� a}M:���}�B����ZŨ�4x��V99���8���ݼ��پ�������e�ء�i}̂�ǹ(,f�c.}�9G�ޞܽ���o:a�Y�'��ak%Q�d�%{u���ߜ�'�s0D�����6�P�h�)3��RښV�;\��U���4)�	 � �5���-�n����ή��k+��K\�9+4�<qK0�Y������ߪm�0�Z�VT�`��*c��J8����	���Fg�ߪ1��مBq�:]�]q�����l^��F�ܿ��G�L������
'_ٽ/\�@�3؟n�[ZGx~'���,`p!����%�Z�rn"Z	�U48�a����[G����e��?�9y�{�B��KS[^Sl�����f>��|ܗrT���C%PѼ�]u���g��}��<t�v���b^?R�j\�e�����t���>+�L�j.�N�#�2������9���ڝP�1[@��y5���(@��,�$3�ŕ�&$~�x뜢��#f�ݖw�խ�� r̝e�xO#��:�i
�d�>d���X���3�ɖZ��n���6�pQy`N�.�}�M��0�w�e��7������V���J�:�����=��4�)^� ��F�5 �j�.��Z��p����-��Ňh:D���IE�"�T�� $��-��N���������X�i$8�e+LQg��ʏ���w���Mf(g䆪=���]��U���/ W�x���X}�?J��55�"��صݢ_&�"OG����΄e�T�0MF�P�5��ؒ� v�F��=���$��){�����@O�,b&)���.��
���[�0�f�g8����q�'�n7a�*�� <��|�ի�7���.����=��ߢ�ER��H���zEkxhC�8M���P�'?@�X�E����bF�br��沾�Ac�����������]���E�s���$���)n��@3�&H
�t�A��&޻�YK>%���W�u.���sµ��`$M�xk��r��˧��<#����w��~}��~���<�ٲ=��v�:��q���;�]�?�q]����L���\��<�I8g�RX�\ث����e�*��0��5��ipT5$����Ov�%�`#�!*���2��=>�߻���8%�U�7�����6F�$o1?�?�>��S<�Bh���؅�
NW ��o�eH�G�=Ɗ��X]u�Pӆ�=W���|�t����!k�?�p�iʰqH�R��>�)ׄ��g�MX6{�0m#JP{�j�DQΥ��viR�`��θL#�M� j�뀰��jOE� �D�3�7�������,�9������\�a�j`��5V;R�Ij�����H�!͎�mz>"13���{�/��7/��뚸.�[�x�#\�4d�8+ƀ�'`�c���{����q F��8����B�VQ��f��Oo?38#�ҟ�3�>Sl�Tt�/� vS-y��2�G���1\b�u����#|4S#�A<Z'���  ۘ��Rg�y�*,M��3�[q���!sY�~qk�hue}綦Ek��.��q�����0!~�q<�l����EFo���<Գ�Nr�SVcZ.�ޥ�H��5;�/o%��sm��gRXRJe
����ߪ~-�a�Ġ Eﱓ�P� ��m��L��k���sϚLj�.4�T���6Q�=	��׮x�&w3R�_��#f[�t��E���}*�j(��ǚG{��l�t�j�����H���m܏���?1���l+���,�̆Of��)�+�/�7�e�YJ�b"�1*A��Z���i��1�1s~/IK�@��ME���_��V��7��>I �(�J��4��O�#�w��l�=gą�^Q��|�U�J�u�B��>��lB5�R+�K��L��Կ���s,��ങ1#�U;/�CqM��r����6N��k�ս�A!^���͚�HUA{����m�H]��j��]�F�i���>�j�L�iAxD`W��۶�W�o[S,<�mūk��G�Y������Q\)�v_�z-r�X�n1��0�](�e�:�*�g���u�E�;�9�p���ˀ4&�B�>��9��aF�;^��SK+�<ŉJxji��;D�_�o���m�F9WPT�:qO?L�Mv�ʺՑ;�.���xa����Lnd,6�7$Ֆj�:��ذޝA���bJi�5�E��1���r���D�a����p�<��Fo.|�H�8���Zug��i`��^��+Ty0�iP�P����ύn���u�K�A�:��W�l��Y$u߷�P�+�V9i�;rPh��S��
����!����K���B�H>|����'�p�\u����g_�60K����T �h��YƗ�7�&vĬ�f;G&���&g[�=�λ�g���G�k\?�s6,틷��?�9ud_b:�\ jE?}�tB�nB�Ք��]͎�E���LA_��JQW��Sڭ�6,N@�"?٥J0D�� 0��3���mZbG銢2v��~���+(�RǁL8B��{���uR	G1FH�8��c�S��u��ZaYa���~�'5u=����I��΂��9�m�$!����Nj���;e(�W�r�M�
�C���s����C�?h�㗰��jE٩M���N��������o�3�yxHO�9*`MgA�f���+!`'\�(�c/4Z��;^����JU��J��<�N�B��;���o�};TO�ї�պZ����i��DīE�T�Oˬ �{*��"H���M�<6�[:�X}i��z�cLY�A��؜��f�k�gXΪcѩ<�(���Ʉ[�,34G���ֻti�O�3���Y��`_0l�^(��"��9��(7�߇ B0uI.��&�~V ��p.����^�=�����F������{�=����}f.c�}R� ��ݩ�(zU�8�=�ebd�U�j�nb��`�~�k�0��'������N��b�?ʙV��(Kv�M���<\�!��Y�K�&��T�L	tyJ�}gusl�ś�����nG����.���ы��,s�b��
��a��-�&�N�������/J�.α�dܰ�Y�%�X�pt�Ì]��#W���	��z�Ҽ�E�������:}uY�������\��L5T
���V�
�M�]!-��U������x�bl����FWz�Rq��a{�KF�;~�yL~=�6-�{c���({Ej]��f��(rB9^����Yh,�Zg�������ȁ_���Ri��^�Y�O���&{����y�qpթ���w=�^a�8-xq�;�7u�j�	m��q	�v49���f�%�O�����e���u�����*�J���C�H�]�>�2�{.鴵�b���!-2z,����!_ 9�*��������^��M��������z�I~SN�H����R4g|�S����lWb�ӕ�N��j���%@~x��>���Ţ�w-	�[3[l