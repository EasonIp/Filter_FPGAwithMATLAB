��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$��\�2����]�Π�p��1:|�Ğ#b�,z?�S��x^ %}����g	ZV�l�	`�+}%ύ���{C�Zx�I��ט/��H�?t�D�-$.3c�����|C�Ð(Sڐs��	"q��yPd]r�\���ŭ��� ��|�gtV��j�vhÞfk�ÿB��ƺ!j��w�B��Ң�j0c�'qI�Pm9)0�^��ZE�s\w"	� q',zEK�rRΒ�i9�J�
���D=�zQ}����h]�
�p��D��3Ux��,M��/�#ـb�WL��
���T\I�`�������=��ݨ�@1�/#s��#���R/�@�R̒�Io�m)�z����`�D�^P5Ax&�a�K\m}���VNz�I�x*��y��Ә/7��LZ�����x���@�<����<�B���2$����p G߉C��F��Q�������{U�|(�\� 6�ڀL�k;:����f̂��H�����M���j_;��SJ���3hI�BA���MN��<w"��a�^�a�<�d?TPX��p��M#H*y��|T��Y���	��W	�3���_@
�uو?��z�����lx�E[o�3��ﺥD<��Ҡ� k�?M����`��A';0�
L��ɾq�T����4�Nh�Hyw�x�}���DC9.螵��������P��2NP�T#X�M�W�]9k�{Vm H�/�e��!Dm �d#{*k�Y��A[��:��4�r�7Ğ����>�*��Ʒ��X��������х������ya*䜏�>^�v�iZ�`�V�S��X+�b�r�V}�ޚ���=$R �,.�(�������K���B�&���A�����"��Z�J�mZi�P�OAY�$��^>e����JD8(�H�6����B�:���T3���8������K�B3������p{N���?�/�Ro�i�����&�x�־v���=75����Cآ��	E�Z�g��)o&�����xeņ�2ed�,�,{��S�7u����t��,
z=�n�N�L��l�v2�!&��q`p��E]�Ii�+Ñ����=�6�lU��h�/%�v ���
F�ǎ@��37�w]���^���	)4�+J����{������&f +�lr�ܟg�4)�=��x���+q�
���v �{����`.���S�Q�*��n �c-TX{(�����Eg�,ᇞ�rt�k�k,��[��'g�j҃�N�A"�K��.���b��~t��GAl6OK���p���m!��=�Ô�҆�/�Y���ܙ�i7�m�a��Q�v(&�I;zJ���y�V�w�U���� F���l�5�D��UT�Ѡ?{tg#�'�enu��=W���E�+�[w7��ҟhh�8]!m f�c
ʿ�̧�;�F-����B��6�Z͜τ�oݫ��N鋂�ir���]X	��+�l1�� #9�,��`]�ϻ,�D)��@��3���sd�M~khaj��6l�/y��Z��0��:aW!>�{��uɢ��>5L�q~c�o���|z�0��@�S��v�`�g��2��L�,�iU�3��SsP�v�=B��L��R<�3	�U���:���Q]ؼs��+��U��H{|�(�i��DD)��%�U{���V�@U����8�!�*�}zeO�LĂ�>��u
6m�#;��
}͎qL�(�oR3�ȡ�nh���7\�a���}]��V��n���Ҹ�����$�q}�*ɷ@xU�jD<�X"&d�~͇&t]���'I��$��g`��^DE�]���`�b$At���i푎 ��)N8.,�Mq�eM��yv6P?����;�eX�:��m9I�c0� ���������̆�!��Hc��44��ǆ�{=z��g�D�KxOw��w����S���I�&Je��I��59ސq�����e���6���%��/O����os�J�����5IE?�8E� A�RT���G ��Mn��3n��#�!R֥qR�H�LOҨ�	#�R�(��)�A8�ho���OpY�0���}�a�l|N��7V��:�9�Ĺ�rʏ^�-�I4?x�����Cu|>p�ܨ��_	���I�C��f���`Uvx�>a/h"��y<L�ྏ�'a��?x]�qBzj�Rܙ�àq�i���a)����4���W��>Y���w�Rk��!�����.m�)�D�:������}�R��(��4�c�YX.l�x�g���:Mp��T����)�^�D�#�J����)Иs�5hr(�Uή5�D�F2²��'��C�d�t�on'���/Gx�|h�ѪAYP���!r��5Ŏ$g�`K��#:��RjR�>�9>Q��Ǒ�ԣ9�9�aU�(Jf��msl�\跹�k�'iTc1@��b/ζ��� Ur_S͛.ѓ��/��V~�=�Y]��Ȟ�(��S�p��	0�~��Ǫ^�vE ��h���ǹ3~��q�
65��a��<DPrc� ���Y։; ><˔�F]<a�>�kM���.O�g��$���k�21��j���{��������|Y���+ꆽ��O�����K#��}���5S�=�屪k}SZ }��jܫ��T�hL����mS�<�{ku8�O���ڤ��|(�̥�ѿwr���;��9Sr.%4�/�R�q�`��"|��Ҡ����Ѓ.�
mm��bY�e�vf͒���bǍ؁��4,j�h�p�r�fY,a��ɫ}����þ=�y$��B6���x�LsC��~�*�y��HTc&@`�F���,��o���O؄z�+I�وj�+ �X��./��B�#�2H��ϊc�UY��]������N���{XH���������O�7�k 2y�����q�G�ܜ������m�������|Y��S�o���	�(�o
`�u)�_����<�#�#u�!<�1L��0o���!�)�T�s��
;u�w!<fȇ�U�8]%J	�B݉�S�ҩ���9%|�2n2�F�-X Fz%������L�*m�����a#F�d?&4^���:&P�Y'�ڰ��|ɜ._��2X���.]��J#Z�p'\%��{S��X҂�05�c��Su�93�r��w�_�����ڑ9��9G*�w(��ͬK��N}��M��)���nE~��^Z�녣�<�����9nx���,����?W3n�1�?����IT�A�*�:A��a��/���2�e��������d�CO^�X��>6�5_������O��;�G��q�X��zV�qK�j��vv���x��=��r�7|g�Ԟ�����+�1{�i��p�(��C�&̡\�hx2���~�xI�A�\��12Q Fw�t�Eq���5@2��2_��E���l
�7���GX�f-6%%0��qg����Z?�C�O�~��d���خ 
S.1�5�弱VE�x�d�� �)@�r�N��qP#�����ç��$ a��j����9˧�f����|%O=82
���ƐcH|a7����1@e�WSIE�D}�Ă�ӷ��%vx�e����~��d]I��|,���F�_��>����.�Jc"��  ���^��h\{�p��^�'����5��M� |�#wx꾦<x�zeJ��9�a��
��PTN�}�<P\$�$�>a�F2�~��ԇ�l�;���d��" Su9u�ܔ��j���2N���T�@�kܟ�S52F��{�I���
�	�P�X��D��񥌚�i�;+r��'Q��Mr�ñ^��x���ˍYl�f�����O�¡��ȱ����j	��M�U#C3�Ԅ�ozx�$۷n
���\r��ڰ�}�u{�:��g?��A����ҹ�k?�0��ie]�tB>!#��۽��*��S��Z�e�19Z�����P�����d:�Y�?Y���9�/v6Q LǊu����@v�We㍷�4[�����}6P� ��lw����4��`xY�Jϛ��H����u]�Q~_L�_$�4-!�y]FC��Z��@��ѱx+�"J4�X�����CກO����D�U�E�PW�8#�"C��è݄Ħu3�TA uF�܌t��I)��V(˜�_G��C��9S	Oo����dO��9]x��>c���?��a�~�N����V����U(�F����� ݢ_D��t�p �����Xzx'�ڄ�|� ʍE6���."�Dq�X��n�����(�3ׂ��a��ia�'e�y�����C`��	����W�l�}��e��L�� ����������:�5 ��hʱ� 	�����/�MK��<'��p��s]��ŗ�hվ�.[�n���+>nn��N�"����y ���zRf�^i�[����]��.t!�7�i͂��<9����9�=o����DX�qJxX���P�ؼ̎\���s.a���e���[�D7�C�U��Eu�r��<>���ԞLkp�:X(�iH�]��E9͚��ֆ��i��t�w�{B�� �ڬ�M�����Ÿ&�4�O�;�	Ԍ�wwY$ݡ�qҟ��l�X�����G� >�@�3!���$��45Onz���)�x�-�&�V�F���f��q4�S=��%� 2�5.��\r7���8k}d���k�;P�N&x���ώ{��}#`��v_݈M��L��'��,S|������r"<��?n�ε�9�����D�f��vu������.��z��d�^�WC�o(���4�=�V���7���@�w��ܧ�%Q'{��N$�4�N��b� �f	�:�{&k��;T��'[�M�p0�F�����-��a�`
��m�4T��Oq�A�L㈑���p}�r�T��-�^`6k	�:��Z�Fe�@�˽�1SB�ѿ2��ǹٛ���7��nU��n�nhY��>~�&�R�jl�0'Uw��G���J���N�@ۇM1"���l�;
\_p��L(�;�Rs�M�t�<�~CINu�[��%m`«�I���r/� c�m�-!1����Nu�9�w�f�����<ȍ�*�����H�~/C�a�0���Z|c���7r̬�r��{�Ҭ��k�-F n1��_7+�d|�T�M\�-���%�9l���g,*���Z����c�#�o���z"��qPY������KG��=��ت�5S��`M:5������b��I����U���&���?�{���!2�/�AWT�hUlb�hc|�gI�Maɬ�7�ӄ�&kqB���&���m2F�*��0���u{W��j�^��"�CB +A�m�!��Ʋ��}
x�lñ�ӹ��{����P��"yE�/=���y���em(���ȱ!�u$l��y�������x��FXv;^M�^�T{����b��W�@�US�g�W�/��e2�=p�ÿ�V�g����(VC���ב���f[AeivE1<�;<=��гӰs=���^[��N�(�̔�}ɅC�u�O0 [�<��F��Jv�M���E(�(ϓ��K�V��h�l��j�4}W-���-��g����rx��������B�h��"U+G���#��2k�mBZ&L��}kX>}Rc�@�)����jǫe!�.���o��R�Ǉ�p)W�&sd�.����?�^�P��-�b�=հ�b\3=b�h�[���ơ]=Y�
)����0�Rq,>��3�su�b��hY�gq���LNN��&u_;����Sz��ig�Z=�8�>ķ�1BSrץ���G�'Mh���X6L�Y�K֕[����aJ�.g�a���=8���_�:��KE�þ^��`�kx/A`(�Ox\�ύ�Y�Lb�;���0�����b%}�oק���樯��,6W0'��L|�R�vp��3�6�$��|��ў?�������y�$�YlwX����)��]�wV�Kuj��kJ�4�l]ڎ��^�gy�4�8�?Z|X����E~*6=�?:M"�w�
�/KRT���@�6� �ׅ�_�!�/�*�#�⧎������.ḥ7�톯z�&����B�Z���
���6�ɑ�B���ݦl&�2�u�f`�8��<'̉H�W.$��e=f�O~�-$]�����`4(ܚx�3R:����}^$�ʁ�-�H�4��A��^#SH�+�z�U:�*���iYdG������
Ai���HD�@�����A4b�����eT��&���Ƿ�1�	{-��xnLk= �H
	..�#�B~P�.�L�\<T�gQ����Y�cf�pE�,4����;�L*`���MV��z"�ܸe�kn,�R�l?�3G����������^K��;�t��y$���������R ���z:Xǜ�X�����_8�U8(�t�W���O�S�����Ē�*=A��{�f�N�B�(L�s�,:M"�1��^�0=�)}�@�sÄ	U-B��w�{�|�!"'��N��?:�C8������xUV��t�b�N���% �;���Mj�M��0�یV�c�6Q�c���.�r8����_/4Č�A��+�����zc繇~��W�G��X(�֞�2o+]4���°�/+4�����J���n)����\���|�beԌ�ȱJ�����Qx���� >�Ĥ�5}�2;�Ø�⋸�Ź�����w�ihPv;�N�wv>41��4�G��ɿ�]��X�7Ik�_%����M	�MaB��v���Yv�{��A�>�p���g�,R�%$Y'y��,�FE̻�v��c�� ,@�'�JmP��O>�!��=�8���ư^z�G�K����S�%�۽����^��Μu�vR�%�?��~����-��3%1�3���*ڇȪB!x��sC��29��'�D%/XV���p�p���7�-�_�������\�d	hP�U��Ά�(|@��9Df�¡D��@���pu�~(�?�������G�=bM��n�P(�2���xDJ�i>��O�(܆�dZ��a��ӷ�x�D�� e�s.Z�3e!��
�xc�$R ����
Bi[��蘌�ki��%�f&2�[;����yzK @7 �U�Vy!=�t8��m��Oi�9URE��O��0���u,T�w<C}����ccV-��@���g�����F�0�ޕ��Y���`jr�/c���H��@�W��H`�YO
�{"2jjS9aV���ף�>�@V�!`z+�P$�,�͞=���X�������]��KaJ�+���ڥ/��1R�g�÷r�W�P'o��0�%�_0�jь2$�Y�������o� ��R����W�y�|��U�mZ-y��H���S���	?��)b��ܣ/�ܰ�t��P���y(�\�+l�����]�;����G���A��2�Da1h�@�pn�cC�	��)�~��Æ��#��F�?�6�Vm]�|��I����RՑ'��z��Bn�=���m�=b�zT���u ���~�E��Y!aĬ&|���X�a�"�~32XB�`�<&�hsj�z�$�ӵP�����iU�e��K�h2��3����
����N�HaT�|C���:��J������!k��q���j��f)r�,�[4�U�A
�s=	n���[�P����[r�k��Ć"tk8��5�64uiN���X��xmG�[��W�9��"&�zÍ47����q�5?�-�v��ћ�\�4�3*O���)��O����n���U�����+�{��O'�"�y�?%{Id-W?�e�<�=��h�MYV�Ǳ<�?nF�<ˀ:xm7Aد����p�_ͬH���4S\:���hfa��W���w[B;�ƟO`D�¦M���%�,��%\�6P�X�n3�f��rW6��"f	4���u3�.�i����lC�X��!��Geiꀱ����S☬��>�")�`�s2��-[>��[3X "�g�����6�*���8��N�O��(�w����:���c�����?�dbIr>�K�m��4��~{��t˱$�	e���CY�ָ{
��� +^�,�Tg�����oé8?�Pu��<����!��h�aY<CڏM�����n��b4h�<6��tZ�V��*4�`��s��2�W�����'��g�X]N�5[�`��<ʑy+�$A<������#Bc
A\p:*I�ױlTu��x�u��M.y�}֭�����\W!K�|�ws�[��9�.�08�#2e�"�k�5q#63�}%hK��x����Li$�EPn�廞%-4����
Grko
)Z�dT�x�G��P�Q�X���OGsb�������B�4;ʙ��7.�ӎ)_
���3���a�3O�16)��[�	3������H�EO�u]�ԭb���/L��٘�M��k0O�R��?�$��T?F�o�X�I_M��h��[��L��� ��ѫj�)lz0�$�I�6��͛��^��A�}����o�}�k�9���͂�#�?}����/-Iq�z�Cp�g����<�Q��ҔC�����|��d� �-N�8OA�>BC����%|b���ϵ{��p�����}b��\�z�� ��
 ���V�;p��9��$
*Xw��Y�d���a��'�k�����s�?�T���ԩ[�;�,�#�f':��n�����d'jVjF%'J(jC�h~��}��u�4�%�����tͶݏ%�nhܔ�Td���c��Z�~�<%�����=�n,W��~��'G�,r�e>ud��f`�����A19A� ����%�G�S.݆��<8�8l�+���P�$���;�8�S���*���9^{�]�"�Hbf��<w˙�7�B?�-7+F�2_<sz�ʺ�T�"A�y�"X��<}�gR����芡���ڌJ��XW;.�F��u�ն��a�*��؟~�]��(
*��x�e�G8/�w��!��I[Fs�q��z(b6;.ϕ�3D-�F��b�J��@Ͱ"֔2��>��)��6��7��?�\��D���G��r#򲐓��������t8I��Ex�����s�����-�)�>#zĺ}b�ʒЄ@pŭq���a��
��b�.d8a@=q����&b��4��"�Y�.|rs-�W- 81$�N����ox��6y�Z,�1 3�R}fI��I��Ԏ��K2���X����#|5�����2�t�B��e7�R�ϰ�S��6�
������UƝwKA B�`���:=Сh�d0�6 ��F��U1�Mh��J9���3�H4{�׾�<W8 ��g��L+�Fo>�t�C���a��4�W�����X��<�\��>���*�:S>�ϴ�aπ�l����{�a����.b|5����f���&������F<yo"��B��d1s�!�ar�~���8�s�K-XXو.>��D���S�>��E.�"�m9�id�Z'��$�K݌�������Do����`���E�
٬�>�8@|�`���G���/�8!T�J�o�|tAalϵ�����ަe75T���I�W:�{&��z𭲾a� \��t���J0����e:"N�3!H���$�橠�g��HgH;�S��\��ܻI�d�t]_&1Z�?F�φ�������!(�b����Or�����R�P!K%ga܏��+���q<9�M>��5l������̔e��Z���3n�a�pwy]�dJ�1+	e�H>�R$�qXW ו �]�	�/�\	r��ɮVg�	�7�f���ހ�{0Wd�?k�6�>pa���{��b@��ž�\E�'lF��5 5ȿ��+��ҥb�6����c�e �#-W\�X�G���[��~Y��M�D^9�y<&�]��c�y����c�4�;�E��Y�T[-��f_f_�o.{�u%A�"�t��O����#T��]����٩�b�����XS��w�JV.�9{��s�O`���'F'��ΡB�'Q�V�ɥ"w���o�����se�/I�~� Npb���l)3I���ւx�&�o^���1֘���n��l��~�'��"��a ���c��?���r�����f��73n�O����х�����C[^��M)H��'5.��h\
����K�~-qwӏS;�S����=� ���f~�g�E��=}(*��"�R᳟C��,AT��>���ZQ��F�b���H�T��4U�Xf�$X)�7���I���N $6�y�u2�U���\�aZg�U< �1J Q�9�9�L!Vj՟E���u]�e/���*��R�&<�2LpF#W�@M�����������8���bg�٥XL�DLF�z�8%
�/.4�P��^�m����B���x�ĵi��r϶��tڦ��n�k��F�3�F�����zU�Y���X䏁AX6:�dJάAх�i������&ȌlҊ�[A�f�
���}����v5H��j8	l2��H�����Z&#�G/S,6�:���Ǯ!�7V;�Q�OtP���cpTn��8<>���c����W8]9V̜��([ɿk��9�wF�;�^}8gR��.3�a6�v	����e�>|�1�~hG��=������7�eɛ���<��)�S���_�ƿn#{ �bڠ<}\���e�|�Ar�?��LW�چ��W�s�d�G�Y��be�N�������,}�1ؘk�@*{c9�%_'M��Lܲ�N��2C.���R�<��&E}�W	J�b�~ܥ� �!��.��W�qR�m�OwR�V;x��K��r�J��zv�K��}VG׭�L:����ЅZc�P	t&D�"6���p��K�15̸κ=��~?�v��qfs7��Uh�(і�綧k�m�� �}�ki�GW�u-E��9�dZ�8X4���@!ero�T�.�e8g"�����e�[bχ��ih������.-����`f��ݘ�KX���r�yr�A��Oc��@��l�a>߼���W��W�+�5n�d�r�T��D��K���k�4�X4x"�<;u̘��`����C`�0VQ�8C��k/#ai������xQ�m>��'���H׏�BԶ�QD>F�(�_,g@F�@�QU�g�)·�1J�:�//AGQ׼�ALo��^C��=����_�Fc�5��U�rc����yY�Κ���[�����������T��_q:��2��~�`���op�2�ʉc�H!6]��z�"�#��?�%��@F�g�s��e��Ӟ�]r�O�:�,�6o�` v]�Z�kgTsg�YR�Ir��}hz��[�Dk�G�|�@ہ���b�ҋ���jp���\R����	ʷZ}�ɳ�6G���5&���Z��v��|�r�.Y�N}~�EB_t�n<z?B��X$ۺ�N�;�ٙO���[��tм��`��O��`���@q/�؆��#��2�8�Bhb�P�`��S�i���]�����k���b�Z�����[f}R�<�l����29����:w.�[�b);^�o@�dE
�
�i�uUFU�zܤAch���#d�6V���8i���D����t��؝�_��K4��5&����[��/$�$��_Ǭ�tU�1n�⺵�B/�ЎU���P=72��[َ��?����~1���pQ'0Aa�+Y�^����t$���;��@`Rh�4����������	���E�B�BJ��%�$8����B��RPV5���4�q,��U�b/0�d���v~/�����3����`��e7D����'���gDM�s(7;��ɕ�,s�֍�x��V����X�Cz
���%��6Bɳ���IЖ�����Yc6�b;�jp� �݉���@jW����i�H=S�CLuI��A�k�Εh�z����ծ�Tl��{�?��c_��7f�t��^��ɽ�t��ȇ\����:4�B��֠&W	Dx(�����y=�a��,}��
�~�3Q�˹��(or�����e ��D��Ԯ;3�^��|�@�yc��/�AP��ંv�g��(2��x�F�pŜ���d�`�)�A��6��P��z�/��
��h�J�����(��H��N�)#�8keI�^�? �N�M�����Q�5m��s҄����yI#U�c�����Œ��˼<��iXs����7�|&W���th�$J_]�P��2^C^)pN�.e�J2:��V�C۔�^��9��˥bC�5(E�ЀcX�����t����\ts>��M�r�̒��v��x	����|��e�k�yxSF����H����t�\sB��+���D����(�V�2�C"����=�2�t��t���Eq��'ܭ�S��L�GaG^�SZ�g��jt�k5u��N*�Xw-U""��?��+��:^7���̩ZUO��c�Z�Q�(�3��`)��������.jO�{	���f��c
�ԝ2�Z���r���{=�M�7��k2N���*$E������y��
��%\®���S�Fn�y��}��,�d��Z��>+6�Y5/��,��w3��O���d[Rm��P��3�uTni�\"��mq
6�W�תer���C�n ��	PMP�V!EC��8�ʊ�n�(@Hl��Ç#��N��oI)�3k~�P�:�6-s��ר]��֤*q�����?�5@�~X���^H��|��_�R��j�<��à>��T�'F�k���B֥�mc��z��m��%|��͗uYx�j��s���޴=&�FZ�A��A3�h�u�T�:���%�V�y4G��\pQar��G�@�hA L�!?(��|�uڸ���С�-�}��9��w�6G��WI�ݑ-��^�7t��^�h�� '3��e�|�σ�ձՀBeH����|l�5x�?o�L�gV���n�	Q�P��`eqg��7J x����ܝ�j}��E�Nb��l�t(�:�����@�	�7�C�u\� !0��S<rψ硣�t��%�)?�L��-e���Njʍ���%�C���QE��y�3͎}�]�:��ehh�yP��Zh�=�_;q�Ub��J�$�ި8<�p;����Y�ެy82d�ٵ�K�,q�#0���.F���e����H_�A]����j�>N�Fю������%�J�FI���Zz�yuFDԴ�@5]�O}P����6C�E�>M��)���� �h]�B�����ۀ����v���&���[�PwP�ۭ�p�F��6X�v�]َ�������$��jN/�K�
	��������-��Uo��Q�����v��$W�Q�T�`$�u�FfG��w%q-�s��3�ҍPu=60�z��I��G�\\�6Tҟ�NFB�'6l�J^��'.��F�!�0��g��^��d��Hn��4|�p��+hⶳ�6g,G����奷y)dW��<�;��� ��1n��f��U�@.�����r{�VQ����V��yw�dϜ�!Л(���,d`�A�p@Mp!�i��2M&�ΰ*���S=:f��걣��[V'9�d�{mp"�񫌺�ɊD�c� �}c�G��cn;C�T���u�3��,�H$t��0T&�5z�y5n%i�^�;�'���8q�}Az�l2z��}��ꉦ�$  �ZQC�x�P~�p��ҕ.֣�Vb�
�E+wr�
`�Q���Y�L.�e$��q\s���>U�h#PE�B�d�=��P��~�O�����U��[J��}����5������rOԷb��V�,�{O�/%�6O��jX-4��41.PQ@�zHK��^�[D���֡Ye��E�_��jh�/c��gb�D*%!ę!�H�}8�?,S����7Qq�>�Fd�m����Z�`W|T���/�.��l���2g^�n�(	��:�>��D��6���wr)�W?�xL�4ܮpʜޝ��ʱ�t[��ٮnW������^)3{+F���3�_�Ģy�#X���q��r���ql�o��G��q/~���O�-^����aү�ԣ��`F���uظѾ��g��\�u������N݁g�n{DY��f���`�Z-Ł�N����y�i��iaK�����STOڦ��ܪ�ƃ�ί�J�1���1�P�x����y���E��Ut���b���	~[��Ľ8�0�����Ԡ������SdQ��V��gyc�R�N���l_�8��ǜ�!����zb��#i#�,�$�O�Υݑ$�׉�
%��x���+�/%aL�OD�BJ�V\'4�O�~��o�Y�PL"ۀ�OLYo����=g:��7"߃��]iB�y��){-Z�A���L��d�)�g�;�b6��>��.�S�lɰ2����wo-�� ���O�!%��G�B����N����BGTv�]Z��z��^�Vy��3.*�ӵ݃ڃ�VT4�����t������/���nNin�.d�f�"��~e�o�\c�Ϝ�b6f�%����0��x���B�8�,MK^ڲ*�]T�t�{DBP6�BW!�Ci�����w���C�DH�sv�En�ECw�҇却��E�h���g�o�W%�ZeT����ߴH��u�$f#��1���}��x��&o]kE��T2�F��V���8a6��B&��Qi{c��Q%��F�_;G�~B�0���n���!9i��H:���/�Vg��#g�N.���49b$v�#~{Yrx�ޒU�HO�$��*�>V[�	ca��7L�HՂf����}e�h�>(hM��d6�0P���V�7��U	%u���a	͉�Ct��M�����t�?"�Ձ�ƥ���Z�p!J �Q� י<��߅��YM�a�3����s)p�Ν��<�4��b�<$P�gى/�\��L�oq�,��<��Ddߔ`��1��_������I�_ d�)3	�/�o�KRE���,��
r(����z��x�a���D>�(��g��(��O;g+s+m[~�x��_l��ds�����Jf;U�� �[�-]�|6hv���i�U���+��R�
�׷0���t9�z>��I�omi��IG��<P1D�~��Ke�#ĳ��^�m��E�m���W����!�p��ސ^'-���8�1�Gޕ@����Q���vi�L�u���zt�.FD H�bb��U�w.(pl�wm�����L�}�}3�e�6dDX��7�% �=#,�Al��!�=|~���y��]����s�o�!Ur�cM����O�wbm���宨���=M��f�Gt�*�`j�)��wQS1A3Y�ȱ���?;�9��y�=,������߾���	� ��z���}E�0����Q�K#PíR����y�3)B3o�[!ꬲ:S,���*��_'I�nKAUNC��-=����՟Im܈S�t�>/��bd���L,[�s�f���$���������7T���[?\�Ph�G�3Z�)?�G�v����O�6�7�C���'�����!�)c?N�Y���6`4#��kܮ�W�Hm���NC� ^W3�Qו:]��!ݱqV��~{Wҩi{������G�%��舞wT<t�c�q�H�h���	���u�G[7�8w��[:���������nP݃�p��fMP�_�Gy�=Z9A1i�٦�����r+�� �59*�i��fA�s_K��1�>r� +��RD�of�}�ص`�θ�ښ�f9
���4�D+�4޶���d�M~��t��3������!��=�DS�����Zu�骼�LԦ�����D��|���*�����M�0�N�8 9��^��!����2��qa���_	^�]NC�BPR�X/�`��5���\/���U�v�.hk�]-��-8��AǠ�9.�ŦO6��X��˃���],�d4m(�g!��wWx�`�W�����΄��9[Ƴ孠�^�̞�]J��Ĉ)Z�~JV�~�PE�Q���� �U���V�x� ���cF��葠�3��P��m0�=��Ђ��ZPQKo��r�%�D��-`��!�NADP�S(A��x�OGL�%���&W�p�K|�`��ST�{>Y���֦�>�\x��}YQ�x��B���n'L��XUo��k.S��)�<����Y���N��-��mt:'�m1޵�]�;��4 $�kW�N������VNH��Ć��n���C=��������W?Z����$.�蠴��:W[Q�1\�S2� S��!�����8�{��^��ݧC��'p\�%A|����y�5��#\�h�.���6p�Uwu�eR����wW~u޾��?'˱t	�ps�dFy%U�˦�?pC�=�S��a����\�1܁�1�0k�Wc�O�-��+~�J��,�	G���r��-,�F��o	����0�t� ~�5�*�͘��+�'Hx���� [�
��Vq}��Xc9:������)�F3$a5�Go�������).�q �	��ȟ�[���Rx����:�Ӭ`(x#��,��?���y��U3µ��+N�����=p�~G�]"?�&�H��o�ĪV�������,�=
��ƽ�J�pו#�:7�#�|2c���������b������r�	
	�bbb���OZś����J��o�J�y8z�om�O��$�bT��}����&�]�:�<��YҠ[u�WhJ	�j��TڦL���͙�	�'�k�E���K�b����?H���� Sv+%qS&���KQ��⥻k6f=F���*Է�3+�]K$�Ŧ��1��h%s�����b%'��K���� �N	��ɟV�7�� �-�����!i�:���A�9h��15�Y�u�h�n�B�L�#��
à߇�B�K��i����2wU�Je:��*�L����7R3>�]8�<Fƶ��|Q�~4��ָ��p���Pc@)��Q�A�(#̃�7rs�xBXg��N�"�`���[��f���.+��J ��Ph!(ڭ"G�[�~.+H:�ٛ��
�p1�Cv0�ZL�	z�n.���Î��v��%V�����<���v��@�+F�|EQt���Zʕn�I���2��)f ^����K��7��+,��
&��+�=�I��o�x\�3�6���0�� �ON����u�)a���d�-X']� � ���vJ|뒖��p�	Vމ5W9�G��c���f�U\�|c����HV�i���N\�7ARi-�qV��/�y�>h'���nLT�{�W�A�i�ۂ
�c�����,�m�-�j����:��9�Ck3���|-�1U����e�"y���,M��weK�{(��Xt�VY�R��Sq�\㋪��Z��������'I���C`|�m��4�w��('+���u��t�}���@�	�2�L��0����ZU�#����:����(:bV�<P=3Ȅ�ɭȮ�eZM`��K�lvH�s�|�n7z�i C�G=�$�=��!� ������ڋ��ț�/>��*�r�>p�����+�t{[�08���L$qJ͛�;]�+�h����6k)¢���] | #9�S�B��0�`.��`V>G�kv��-x���L&̜h~�?����g��� ����ԆH��5B-iEV=���h/"�(5{���V>S�씾�0�Ƙ��l��@�R�lΧ�|�_N�j����c���_�+�^����٘EFe�_i�R�T=۞����6'���}�_J�(����5�������k����u����d�R�'|~����OU$���������<�ծ��5`Ͱa��t�/����{D���Q���8b��|���6��m�G&cL����O���c�w�E����3�0|O�����@E��3d�&�d�G�&��Gfo��Tjf$9�cEֺ�Ф��#�2/IQ"&�Ek��/<3��˦E�X����Gc��٘�h���|c;�g^�9����]�Y��!%Z������y?`�(7<i(H&B|��e��dַ�-�xy�ѢOu-�#x/����TXa�Dyay�zL���1Ո��Fc�=�k�@��� ��ľ�O�-%��S䳘S �NbƯ�
ד����2:cr��*�bӊ�^6T(�(0?�+�(^ycR�9E3Ð�G9X�%��x?��F�"�`i�mо86X�% Ƴ_�T��щ�jCvr�E~No��b�|`��m8�,����,5{���W{����0�"k��S<S�B-V����c� ���?+���);p}���B��m̓�kQ���=��Կ��λ�
�N�Ď�&[���{\�!u�=��5�x�)IY&��?koM[ƤC�.%�续}�џsZ���<���J�2�OC��5`�y ��]�~���Q�
��t`B��k�B�i��/f���H���n�瑐L5�&�c#�NYLz!������O��kK��&��
raǤm�nIB)p�ÿ�]���u�ݩܖԇ柦 � Tf0�8���9۟g��NM�q۹��g��[���Qd�N9 �1�'�p>���t�����D鰓a���cl!�iRD\�F����rq��X�8�4'��s�s�]�ΐ[G1�
UMjm��(Y\ˡ�Eb�{@ۋEL�A�vkb?���������W�7��v<�Y��닯���e����6i�ݜ)���<�K�����ic��Q�e*��7�ٰ�8�)O�Y�3C�u%�Z�X���̰���4w\�=�裿� ��͓[�ߊ�W�).���l���h���<�R�ih։�t�4շ��/p��Ѭ.I\J�ry%�W�2ȋ���/�RT�9�J���x�s�ޚf$?!�]�Ɛ����Gצ�a+_���p%>��*�� 1��g�������\>�.�>?ʩX���ԍ�,����mҥ��k���f>���׺h�KV�pܟ��z�z�?h���(sQk���p���Ǌ��E�M��P����|WTS?��ɂ}��sE�N����&]0��n#Cj�l�D�8x�A��*��_�r���?!�Z��?��uPǑs}�y��3�#=Y$�p6*�*m�hu��H�\T�qj-'\l˔�qyEQ��:���uj����������2lZn�����쩖'mR$�*,jY��,�Ɖq!ˣl�,d�w5ʒ��\CZ�M�2���	�\���X��g��~������I�Z{~��.C8H_�G�eVJH*�kPkA9#<���KsA�u���
>�,ܢ�A����Ucf�<����M���Ʈ5�:��hTQf��d�L�sq)��v���],��)8j���4Q]��튔{��+���ٍ�C9*�$�;a�Y�����'�.����-��&�W�����O=�c��c�W]�	�ƼLո�K���C����%2�!m��D�V�$���`�+V����-r+��c2ՏK fD�+t�ĬV�N��GB�m�䵹�̚�1'It0a����֡�i���X8����u���h�����hG;�i�B*�#
��4�ʡ7	�F"/�;,���lv���_��Z�@�E�{e��<�C����|�8����G-CQB�n<_
�k<��Ň����N�~�J����/�ً8$Qݟ(���)��w�L�oոnC���UQMEO�U���XL'�s�>�0h]�$��Nq�R���,��,�+�@YM5<�}夀mB�����U�i
l6;�(L�0(����Ѓ*d2��o����B/<{."���)Y�aȀM8�l!f�
}-���8"�nJꄮ��̀��=�1]Z8^�N��f�w�އ�@����E+����G��S"����{!
�&�vE��ܟ1U���F;�-�b����#��CFH�s�o����w�.fJN��6�Ĩ����**���m��:t��?�L1w�Αy�"�P;�q\���*C"lL?��q	^B�!"���88?���mM�����Rʉ¥tl�n���Ծ�Z~:��e��!�{��a^�	�����+���;����-#��v��W8��z�"h��8Q��*\v��޳>�1y �V��K��������P�c���]yl���r�c���>Xp�քk�,>@&)�D�~E[�؂���-�m� ���GP����W���Y�J[%sL:%b��rI��ؓ���|�Y��*m���ˌM^�[0���Qj7�:���F׻%5���Vi����r�ղ���"';������l��Q9]��L��X�T�|��F#�p�U��a��>2vN�a7Kt	�Ę~����|��kuQ�^�i������J���鴭mtI����t&o�ԟ�u�2h��P��A���GM-��gN�*����M��Xފ�m��m�!0�R�I���D�"i-O�|�<�i�7�zM	��}���$}��L��}�էu�YKk�ǹ~i�02\yWgH�$L�ޒ #䗴�2�K���k�݈*��T>��v7W�P>��c�	2�s?��9[��&�rč��D�T�.���<����CQ��M���`g���H Z�m��xc��ؼ��R�����jM6z5B��H!J�dΖ�v$���-ﯬ?=��Mo������=�%�Mu�w�G�����1��&����9M�1(<-� �?��x�GXM���1H��0Ɓ�E�z5��-ʽ�`�a��NP}H�@�;M�/�>���"�=�l����e[\�O��Wk��	��TȩR�I�@�f��7��жug��z;2]�~���D�ͽ(E�	��5�Q��lxF`�.t-��,+I�6��<�ظ&���iYr+e�z�pI=i���,<��%wDp���5k�y'Z��d�Vp��<���죽$� �ܣu�Ŵ��>tkb#���&A�ˇ�?䷸�01��a��~�y�d1��NO��M�	��M#W4��G(��ח?�W�Q���!����I�.O�l�l��d>���գ����Xė������_������BK�p֋�o��*_�-�߃eK��Z�Ǟn�5��b��qv·���������PVntbf��3�:�!�d�s)B�(u��"2���$�&���]����vI������;7�w������y�����H�[��S�� #l%'��F^�8S�B]11$�%��O����NGR|���`��=��`�����P��{ �ڒ"��19!�!+�2�~�E`�����W�)�՞�-<˳�Vd)��m���W�i�y�j�/�����J�7F����۳?P��ۦ�W_-�2���Dx�|���n����]�t��ک�"�p��H���%�\Esd�+��1A�/�
�<�Tݻ8Gx�w֔�C"�t^�'�T�d"`�J�Q� �Ve7V��ԥ��[�ҙ�&���{[�}4�sW딦r�}�pFa؛$�mO%�*E�3�eՠ���l8�>0�g3�h\¦wm��$P巑�k "x&�PI-��G��I���>f�'�e�Wk
��~
r�����T�P�黪�ı'�^��$[I��!?�Ar��#�"� |��Au���&�Aa�է�X<x��B�u#� f�{!"��ܭ#2��4� u��O 6�^8��,E2�'X�q0�.?����L�g�z��4|�S;�8ҳƕ]�� kW6<��ʆ�s1��(���t��U:�F̂ҧ�dN�-s
A��y�EP֚��υ,��N�BNq��d���z���/��2v��_�K�+C	����O�	vұ�l�񧨜�<�0U�A榺V�������k���J��d�l���p��r�O�F�Z1q����'�}7�Ik�1�J֠0��$J&!Za�3��Dg�-H&�8�i�+_�8��U���$;�����׃�q%/M�HoF���zy��ܭ�ė�_�M���r|@i	RMܑ��Hw���g�(+�΄q��hU�[�������`��Ii/���V�3Z�ཉD"�w���
Y����Qox���s�.3~R�t�fb*�A��|��G��
�3���o����F��A�w�����K��i� ����Bz����OE�a|�G�A�E��IȀ��LH��E��҆��9��S1/D��ra��C-���V�9.����Q6��/fg��?3Q��{��e|4F�-뜍(���H�9�k����{����6�E[�%YEW�(_���V[M���lh�t}m-$"p<%��%������g�:�9]�e�V흎\���,KP��$*�*η05�����	���n��>�8�֒Q�iz\���� �j��dw��}��xi�f�����S�`f<��f�H�������hC0ϫ�:�jTt���-E�'q`�#-ǻ#�{���N�:���\�l�݆�f���GoA��К�N
�0s��e#w1K�2�XR�&�W%ӟ[�����~����d����5>WDg��7mJ��~��Z�k.��ḇ%��wG�K��+ �ӝ4�DA�P���R���j���TO�\�7��8��>X�D�̲�|�C�>�LJ7*.��1�z���(c\HWNٻ��{�����������OE�M��a�Hަ�c�+���L�t��, ��h�N��j�>b�M?�'�h�G͆��}��}����������	?�s�kѳ��ʓW�j�^]3E�	�,����ѓ�^3���2���.e�������B���j�/h��V(�-���y��N17�wE��N��5�	7�7��[��GX]��s��>Xt� �>�������	sڹ[�_\���y�a1���ɔD|X��R�w�\8m��8�����-��r(�"��'����&�� ���3&[���a ��>O25 ������>�th����Q��lJ�08�;�D�B��09�;(��}��?�ѹ�%!��`v+�џm� ��%�3���Iu��
�Ő�P�T?��U8.�ht�_Z�⨝:Ю�,�KR�Ɂm;X\H?����5�9ۉ�R�v����m̶4�>�5�}��R����_� کwm*3΋�%,t����C�*�{�8}ɫ�N��~��U��w�F���զ��D
W�Z�\�yr#x`���[�fc	�#�y!���6�t�?3����LО\v�m��igr�����B�[o��,I��f��%��A���X"~�(W�ʲ8FĴ��0f9~ɵ�����i�*VH��h��#�-�ϯ	�O�&T��,7~����AlT��^_�E'�֋������3���l�WZڄ��ͥh� �u�D0���k"Z���B�����7zH2��,.Y�w�)˲��u|��t=�}���e��vBx��]oյ�9�H:�Z+��N��I� �mZ�աl}|%����=H��!<����[Vl�S���ɍ��5y�Uyp�"��x�R_. t�E{�͊c��_OԎ��;<�`��� �r坞��	�s��J\4��o���^���S��	�Ǿ*�3�l��L��V2�9y�!҆v�+�[I1�z��ݘ(]��)6�Ň6@�c���䅢 ��֟�4
��'Q<<3�^*kDY��$:H��w�a�^ժM>_ ��|��Lh�sE<���v��.��#��
?z�L�hyވ��D��=w�C�(2wc�T��\������i�,���@���u|)}0dt�[��n��i�ړuI��qcw��1�,s�?�(���bx��Ћ�Y5��=��}��������i9��o�[.���,Nq�#YG?���[��)8S��U��%��Dx�%x~�I�O�y�	�ʀkC���-3xN�=�_{t^�4�
�v F+4�+�D����F��Vꘞtb֡?u�V�U5�\��!���\EV
�j[��� z�?�oC'��2��dV���""	��_���MJ�_AhI>"�k9DPh�T3�� ��'��ۥ=Q��TMl!'�����r_��r��T.����2�O�DX��Wlכ�%��I��,C����a�{��5���B�LL|�Oo:�o��-= z����1c\���u����c��O��C��U�E3��K	Y��i]Y�E���L�I�U��uSK�*t#��\�U
]q^	p+�����;H�y�y�g���3��dYL��e�/��Pzm�?J��'x���Ԧ�s��]�2.�N���` ~��wz��)Ho��(C-�I���Ǝ��Nە�b4���rX
�(n.k
-
���`C�����j�����H��.�����nB=�R���MY
�O�tm�����������H�8�W�˜�B ݾ-Y ^T%m�/N�i�|D���IVb}�8B�+��%>���ͳ���o��÷e�O �@5���u��H��Y�0����� �E�3�-I�(&�p.(�B�GG'�%�m�"|e���<����$�F�
Z�b�#�(+�x;96=��c��+O
�P� ���}������R���ѸmPi�'��f�E���lo�2ψCM����O�v���L�h��u���h�����n�m]_D�8����~�PU�eDR�ly�Ƭ�ѭ9�c��e1��ұ���;ޝ�ز��TKȏ�n���q�$�f���-���A';�J9�\������1��ES��"�
��{��N
��(��@�zN�}��"�l���ū�QamX��v~���� ���SL���s��H�9Kce��Y�=�<�2v��	ı��!
��`:8F�*np���_X��0�GI֞@���sǛ`�4��qV��RKN&n�j��j�F�X=__�����Ѫ�����-��� ;��꜅�Xg�v�ľ���3\P�[b�]��_q���.�`�������
Um<s-cN�Pϰ1o),�E��{�\ʺ��o퓮$�����V��g����|+]�p���S
�J���7�N��vۼ���Ʒ?Ap�2�_�L�e�Dy�Η�#'͡Y":/!)Yӽ�z�����ytP�õuC�6���@֏ǝ,U���$�����9�
���S����(� �P���O�_T3��τ��;��%�"a�����*'��Y�$7��-i�K�Җ�����!tB�8�f���%z�璇�xQ:7�ky�w��nʃ�N���M�|�IߵY��C�:�b��Y�a��3Y�X�����@�SK+���� ��Ƌ��*�6�T��T�4����/G�k��Kz�K�,��������jh���� c!�p�昨�#1+��W,� X������20����ܶ�� K�k�oR��l�v<2��<��Y@�o��ls
^�F�.Fì�^9�G"Nйsӱｅ����H����i�0�K���0�T�?�:{'������<��( ��ڙ��~_�C�#�߸��TMӣ�Nj�b�;!3qF(�ڔ�_:��y�����eB�3t�s��:��~��d�@�(�H�bov�� R�d��y��Ajn_��Z�����Iߗ��~-kUP� ɴ� �܂GX3q��� ;Kȍ Pp�\Ѧa�� �mh0W��]]֪iYĮ�ʁ��gI9,�
rU=�
	��)M�-Z���s\��˧%Ѽh��ʃ��@߯��g��G�ASm�4v#y�L#�&�J��\�=�H�xN�VQ+y��H�׮�C/���Y{&OuG�Ptb|&4p�b00�4�6Ý�M�S,�)m�����'R_�2:�@�Kג�&�U���7��jKΓ�	�C2[:��#���Oe04^<��pȼM'��m��H�$=���v�ӝu���ju�a^����@��b�?���X�՝t����_H����7��K�a���o�/z@�8���G�8�'��\��S�@;[�B;��(��1��~J��{?��HӤy�И!�f#Q����(���^i�%Z����R���ުb]I���S��������[�4|���QU4��(��8d5ǈ�.#�4��Y�c�Q�ݸ�0|��jb0�=�<���z_�1)
fL�G�ʛ�k%+x.8N��l`�}��C;����fD@�-�R�|}�R�*
�Q���7�g��X]G(��i1�I���oe��P]�TwR��+e 8��;�SV< 1���&�5������W?��Y��	�ޚOy��٦tƋ!��U�V^���4��ƫ7a��+���<H���0�Wh0�8��Wy�O�Gq������� ��0�'U�[_3�ܮ��**Ek�S���-~���sQ�jg#����NH�?�Ƭ	W���/��薮�a��6�s<e�쇄iw�xdG��� �`�z�,9Oe��"镡�5e�2W��)�=z0���q���et�T���}ȥ�B2�
��ϳ^����� IX�4y��nO9p�]�9c���R�c���2(k��;S,񘔛zG/#:�T/�̅MD�PQ��=&��?''4zU-A��#����#Z����7z�5���k2��t���?�uk����dӫYR��-�������M�r �����ϟ��h��Ĩ��l�YΎwF/Q�1DR�
�|V�^������X�'`vg��77x��J���D�������
h$#'Gc�C�pA����2�^w"�Ѽ�&���9R���B[C��k�.K��Ci`��|˾��3��(l5O��kW'�Ԥp�a.J	�{��"_5����x��P`���5���^&��Mz��� dU�7��w��ǆܚ�zq�e�2 Y8���#��=� rҨƽ��z�L���>4�"@�JA.�w�ݳ�\��
���3�F���j�~j��%r��y��wn��"��t���#�nj�b��ed,�q�CR-�06�}	N�/�Y��$X#��h`�����*�Ǐx�e��g_�58���[{�E��>�"�Y�B��8V��/y�e�vJ�f*���
2�)�@�'�"fB�P��s�$n�N^���/�]r���(Ienz�2�ݘ��h:��d��]�~ҝ�|�cڧ���(��j�����Qu��u���xGJ���$�S�d�*F����so�$����w��� �Ĥ��6�~�+��c�#��$b�(��L��=�m�X��)��XϷ] D�=��v�8.4�.�%���/�Ru���sb��3tT%�j���C~��ˍ�"9���`+��d(�GIr���{
��mT���H_h��9_׾��`]Ʋ��dG{J;�L&����n�S�r �m_�Q�F;�"L�)RlI}�L�����i~��r�Q
��A�>(��O��vUy�n��āU,��F7�zh���X�HCQX'�z�2��,̓e�sws�-�mZ��*h���֕�&D�<4E�'oQ��O��X
S�����m6Z-� (@o#MэTI"�-DK��s 1�,T����6���J��D1�Q��KU�qӳ�׈vu��+�(_8#kȊn��z
��,b��";���`7� 9����Ӯ���2�i:���ݞb�}���ڑ����q[�*_�W��rU2߳Mn'o�>������?2\،�3�!Z�K�ZP�$��a�p�D# L�.z��=QX���)k�1s�(��k����~Ȓ:��u�]���b��j0;��Òo|�a��㚪 jD)x/����jMq :I�_/�����%X���h�`ۦ*hU�I	6չ	h�@`���Ю�"�R�o	���&��'-�U���_$��?D�d9P�a9�����1w`A���_(�`p�����om��5� �Q��U��\�w��{�칳�I�ޒx; ^��d�:��8'��6��^�����Eȳ|�CXpZe ;L�"bu*�)��˱,��zȬ���E'����h�J={�r�|`����v�^��~���ܚ�Tf�8p��`6H�qB#@4�>ڠڴ0ޖ����� ��a��Ρm� (q�`g�����L��N�l�T+��"S�ċ#�*����ʦ��O�qq���6�z6��ʄMV����g�����]�G�!�%;Ƽ�vz"��n�Q�0UI1����H r�����Jz鲮9�������\���`jCr'%�u����Z��E��������P(�i"��z��Ηf^��׊�̞[V� �$��u�Lu�Eh��=1%�] ��V�G����JH��J2˾M��r3#��Ft �}CVu��CLh��T}�!��Rx���y.L1M��	�lF&4�y�h�+,\�t��g![� �9�+�m_��.0ҵm�X�}��ڛ�M�3���w���W�%c��+R��U����')��],��i�K_����Ob�a����ڒ�G7���M,�������v�,-MbI\�-m�a^� �ǖ3%�[֨s3��{�I#����ҫ�Pг���W���c?��r��*��[��������F����e�T
a�+���!�є�jzbӎ�zƤ�rq��1G@g��G�d��ӿ��f
;�=��`Po�G�} $U��
���{����2��&�4���A�-���>p����}y��/�f�R����h��^��d����	,��;ݘ�
�!��w�ۜ��柯�֩��ہ,�%10t�:%�ĕ����V9���|��X�b�n��z��CP�#������ n��La 㡴�% �bU�F�W�jv��p�g��N9�ZR�P, ��>P.�RUd�G�p+;q�
�����@�BA�*�.<��ZB���W׳�9��BC
tU�"Ã�d��F�ƪ�c*?��㇨��U>���qY�.�WN0����c��-b�~���@������ 57gP�M�����o�ʗ���5������]=z�m��	j��\������H �!�̀5�b�=I�a���8� ������*Z�̗ ����+?�Tw��6�W����M��	.]9�=}P@�o�����b"m���*���;��E��!��e�1�H�Q��cD�ab����/)Y�S�z�
o�"���� FVI~�}~y�;�G-jSs�b�3��N�ր�M�������W�C���x0ރ}ˌe�S�TF��T���:ı�hfd���&����������-��;JF�y��\y�)}/-c��xo	\+[��Lz��g�3��җ0H.����^�MA�>X�Tk�h_��oK���<��lp���z��F"���
N%��ʜ�-ٔۥ�9&�Eiq�gX�q�fi��B�Ͻ-�b쑓`���lʅ:�ן�:�?�Z=�T�2�CMY��@sS�%��*��	��ʽ�a��ۆy�aT���46�qpjx`�����gN-[�G&xW5s'E3���ผ �w���c.�0��:�H(j��^A5[(�7��A���k���cHu�i�晋c�Բ��]$����@���xj&ыw<^�eϴS��2��V����
���J�2R�O/|.�:���h+��u=�he��uQ�H:��⪧�zX6̍�uc��ڶ�d#q@zጧ7�7�Y檵*�:F�+90p��~�6_\�ֺ�p7\Z����蟫),��uļ������:C�,̸�m�R����K���1��oq�I�c#��?�
¢��(���)��a�b�Ρ�<sE`����1�O�ݎ�+ސ�Fq	Vl7��d�Z��-{���I��S9�N6+<[M����U!���Dv��D�|�1��#U���]�q�Z��⚷ʖ	���� ����$d�t�qp|/���~MM*#�Q��	:�"�H� P���Ru�4�҃�#W��@u \>�ٟ<��.�&�F9�oa��*kt��=w��&��;���.`���a���hj�G��	}��Mg~8��6�����(�`is���B�步���o���{��<�4����E4�#{ӡ�����+����q�l���`�U	S(�7�4�����WK�	?�5�AiK�.`�����C`�fN�Ȼ�qq�t��C�fݰ��NS:�8ڮ2����<X��H�*�L�ꙩ�F K��C%GT��x�g��z
"�^�Ѧ�� �C�)�Y�Q��:�cP�P��S��.�����,�ۆE�J{p�h��.��O7#$�_mY]'0�N��
�%���v�;�`3��# �F!�4.ݸwo����|���������%� �um��8�V$j�@�&��#� ��1��o�sz���a̦�Y���e�޶�{Pw��RK·�q��b����[�����'6K��v.�����)���C}%q��������D~QFλ�.q�J��sLdh'.�F��T �	�1��v���r��N�,$��l�ս�5/s*�5�ɽ��@���1�lx)k��GL�̗�?�2��0�#�P�W�s�}��e�zP�p��k |��3���O����	*���X�]<���� X���m5ݹ���9x�o~�>��F+�dR�
 �5;t��Ev��6����g�*����vJ�=���%%ﳈ�N1B{'������X���:�}�SK}��K�S��噌�L�p`��aND� ��댸(��*��I���yŤ���,�H���!%��X���Z���n@�M7��є9ĢHÙ�+��8H����,)i�4ᘗ.C�t�� ���M�X�a���e>tl;��F<b�S	�B�됯" �ff���Nu�.�v&͊��E7��t�r��xM���<I���+�M>~n^]�I�Atn�����t7��q�g`���3���D���n�����޿�W�N+ű*�N����2
�~Ѿ�"QXӑ�i�&���f(�'�[rs�)a��������$)�2�b��3��^Z9��>
�����I0��F���f�W�9!w)㩞
(fF����Z�Ips2
Y>����14!��a�!Fo�ug�I�8�..պ�N�?��� �m�����!�\�.!�1�ŵ%�1!�Gi <m�8�;��6a�]�(Dg�^��:���,��?��5������O(1�N���}T�޺�.�?���o� ��r*$�Y�3:���@���7�H��9ZӉh'k�f3�<>*��bL��9�q�ز��yz+CvT�s�E:} kc�_�n��)	E��˝�p�C���ZM���@�<�&(M:�E���p�G },ߞQ"eղa�W;a��)
p1�m�}����L�Ds�}Q����0x]�+=G7��Y:=�`:8�e!�zI2���E�U����r�Ț9�@��S����I)\�X�y�����yo�B�F#n�%�x�SzI�{�R�5������k'ǣ����khA��H�9!�v��l�<~>��إ|&�����kl7U<�"R�h
Ml,�/B}� ��B�K�HX��t:�0�ɒ��+c�0�U���4�|��6r��즡���e���=B;m�m�4tT�ƫ�d�R݌��r7����G�*P'�
C�S$����/KC��Ï�EZ'Q�.�'34��,1����������g�B"�v�����|4(�B;�n�ڧ_3A��#'�p2F�c�Mx�7d!a�=Np-6YEifC�I��K�M���3���רs.:r� �%uH�'�A��ؾ��}p����������J�����W��'�4��u�����Bi�x������FP[���0u\���OX:i�'���϶�����6���?Dˠ���Visx9]kk���k��)
�7��\G�'9Ap�_&�m������i�L�h��1�HsQN|�6f�38o��)3?���{��������U��"���j�H�IF��1�m�{R�#n��y�G�I�"0��g�m��Κ�@�rkc��ԺL���g�1�v�&���������jw-�2��~rXŊ#��)[���i�|���9x�y*{�&ᾋ�b/ǝ�} QߚiY8�GfRt�3��啓E|��0��2�2����*n�'��꓆�j���}4?��a3u������V��Mf]A�Ql��m�rP�9^���k��?{�H�����Jj��zr�tq�����8(�����7�y5�C�ϐ�!�TG����~8��AFDs����
Kr=��瑾r����(�x��?�e�4zl$��6�=��5�`��L>f����Ƙu�*����@9���"��N#�Y[MFQ!�,|��0/�L0�
8���*|�jk�R���̒`IB�1@Ay�Lw��)������(��!f��e�k��'&1�K�� t2:#ȱ��|��#� NYS>'��3H�+P8��K3%� g^�(8���n�#��ǺY/ ��=�3䤚����0Z8�o�b�[�&�j�=�'O�3���	�?O�p�-�Q����C�����%�����,#'��wOd����ϥe�!���Y)$G�e��i
�A_[y�ߘ/@��?�(���J7�ߕ��Z;b+���bKM��1��(��>ZE=Q^t����ږG���'�뙊��{,Ҿ�ĝ���z��Er®[�.a��0W��<:�U���ڨXgĵ�x�&�m��'_Ow��!��2+5w���������&�KZHr����i���m:2XFyRs�Yٮ�:'_H�ۖ:f�gu��1����rJz$s����5���N�B/�b���Eá4�@���d���*.Ȕ"t%�j�
X�wo�Ǩ��G0ƣ:S� �{$ �N8O�Jl��d9�F�N����G��C�D��&�&97>�q��g��g�p7q���<)�)����s_�]��I�l��-V={��̡�������vA9-��]�n,������[���W'�D^����r��	�y=��S� T�#��w6����b8c�@$��!6�w�ݔֺ.8GM s���ϲ��9�d�kJ�aY��a�!��"uj̫uَ���X�d��H�?֎���Yl�
hV��ܧ>�oh�#�?���7��?��h;@��W
~!d�
-\�Hv�~I_�q���;���D���~&H��A�)ўǅ�P�*�""!�n���f|m���_n����fOrk�A�}���]�d�&�e��zm>��� �:���-k0��`�Y�$�n�������q��g�P�	3�\D7��&�k	X�v#>h��h����
�z�{WׯY"�9,.<Mu�=�}8�ڊ�-���	�|���t���޸�G1X@t������pg���@}�/"�((_�r0�4z4f�������Þ�ns~@�%tt��㩛�D�0H6a�}�2ty6t1��&��6�p($u;����X��_VxIt���p���n���I�C�-U�'�Ƶ^�ybᲑ��4C��  ��*C=��AZr���u$�{���}9��(�.�R����͸��Y���R��SѽoN��ק�e�d>�v���C��2�lvۀ ��xc�5��W�Y�����gE`9��*Hh?1²�f#�֋���P��s�P��ڱ6�����Y�c6��!�g_�/�S����)�0L�E���&����d6c$1%������/R7N�>E��[����:n�us�kz�J�ũ�\0lK�K��$�$=sHt����.9�w����z�#���V���F�Fϯ��r����)�� D�n�u0���Q_�� ���č'[��M���&zFbl"�#�`���)ȍ����7�\��յ��0��"�oC"�J� �&����\[ͮ70l������
���3$��<dhU~E6������P���W3Q��[�A�V�Y=ƒ�%U��1o���iQg0
c�	@�FZ6������K���Cy��&����0�Yf ���Nr��7_O]u�5B���<A�KX�'$� I�g���NYZ�(�`֩kk�a?U��tN�Kf�cJ��+�N�g��IDNv�baR���	��TCDl�%܃ǶH���*Z�&�]����`��S�B��ÕM�y��R��'����w��]���<��j�4�Y����L[F
9k��Ѝ�Eiп�Q��j�Y^V�'�s�/�%肔���$}S���������%`�� 7�Y�KƁ���7�w�
�T��N�W�;,�:�gao��v={����Ƣ~�f�@H"��A�ٴ|p<*q"]�ɭ��T���Ξ<2��N�h�����%�+��/|�59�ok�"7S]F�N1b��aB����m����r���]��/���/����;��A�Jx��6[�C�t	n1��8ڡ�h�׬����q�i��!��qNIH0*oWz�-]$F���w�솂��"�(�<S�&��oD�b?L�ԯ�+E�~J�)D�%[hi̙yf}��;xԠ��v�m�o3��o���u������J��4O�`���R�R?l�ZuU�f���X �d�)G�k0����4}���l���
�=��� :XS!�N�e���Jm�re�8��{&���!A}�P)�	����ї��xk�ܝ�ʁ�ha�B3�]�T��
 ND�oj�P�v�; &����Ѷ�,����7� �~*�PX�d	�0�r�k��p"ޯNjk)��r�xiG[�|�b�!Px���*8km�%�q��Wk��/�ku׷F�.��`�]ݭ��ř����*�K��4��q��Ĕ�(�I��;��٘,��5�]zY�������g�ܔNC�&�je��z������!̏���`�ņ���
B�2hL�u �嵅�7��kq��MQ�#aB������KW�6��IK�=�u#���>u~�ݖ�����V]��c�,�y�kB���zG� �.�P��L�	#����B�\!�փq¡ *�
\����t���ҽKO[�ҲE���y��ueW�9D{�o��}��� ��1$�O�oUcQ
6�^�yk�{�TڂD��O${c	��	?�9%p.�3�`¢��՚�Iǘd�mt�%��r��K�>���Hf��nө��I�G�x����;���(%�%W�8_��I�_�9^�^���K�4ē\���,"�;ҋˉc����c���9 }bV�}������	�q~�]�f�Q�X>ṋ���0���1�Z�pȨ��V��⎬�R��s�����=��#1qTP�wha��n���T��Wӌ�+�&I���1���L$(w�e 9x7�[!RB.v�����l`z��&�?�Y��1'xPp[�v�'4nDB�m�����!�au�nM8F��V7�u���D�5�&�fH4��z&Kk4כ�.�:w��lEm߷���f�6x:�wg�$�Tφ�b���,��i��g9ܜÎ�ၴ��)Twg����܂���
pC(�j,�q�<��T��S��{4��cnN;��&3�7E7l����f���	����z�F��j�<J����WV�(r�>�XX��Cw��;��}N�3�y�����)I/������~]A�ŵ��� 7_%{�P�uj�<PT��i���2��\\EFL�E��ƿ5;E-85Vq��,N��{;��K�Y�Zq��-٦���WO�ڣ>�׹ �b/,8��w��Y��֯Ғ�Ò��*�Kn�xJ5i֟`P=�a�S�/�aă߫�Y�Kk��0�sL)�9�u�^�f���㥚���(��ч��H���ݬ� ��� ܄�Y֝r��_�siߣ|�G5�χ��e��.O2w�Cb��wm� Yop-u5ҳ�s�i��7�17�N�p,��>�0�8"�����
EZ7�;c3�c��PD���v��L��\������n�,�+��L�V����m�D��m4a%T�
/ Z�d�@�y�*42@���f�୻�Ψ��䜩��9IW��|��Rg=��B_���iLn�Gl��yR�`9/���"��&�w{Ԟ������^�9���<���'���u��jO(����ؓ��#׋���`p�=��|�,M�.$E�;���xjD7$��- �;����;Hh$٘L�K����h�V,�B2��QK��\���C��Cy�ml�Q���Tt����"���tj�Y�w7e>_���0� Uuh����p�7�n��}���,�� �����+�v���v��m�#�1m�qz���@y����ox<�������������ئ���3�$���F��d��2�`!��;��Z ��ϻ�{Ăx�<�=����R���>�o�LifD ����f>m�o��m�
I�DѢ���.�N���ǤA0��'��:��xUYPK��QC�5,q����E��\��\-�~fi��ae[�����{�\J`�ˡ��A�ެ�˟)OKH�]3?��ˇg/��dεf��ۀ^"��~�U���Th�V~)�_�.��P��u�f����ԥ�6��~$���M�DE`�;�>���N.�Y�]J�%��vMA�r��%��/��ٕt�ş�b�A�{1�D;��\��}+G����. D{��Ie�Xɱ�3��u��(���t�Cn0��:z�6w_b�]����1���{`% �@7L�O���*g� r=���q�P���h��9
��T���{/�Vk�Z@�lƽ��6���eY�����EW_��{4�����F�'y�t�-f'���aA�lt�5�]�5�1�XHu�2g3'�!¥�*ќ�D�U�m,"����}%����"]A_ߚ?1��˖�󕕳���ȣ&+�>��B̚,���ޙ?�"����������L�(�y��u�s�E�C�XΩk����H����N�Hn2+����0-�0����/n伂��y�um���Eg�oun6ء�`�8�]sحF��֖�R(�� ��\�gmQ�#���U��M�x�渗���C_��x�c��"/�"$`Be��Oɽ�>B ��:юZ��K�]ۘ�,_��)���id��Qf#6&���VX�y���g��n(�oo�c��ڧ̀���$t-��SfҪ�X� 0"�6��d��u���rFƟ�I�''0njC�^�����	�汷��գD��{x���
��e�#h'��J�,��-.�Ad�3v#w�x¬�'�966�s8.�uk<̓��_�1����ю0�1eeq������\А�R�A�#��
��hk*k��2 r��䙾j�G;�H/B�F+o�΋'�EW�
ݠc�55L�?�f�짩!�C�7*Y�z�n��il��^���T0
1+/��*LS��פd+|�^|�x������]�=�hV�ڍOvB����P�u��;1̧m����ʅ�3<�Hu���8���g��=�x��R�R�/�+[�7.#5�0mV�ò�n���
d8)�r�S��"`ҵe#Եm#[�>�?�@7�w�eBc�ר	 ˼[�?ڐ伶IN�~�ճ��X�	�"z�C_'*��EAtx� )�s���@�T�LʚZ��"}dox�{a�\�q������F)+���5Ƣ��-p`��a��E���Z�M�����c|ρ�J�s1YA�:1�!� ���ޚ7WR.�H{4���S��㶈/7[������pfB�L����7���:Y�!NP�c��ڌ���I�RA"O ������?%(���܍l�͌�6p8j�!���0�}���v�	g���fz���5��^�pJ��ߚE�_�,�"c�nT+�ʇ�z������*�8����X���^)D�]5��p;�a|�%�5
��>�}A�d�����K9f�6�0W�����x��X���r�,J��'�f�f�;�
Tc� �v�-k�&rj���~ہ����?(
:��� � ��D�Y� 3���p�^�gf���r�͘��"/�5�g�5��Jk����ez��'����+q�N������� 7!=B�T;�n�����H/��VŠ=����0ı]I�?'�칔��,	�o-�������U2��gv����u���.(�yЅY�1�An���}���A� 撔�F,<!���ٹ���XX�
~�!�Wj�G���i4k����$��]�Uh�MrC���m�>��q ��3;�5�П޸��l�Tж�L� ���rl0)yk�W�=1�����4�����5ӌ�_���2�g�	8B����[�
)���u-xɱ�s�c�\7P���N��?0�vO��_�]x�p&h���4sV���u�	\#:,	j�_�]�>	~���:��[�L���=]pRD|@}X}����3�f�6��P���_h0����*�Х�XU���R�_�N/��P�55/_�����|4��\$l���KK��$NL�?C��`�T[j���6� L̐�ӋV�a?�0�8��̊kߠk�Z�2�' �<��!8��A�\-�Jc=v�뛜1CW��d�*��&5d��EJ���H�L�Ə�1���Ҵ��,%k+� VI
+��,jDV�:��F�L�����X�h�~gcQ9��K�?�މ��ݏu�L@��=>4S�B����\c��Y��@^U��s�]|h�P�,Nm�*�D;tY=��ZR �)��b�0d�1�����k����ߑ�b��C��v��[�ر��ᆓ��UQ̠�kh0"݄-�s���K�WոJ�� �0;~�ц���`�O�2/��Q���%^5R��9�x���=�rEb�����W�@D�1c"��/2���G��;�8�����xIN|x���߮�.��T(�O�G6(x�$Ͱ���Þ��iq��}�k�d�$��ݩ�.��˧��Ny�7:È�M�o7؃�mW�
QQ���Fa�e]�n$�=���IZ����r5|}�_LC�x���� y&�܁�4�ZgT�-��]��iZ-X����U�)�)�Eϗ#G~���h;]���oEJ��}��_��wj���=�l���G)�)��6��R�����G�2U�F遲�G��C �9�[��p9k6�c���=�3��AR�~��"�z�e%	|�N{�8W�º�w��uN�8���N����p�?K�!�[�KVG4N���E�S�j�@�eBi�!��Q�q�xL�#��JJq:4Anr���9���*�@`������2pJ��<�w�R��v���RDnM��^��i�,e\�����s�k������ɶ�R�u	Z3�L���s3����x�A�l�A�����cj��;���Sz�XaK7��=(�>��=N�4þ�}���
βh�+�p*���r%�4���nB�ћu�3o<Yਃ�Fh�V�/�h���B�=k! �����-a�J�����X���sF;�{l�q�� <�^Dq�ػ!�L��
C7Ժ�@	��oٟ�j��}�<���by����c7Kf��V�}�����j���+����	y	x��J4m��16fY��ހf�A&{��1|��F;j���\�V�5xYd��f�Դ\6It��Be���x۟
�����&7�hԧ�Д5X(� 0��8�qu<����
���b�;q�՛�S��NK�&jG����}�:]�ñ�I���R\���	���b�S+Fw N�S���7���7����F0����R6
Tm��\S_��ª�=i r���F����hH.��.e%���4-�-��uQ"��ΥZ��w�fBLvLjdk;(�3t	��σS0=?jE	6������ގ{�.,�6H�o"�� 7�	�����:����bSl݄9�W���){-%@c2;���x��FP��/O�I��<^��x �%�)�,����hOΓ��.��g_���"�vl�<U����!/�
R7 ��Ñr�n�ɧ9�H��R'��E�$��4���y�Q�gOlUOݲ�k�������<��Y�|d�I�����k&+!g���(N����'���(���:�t���Y8��:#:#kA��cZ�V`H]�^�=S/)l"MH��Z"_\_|��|��.�a������~�`�����\L�㹺��B!Iq��褮��,����^4�p��Ҫ�~�L�����i���P��8�p�;p��!&>1?�3L-H��'�
�U�8��\ �f��w�kS�0ޅ����=��$- �y��2f>��5������X�`}��Q���	�v�87�v���#~y�\������<#R��>������%��a~z�ƲU����r�/jc�M!B�S_���2�>��"��xԡ I
}Z������<�&0�ޠS�,4���
�?� :̘G�"ܰ6�f�S�p?�(���|��MB��}W�%��{3a��5#T�Q��I�٩Ln+,�����F��3��1����*��I}ɼ���0$������Qj�� ��H��F�k]Ǆ��LVc��d�k��jc�S���w��9k�;]�χC�=���a���Jb?�*'�X���������P�}L����_>Z��ك�Gc��W}���-k
��N }�&�}�I����L��=甂Ȟɵg��JN>�⊴�������x��&_��2�`��V�8Z�l�3����t�w��e�Y�#��#CP4�6���;w��+Lw�ev�2��"�q���9)B%G��Z���v�6$�P6SY�h�	3�ٛ���{����˳v��O���0���1�t�G;[Mr�8� ��C�=Q+�&°�Ʀ�Q����fmz�y� �78j�at"�N���Hd�/+t���&�73a�ml8Jt;��X�ۡ���$�W��.R��j�0Z��M�<�5��r.�~E^����&�-'������h3KK�F���������/%����Z`I����y$l�o13Rb"�L�(��#/�C�����E��Q4	�$Ω�N�������0z�	a���i���$>��w_�?2n�~�'qDa7�2�]��T)
�5<^�K��+R<]��#��
� ��'��OSg)�� 5J�=��>�/�)υ�������~�3*7{.���[�R���y������N��l�C���ER�� ��(<�z��P�O䛨��<����*a�`� �0c�ަ�[��Z��3��56�6Z����-+��h0��T�چu�g}E�˴ٱ�r�)�c�)�}�%����W)C��|��Q�Tڢ�]�7ߔ�
r�U �;>/h��[�J��=z��<js��a��SF_�́6�����oB >�Fi���:��i�B�}�\�����u�#�^x*a������%��N�_BzC�[�f��Ғ�4zO$��i��/Hi���g�'���fN
lRŊ�`ؿ��x;�����g�e��~�Eh�5�� I���{}�� �~ÿ�����U��M���e����Xt|f	�(�~M�����r�Cpk"���!R����/�1��S�I7����*�he�ZPCfn�ͽ2۰;���{�۸���"z�r��n(��"3�:e=�S ��O~�߼�|�9����V�;^�sA��L%�Vۑ`��@�{Y���R{ʜ�OA8 ��1��;�ܭ�/�E�?��?��y��{��;Z���!��t9�L�*ow�֤)k �o�̈��&pl�����P�*&�����a>(ݢ�_���{{��6�������<ܒWg��v���x��8#�_e�����E�J�䐣{
��,�'��̀�C�=a��IŔ� ��!�Iز��l�L��U����}��ll�6�GW�y|Ҋ�� �\?�=�ى	���#Y2{�c��n>�o�,���|{������\�Ȍq�1^�p��6!C���g���8\���AkJ���YQ�jK����5�OD�M㊁�Vք���zg} ���SGL�+ZE����KQ���˩6���Ƙȱ\����T�_�h(���Ը�Wc#��7�0'.q��A{xl ;�a
F1���e�O3���)d��]w lQ�/7��	Cm�߮�������(�ZM�cE'c��B���o�uA?�'H͸�P���Ls���6ܪ�d�kq}2(�J�-�P@l�%�fg
�@�L7V�y-��#7Ϩ꯸"x�.!l�!��m�
0P���v�o��p*6g����8��6��� �c��/���a:|����FypqkK	R�\��@�LOD�����'b�םZ߿�Y��:�����h��Z5>j�r\j\���l��W<I��m�������'�,��F��We��'�l��2��l� ����q�锲Ff�"�����]���0a
�tFK����5x�q+HǜJ�	%A��XR���WM>$��:=�b�.;.����V��q6�ț�P�s�֟�*ڠ���.�-�CFl�͂�;�7��9�����ڹ��d�6����i��T�<=C��3�w��T�H�jx}��}aY��.�p�l&Ǐ\G���<B�r �Y�q"Z�xC8s���ʿŇX��:��$�L��=��g�GW�n<�\��4ı�~K�Xܞ+�3�@��U�#fMcy'C ��-��1���5>���,�D�G�:ܿ@?a���WKV�~_��[�9�^JcFiFH���(�f����7ed,ZQ/����{h���#.���5�"�ԏ�B�"bB�TȮ�==N����e��[��� S1G�9����c�!-`�v���"�w�&g�Xi'!�Vx�(�Į\��'4����AQ�a��������wz�5 �7?ؕ�pr5w.Pt��G�=�����;SAy6˗�v3�(�8^�^(����n��R�&��ڰ��Xz��}�(�O�I�!�xH^8�1>E�WMZ!��\^�sZ��ժ<�'�����n(����7��}����� I����X��F�QG*��M��}�ٛF�&F�������s4c�i�U�8/en��q.z��&T�j�"Z����WO8$�ň!��[�O.��툲@.&�?>�҄ȅ�AOz�{K#���$��!6"iuX�'�'6�L1�ӺVl��iɋ���L�U��fوJ��{�7$NH�^��� l�%��ʣ�z�D��>;��C�w ���	^�Ʈf �9����_���G�
Vų���`����k�̦oQ�"/^1e�â5�J��ư�:�O:�A�&9�I
�ll�e��3ƍ&��S�_��Y6]?`4���)�7#�>^�#w�oO,�]����,��	{��'bg����Շ�h*�W�f�.��[7�M�3������2H,���K�XjEG�î��gݡ�yX�����Py9Ʒ�H����T0g���%��YQ������|>�6p���sNɒ�8`iֳB�	�v��Z�t��M��-��=h���C��أZ�����<��B�Ǟ�:�D�����@\�����D���f�ȝz��S�coN�r���P�( L�a\r�A�
ʷߑ�Mo�2�J��V����TM0�s=:]���Vc~Ya��$k� ӿ���a����fy`�b��nҏq=��:')s�[��#%����űx|�+�`ddMQiJ�
��P��eSn����&w��6��_f�l����L��xbζ	�e�\�K��jEC�{��fr�`���
�k6!R87ѿ���W�8I��%�0J��U���=���d�|�}.�Ԣ��-��]�7�:`k/4������Q���JmBs���Gٍ	�.$�Bdq�ޯ�n�Ew���_��m�S'[���ZV3�~�l���Y����`OFX|��S��v2�G�a�m̻+���n-��Pf�e����{����8��hP������X��\����Tv��N����0�.FW��(�u��7Sh�QGX	OB�/vzх�1'H�Ryj���g�&����w��Ҫ�t�~�j]ſN���MH.]�VV�ռ	0	f�D��`,��H�Y��L���R�ޭ�D.52L�m�)���Tf�Ǝ�;W[�|�TM<���M�je�E��c�!2��/�B��}�A;�,�( ÿF����ZI���,+��|�Nk���_|�aT;v}�s/W�EI�g�4�Yx�t�mۆ?{�
�|Iݥ�i��Y�@����Q�ck��̸.�TRs�Hi:����� �j[��K�%�`��ڡ<��LK�aY����L�ix�˷MĈ7�?(��f��z`�>�_���Ro��$L��V�^�������P�pu�Lx"Y��{�����{��j/E2K^��婳���V��כ���rߔ#����(h��&���ĭ�)�2�14qS��Q8�I8�l�g�H�����UF�C��Љ��� QĲ�c??����̟(�KV������ITx�;͙���3�����p{t<5��9�l�	߰�(������馶%�>�E� 0[a����AXMZ��
�A������r��q�u��"���^��H�N�]�����7�ir��-U�@,G�$c�E�p�&��!kĲ��PA�֭V;�zC�*vm��'�,����{?Z���r��X���I.�����/�.���ap��l��UޱR��.ׅ'Q��t5�h�47D�K�v�#�Ɍ7�#n�r��k;�uDK{V5.A鍨�i!��w%�����I��R�*mbLkl\�k�Y��G��DSH9pqw��4Cf���M�ª��y/�ε�'^Ծ�a���f&��Q�aP��p�.جb_�~<����U��Єh�Eg�P��t�+��ڐ�t(�������9E�G��T��͙qq���m�P�M��z�|!����8	��,�I�;:	�$0y?��.Ȁ�@S髇T���S��?ZzZ@m+��n	F�H�\d�+%t!l��� jU��rKF�G,G���E��;��4�m�|e6���b �k{N8��&�J?jz�%�N���6��W�k`ܹ�/j\ �t?���E-7���2�Og0Ɖ����}Z�S��Ql���r�C��2�B�͐V�{~b�!��<P�~8�%��J6vl18��{���ӯx�� ⟊�<���B� r���c]v���\��C|}�H]�Ӕ��or�X}+0���u�U��� RY�����K��?O��[�}����?�8jz �C����_-��N���~~�>��u�ՙF�uyK�\��{,�"�֕�Y�����?����܀챻�X�uKǰ�a������.�e��{�a�^���倣�L������f2�² �Ί(�<�I+t��^�����Q��W}�E1���G.*uw�)�hq�
��%�yQ������\x�ű3�
*`���ے8Z���?�	<,Y È%���{2�;�y	o0i=�m���[��;�HdP� #n�_�=E<'oq�� ����&J��j���	g��,�~yl^���W�Ij޶�A���h��Tk
�E�b��e�VT�u�1I�g��˲���ZM]Bj��g��P�W����{о�U�b�F�To�lC��FR+��\�5W�f	�e3��UU���^�8��/��U�a+��ӊgC�e>��EWf����*( 5b���v� �e&����sZ�㌛3��<�NXX�*�/��"�T��1�$��V��{_*7���zD/�-���MOwI:yO�̪`������3xr_�X�/���-�ͣ�HE��8��(��DU�S�鴐�L�r4]�"�U����V��Hv" =�e���m1"`���)'i_�0�l/*,4��a!�(�p�˂���b��k�ݶ'1������x�[*�6���bS=������౼� 3�zF��ׯ�w��`��#7�F���?�Ϙ����r���N��ߜ9_RDù���|Y�B��o���q�hƴn�8;��`=�I#�z����� ޵8�-ڵ����Bv�H���c���[p2�H����(�@��E�ֻ�f���(�>�k�k�ؾ��f���"�u膜�>�� q���7�h��:KY��h�&�ᰮۃF�61����w9��|���*���÷�R`�D��gO�JD���>D������+�!��.�"/ZZ �rD�B�X��o�񼨟��B�� -\��	٨����*�Yh��g���F5?i�@��\�> |�;1f�^T��X��TL��а �M��\D}�u�\�9���w��JC���ӾH��VwM	M��,!�}�8$�Xu���N��6�]��US��#���Z�<��Fa-�F��K��Y��+.�眕b�tT���iV�/%���-��}����n�J-�����J�M���AhW?��V�P��/w�>y��sz����T�ghN�+]������DGo����s��c�j��J8 �a�~��m�B����=h|��=V�o1P��e]웈�i�N�RACU�>8�t;ZO�Y,������.�T� �xuo�І����Z��[w���"(:�����,P_��tn6�^'uQ�x�:A��;:,���{y�,t�j@�8���mu��c�nY���+e���ԡic녤�^K��b�=�7����mF.��D$�W�PŸ�S1R��;Y���d$���|O�i�K����Uv�^=Y�Rw�>Sp[�"�L��XX#˷	���/�S�_][G���ܣ��'�Eof��uk|Fֻ�O~'�/�`vKY��rP|�j�ŇQ9]� x�	�����2j[���F�+�̄�}��ֹ����ݑ��m���ՅS�!fL��1���E����:^a9��[ш��RŶ��'2&��u��	���&��{��x�#����z��X�kH�>��͎T������Ehۺ��E�{�����dd!|�ĝk(��l+f�`�Uw���U�)�L�$Q� �E=q] v�o�����r�⮯4ƌ�D̠m�*���2{e���:'VkB��YJ�\PD�>r&4jݸ����}�)����!Dd�s��\����N���o�w�͛+O�U��Ӭ�#������xm-��'�d��hGxLm���c��yO@��K��j���z������t^��W�0�
K��cп���Y�#r��z���*���أh�L�h�}�����CiRMYi��0Hs����YZ785B*|ֻ����M���qv˫�Ne��)4QG�Mׇj��:̭Fd�]{:+�ýw��TJ8���dĳV� :J^X�1D�� ��sao��
�J^�~�$�Q�	j�:���C��t���`�gk.�B L���0Z��y:]5�B��/����P>+�R�E��X�%��X����8g�o\��J��o�̮�+�DJ�o�zO����� M��t�%��k�O�J��I��_�F���kN6wI����BW��;_�䧆�!z3����$@�Y��݉�[L0���\�s��P�ROe�L���Z�{���ĸ�.�g��\KH�G��&G"Y�ʭ��I�'��h����-�QJ�z�J����B��gnr��x	z�	qfF>���׹>��Ĩ�n����)L��byG���
(l�O��e��)'k�tY��VAn���P&��}�L�M�����	7Ȯ"w^��m�*�Q�#y�ߚ�S=���Q�?Y륥��Ҁ�K���c֋���RL��&<gRhQ��2�c7�e*��i��T�3@�!����{�i}��!*@g*�wj:wݭ���4�(x6Χ�M��m�Y]Y�=e<iӜ�n�I'��}[K�s����i��t�T�Uĉ��F��1Y��HM&�yoHx�<l}aW�{[�Cf���˦J�����0&�6jti\�Я��YЌ�,��G��	�	f�#����A�Y�Fq)���z(�F��8��骛�u+:b-���$��2��9bx?�H�C6�T,�@�t��ե̍M�����ur!#K������P"��tM�i?���SV�r!3�I6��KO�g�K�ɰ����6�k�DRr��E.��У�u�+X�Ϲ��1���t��Bg�>��"6���|-F��u>�z���[�~P�'0�����0�]�͌%����L6�#v�3k�a��Hp��/����\3��g��ۇ�sҮ�0��<�p���MZJ�q��ILOig�1AH.1m�HgIã1��oJ{Ƣ�G�-�P�H��Y�y��*�wm�S�*Fv��
��u��$@�]��=����斟b O?4��J�C���#��K�h��I��>�%b,���t��A�����zٛ`?K@�H�e#���~K��mh�8����Q|O�Xq2�*e?�B53or���aC�
�hTg*׀���fή`RDB/xX�#��X�2� ��%{$_	2kCc@�r�M��fĂ�Q����<2=�,�ފWs���0Ez;s�o]XG̊��﹨a͚n����}�>83�c�}�Eܬ�b��#a�����#���Xs8rˑ�ʞ��W`0y�̤u"���sO����o���iА�݁�F��$�d?�5�F�D}�D���׸������]�8���J3W��L\���ߩ#���P�X˶C8I���rl�	�� ����{jAa���ѵ�2�,�axK��ڋ��t��WLV�*=
>�6�c��z*u|"X��sF�!u�� �.yWG=�;�!
���(��@�N��H��tn'�E9�8jy�x�K�þ�t'����b"7/z�7�>�ڤ��cܐ��`*R7��Ry��(J� ��}h�榚�����ȕ(��<��t��A|9Sq�|TU�[�O��ϩ�uv�`c9�idC��X�i֪��A�A�vm�� ��	�&��D�ܮ��#�YOzr���q=Y"�h��Z�M�HLi�?����q��YA)ֳhk�W���E��1$;���Ze���,$B�t}�|��-��ܖy�zˬ){����j��� y�,(����͂��=�&�ژ췀��]��������fZ�	 4*�>4���iBƘh�Pj��
��:T/멹��m�ڍ̗���m_@J��e�$L�95���������ހ��y���+ñPj�3W�������0���O�H	�
D��$a�T�5h,�;YH�i���+�����\��p^��8�q��b����������ʸ�������������6��y�v�AP���K=^ꢸ��6�{W6�7�ƫ��v��`{�V�w��d-��vkN&[²	����8�/cYL���
�@�Y�^r��B�� N2�("�����=�56�U<�GC��ז�ӃV1&M�� ֙��ac��K�.@��}����l���z�u�J!A"
�����E}�?J�v�yL �A(�?�o8�@ϾoRt���+�����Cg�Dm���rnN4�6�,0
�5I�Ѡz��#D�]f�=�G%~i�g�ɳ�	�y?�3�#��Mn��L,���������R ��.��P��A��)T:�\)�b��E�Z�d���#�>X�X\���~#�.6l}�L���c����V��y��D�%����C�i0O ;��5�c^��{b�k������D#��*C�v06���j`�8���,)�.r�u�-��~�6��8(�-�<� a�;r�ʿ(�\��r͐����N�Qy紟�hU���5s]��,��ȯ��FwN8G��T�g��l�����:�7�NWs�b��h�����<+����
2Ls�����e�ȧ�F��B�\�h������qI��=�gۊ
s�@��C����/5+~�`@X�L��@}CSfq���l0�a����9���ʹ�O�0�+Ga�>�N���K��\?>_D���c3C���!Pvߝ=��3����B�-d��6a֛&��X���|�J�y��d���Db�4�bP9~#��ݮ��E�R]�?���)0=�W�L���đ��͏���j�$���Ce��q#���?���~��������t�����d8��W��Da]+��A�I�;k�F�9�eW7�<&��#LXZa�	AΎۓco��5I��d��!��#�����&���5��
,c�s=S�R�Z��'��d��^t=c	��+�]��o��y�-��u�� �T�]������fFt�"U�9�0Z���5g��¯���:�"��X�8&_4���-~k�F��){i����5*m �kk�6����1�f8��P: ��d����}�G�����wO-_��HI����j���L�A��sτ迉pSo�J[I�dU1�v�DZ��9��� ��m6�c������:�^}�����Bi�^Ѿ�=�����������v�������z{���7GQ��t�� rC&���ԹX�8A)��I���fg)g�n��j��e��V$ @J������<�A�b��|T:Z*��ݭ;�Wz�[��R�0MCۂ}�}Q�#s���2�*2�-�Y���S}l�D��G�0#YŐL�*�W@�ԏT�ќo0�O�~���q5�[�̢z޽C�P�X-��[B
4`�Y���zb�L!R����ot���{���Tn٫I,K�uzI��#���	m�R�)|�i��i��YU�,��+]��C_%J�"���ۑb�Q�f4�M ���=:�x^s�u5�o����4���>))����*Ss��٧4O�q&@�ې�˗��^��L�#�
u���̥�u;J����q{f���mv�C 7G�e��`�lp��c�CƄ��+ɠ��\��^!fQuDjFz9�����h����/�V�.ilcR)��C�0�����wnD�ޞlB��h7.�4�̅�u��޶����b�	9�8#t&�Öc�_ �lsFcD�����r�]Aea�V:�"�#��@ݮ J�$�n�9�>F�Й@���Y5�DNu%��U ��A8�RP�����W�-�:V8`���n�<�k�x���}��㧔�Y�k�+6A��#��܁Ο�m�D�ڞaC�ҙ�>�F��z�YK[N��~�a����BE̦��ު?�%q}Uj�N����O��������L��F�D�4G�^!�8p��jvS5+�Y����f��N�'Į8&�s�q�:���K��$���Ѹܙ�M��Ȁn��-���t�S�eS+/�]n�\���O�kü�]�N��'DO��r�*�X��"&�J�	���ZFT ���X�H���ԧZ�<����#��D�a�%4�+����Z	B�R���1�&}7�œz�C����80�L�������w��iaT~u�(S�m*N�Ԑ6|3��^���¿�k՜��nb�1������"=*�\�����Xu锖��k����gaC����^���$vF�>V��nl�09q�� ����V*�˨�*���i�p�qyTB8�C�ґL�M c{!��p��$7^�3R��
Y�V����;�k�2�zV �|�����]U����&r������A�/K����R���V�\����-�9�PV��n聻Lkz��F� 2���[��e��z�}��H�v�1&=Gc�?�-����~��51�B�r�E��O��m����%ٵ2���	̠�wDO�����^9j�݌Q�9���tP�ofM~n���T���R���3	G��b�p��� 5��~�u�AK�6E��$7��\�N���tQ�ɐ`S�P�t���Pè5�g����D��������a��a|���}�1���G�ĝC�m0���]H�)=��-�Wlå�vkI�ϙzK�+�� �y��ጲ�М��R�4\24䆴:�}�b��̶�HŶ��������r	���FXT���C3��J	%{.�s�U���'�/����)v����<2��^R�ҫv�k���k�i�GYS�'��R/�F�VDVf� ��I�W;	R+�x�,�WyI��fx�>��I�o\T���'�N�+�g��>�x�v�v���`U(�U�H�	 >":��G�6&��v�F�.����I*b�X�/���um�a࿟�8�"������f�v�z�
1�O����i*A1�3-�t��G�IZ*e��eD(�!n�#-\��Ϯ�]�����8��-o0���A4�J6?O��s}]�:c�_~����Us�]��koǢ\0���v"-��vn�r�j�U���[C�c���Hϡn��"eֻ��*ʿ�7�C:WKq�dŦiξO���A�C�RO%#�h%�t�\7� �c^�c�O�KҌ���O7�@A�樎��ѵ@Y�p����k��F�n��	��w�����"̩�HJY��Qi�F��L�jg�Odn�VT�V��u���X]!Q��?Q8�xp-�繈�]��ml�<�.�jRM��m�?<��w��E�׿2_C:2��M�\Wfx��/�ҵ��:����܆ AG�ǣ��r@��zj��W����q;���86�Lfɮ�q�/�y�5abGv�#k���$��
V���P�m���Ac�l����Md�O(����{U{T�S���m�O�� ������#���4��1�%p5ݛF�HW��ȍ���m���hf�Y��gPo.}�[���:xU��V�e�@X�����=�+���86�U�ݳ��i�}�{CH9���ګc��jA��Y2x�;���Wm�YG뙽����\�1�&���MX\�.������t�9�`j`@�X�҅�kJ��"�b��2H��Ǥ\`Q%+��E�������	����t�B�p��κw���Ί|?�����A���S����'6��?5��AcGT�s�m��/'8�&MO�2���K"~��O��L��Sν,���QHΠpȞRY��x���a.&n[�?�W;"�kSz�?�>���
����hT������w/b�1����f��!Iy--�Aa ��;�m�+����Ưێ�a@�PG2��,e�^I��AAC[Q�QA���񶊶�e���&@��ֺ�g#����L^ ���M>���䤳%������.�(�����B2S��E�u�r����O�"�bI�������;�@<���r�LLB$|���@3���W�t� D�?�
���O�M1�H����PcDh?��A�\1P��ǻ-D�)�OK����]�p~a��2���<n��#C�Xg��_��z4xq�*?�Wo�@���ԹH�] ��O	�u)o�o'o����I-��B|+�Z��Ps�5*��3��R�E�=�t\�vDFM��t�u�	�ʀh!�:����_@=u��l��w��/A�l"����:�+萆�f�ɽ7OXD��5d8��W��y���}����HT�{�m�N�A�6�转�4���F{.M�+&�=���tp��U҄#�F�Ա�WJ�|�j�[�O��z2�5-��[x���Xsu���?�<�\VzԚP��-R�<��컩1׽��ۚ��t��x�GG�/����4VH�Q���O	��̙!y� ��pj�ʹ�)NRo,'_��r[���((��[�Y��J�!�a����Y;�wX&d�a�H;rC#��q���f�G�m7�pDۢZ �P�Pv/��rM���T�M22C�`�o����zº��PGv��"
�{?Q�	=��Yu��~�5"$��Q��Ⱥ�}N?@�Q�[�Q����grrH��
>��8�h��*n}kg̼�\�h)#"�H?�R,����+�@��Ʉ{���^�ҙ����/ӡQ�Ն6�����r)�v&ǵS������J~E�]k�٣9ԓ��ߌ*�s�s�@D�(�����m��vZ5�6ɭ]!})�[���T%�����&����?;[���!�'m0\,�^�}��)�1S�[mr�ΰ�.<�*�:�փ�\6m�*�Tf�J͆���@���Ȏ���Q(�6�«~�eB�ʑg[Μ3ʝp�t=�.�y���=׊�^����g=��qe7'��dx��]#4 �I�]$B�b�s�@��dn`����[����W���t\=ߗ\[5"*?/%��1K�}A�5���P۷�ڂ�adΐ��p��D;U�w�&�X?�&�Gov6����#��(���/쭳��B�?�ҍTE�*O��)�ͦ4A�-/Ӏ2m���<�l���k�z�*=�ﰝ���t9*�+����cw��n+Z}��L�zɠb[����;p��4��J��D^�G�D�܎Z�X��<�`�$��,���]��%,d�i����yq	������c�ǘ@g�h�sʦ���Ky*�2P�R����'x�7���aL��6&���_�2��+ Є���]���
��E$b�i�P�$�d^�zu�>�R�#&��ώ�~����Sd�3�Z�7gvS� *]E�Ne6�1���ג�o��<K��X�'�x*�B����OŇʖ೩��סETh%�zu�� �˜3T�R����ER����x4����񬥼��]�_���x٭rck�MZr>B[]��g�f�W:����,k &��>�)saSAPd3DK�g{Od�KG~?�^;�-X����<r$�K��+�ˢ��r#�?��8u�s=��慍Ҍ�]�A}Xp�*O"��	t�{�*-c�#�1U ]&29���Оg���л�:e��ٟ�핢�eQ�a���ͦ&���Jn��t�p��o'�w�����&{�ǽ��=t>��Z#�_6�+�Oɨ+�r��d�T�[���{��æ	ͧ�f��3Si��p=���Ym�٩t�(�l��3̦�2>�(�]�"�e��=��è�A���B���z�j�����O�Z5��S�yLw��ޔ�������b~鷭����]�	�u���t���I�l�&T���]�$���
���`��XP�}L��w0�Xd^�$z�!�PWZ��B;�t[E�	�6v��������IΨ�@�x�&q�;��X��(/����_���;#��ϳރ�!~�,�{'>kƐ�����0�P�U;x�&���1�2Z�v�E�6���6�L�;91O�����ץ���o!5[Y���RQ�^?�/)��bN}�@?1Rv~3�8�z����o;d�W�UY�l"8�� ���
k�K���2�b5ă��@o�y�����~}�?�*/�<}�q����y�#Mo�̽!���~�2��M^�K߅iӆ��(V	�5ξ+t7#�ab�q�o��g���(�4 �Z��Q�K��TD�Ju7�ܱ��3.I,UZ��7f�1�G���Gvk^T)1u�$9�A2 ����_�����3���ګ�������*�v`fDE�|���wP#�ܻ��(���a�d^5a嶏���QR�N�5���%����?�(�h�}����_M�Eg]�y1�؂��7��)���m��UI�s����[��N�	�X��&B*��Y�T��r����˛�{���i1�}x���+�q�912F�;���ZÍo��x��K���L:t���mDS�o�rq$F~z�B`��g�����ӑvwl���	���(sE�ʵ��C�k",�����6ZP�*"�)��-e��C�@����	�[ò+!Cy��zB��U��+��Y�E��]+.�'� ���m���T�Ҙl��wZ!�K��V����(L�
K��n=Ǆ�*O�~����Uk)�u76k�y4%� 2^�),�r�e�n���D����`lK`���A���;"��p?z�d�y1y�M�Q�ۈ��x|Qz�n"�J��q��"��V�G�.� l���"��u�Ӯ�|3"�=�!���;a�E	0s�j`��T�~V���jic֘��Ո�$�_��%w�T8�2��0@,��I�����˼�+صbk���v7ľ?�4>�Coj(;����t�0*�6+m���������NV@�>Z��/+��K���ѓ���@��J��i|��V,��zJ\���n��넩,�6������;+G�(��"��1���r�'e� z�d��V���3Q��M5Bp�4��M>�Ēk�r>&T���B��-nm�ܸ0ϗ`����S�gN��O(�l����1whu&�S\���zs�,f�pGI��d�����A�6�pY긵Ԙ\VWՊ3(S!� �;K� ��X᠀��# Qm��u�G�Bi`x�NΖ���4^n4���2�@H��8t��~GcPX].3W�?��y�̖峅����.��k��WL�|�c��1X�@�	��A8�em��39?41^K�؄���Vz�|�.l�D��,֨�o��G��r�*
���lqTl���0����.V��HBRLV��.��10�C��N2r���1���~��@�[���p�z��Q�2���A�KwX
���zN�s�{��Åu� ܣ &��w���$D�xz�JX�̧؏���FD7-`�uH%c䍑��a)5�i�x �b�e�z:>�5=G����!h{aI��#���2s=�2k�d��\�ުx#�e�����;[�¤qD���S�q�^K�e���*|�Km֬B�9��£��{�CΥ3��W��\N�[:Ds��,��� ~,<����3�D�pz������+�ͤ�u:���K;Lh��h�R���@�]���.�����v����bA!p���.�GR7`sQ���$�CG�hw�|�G�Ҕ�\�?�0�Dd ��Z��^k]��>Jȥ��.qgvb=�Mi��!�_s)/���;,efj"%�rmpx"�.�W0M�� w=�'�2qU?�!�R8IU�,���G�s?D�a�ß��u�IW�;�܁���p���S�tJB2,��+ A�Όm0�(De��f�³�ǖ��h���s��rH��kh?B�D89��Bun�Zy��p��
7C��܄PO��$ޙ�6p;r�����L?��}���s���q�� -J�!�&:2�� 6*�A�������k۾h��2����Jk�9�� �|d�F�â�eN��.�3D6]��x����^�B���b=�(��z8�˥2#�#���Ȩ۾:m|Y����Xwi �C�x��,� ���<���2��a�?�� ��>���O!ռ�~�saXN���,��gc�Sp�P>�%J5z\yȎ k�0!=7���8~�5	��m�Ps�v�߁O�%�F�?��ɻ�^�_~ꤥ7`y��,��zx����8n�X3�t7��K�L'>{]�X�W`�%�vа���【�4Mw�;v�jUWn�He����*����*�cur�i(�4�j T��0$l[��ZV	��V��!�^VNv��@O/�5�.�d{�O�0�t��h���~�a�c5s��v����I��v�#*��٧p2Zz�]�gb|6	�7}�����n�/�8���@�!��P��Ś���,?��~j��o/��(�������U��x|?z������)�]!��1��.�X��BD�	]UznҦ-N��] HK�$�	5����锑oO�se�U������e9�^�������������E�BE�ϊ�JQ4�\0L�Oa�p^���`$�e��ߥj_L9 ���
,�Qn�L����F��r~$�>�Yl����\����)&CHE�OG�Џ�`������Ô3�ütɂ
<= �)1}�֔Rh�!ӛ�Mᖥ6N� El`w�g��1ϧ�.���� ����SbM6�7|��t:<�[�G�'6y8��2w�y~e<FY��o��;@����wX���q�a�-�s9��	?�mj��{l��b� �]��������l𖥨�V��X5����5�zK׏�Hi���"����2�����!D^t�K���G<������P���֞�8�2��&],����i��{DH��F����y��b>	�i�^ˍ�3~E�ܡ�A���[G 7Fz0m��@�o��|7�S��L�+��q
����ԈD�]����zC~&L� 8�55 m�
�K������ܚ&i�B}������`�W�M���
3���g�!5��.nj���K�i�ԉę��������D����lW߉�mm ��o�MD��|Y �w��U��D�tŐ���FXA4�\��qX�Q�eO��y��0`��3M�<
w`�߬��%��n�:�wE���Jn�h�16�=gC�m���e�Aɖ���T��$Y�2v(��RS5l8��o�Y��Mk���S���
�ɧ]��r��"���F�������¢�5�	�H�pW��l�^����ؼ9	�r&�]y].�����=��f���aօ����Y�8��a5��v@��S�2GA��F�5/�}c���pݖ��'���Μ�r%���`s�RS�?5�~�@30RKs�����!`�'�sR��a�U��6�r����!�o*�����h���T�N���ZZ�DJ��7��Zsu��=~3��}{����b�$�U�˦���^�"~@o�+'��v�7�na�t�qfl��R�	�[���HJ������D{���\����\�V���D���fr�8N����9�O���힍��?�m�F���2�97�1��hI��P��-��Lq����?)'��a��z����"Y�ˉ-?��Z��xfh����!�8֬�}7�0���`ؖ��P��������I��1u
/��;�0^��d�������Yr@�W��������1+#�n�st�"���E[�!l�ZC�1P�U �;I��A� N��q��?£�A�
\w|�*��vb��|s�r�Ӂ�믮�k�x�e'l8��vM�����AJ�oZf1�۰�D��Z��0��}�_4@x
#�v��(#Q���x�Ch~�s'�u�O�^�^�g��
W�l�lM�-@6w��Q��B ���V{R1>$�WъJ�OD�X���ů�w�Ҭx�<4j����X0R����q�A���q-4=/t��jnjZ�a�˷��!,j��+z9���?���/\)o�v�B�}�s*��f�?H��oЏMN��m/�5>�W4x9�Q��A��a�xbqq���)7� �dp1r�?��{s��0y���,#�9�f���XӾek>�����+^ar�������ڕ��ÝA|��,��ů�h�C�|u�V.r���܉'��� �k�Z�vL�'��w`��߷v�P�٨h��7���D[f�.��a,���wC���%��&G�Y&Enw���^G�˱�kP��"�'I�̍7^�a��?�γu	��>������T�#^�`��Eܯq�6����R&5�y���wq����r1\I	�FB,}R�.�T�=?�C��)��팗E�Ug� �O��俛�LZH0�}L��3�o����9dg���]4�1�M�3!^b���g��?��/���ot^�T��ɛ9,GՏ>-7�����X��_V�?���3*��8`�R���
z�UQ�=���ҳ���G.�!��͞M�d^hax�
<^�j��?f��*g� \/d�bצ�w�v� x�2$:�����r9�ؔ�3<��񡍠���p��d�[�&��}!�D1Jc��ˁ�GQB�(7����(*K���)溥��=B.��?��R�ǽ���S�>ky�%�s��x]H�Z����~��b��ƛ.�b�x�����2)ɖ�w��\��a:�'9���>��d0���)�;]��$���ȏ�u"Ój��%�� ���8ȓ-�u��Do�N̸vHYr�ڡ.�xϝQ� ��E�M�~g*�e^��xt�Ō���J��I/
����k	-��*f����"Q���tA���� �n������5QUb"�"�`\}7^ͧ�"��w�4�� Kݢ	��W|�;	�lG`����)0hX	��_\��%G�{��C/�tCܻ������t&�"R��������uޮ=��D����{�A#�9��s���'
[z̙�g�L��h�
7�
ŏ���[M$I^��5ߙ��R'�XC���C�"׸<�	�F��8jaK�q6�ZB
Q!=����>᢮�	�X�ӭPNyn���l��O�8SYg!+(�:]AUd���8U~��a������C���pP%,ù����<�=�n�*3"!.+��mx� ����ҳcw6Fu9�"����K�)��q�/�np����M�8�� �M�%�S=Y���`�~4GA"�s����J�3`�,�u�\caS�$�pP�+&�J��w���mwx��T�� IT��?�(̄F�OJ���9��K��� ��z�RL|� ��/Z>&�����յ��6��@N{SaHo�b�ŝh.cD���&�#��M����"S�R�R���9q�r#��J1$ʧH�w]�(��q���.ޜ	7Ɛ��4P�[�Ƀ��z�k�y�B}NZ�C�A_}���\ҏp�C�p�2�Ĕ��5�Յ�ָăiTp��vo������,Cl�J���RW���P���M2�Z�����*����B&>}��"��%Pdw�Np>ƱV8�/͹Һ�Zg#T+�$�J�g�6�)���"ݵ�rT\�^��ͦ�%Z�u���Xs�w��`�Y�A oLCY'&:��@�C��qgC֠㭓��o8�[=$rN�:�D���a�N��;0
��բ��*�0�;sɢ�m,�2�B*����5ѝ/��Ԣ�H�E����v0@��3(�sy�q�o��X�M=��L���6z����;�W:��>!���*J"_U�gyS�O	�?FXQb�Ǳ b�w�P����C�GvO��TFi �	�~B��01�o	�<+v���4{"M���2B��yѕfX�t=�5���noMk�t����:£���utLL���T����R8ܿ�)��L3�8�:o��>����j:�&��+s��J�/��J�	�\̍�P�P\a���<U�Kx�7Idؓ@Z��}�L�Y�s�B4�Y��tq�Jfp�\0"B���Q� ��L5�#<yZ<Fe�~	���v�.�ɚDOQ�z�77ݸ�lz{��W�n�I�W�6K�.��~����2�mEϝ�Ch�-}�q.*\\!��	$適�� �}�{4b��{́�}�w�g#W�|��st�M�jҵGR�'�I����p�?�9�B�g��{�LpӘL�������i�
.��:2�Y%~���],b���N8���ؐe	��mk�n�h�]��Hk{ɷiu�S��m,�Xj�U[f>�.vl��!3P��.��1��n=�S���X��?P+��s���v��L��b2ݨfw�������<�N��gw�K�%k���zX7a�0#�־޵��֒�)7������?A�݊�[/�UP�����E� ��o���vɒ�d��~�����C�Ig�<��E8�
�o��!p���,E�h���H�_�z$�+~���>V��f?��Rr�1������ѧ�-��y�C-�l����v;�3���U+k:7nFM�,%��>^󞳩W���0�M�0��˹^&��c�;��Ry0��Ɨ���HҢ�� ����z�`��',��?�����g��� �6��O��y/�.(�����#�{�4^�!�� ���32&;!�]~jҗ�'���xu�gNZz&'e>_.n�u`QC�� &i�#���|Ob��+�R���/b
�H��	C��i��G���b�-�����.��ᰲ��Z��r ߀d�`�KNV�T͂Hґ9-Q���e�>C���*xoF�=�4��K��Ӛr�~Ceή�&�-����~���쟾���̲p�F�8�����$9xO�~����'���
4�քx��|���{u���C������[Et�a�[��E����4���96�ly�jI�h2��.d[��B�o��x�k� �<C_�7 ����Uu�X����3^�I�L,yQ��{b� ١��2��m��K0D�m̧�'[��b�U����R����Y*�� ���r�Ij�>�]B�r��&�oZi������B�;v�sr/�����4e�X�ч?s�2�ob��
Tts����>�D��#H:��e�6I��=
;q�N��|m/�q�)�)�4t}Kj�����<~U=_�V6!�X�P����?�085�i���$AS��^�+[�~����pI�MdW�ƔƼD�r'���ϛ�I�7�zO�>(���^�eO��������Ms	|W��=�_�%|a�Y�B�=�W(�av<IE���O�R,8�<Z��S�XS?O&VNg��a��fk|�AYG<Á4f�8l�<
J��Ns���RŎ�����L�8�����鴍G�i��߄�1�?�gZ'�mB6y�1��դ�ų�����Sg*V3@��ړY`��{�)Ḱ�?�2�%P�E�9�sϮU���0+�&
QM6���Z��c�Ԃ��k�hO�����wr�<�}�4Qe.��z<Z�ߧDQE��1��!4	��򹭽�T���Q�m�M*�n�%[����j�2Ls2�yNB�����7���:�����*���k���N��NgԖ�\��C�0KbWS�;Ӵ!�����/�D�),͎�xM͔W��bL��+�!��B�[ܰ���{�m�#��哨�&\߇pz�=6̛n�]^����v��r�L$�(��Q��r�cGu��{�[�!�|����O�J��FJ6�� "����Q3���%k0�|�:M���,{@;g%D������m5ց�kqZQ6˦��c䑟���(��a� ���q�~N |�I�l�ۃ�����T7�Ԕ��� ݚZ��h�յ�C�ז�L�M� #UoW�z�\��Ǵ8�����s� ߭�?9�}*�����tm�G���W���N���)8)h�2/B��+f���䀮#LH���!�snJ�RrY�|T9�W���G�v;�>I�5�wHV��� JN�rw��7n��^+�Cߑ����S��lE�O?����O`��������w1v�̰�=!�4S�oh^��z�Y�����9�0��:��H��������G���.
ar/���e}�k�/>f��p$m����G7�]�S���oy�3�r\��Z�� �W\�i���z�zN��<�8dF��1�<paE�"�ZKɗ av)I� OS�����P`�
ie����5�O(��ւ �L�[���Po6�YSk�̜C-w�=��=\��`��0�Dw;9p[�C�r3vp����~R�f�LvX�,��Ja���"�)��b~QG2�A͍b�L�Ef}$���D5�?
�-�P�/�T��9�l��GM��K�Ts�H����F��_�z�=P�{J��a%zZ���4xa�t�Yo�f@q�M�z(V�P��L������z@��x��V��OТg�d�����T:�RW�x���Ї� �ٶ?�%4�ZG��<ܲ�d5�1�*zt{:�B���uB�R�N��9J���ܜ)7H(�1!����V�0zPEČS�}���Y˥�pt����*P�ޒ!A��>C	�0t|3��&gK)����<ӭ-��&z����������A�Lo�BZ'��3E�Crq���X�hȫ@"J�q�����J�{��(샙��`�fmBC��p���u�k��Y�@�$h�h�E�4��m1����g;#qF��V+h=*V����N�זj��>z�#��.���>��)A:�I>!����us)�����B�[�'���[�]gȄ��)SB`+_������\��Cޗ:��:VZP�$�i�����m�ďbG�QH��s��K�a�E�UVN�;����p��@�<I��=�\�?����(_i5���wf����wޝ�z��!���e��?�ҏE����)������M�l�w�e�Ƒ�v[�g+�HiM��釂��О����6΄�#����S���1l:���3v��RΑviH���~�Ż�^\7��eqs���B|�
^�zoC�~1��~����]<������
U�2��s=]�f8V���SI�L�p���~��[@��r	Zޯ�?u����֍��4wR=�O��E��v�Y���n��<<� �Y�M ��;Aiq��է]Q�81Y��!M�f��5꒠y�E]ϣ����vO�ؒ�Y���׮�T�3{�[�I�d������a���[5��sgx� }ha�"��p>�B�>Xe�E��<��z_LP���fS���#`�,l�tO|�S�yAWm��ĔYO����6U"��\d�����|���߽�o���&��B���쥺 ���"������,V%�',}Tz)Q�["�J����]�W���w�W���%���d��=k�\�c:M�K���\��F�/Ö��0��+bi�c�a����������"*!P{�h���P����܁M������a�c���t�T��BcLo�ym��f.�N�k�Ug̔�q���Z!���?c+bj�|��>�?��D1�;�`��)F�a|H�KJ��[��#���b�éH,o�4ae�h;R��i���ef����ė+?�z����1# H7Ǘș������۔�@)��,�enll~����m�.q�h��K>~�O|q�Hm�k���{,�Ք�΃�*
���X#�[�~Ky43���_�����p �LQ]M��VeY�Mͺ�&�6����@�q2@�G��G�7����j�b~��z�s*5��Fu~a�ܦ,n�|�<lǸܞ�����AW�o���<�ʗ&�hߣ�#� ;J�V�v�5�VohᄰW�j=�=P>�ۋ����#���-�"��]�p���ѭ��2�ݐ`<�;4H�Y�X�U�V��%ZY��W@��S�9�g.�	�J~��V�� ���TifM؊��U�3yn8VI��g�:q��5ͼfЦ����M_*�I��$ؼW#���1l��}qE��¬�J��W�VӜ�oFTa�=�<��1	���$P��sP���z������z?y<�'�$��7$������$qw���&�w�ϗ���&'N/~3��_���@%s�LT̏l�0ﲿ4ⴄ�fxF��n�P�*��`�^V�t���d̉~�y��� ��2ù2O��S�.Q&�I}0OV�A�`M,�\�OV�mŢ���=-6��P;�ql����6�}:}�/7'�סT_���\n��E��y�V7�pS�~a��Ra�G'�}w�ӵ�z���H �l��Y�S]�Kj@�8�lL,D\l��,�]bde>�dB�I.�bqe���F<�4�}��WܰTc��U���ǭ˫�~���t:�}�4q�LS٪{Z���\�r�x�S
q=0=HN������+�8uZ�'odOV����r~��6{c_U-�'�M�Fפ���ʌ��|[8䠽i�D��ұ� h#�:B�=���/�[�S,q�+�����>A�Ӈ\:4 ��~����ɖ�y�ھe�ѣ��]���`��0/2�Q �V?o��{��ҹ�#��r����7�D+@�0׌g�ț��? s��b@�{��f�T97>�%��<y��Q�1�wd�v� ������f��Px�� �-|b�=�>P�%�b���5 ���e��{�Y���m鶊��1���]{Y*[rv�'4|�6G�᳜��� ��c�Y>�Ik]J���jP�k�D�����(:�"����L�������"����:,�%<�[kE� ��&F��q����P|ժ�QSd�+�c�HL���r�a��'|��8G| r	~�:��
G895 �,p�0�j�ض��y`lwU1Uxq��5�,��JQ�Q�.���l�[�c������lG��
�yu�hE��$�e��S�|e��ģ�z��uyVL�p�����R.܎�o�^aL^?�LN`���f?x2�p%��5��ϱ��O�k�}]�i_jy�#g*6U4��x�;G�fp<�����Kioc�{t��;��~h�IZ�sV�꘠�غ��E�Ŋ\���7.Bڧ���qӯ��.�^q��~,T�&�(���R�I)^�����|����O	��_,�x���'�.�CG�Y��Ib�9�X�Q����O�� [�j��� ;ݕ#D�@j-Z� z�fÅV��n��W&�7���F��r�5K�apm�kj�����R�M�Š�}�JgC�2��^Ttb�&
��{����߻���N�z���ZRPy��Z-�������'����H��m����qᏣ��ϠЌ���*�Oo ��%��~V�_%�H/���G�d�#S,�2A[�gG'��˷s��u��]GaJd���J�[��n��l
[Ĝ�2��0��!�%�i�M�@^��s�aV�Z�%��48I��$�!�9���n��C���������5��۾��I��MK�|��_ZZ%�9�$YY�t�����PΜ�P�2�3i�����xx�t|�or@
��»���񬾈�FSn鿒�#p%(��ly���ޭ �CJUuA���n�#��*+���V�&���d�<R�]��m�!�a3�qw����8D� v��N�j�b��Y����&ɌJ�ٟ����	�<��� 	p�R��/%��.CR۾q#�`a;�#��������$Al�xZxL�[	e�_�G1�o�c5�bo���b���V4q'ϥ0�8Kpx'��0�X��_B�E!���jfT��}�ۭ2��E�g^1����L+�ɞ@
�e<�cLG�s�\w��f��~ٓ=��U��X�n2ƪȑ([(C�cY `[袉�C��X}t�Q��oB���W*q�1s���(������.%˃u��2�=�����MW�zs����U�1�����]��U�YR��#%"�
�q=��Q�
B
D�7)K��m�H�8yi�a�؞�s����7��,���:�.6��:}��X	�&�r�$zU2��@H�WCu���{�'�=�4����	��*#]Uw5�W�zD)��8����6 ͻ_S��q�:� ԣ��%Jtop�1�Uԉ��`�D��[��68����A'B�a����D6J��A�-�F�f3(a�ȑ�3�xr�؏z=�W�IA�Ȯ'�a���P����� q�Xv\��E�)��H�u&b!�a�,����s��2q�k����}�S�P��]ȲG����9��=���;s/c`厲t������E	��M`������Db6�r�Jo�l�d6[��ͣztiW�(�� T|�������)�QLye����w�P�v�xD��V�����a��U�tFXv �ucw�q_�՛��rv�ڪ�J�"�<���8ݾIh�Ƭ���>��b�8�{�I._5"5^��x�{�#�,��_�_�|���f��\n�K��oy��q RA&�c����cZ���K5�u���*%�7�4��*E�5���[T�����?�����eU2=cn��@+mf���=\�
۳/�c�*�%,��|a�w$�@���9`8F��u�;��[ط��ma��^µP.|�PH�����	dڱD�c	{3H�+�
N�˴���M,��ǔ/ ������5��)�����&�a�/�^�Zs�כ�]aM�fg:P,1(+%�Enk���k����;2L���tֱ���*�;�da�pes�ކp�������K�\(��)cZv�`��|��+T������[1�(�z�G��9���:�Um=�.B�ZpNh���ç�d*X��y���1l{���}v}Yg�}*��S�	�D�.u�)�����mǒɠM���>�,�?!�����{���k[(/�\>@�Z)]}�C3�
q����l���x&B�%`n�7-�E͗i�3� �X����A�7��{<�')��Њ4�W
X�ۅt�<f�|-�r�z���'߉c�K�%6�x��H��ѦQϛ۴u1��UVr��=��<�)E�ߔ!�^mS};$)P`-�p���Ԋ���(��Ԡg�2��7=T�.�=_:k��(լ�����s�e	��-�	�[�F�LF��Z7�=a��j�2SS3c�oy�\��C�sl�������<d�Bި�W$�qx��y����H�����(.�>��e�gm��4�Y_g���(6;���1wܑ�8ᴂ(Z��˝'�W%0޺��zO�G�1Ҋh��Q!E�QǦ������;���
<�8�rS�/M�^���&��������*�H�{i�8{� �@�!;�v7W�u2=M�9�v֊XH���B�$�o͌�`�+��s��¸:����
l��w+FO`��5������Y��l����a�=Aʉ�$O�@�P7@��Ԗٵ���2����ehl,V0��Q�]��(]��%��/����n�3�t��0���$�O�2|=�6C�M���α�"( n��	�o,�9)��ؤb��{��/>�B�����B����|��p�7m�qy��@6GI�/$J��i��^���)�����'K�����-燐n�7���+%��9}Qm@S�b&�O�)���N/��1�Y����f�]����� ��ҳI뤵_�`��Il�xzEq�`�j�sdA#���Z��77%��<�N��"C&=q,Y�Y���8�����Y2�7�둩4�ȵ�v�3�kl@>�%�eh�6Q4��ί.����8z� |�H��g��RsM�آ캒z�y�����p���
Iy�ڤJ�N(A�Sw��Q$+a
�}[�G�I�O1�!�A��Y`%��y�H��_�#x��LdR8��cV�b��т �2_�+G���٤Rm^�Ҹ�o�ҫЯ0T�n,  �o�0�Ѩ�*��[��n���}�
<2n�S�M�{�]�P�����A�����q��Q6�C l"���5�� �%�8:]2!���$����=�Z&�}\�أ�w�G�$�C��{�啖m.���,9z*{�տ�[�'�e�� Ȍ���r���i샅A�F��LߨA�r3�j)c��g�LMB�^^&i���a���6WQ��@���xs�ᖫH�n<C5%����a��fJ��OZ`�y���g]�-�\��f�5�Krs�?(�\��j\��O`����cz:�*� Xc:���}�H����y�P'�$5�:��_�39�y�Bz���2C��*ݧ�U���Qӏ�(/w͛Hj�gN�!G����ʼ�A���Tc{9������-}᢭	�1|I���AQ��!�&��ⱰV,���A|��8�ӭ)�}��~��C вD���jSK1�X�i�_D����еp����B�����&�(/��V*��߽�ԃ�4&'�D�v��uգ�9���.0���.ĕ����Ǐ9+��D�W�3���}Y�C�`S��}o����ۑ?�G������v5IҘ��]�1&��x��/�$�w�
(���䴔A�N��5dc[_]�Ut V�0��Q��O�|���� H�c��)�
�;��y�Ƈ�
j�{c�6St����6|��=��D���~oS�c�,WX��u�A��V���,0C��0T��������qFGD߄U�c����a��$q���X���$�q�fe?���*"�pC������qx%qm?*�*���7����e�I�j�oBc��+ۅ޽�O8myl���<5�<��h�5T���E��>5�������v�)���z��tV���%������6�����n)9�^'�(���c�m���8���Ɛ��J~�A��@P����NH��ӟ��^닖�d��˅�@L&�kV��-:�Up�p�m�zmBN>�'�Q����T�[�\Ё�	��n��aӛ�z�x�Ƚ����v��J�럑��2J��:��U���D�G�����`�{�JK9
�r��b�u\�W���g���mqb�Ъ�r��J�)��gO��ɲ=W���4l�W>���Q'���Ah�R_�_�T�'�kjn_;5����ż�I�'�Z�fS�"�O|���G�V&���ݓ�-w�zܤ��uh�����*�s��غ�V�۸�Xp� ^�w,u�;d��ur��m�#{n�?}�`s�:AU�/���mA�P�m{�n ���2�?6y�>?��
.24�Iz�5�G�$0!C<I] �EnL����!��YUD�=Y�������آ9`����Qօ�?��y��V����1��y@RuSZ,�"Ok���J�*6��G�*��������f�k	��F�#���:܈�5`1�Nح@l�ˤ{1aꜾ�R�vt`���DjQ�L�h����M��f�S ܶ���hn`��A�!��.��z��09�l}I����M(�����@r���J�I{�h��ߴ���e~\�(4��bd�����t�{���-P�1�	+<���m������Z��G������j�.�[_nB��;\\�{�-*�ӆ��@s`g�"ډnC��X���1E[D�`�X9'e�Upc9�"�hw�e�G�G_�9U"#���'���q�5�K8���}��u���<G�3�gK�����~�`^���<y�>�g\T��A9����bqI�F�� n���;����~�r^��c��p���_�AJ�)�ƂK}��v��o� ׾3~!`7�� '�S��+ɷ���A���]�t���x�M�[�U�eJ�m��#�-_���R�g�խx�I��vs ���`�-  ���Lo��}-�",l�zcu-��,���>n��x�Z��k3�dԅ�x����)j�*-z�w���k�lPP�'v�n�a��H�w�����w�� ��	th3A�}�0m$������4{��̺�"�����.�@�j߀�lWN��[{�+�	�pQ�� L��q�JH��fn���#݇P(/��d��Vn����H�zuϧ(�E�
��(V�afV,z�J0�:�P��Uz���Ka�G3�D(/�u���.�٣��0�}�����W���ep�B��O�`4��H߰p.��������֙�Jw�Ix)�5Zd"�e^^�Ǫ���o����bT]n�~�i�;bֽ�f� �6��A��Jё"��ƪFQ�.��N���d�[��F�A��$ �r��I�X�z��4�;�z���L�w�5���b��A�P[U��OR̃�����߲�::*��t��g5Ź���+@8�P�$m�〩�fv~?z{�����D͑�E'����r��f �C��/-RP�F�DǘX�(P�8�eV�ލ�R/8B�m	oD��GG��i��Y�$��O��_�`�{/��;�� 7�u>P�V��S����#YO�8��RX5�.3W[���]dP��d�4�O͢��0�e�ΎȒd��g��� f�UGgQ�;��NmI5.�z@�ytZ�H��o�Sb�\�Z�P>�r���D0����#��0��#�+��x��_��㇙͖�Ce�������սi��0#����Y�rg����4۽���8>��Gp$���[#v_��#Rx:��$�00��U�$�4�/<�{��5�*���Ʈ�kļ�כb���R[�j
kw��$:\{;��?,�b��X��6*���� n�X��v�f>��W��n��X��#6����b�Y[X�.�W(Z����SmS!t�/�-�����S}.癫Ф n�)e�� ��	����^��J�����Zz�CUXg���[ꐺ
�����T̺N�j�b�`
��j:�}�� հ;��Iv��A�n�i�f9��4N��Xt�����(�{�F^V^��6Ƭ�n���FTO�jnk.��[C"Ii\�==�aN���(e��4:+\�o�E��Î� ���3^�K�*G3-Q���R��j�[������q���릮�T����&MC(&؁���,�A������M6�Pp�j ����F-xUml�<���?ɤA"X-�Ŕ%�3����s��B}�$�����l�u�2'j�1 �,����:
x����#��w[:ǩ�0*G�.E���c♙@K�=�#�l"�Q�wn�,����{+J���c_t`E?�.�J�9��7��I^��#�%�Y�>B����w�Fo�P9�Yp��C�SK���(�&�3Dv��Q*��L�Ĥe����#w��I��oi&��)w�[2����V�[�:m�4G�&D�V(*�Q��t��>βqyx�T|pZ[�Ы|@#���#lF+6�v��!�3.�|�̨a(Z)4�~BEg�J��K��CJ�#@�t$��Wm��YIq"��V�ae���uY�h���������f�Jw���9z�K�D�5�;����B��� S�H��p�\l�U.����a�k�zKo9�휞h�A�N�D�GNy�
p�=!<I8��4�����!κ�N߉
��ءD|2Ң~���r'�$��$:�/�|P����
LX���`���x&�9�V��;�1nt�U�Y!W���*�\'=+�`����*��ЬG�-C� ���-U�����!!H�.1+A�Ӱ�J�%���zr�S�b�6���Iw��R�uq^�p����������Z?d�r%��0M)x���D�ӯ�_�@�_$ f��>28�%[�1ۻ�z].�N����a��5�J'I5x�/��o���G�5�N�!�B;�a3D8-{�_w��e�>��D�0 u�ٓ�x{I�9�����E���rr��4n��W��5p��!q��i��T�Kw;�]�������,���ML�Ό���c�F�t0,��V��}���
��3)�p.%|�˶'���2�!X|�]�JI����� T��H���}Bҵ�.�Zr������<TQe�qƂt_E���X�6�z���dA����� A�=�6@qDV|y��-��n�K�qڱ��H�aO|�'P��q� �݂$]X��2�"0�ڹ
ܬ�s5\���$���g�u}�d�O�P�^�m��<x�R�
}�@hV����NK�Am�E�q8������A�����ܥpjc�-��4���vW�M����q��w��ܮeO�/�6Ф�����aB�h��b�$.}|?06��v[oJ��Le��YG!\�� <ߵ�	ُ�V4�	�*���=�[ַC�
��q'=��X&gw�BфhygJ7:&�8����e1�-�'���������-�����9�����g�5GS�si"iŴ�%v�DI��H�\s�d�x����P�o�w7���]��g�
el����~��$����������W��`>��1�����I{������*�4�,���b�����Q	� ѷ_F�=&Nm鐙v�`y8Y�&����{��=-G��*�Q]�� �F=������bo�M.��yJCu�࿜��ŋ�Q[a8$*"�����\@4K���E���'���A�]�a���Xz��=7y�w����H�v��{�}|x���K�3�qj��I"���Z�O�����B�?�8�;ϛ��j:����D�Zc��l�,�C&|�5��Ճ^l�jܴ�C�P����Fpp��t��=LS��<}6�2�Z����~�!!����1�*�\��_Z~P*���[K��T�'�z��`��Cc5��W�z����k���)��.��=���<��kÞ(2K�)!�T�\��R=�$����,F':o�1�:{K9]�4{P��a��NW�Z���Ap�zo6ӠPÈ^�Co��ь���ٳ^��d��\�M%�F��V��J����N����I-�ΠnuR�J�N�� ��Ml0�ӥĸr�FK.�Sk��@�3�iOV0|�.>�)1����y��D7�~�+0Q /x?!UF��ӗ9Bԣ+�AN2��߱��Wڵ�'�W�B�rs�/�k����G��G;j��0�wn0:O���t��{jx��G��d�#�̶�<��N���[�19L��|kXP����%�ɺ��v��7�o!���8�V�	[�?������TX���mwy5�+���i�Y��b�pK�H�H��ݿ� C7B�R��1�u"B�T��%SV�;s
E�N�`D�do'ګ����^��2�Gv�Q~:���ٙ��z0����_�P���"��F�>Ӱu��Mmp�B�9}yoEk��-Q�c���G��8����
�+	����C��;�i���y]���Ҧ1�i���R[d<y��oj��Oץ/h��dǝ�Y�6���|q>0s���T��g }��G!�����{CZ���q���w�����5���5i���\������mG�^&�Dsm�k�ja?��c�������?n613��F��H� �2,Gw	[��9�w�Bŗ<~K���u?=�2'�'�H��H����\>̏P��7�*3�9�������U���L_K�F�FJ�C���@.�3����>ҿ�=m��L��K��Z�M2J���8]�D��j7�pI�%8�\a��\�"G��PW�Wq���G0�H6���9�z OF{f7�Z�R|J��O�!�~���4�����W� �lL��d�P,��Ѿ��ԋ�'~�Y�hc��f����ێ��-�h���7!4�(���Evy�1O&�'���������֭��E���u�fI>/��u�4������V5��D�M:�oUS]S�chr����)K@��d�l_�T,�?o�
�:�6�����{���Ie�qJ�I���L�A�V�Q"�Ť�.0r���spM����ڊ��JoJ��㚔�N���U���wl�"��6ȧ1�)��Q�5Q�Y-)����7�ݻE|`��3�x&�_�Q�4�Hk@S[�9�6�o��s*�&e�T�]�5��/n8���U����.�����G���9�����C��@} n&(�C�}w��j�d��?qڎpcmc���@C�@��3Fn�U$A�M��;�L�-y�r����i��u,S��!����$i���q�_nM�籫�B��'��;�95�����m�Ա�v#��5Q+�z���Ly]%��C�ϲ�M�ӄ�-h�~-X�R���	!��p,�q�\�Jq��څ������)	짽3�
=�\�Ө25�e����H��3���~�B3S����T��1���,%(hɒ�Zy�̬\^<�?a�b�߮��t~A�㲀3]Ɇ�>��Ha���/�'�	Q��-�t�	�U�(um��d����<4�{����g)��*�I������W���mD9����e+-�8�H{��n�-jso8��j�Igt�ڣ��Sp�?a�pZ�W�/��f~,���-x�g{!�̇���ӊ
�Π�G��_PFxG��`�2�%{!9$ׯ�%�P��  Z�W�s��9�Ғ Za=�|�'7�H}�V�nr��X]�#���Vc׬�
�2�F���$3�]�����b����[I�2�[����Ʒ�E��0ue?���I�5N�I?��>��Yp�h�^��ċ��ȑYӉ���nuTK�y\v�
I��\��UЁc��żf9�s����Z?K��B�W5��i%{�2}�}��).��4w�G���H]���L�ơ���nɗ&]��s�Hd�1�c���-
�"����ۖ�s`$6�f��fe&?9+�� #���~���;�b�#�ڋ����+�t�&�Y�O=|��?�2��g���'6��~ø?<���K�Yj,�ԉ�:��b�9?������^��6G�l���&&wȊd�7��c��4p�!L|Y��'3��Ib��}�7 /�f;�*�R�b�@D{��=�^2麪=�w��+�Z�3Ԉ��
Ź0hvPR3J���$}���5@���r[�GRϼ	���<N��vx�9�O����!�hӨ�(�&�W�(h~E�Ĥ���"� �)Y�V��l"����
���B,���?�Rxǁ[b�J?za���;r^I����r�Oѳ�ckk*����#�O��p��Ni�1y)�V���Ċ�&ɑ�@�-US��q֊R%�?��g��c�����)�1;���Ș�M������;rl�u�O9��?�Q��ca�c�a�R�Y�?u��
>���_�k����j�����?��|����(���6r�0�p�l�hv�ٚ����S��*R��:��������^?:��Y;��.�v�h������!��	�:"x
&S�HG�C^'%��M[������`�8�'��Q-����Kn����2��@���e�Đӥ�]�Ѵf5�-�3{��R��T���/5�����
>���7�a�����2l�q��x����.�r,�1�vh@#���M!�]���e��k^_N��C<�XB�鼣��V�g���}aO�e9l��/zk�vG��]��O<�S�b��ieh����s���!��7��^H����<���o͚#z��7"o�����	`�IF?�c;�����ѝ�[t���Z0l���i���V �� Q:](��?H�?	�
��xvp�����3��o
�+���Ģv��.�YyK��ïv��������F3z�r�pth�q�)7e�35C��Í�]Urx|��DKs���+UZ��1����}���ƃ�8B���?^ ��N�F�K�S�Am5/ȏ"�Ƒ�}�9�R���v$�U�r���i<�4�A�Ü��a,jۑ����=d�.C��7�}������BUϼ�\n��d���9Еw�B6�q#���}�I~/�]g~�Ϭ%�fy�Q�}�,v%���]�A������@��m�h ���,��_,�������hyC���>N ]��d�f)n���Ut��htL$5m��g�F���܈���?XdJ\L�0��M���Al�7_l4�7�K����[��ˊ�Ê������+���	|fwD�7Q���o<����:�}�����p~���HK�To��Y��rvyc�u)�]1�#k�W;���S��#�le��a'�^(e�$�&��B���b�o�8�����q�:����?4|���Β.d��n�'�d��uuL#}�����9�B��u�2.�P��~���|e|�x٘����ʨd�J'�JtV���I1�H�������|�c���Z�����5/R�P7�c ���4k�pu���2��`��Ŋ �Oѐ4'��C	1�K�Dh��35�E2D� ��[��n#X8���'f2s���|��r��"܅��2�"͓�dZ�h-���4@���{D)��\�H3��F�OL�4��+IN/��D�d�W0��Cqv�ϴ�ju���{�/P(�Ji´V�`+�H)	Z�dY���2�y��6�϶�X?��L�����,�+�*�\lq��c�*���L�I>ΝB�]GG���x��e���@�V��>m4�W�Z�����q�c�2��I'�7��reL�K�c�V�*��5k�|N{��"!�̲�PSF4�s��v]��N��YUN��i���p�v� �m,�1�g�UQ������ג�}�f箊�w,d�;|�B���L�}V�x���(���	����qf`5zo���� Π���S��Qv��s�<�:�DE3�m�Ȟ��!��I�O�x)=wb���˴&�t�H���<��2����d趘��q�Rs����댋zEƸh�r��i!��.N`�=��~%�9��D�n�b�����
vf�Yx]5�0�Ss˼,���;F:r������Ō���d��1z�9��p���UILl��������ǁ�}	���d�\/h��#��$��S�~���F�tJ��t�c1��1�,-���^����稆��o����1�x�s�{}�{�$2NZ�/i!0���KZ�˯���؆�-]��2�M��XZ3� ���Pb�%�ң�y��!��Y�.�	�[��+�6�\X������sSu��B�z}���=�q�U��v3��tR�3)
&���b<��L0p��d���)w3� 6�*Y@P�����,Gۣ|�jҵd���D���ՠ�h�Y�A+ �is��#n��9<.�{��q��1���s�8�����Mp#��l�X+t�icb^�����<a�?�_�aD?��N��ϕ@��&�������t���F��.��ac�~�͐0�]߲	y��-�8B��<�s�O�+K6E���;�V9=w�coS#�"������O�����$U�MYR~��ŹS�˓�˹Z�.&Ť�퍢R5�z�`_NJ2�Ϩ2�yfQ;�=c�*�:s����3W��5iQWD>���	Oݿ�m3֌�)f4y߹�.��y�(<�8p�@m�#�Ģ�6�y�Vﮍ���%D���[��1h���}o'k�(��K���h �h�b�*d�y��%*8~"��%�K��Mʜ;,�(+h�P�vN<�DƤ&E�8x4�V��-��A�3n��N���?o����n	2Cl{� iD���
Gql�Ú�9�oͨ�a��#�ש������`���?��"a�=
��[�=`&(�~)�˾�0E�څ����h��w��޵<s��h�{����&��;�vw�3I�j�Dvޑ��G� ޻��g��Jd�5�����-0Dї�r�ǖ3`��k4C��N��P�W����)�|_&s
o�z,8�"Zue�M�u�Z�8qB�(���P1�t��"�j�;�e�C/�v�Tt��A�4<�6:�K���4w1Y�^��5K=f�	���x���i3b���{-0ʆ`�$*�uMm̜��Ig�P��#���Vd�r��`6�[G��}�lkhB~6]�7M���G�(�d�Avm��3�"�8���и�s&�	z�:�l��$E��f�CJW3�qMF���������0��%��(6�0�@�>�~C�H(�[u�E9�iEՏ�;�M�`R��G��
}jZRq�9����������,��w#D����KeS�0��jp�V�#k#~0��hwc��"'��h4�s�����g�]ͺ��`)��Wt+s�Y�:1E�b��8��"[j��!����g����;@i�`��{�b{!S�W�A	و��Q��s��N#a�m)O��{<q!D�sC�AJ� E+b@�؅fF��Z�g5�y��i�C�"��i�Q)7�kߛ��gj:!��, Nj�)1؜��y�5[δ�)�J<�<��^�Eևm���p��j!��sÄf�f?I��[}w��ò�֢("���~m���w_}���)�i˥;�M�t(5��Ī�
Ӂ ���j�4��Q%�i���\�\�X^�Q���;����DŶ��T�s~6py��dq������zg�3�
J�l11ؙv�����S{���͂�-M�Q+�5r��V_Ēh!�'�a����H́H�.j!Z1QKK�;��g߸N�2����e;��ݓ���Z�r���'_L�Rg-d��Qv���z�;�@���V�q		�Y��;H���|p�K%��*�5�P��I�)�	��<TwY�
�����O�k<PWT#/�	*�-�u�M�:yn� Ĩ:��S燴t�.���~�jM�����k�u�Q�+�o���l*��T�i�I��cYѫ	��=�O�@4�dp�d6"���ę2���z���)�I�*�X%����(���������Ň�j�F_Ҩ1v�3����(?9����=?QڕXk<K����"����M+'4 �u�J(Ls�:8ggq���,2Χ�G��'d6�h��bU��r9N)�Y��c;~�ٔ�{�/A["�˿@1Q#0�4�����b���Qs(��f`�\�0�b� 9[�Di�ֆ���}�?�H|�J@�p�ܽ�:B��x�_�V��/[�g}��3��
���6�����{�]G� ��Xu�C0��2�}G�Z���u��i�i]�-���x��#B��Y$F �N��L�9 Z����U{R�p�Gڕݳ��.>g//ߖqH�t#�?�GK�c�!54�|-��ȧ!N�;	ά�m�m���	��v¿4!�����ϔ�4i~����3ĸ���~CG���xJ��y��5Г9����f�"��Yb���(!ԉ�P����]l�~���7���:����#maеEO�r>?�k���Q��p
��b'_mQ��,9�ވo;#�Sx�op��1[6i���O�Ъ�=]��<�/��a��n�.u`y ��S��Īh �D�Q����S����1J���Ě� �^�D�.v��G���T}����16`�+���,�u���q��YL���k9#�C�M�X�j7�i�~\��W�s����	Ä���x���SY�*�^�ؕ�>����tDn���ּ�.��_�V�PO1��qD	�ٝt�]�Pn}���/�����F9��{���XH��B��cUfrl�y�܊1:����>��T��kh8d�;��y2_���f�
�W"�� �)�&�F64��x��1��*� Fѝ�8\�.QX�g�����d�6�Ly �]���Q���wHDc��%��e&���-����=%CG |�B���?�1fS9�s$��W����t��UG)����0�Q��Ն}��A����A��eB���KwK���d��k��.��")T[(C�>��?H o�S���CU�1z���c
�������&��b�+8��ֽ1�L]��r	^�gc���u;$�hT�b�*���[yx�	Lp��<եӛίYҐS���j�n	�R3����%ړwO�sﭥ�t!�X�皶>��$�P6��lr���u����_��i�-:�oH"����Q�찯\����X����m&#���k{㊐}�\uv��Ɋ��,���%Slgv�%kF;�Ү����;l��i[C�.~�`*�C����taVt���S�� �nM�ʧ�O*Ù��
.uV�JJ���/��$���S�Fᒥ�o%���4k�|u���A���LNy�<f���_;}a�|��NJYZ��َ��ڥ�a�I��T�$mO7��&�o{v�;���!�T�[Ϡ\9ʑUy��d��J�������oՕ���
@|~�R�/d��p���
�H V��7�.R so$Cˆ��|�y1Lh�����-&)�=+>�i�h���w���1���?Ool�{oûe��x��#~�BŸNw1W�iwGxZ�|j1��#��T(Z�e��|`N��$�g����<t�e?�#Fx�&�Z��$����������J��@��0n�9����o��ƒ���gM=��� �>�y4������#ޫ�c��)-x�ϙ����z�T�s��K�4�g��%b�g2��甾�$e@q�CT�ls>wwC�o�����{�,�����f�3��ϕ�c��h�FlVU��SI:u�FH]$Faz�Z{���A(U�>�d��>�#s����`@&�޾���<�3�b*'RF!�3�be���2�a��i鸐dCT��w��x�~F���dqBX*���b��w�F��}����b���<RufI�k��	��9���5�Ğ���2g��l���8��%g��2 �"D�p���f��V};�W��iF�]t���6�x'0����
?j�Q됼��#��ׯ������0vI��9�`_`���4r�+�P�L��:�4ܵ�\(_e^܍r�|ln�����,�z���`�~��0�Z�,��x©e��n�5�ȼu�L�[JH�Ç��n�������oM��N�)��I�||��5L �(��QQ98R@�`A��4��co,�a%tS!"΍��- u��u��dav��߅w;e������v4�U��StC�b<�A�{�X���=mՒ�1"��η�W��y�mpk��7�=��p<�9\������>��j�F���Y�hh�yH�u�a�"���ZB�MXl�_'F�*Sc��\(�ҕL�����q٠�<�s�u�z��e?N˼�/>���7t���9	��ߧk�h�M|E.-jWH�@��],��}1ry��O짉�	,@4�1�`gB�o�q���@�B�Hkc��]H�^���O6���'ŭޡ�8Z1����t4���ᶭ�ǎIx��o	���� ��6c#������^r������yإ4q,�U�.Δ����=�v�����l�T����)M��
F.�3�#����a��;\�����L�faj^K�q�p[ޚq�r�^�|��\H�o��c��kU2}ȡm"�ZM���%{&B�P�ڿ¯3�a6du!�x&�V����&%$��"��ĕ<㮍ǺZo-�X��橦��>̔��|X~�4&�"P����f�㝂�nS�<�Sn\���L?|������z���#��Q,t��S��M�^�Ov~_~t:U[�NSўܳ��طø"(���)�GbV6� J��10��n�8H!�D��j��?t`$_�ϳ��>�����%�"H��w /������������ٯ�Ish�v��WĻeGTg���o���JR͝U����������K�E���_�"2�������������K�y�jk�ܺU=y1f������|��}���+���LPx�v�%�L>4OV���%{�W]ؠY0M{�0�G��9xA���@,)�$�
oC�1G�lcR^FҋE��˟M
�_�6^I���қ�73���1j���#[�&�kn�mT�ʈ������Kuٴ�@�������q������h�J/0��mꠙ}~K��ѲƮP��u� �_�0�V�Cgb�kv�݇�����󭝣w�)�������E��]��zz���}�<�-�t�!�t�'O���V���������Ń
����o��Yb_�q	QI�R^ȟ�P�}�/�=z���-�>^�|/�D�U�=F�Lw�D�,��%c�<�;C쮦�5;��&Zd�8%F��.h��@��f+��O>6OM[5#B+�8�����	.��V���X�մs���{��A�7�{�}�x�&�v���|H���!G#F#9����܅�	�,)�*�~r�+@��V�ꥧ"\���g^�{V�Q%�(��ۭ��;��ꖚ��d��;���-�W;1!G����}�ÜU�t�����f��s^2�L�E�>���!҈�D����֘�}�bh����g���g�܎��1�4�e��[%&��,!���� �گvhP`p�"�{���o�{%�"�������yU� � Hס�%�

��(��Q7�J�
�F��"��7,�7/Jٴ�x:���]��wp�CZM:�ǐ�P�l�H��f}d�(��0G	�}o~UW������N�&O5����gΉ��a��j��?Q�=A��+S"�j�7����kd"�Z�c���tt�>ɏC���8}B�=�^6# "������M�6D�a�E���`�'�!N��k59�+A�ݐxV*�y��>���\�т�V�]Q�3���H���$�i��4��eh1A{	Ȳ�#�Tʮ{��S���%���R�Ԅ��ȹ5B	��rqt��j�PTS��� �*Hf���:�̏�佖U�<�^o��;�қK��-�K��v�"wuT�7�8\��<��tK	����汇�^�C��E~�$a��A���д�����頵�ؘ�VFe�*V���@8�_��A �Ʉt�oD�YYB��b��Ff �}M��:��Mc �}V�Zk�-�|��O�����GJ��lࣱ�ߐQB�e7���nyr�V�@��D%ڒUf!�X��	�a<�;��/�uD���ǥ$žK��O��BiE��X2��$7_�o8@� �7ó��%k~0@4�i�R1�i2O}ϔ~�i{�U�K;~�۵�I���F�]f����Կ~�z��{ r5�S��R��%cǝ.[Ӣp�oG:�?0�.[��0�VP�w��<��OZ�Ҽ
ɏ�{�:�-�n�_?ʁ��u\1��mq��u%�ǌ����ޚ���M��Ru�>7Y{E:�d6�(^���_Y]2�xn~�����mn>m>!jDL�|[���49r1?�Z��o���]��P��=�M��)�7�$��{y��2��I���7@��$(p������81:���H�v(�#S`U��ڌv�j�-�>��<���TϜW*�J�5�U��3<c.��7ӫU6��,�(�7r}�.�����8uژ$�>Gr�n��[Ȼ��������rj@�ntu^��-����b�2���U�>�jr!fj�����=�Z�����@`r����!^��e��v�w��W�1;n
�J�kP#_��J�Z5�nd]��*'x���JX`,m�-u�J{��fu����9�=��&��U��W��9��ޯ
ɲ�7<Wᩏq�V�u���y�Q!�y��Ś��s�ʌ�׆f�i=E/�p�`��2l�����$��,���d����]a������vrx��>�6viR�~�[���r�·	�&k-��;lN�B^�$J3�@7��?��(��·@`|I��b2�`1o��/hN��%-����2r��N�?*	�S��k����;�a\�{�prRxH���הշY ��G59|knjt���t�l߂�|y��	��6�)��K���K�|Z��}�,߼���xM~��l�Aj1��$���9R����S��9o�j9C��L��ķIHWn�iqrN$2�J>q8���F�-��j��ָ��o�e	J�Lڻ��Y�����:f��-�6�ޚ�H:QU�p(O%X3��'ڇr��+��_�r���s4.to���cC⁹�|_�������0��N�V�b~�! �M����4�4u,�mӂ�D��3V�eqnH\a�̷��'bv1�d��E_����+�<K�[����,�%m!�����5�6Z ,��l
r���dQ[�����Γ�̣$�P�04æ��O�F�������я+�)TX,\0�����~4�����r	����ΈL��g2{��	���^�OXk@�~�7� ��'n�$EZ�]��O��(N�A�;��IGP9���	��FUd;2��7�&D_�_S ���wn�N�o����.>�)�#�\r��7'K7fjx��NZ.��:H���o��F����{Ν����r��N�)����4И6�z�1T�?sD��C'�����o�)�a�!�1�;���+Mח� a������IyZѢE�cR�ɦ�\���h�g8��Y�/j 53�,>���GB�e�-�,�sx�߬!���Y���1��a�ds�mw���d��t�3��<\�� q��R��t@>d���һ��h
5Q�Y�G�������$����ۓW�-��2;>V~�%f�G$�����j}�}h�[��k)�U/N�U�-�}0���T?ClI��֌��y�\Vx]T�f��;'�2��V8��"���^��1�����F�戵O曬A��q���H���J���VrF���\?��f��3���Ń����:|����M��	dc�8$*1^5@����(+W���U�C��T��&��V������lx��������ݘ���5F^���u�(�Rv�y�Ϩ��.tԭs�5����]�s%i����`� x���tޥV�6�U���z��q������J�O�Î��5�JU�/'�ݯXg�u��7nZOdS��σ�:ߙ���	��Y�f���<�z��vO�����b@��W�
X�-���A���_!�B|L�L⨕'4�ƞ̺pKC�i��.y�`՘�v2�oP�)L�꼏=~JR6ݎM��h����Z��icˍ�"ཆ��b#8K��R��Y_i�V��\<A>���H�9��^*�aj�fŠ�{5��XN	��fm�T4҉�'�h5��ԯP����z�>y۔'��JR�4������~�\+A���%�rY��l�ו��~��:�_��4=�UE�������@
z߂x���	��d��9��e��-��KmF�P���&4k	�+�j�W������Q�O�=�v ��XC��y�;���U�̶NP#RX�&�m�
��'ش��dx�Kw��b)�Eo�5�a�^�p�?���a�ĝ�c!2a�T�oyɀ@��5Ƹ2��\YL�
����P�\�ޏ�E#�5�f�N���;\�}j��L_7ђ�u���o7}YPK˃Y�Aggc���6���T�2il������ A,������b}�+K�;#�p�g�]8�l�g_&#� :��T�u}=O�*���X�)yqa���=���vS��-����2�\t������������$����c3��[6�ߐ1�p	�8����[�Abm������{�����u�&>�ԭ�fc��|J�%fnp��\�����j���B�_K�"Yp�0Ϡ�Q� �Ս�2j��cAةE��Z�3�t�L�-�Y����+��:���P�TTi
�aVG����<�°�>�H�b��B�z�֑�[������Y�,�I4�J�b+�q�sJZ�d]��n]�J�� �t�$15�2�vx+�F��&D��)l�P�G�%���$9��ګ$3l�l���!0=����z�S-��쏤pv�@}�('����E�+��Mp���]jG��i�;D�r�s
�IH��e'67��Pu����E�%��g�0<�� :_#��#�e�7��a_M�w[�:{w+�l��/�KCi�$��v$p�P/k����"�cv���ӡ?Q���4��s_�YW�i0�c����bfqV26m������*�ŒO�]X��x���z8��h0��f���0�6v,q�/��n��k0�*=Yt�g�F��j"���5qbG9}� ���(yД��D�<����Q�;G�ֻ��7 F=���&�_g&Y8����p��/��h��}�`�<Hڡ�ZKo�Q���D����_���mv�(J���r��ӝJ]r5�:�-6�����ZSZ'N��)��w�z��U��f����+�T�)E�DOT�<�e>z�G�$�-�����+^���^�7hs�xVvl�a��\�:�m�l"Ԛ�4vB*੅����!�J���e�i�������m��KNnvT�ʌ���2�(r p���i#�M�� �����`1wDV��O?��^��]�N�N���f�E�Q�嶑��7ƬF����U���IWGu'o�p������D�0U�2�l�$�b�Y&A`��5����i��;^�[wWd�+W�5٣؅:�����$�T>�-YQ�oY&M����x
�r���b�7�E�7�w6���¤��Oz��Z�c��4�Kda��5#���:��	.��(��!	�i�/-��h�X%����������LL��������m��-o������;�M��8���Oj^(t߿�]4!M�o �<�� ,����rU7��q�oۋd6y��k{�j����HH[@����ߍ�����y"a�HE�-p�^ދ��&I�z�\�3S�ւR&$:��M�ʒl��D��&c�2�����9��7�=M6��>�`0W�;Hۼ���ol@blr���:���͠K�U,eO�����Ej�95z.U�ԁ~*(Y߆j�[�<����k+� qb�H3�%�&tsC���f��c�P����o|���	99MY�v�l5%
ļ3pkߨ��d�`�F���ܸ����mydZmD%ʞٺ�Q�H��
H����x��T0,s~���K5k����Y� tXA��,	�]���v�e��o��#%���`熆lQ���\���)�9�l!G���.��#h�'Etd��N]y�|nȉ|��N�m�x%"|� �Ѕ\W\cg��5�V���V325A����^�o�*w��qfˑ�a���������MB�I��)H!�8�5��&�T�@�;��;y�u�ZQ���M�aJv�0'���͇��;ήZ-���ae}蹕~(ue�
���3zr|�A�[�\�����Fs�gҾ.�;J�Ʉ��'��
*�ply�����dh&�G ���k�]�GѤ"��c�f!"93� ����_�q�4��,�S��}�w�K=��z3�g�ӄ�
t��:�턊����hZ���KwȂE�F���sX	b��17�p+l�f׶�0�����VK|+cc���?6xCZ�# ����"Hx�iX���Xȡ׊O�!"4�ܘW�csľ�p���l�2�i���U�	���>�u�F�7��[j���J%�S����;h�����s�y):!�����bQ�������Js��r�[~ ��'�eE�SJ��$�|�5�:�X��b�7���u��N_v�]T�Di��.sۺk��Bе���� T�G�smj�aV� �S,(��z �ʾ�7������R�B��E���	�3��<��
o0`�����M����ؗ�7���"�y����7�H�9~��O��GT���돟X4Q=z}{`��'��,	��Ux��Q��Ɛs����W�߇Lr�ƨ�VƑ��6��BB�h @��D,3^u����r�������RfN�}W>��s� Ⓓ��*����rV�Ԕ�J"'F7K�Uh�h���7g���!6
��%�F8�O�@!9� V�Fo¶>#V�-�]ZQ���,(��2��HZ\w�f� �P-@�7?��ڝB�����m*@���h�kk���D*O����w���#�9��5l�AD�i��̴] ��]g�+��֒`���%�+��ZG�@���P|�;�8+1R]�j��-��f��ЇC2��5�¤��>��zK1�9x�n��+�' ��uޑq����&�S)��Qaȋ'��AG6���s�u���|�sm?H�nY�u�&~��x��L���@���}�� K��kt��t�e�*�$An�]x9ņ_�cüFB:ڊ��
L_.�ʢ�zk�oM�*�ʦ�41��Vw)�,w�la�,svY����P}��עQ9&�����VşE�w,���M��ǲ@;Cɫv�6�_~�m�8�1��Cĵ�?�W�˦1(��J9�iQuv':5nj����K�q�S����f��`�۸�^�6س����U=_�\�<���@�\ހᲵ�G`�8;����E�ȭ��w��b�q~�vV�	�3!�+�?Q2m��0��-s��`$���18��qR�������Np�\�K�n���,q�}Td���|�sJ��XP���T[� C����������-y� �G��0�}I�A�Ҕ����0�j���|�8�d9�����]����W�`n��s�r$2��N(}`���HI������3�Q�gKF���U�#ގ��|z+������0I�fb��Ɣ�,�������ꒀ2�U�����l3�0m(�&'��n��3�뽴���'�����ko2���|�h|��}���n�g$k�l;1��#��5Y�: �YlO�w�\y�&�3AQ�zM���c��a��d�P�>apn���Wl�����!E��0�B��E�B�Bu�~�2�W�-e@b����3K�p@�뢨lG:s��(w�덕:t�H$)^��������U�⶞��-�\49_s�+��X�͂To�D0j/..�yG9�Ȋ�9%���~	������?�%�d�����?�J�-���6�	�Ia.N�L�*����*4��t��3�c0G��g���"��N��Ԉ�V����[���F�)W'9�>��o���t��Y���o�n���	O�8p2���g��@(p�&/���>�_���ϥ��۵��ٚ^�	��D��=_5�^�_�ڀ7t������2�XR3ʿ�n�;t9u��gv�ۈ皚sOB5{��6�D�I~kp�Bk�U��6)�w�g����ҥ���H ��wۓ&��Dc�J��F�e&�B�fP튝�cgڊ�5� �v*�Q*�|�F��m;��O��5��\?t�r�c��u�d�a��=�Ͳz�b�X2<�<F���i��J��x��9�:d�@�R��W�PU�*�I��@�W��,�.��ƽ}/+HI�|�J��A�M�$�2���ZQx���� 	�~��(N���>�C�/������ǉw���4I=���K�I�ňK�Fs�i�q�����ieL���б��}z��62�]��FGcF�bJ\���Zo�Xp����}_�+����[����>�o+��&�*jt�s9
X�(,�c��w�&m��$���vc;�l�b�ԥ<Q�w��zY������ ��x�79�n����-0�~�y��/�A�%�G�ęM���0�;k��X��g�k��� ���� .3�+�a���+�~�{�Vԭ��le�;m�����$�%I6�0�g��1�i�&���S'�;EJ�{���z���W^Y�~D�_��N��n�� ˸�44�+���eOHƸv����~g���f�k<���aÏ�J�b��O��
1Q*�|*I���9��}M������V�!qo�����Ȧ-���ѓ2�8�t=ͻ�$�%��RF��);�g#�ۓ�5O�ea����}n�#u���b��2�A�����V�.���Ǖ�/y�s���s��[�~��J6"ؐ���Xʹ�,2�����G�{�.�o�7�5A	١�%��!5��u�;%�1�Y��ߝ��E�F^��/	�b[Cc���k�U7S��9*��n�!��,3�m�H���&�O��I[0��E�e�@�0ay�i�(����0�����犄�T�=36�m�o8�M��`$�Ӄs$�+�^�.�y�s�Lۙ���F9��~�EC�m�֑*��;�,�}��P��CU�D�=7�f� f����Q�ē0�������`�"�>;6�%PJ���Ol�w�~\.�����C ��э����Z>�h���&�kN|�ٺ���|���qy\â���5%�*� dG��L�D�t��:��#���C9-���&�ĐՄ7�b�69ec�I�Gr���!%}�qN�5m6�<P��v�g3�����SK�f���Vi\�`�rf�W����m3�f��\L��q^2N ��8G�ER�~���K0P�}r鮯�VE"�KE�Xo�,!�U#k����E�7��8ދÀ.�!7)`�aZ�;�:�Sd"�K+=X��������;o�p�^���}^��:�)���	&�u2�Cv��g�2�:Uo��
��G���ȩ� ,��0Q#�I�(_��R�w���%��H_��4��y�G�Q�n��ۜ�Z+�%~������B;�.Nzv����9��d��[*�Mn���=����������4�a�Lo��_6�뭣��q_O� ��nsFW$=�F�obs���^SSc�zx�!R��Z)u�Z���9T6�������ӑ��sjm)9�/����_�^�׍6�%>0�n��Ʋ�N-jE�)$��WUҙ�xՒ8�Xr�a' �܋h����F]��@��
�O�ꌅ!��Ϯ�\��9p�9R�ä
�pS�̂���Do���J^-F����S�,��լx��K��ʤ��y�<�Z��vUyn��/���vܵM�l��&���� �dd|��˪t�{AL)3�zE�d��{�4M>JsW����7C�ȼ����IL|�'�]�v�l"#��L#��Ń���h�E{��)t���?ƃ�� �/�&'w��d���\~����f�̕{kgję_?0��a��iӾ�j�xfj�,����\�Q��,�����6r��v�	4�z��i���C2�p��� p"�)�\������>_�ʃ��;�/	%QS\�t�[#������?%�W)ݳ��Y�K��ͬ�34R���/�Q��3I�ɫF)��zo����Ќ���A=��\D�2A�A󢿚ۓ���BHkC �Ch��hX9<p�[ԣ�#갤+$��F9�4������lu��ס��yK���3v��h�HMX|L֡���]qg��<�z��>`H�ˬ�)w��%����as�Wh	��:ѭ��jZ���FM�) &�)�O�Mj�1��Ft��- �zS���L��6���_�u��o�̸��FF73�[{TVN��������]����$��]��^���+~[?M:�>C�&���i�~�/�L]��>6���R]�*ܴ������fM?ߚ ��a�KZ�+f��8�`)��#�X�|T���7�K �P���w(��P�*�
'��?��Uҋfx&B�b��Z���G	�ok_�i�j�pE�}�?�j8#�D�$��˰�j��Nb�E���x���74��D��"5I�e#�J� �Rq��g1��,�[Q�����)���%:*�dC�z���/��ntG��HV�(XU�V�*�@��x(	�O-	��rʷ��(�+^�/��|���^�3��ǉE�������E���`��k%�71�M��&�}U��_��8w>c��y�y�������E�"䍾c4���$3M(��_�@�Dm����u�v��'R�4U��k+��&7-����o��n����D~�_o ���ЄI��������˲>�Eήp/�}Id�� �ϙnf�����:��
���8bD�����d��Ӵ��+,�_�\�L��bI�����<�lg���?z�v1X(���o��褽t��AXA�x3 �b^����h�ɭ�b�u���ZA�G�P�Mc�U[3Ӧ�cۇ�gI��n�9��p��;*]���'� D8��wD��ֱ�vN��	�SJ�7�5ǡ�.oaV�Y��i*h�z�F��N���;tGw��M�]��x+�/j���c��7����X��[����[�R���e�SW�����ɨU���ݙ˗T+���?�K�u��m3��������
�����a�P�|�.�Ί,97�}�,� u�]��<�Q�c��f�c�2��.~A*����=�@7�y�Ѓy�b�2Yۺ��KN�"&��Z�B�S�wx ߓ!i������z{5'���+��f��b\O��RVvF�WK�'s�u�}ɍo�(SԂ;l�7��9Qшp1ht��G�7BP� �˪��m�j*�0�˻l�{vIM�ޕ�)��S���y+���ox�i��&[�^ˤ���WpF�
��}�������<!;8���L\~�):�%8�U�R��E�t�v�҈��2�7I���Q>=��}Cʝ�+��Cq��Ru��������7o�E��恀7��m���Zy�}��p�_��5 I�p�TN�=��a��ҏ'Z��	���7�%M���TB��e����$��a�~�xh23�����W,�d��x���23�a,	Y���i�>yarO`Q<�����Z��"|P��0�1΍��$1-�?$�q^����� �gV�!�эxA���[v��ḳ���ӳ�Ҍ-�4G��e���m���.�Y����b_�.���r���x'��K�C��L�:$rx�x�ΛH����(�Z���J���ݞ����8��p�89f���m���%��;��G�Grwg3$�^��u�vo�'w�l�>���xz�?��lY̖��^���RR��#�dqP7|�����m���}jH�,��O~�cs ��(&#�"ʫ
^��3"X@����-y���l�ڥ�j@B̓/�Hм�
Hʟu���3�����j�N��/�d0�rY�Ξ��~��a�hnE��ͧ3��?�vs@
14T�
�B��.��uH,�-~R$�M*8�� D�*G��V�3Wvx�q����qP�b��A#^�x���J\�<��e�n��,	���oz'Vܩ���D^���N��ʧ��%�X��,_�y$Θ�����z�G�|=���b�T�n��Y�!*�`�������s���sN�T����Q�b��#q�6�X�����������[�KF����e)qLw6鳅�V7�n�Y������#%pƁm�f4�"�J`#9����I�l���G�E�m j:B���.��uNWQG�V=hy��t]�1h,z���$��N*�`�#/ր4(�J	ӳo,~bid~��i{G�57�2��ȯ{GJ�.���Qf�V���%aF@�\��)�Π+�Lj�u�4�D���13u�)Zլg _�� ��?�?�62/��߇{��1�)�)?��n=[�J���v{��DҕW.#�T��.f�M�e=�&s��PC�ш��v�����$z٩�DwS����ӑy���}���^�?	5��1���H��S(QO�<��4"����h�@h��}@2%�i/`�h�0r����d�����j��v����[O�hn�\P�x_1�Z��;!���_���G�g���0�ƺ��dOEԬtS��a�J�)����咢�+�s�QLv��F�\�������睌��),��.{�������Sޒ��md����0Km3�5I�}���X��k��	����as3�;���\P��=сH�ݑ�^81ۡ�  n�=+��U�/}]�P��A�Î�3��j�*��BK���|�gf9�T,�n{<o�8�P!�5�5�Le���L�u#ʕE�C��~i�h����m�!�@e[��R����`)��O�U�h�Tm%���ӧ�c3�^|I]�X>�
{�
�z%�� �9˄��fp�ў�g��5;�����@Ê7�6\dW�{n�Ɋ>�c�.�`H�>;�J�=І�rj�p�!:fæ�Nu(�o]�������l�\�b��X���W��H�ո�d����JBj�6�hw#�+ۋ��,@3>�����(�U���x������AN=���/�\;��'�������v��P�l��.#2��R?냬�(i�}.s��N��h1�VŊ�	)o`��d�C�� 5`�J�������2I�{��R�q�\&C��o~�}.���F���SL��y�h�`*��Ϥ�J`ܻ�˿�}���ݸ9%zz;m|���S� �L��+���I��N���
Ux�Mb�SOG�S�k�F���-S�y����CR� ���#� ۇD��oT���5 !�"��ԣ�zЂ	A�'W�J���3��"~d�������8!�F�V�SX��8�*>GJ�
�u�����:����t�"��a����$J޾?������0�vƇ&�m������#�jt
g����H�i>L��9�g9�|��,��v���/h�����!�q�DR ����s�I}��2�#yZ���6M>�M������}9�Q4bF'��qv܇5�`H򌻲��mhm�z'�Y.-���b�ٿ2��|i��QĲQ���؞�����_?՘���/��E�:���	,���@�p�QM}�r�)�͝����$տ�܄�� :�ܢ��B���$�{�u�H~�v�[�9����h�0��1��n� 
�e/bֱ��G-jeDT� �ѻT�ʴY���n�DV��ݍ�7���5c���h�WK�Ô���%���EPX�c�<��|�,��K�zp<�+.X��k����n����c�#��ۙ�5j�ow��� e������ ��Rj^D���v�� ��w@I�@�E�D^��{ �˭=B;�y�y�DǕ�X����;��C�'����鞲3��~L-٬W�9������@�ǫF��X�n� ����eʃ�y��ײ��hagY�8�� XL�g��zg�-S�A#Y8��`\!��n��TթI+�0�42��j���=|9���5�#�n�;G|&U&���Cd��Q�;��5В��J5���n������dV�S�� �,>��֡�XQ~b]�-i��#{�a�k��m��3�3Щ~ݹ�]�6X�^���E�C�j��Qz"D����?#������h�Ɨ�q�ܲ3T���s�K!B^��ř�b���R����Z"ΙR���z��h�ۜ����̜_ZV�:;��P_]���Dx�7;�,9��n��ײ�y���[!�BNʱ����T�[f����w�e�\j�c��zi-˵b�,@9p����N���aW"�E>�'0Үe��nPg!�E6@`@��D�F�RP8Ə5���X'�(��t���?���ٟ�#�̐�N�_�\"�7B���Cᬄ�>�\O�7����������2�,n�*5�<r����z�y�PT:V
?ǲ�c�C�O(cg�����C(3P�ő�H$䃻����ZJ���##wQ*o�[�Cmݙ�ᐥA$Y����kxG�//��!g���CM݉�b��v��\�G�X��4���aP����>�GkY§�ﾽ��;4�_�8S �(��!��
%?%B\M6z�H��I#�ņ�>:��u�f�^��d-C��]�^ӏ��M��&���`�}�V��R����u�g�<_��v��y���АP�x�UZh<G۽���/4|�\��SY���"�Y�}'54vҲ�[2��b�X�}[�;�}^n���>Slw+��~{�+"Q������1�Z�'D"�����������x��{���?ۓ�f �q|;{���d"���*R}��? Kv�
,��`�["A��y|�(J������/G��qz��?:2s�\��2�-�.5��e��\��o�jJ�C�~�P������^�Ư�_������^t��Ie�l32�*���u)�iN#�<��Z��=h�;��5������?C��$���ßl��#�8�2<���H�´�WнAVgc$�;��i{q|��lp�;O['����~n���uBZ� �?Z���K�,��?�Ls0����'.�'����7���<���/��8�����eH<p,2���c$b�rgx�gvH;���#X������8��;%/�ۛ2�Ј�T��=pt�Y��U&ZCP� i�� 7�R1.�&�EW�����(��%���g�6� :�!@1fD�x��7�TI
��������5���E��'F���e,6d�i$p� _I���X�i�ѭ�'4��s���+%C��c������2��^㻌Ѕ�oG|{n��K����z$h�s��T�o�r�)Wh71��5*�p����P�������	��c���U_Fۼ^�y��%W&�j���E�����Bpc�q��VK�rӁ4	j��	�l2B6��}�U�������?0?���펏h�#r}�Q�_aj�MQM]ccK !��8�R*2��ON�T���4���u�Ns1�+�t?އ��j"?�e�)Y��ll�c��z�` $,����D�fh4�t�5�+v�\�4��ʨ��I�F�)�����^�SϢ6ki&�B�֒��,!Ycq�5�f��t�� ؗ{��~�sFr�H9	�q*/M2f��.��H������Dʄ�S�rCcھ?����)^�%�Cb5�ˣ���N�_U����(�,+T��"�bٝ�1"����YcW�B��Cf���竂�,Y>,���A�ֻ���=3��3)Ӂ=���/�ޠ�J�A"��P1K��2�B�˕���s��2�:��1F94<g���@O>A �	D �,��geZh1.]g�3����n9��
W�
�)��dr�@��HY�`\m��\�T24e���,9�`�)�.]M&�c����Xy�9+k�kg��H� ������e���ޤ�}���9�Lr��d�9xBpm3͐�s��i�RL���|�m[&�P����I��<y'"c�toH�ڱ��瑓$�q5����,[ɟ�N�u֋Ƹ�G$�d�6����SM��j���]yo	I2�k�]~�6�z;�l[�8E���UЩ�c�����K,������C���l��GC9Ɔ���L�-�ǐ�T_䣕���Dx���0��e��>�8���@������7�y� �6���aUN��ZX@g���K����ݫҴQi?�}}���d�V�f�PR�U|�D��3QVvMc�=�k_�}0�V�w��v/�^���*���e�U�tl�*ɷ�kv�Q��mՍ�0���?�R���%%���B=�P5�a~�Nn��ȭ|�uK��)\V�!l�f>��0�d �W�j�!�"Y�ۑ�;%!H��PW{��
6Y4*6�&����4� 0�3��2�s�3�Ck�9�]Zt��O;"�1o���r	�@�GP�$���B
�����"A��T��HP2�\��C^���?�M���ζg��`V)HLwܭk40��D�����b�dm'�4i�a#66����+�Ǹ ���_WO �j�K1?a�˹�EB,�nDV:�#����xJ�3��q�i��-��t��jJ���J�`�SZ���'<���$-F�n�[l���\�'��J)�MD$��ߊ�,#�{�1\��\����,/��k��R}�f���j���������)�,�GG�1t��'%ۨ]E� �
ʔ�t,� m� FD�� '�KM��������
R�-9����u���sD���%z��U.�+�D�^��Hb%����Кn�wgf�s�B��RP�g�	zzw�����s^e'�=
�)(�.�Zqt���d[���(�#�B���s{>
���3�]���d9_6*N�N��&w�%����� �7!��Ҵ�E�)�l���U)D4��
h<���l�5�K�� j:��@�\4�!>@7������"@�2 u�a=w�~�If��!��%T�l,PQW�~�cP���nH�$���𫗺}z�]W�4��n��Ή��05��f4���t��_���M9�����t�!��RI0��Y}xs^�ݦ��M&w�Q�^#�?�gU��+��A�%���K�YLy&%������9V�Yو��M�d�߂���ξh`Z�!��O�XQ�s�6|���'	�d�}������Y�*���jhj"��?�[�	��=���@;�^�'�#�*����[�G'Nj�ip-yܴ���.��H�'L��1��xq"��K(lǃ�zkm�ca�A�2U&���u���Y������NΊR�K]*��u��-ͩu���tַ��x^��)� �}�`o��Cm�̣nz�h�p���)������j�
�#!
(�NJ����Jp=��/4�v�W�n�H<��d�W�� �_�CJK�f��fٞl�У%l������v���P�%�E���ܑg��Б�9]0TH�S�+�p\��\���iot���kl������r���ә���Џ9��ߋ4�bgj���/�)�i�*����O��2�0�)��a�y@���8��<����Z����b�G8�	Ȃ
{ t\������m��+9xī����*f �	,��]#��PY�������_�S���v�LzL���w��$k�"�����B���4���n=p�Np�T�$��bi�`I�6_���%�<����������͙�hfX��b�'��0��-�cg�Q�}QE� ����"�Uo�f!��؃��b�+����o�@k)��\�>�KV��Ps�+̓�Zc߁ݍ�X�����
G�G-�;m�h���2�:�h 0Lx�:��"͠w!#Z��W�"����V28�؊{n_�Dh'�������"E��Fgz��~�s+,nE����8}①T�����n���G��D��]m��Y�M
�VJW���} ƍF������<�������V�2Oʹ'�kv������0��7�1��M�*vM�,*e-l�Y�%�$')�CLK��Q�u����e���!�Z�^A�i��`�w�op�<@�����K�7[��LeLP
�����ՔǇF����o1<7���ap7}[���`t{�r��l�~����Jo���|Z���M�&�u�U 5�|d��,��ؚxa�~���}#��AG���_�kgU$ #H�	�j
y�J��~��Rc𦟛:��`����jݗ�} ̩�7*�~�����R}V��5&a�C�׊����5�"��[�I4^�"���g�����M.y
����cDѡR��x�e{���O�nhq��b��[�a��K���kX��	�ktƝQY~b�}d�i�,8�MD��X�j���8ӭ��oװ�,e�=_�x+M�=�d�0�㋡)eK��6�V�*/J��l����g��<�����1�enhЇL-Q{'\t��{���)zׇ�X$Lk��iqskqFVDz]�Y"i����.�*�)z�9S�V�?kJឮ�Բ�}��h�Y^�;�w��|�`������%A�"{���Ue�ȶ��}�O��{F{N�N��
c>(���qK7}Z���B�?�S�fTf�.B{M�
��@и���T˵z}��~�P(/�w8q5KL����Ū��	0�8k��`K�Κ�RC�TT:U:��>����-�%��?F�/�٪�-_z����2�ϷE��B^�쓌̅iY�Bd�����N�^t�U`�n��	�>A�g,+��ę��K��2�7!h��m�o����Q&�(J*���!���/-���C�*����9 ��<��������߆����_5���{��#/�Of]�<�RjT�r�v+d���7�ظj�����sY�Rѩk�J'�%��뚅�D罄��]ӁTe8��/"�bL�����Gҽ�����dv<a�6�T�|U9��.�n?�u^���"�vY²Gi a�P����[c�pלo>=D:��i��6��8�*!���Ф�9��j��u$��{��XC`�����8Y��lFL��c��� 2d.�߆���K�lm(�]�o�����RXM�M�ɔ��For��q�b�%��Lr�O�g����i���n�_�*�&���͊�z��3��㦅����Wi�.Q2�"�oA��8-ý[�t_��s��oMTY
�%J���k�w-`]�5��Uh9!9�g���>ލjt��ǵ���N��*�OW�x�XsޢƗ��)ﵬ�	�0�U ����p�D�ܦT���aI�5k�V��.#ށo�j`� ьe-���!w��7��v��BZ�%�#;���Nٻ$�M��_'���it,t��� �{�t26a^^��S"���Dd"��,"�H�~��Ӌ�����JZ����x�mzjx��:P�ٹ)��h��tp{��K�4��N��'�Zo��ҩr��zƦH}���.��)YQ�H���:���j��\���_36����D�*t�LF��x��u�D
e~_z4�gk�����L� ��I�٤*Ѡ�M,�8M�1ce�(�Wϧ�-N��ث;��?��+��TǤ֜{j-�lxj�s�	���$\*���*��2����Y+�V���	��KS�vP��ҤON��aE``A��ʵynr��ѱ熎�#�Y�#�B%��kΟ� ~4�A�a��YR8�s�� *��m-�z��*��\w�ݡ����ȵ)ǲ�+�ʍv�/vR���Pz�)R�k�g����/= p>ʎ�<ⷉ����'V#ǵ��������B#%��� �3�aS�u��<��e+N�$YZ;�J�$Ed��`l��AH���%� ^v����x	�W���&�ۡ,I��iG���W��i� X|��:6g<�yDRA��Ul���1 k��g`/�no��=Zmj���4EU��H@�Dp��=Y�e,v�g�t��.V�Ej��Il�q=I�/��;2H^}\�?�I��c�m��7�C���ڍ@m�����&��ؙ�����5��!r�a�?�4�&���7��.�x�T�ה������V�00����R�k�L�M��s�٨Zd�|�`_�t�c뱇1��^J�^'�_��9�F6����$���d�3���7�Y�P��MʙG�X�J��FDX�/�c�؀}R!Z�_��X�8La�m�
�͏s�8�#Hf���=u'��r4�sf\8g�*��Mw�]�p�a��lo���G`�1!�����c?cG3�Rɩ�}�z��9Ȭ0�&�w�;n�cG�I�C�cC�u�o�� �m�eg��a�����5�--X�6!�����~{�K}�@}jr�� W�E�:r�O�.W�'R�#��T���[&eb�O ɣ��eh�:�Y�
�QVm%�YO�z���.��Uv�G,
�+����?�Mz!]U��4���G��S���b�5��*�'�\mU>7cq��_�i7DF�l9����=˱�xP�
�ʋ�ʚ�Ҁ3V&l7������~�f��C(0���S 8}
�L+��2��$4�"z�JJҰo	nj���}9i��,bFpp���l�Z}P*B��_���߷F�aY���C/^��� �jU�
`��5(��-Q��Ԅ��7r8}�y��t˄S���y���9����j���t���~MrB��$�'���|:�[�I?�U&K�9p��U_�<��\�g�`�M%E�^��3��x�����5jK�������]���F����
]x���,�`�/�L=4q�㑂���� ���<�	���f�Y���=��������tu!nC��*ӏ�N�G}�O[��3��>������ĩ0�CyΠ�8��j��eƷO��L@˦I�vѪ��Ģ3���mӡ�5\���p��Hi�k�ͅ�����MK���]B�F]͂�雞�q����2��JA��Q�Jy,Z4gE���7���t�}cOp3
����Pz��n��v�Q���Y�Wm	�8J�5N�Q)�[�~þ_a#�.���U��-�)1D
\�5!�~�w�1���3�D����S�t|C3�O�T����R�ww;�����؜Dy`Xzj7��5�́$ƅ�
��\�"���-�ku�{`���zFӔ�����
�`-�!� �N�V���N" .�jI'_b��ɵ�ׯ���2a;�l��R+9��!��[g�D��l�j�h�G	|�P�sg�"rn��跍�o4�Z�k.�J_�^"}#���Zl��F�&����AjMmp.ş�st� ��&� ��e� ��)Wv�/2�[���+7,*@�)���g9�1��u%����n{�>�x�|�����cC�T 7JTJZh����
E�'s��˫e|�F�S������0�����;)Fl/P�]WR�hfk�a��s�Ud �6.��F:����b.[�Zdtb�jQyI� ��(E��/X����J�Զ�n �O �ba���؝���H��ze��\r�E�'�v9x��u6�fϬ���Bz}������(��z~��5�<�DVH:�&J*<߂�S�N���D����� ���ϰn89�ޤ� ��1d ��~.k�U�+@y����1���l�W�{�˗��0Y����\ӹ@�\�v/\����/9�PF���X*�A��ѵJR�jP��a~��sR�IvU)�9:[)g?Ζ�
>#Y͞^B�B-�JC�y9i�����+���q�³&�G��A2�e�`�,�J��Nn��t�R��+���ǯ�6�a��a ee��1`� ����揵W�8��)�Dx�N'w^*c����Vm�y��CT���舩BR����@��˳��:/{�kgA�t/QG�w{sr���^��瑩/+��X!�_����S�����v�t��	�#��x�މU�Ͱ4u�����S��@"IA�X������ѩF1�;L��O�k�/D	Uǳ��;��ڮEv~G�b;�M<�@�*�P�⭟�����bcLds�*M��	E�'�48���?����j��ρ���#W��+�gh�o&�F�8�\���u��#@��^Ӌ!���]l:���^
�x@���B�	ϝ��%�{�l���<BC#�U��͗���h��!���(�%j�B��vdz3�	#V
j�E ��7�v�:�n��n0j�~>Q-~nq{�Ώ.�0��Y�J(w/H�M��c�=����ׂ�=�2��3&N�Oߠ^�C5u}I�4
-Gg��9vڥ� f�c��[���B2���m{Oe�Fg@��)��5��< �O�?�s�:�g�������%��8Dk����{ ���2Z��g��<i�7��Q�>�YF�S�ܵ8�O���e���c���bhC�_�ద1��6@��f���d⑒�9z��q��K�l��o���g�"�/�m)���p�>󬻄KFJG[�L���[�� K�>�'��+��2��4������&zɼ�j���N)�n�)��?����U=z"(ʉ����s�)���\�*J�c�8�Ī�i�TN���y����K�,�������Y*�{��r�
�-Pm��P���V�m?* ��TH�����e@�c$6���,�+��H&���r0�I�-���8ˮn.!�7,���5EH������t{�9�����	o��3�ʭ#��S�Ӷ ���h�j�D���v���Ȩb6�'���X��b�HWt���U���N߶��u�a���IĪ#q�=N�y�2C6G��Fp�%�.���C��s�ȣ�宇�P��S$]�#v�����G�����D�`t��Q@�8b����A��p��P���v����!������_~����@����X��߯g��u N�3�@��}�Gc�-H!���:����fa�{v�>w	��U�=7e�2� ZX�j�z�,����Y�?�3�a��Q"`������\bJ4%�����[f��!|*	�v�g�)��&�;ɜR��n�0�] ��2��,��N^8d�5jبo%��Y)�3�\��޽���0Kч���q�ߘ����^X}�.���E�: ��N���T���d��E�iGgǬ�����{�*J�C������з#QLsh�|f��?r�t9�:�=����8f�.f[�>0��hH�B1<&G����� h#A��&U�O��a7.*�p���@g�$%�X��2,��dx.*��ou��lS�ީ���9nv������:sa����Xl�cM�ئ��7�������d_��7��h!K�)�qy]�Kn%�z����zg9VqIY��.�û�=���;i�Ӆr�cjC����8[�F����9|���0�Nt������`�q�2���t�ŗay��4��	��S7'N�GÅchK]��,L����A�1]i�:�d����R�M5E�2�{,��9�OZ�^f�NZ��]Dp[�TX�J���eav,ZQ��U{ �a3ӄ�!�fǶ�DR�E����n�ƓxSI��-Q����pE$�#y������E��g�8)�)@�ư�"��]�#��;�N�m�&���g�L���\,8�U������D���]x3@��$|Zv��
�L��.��⊿�p�|��ze���`F�=G7�i���
�K��xb�K���L�	l��Š�6�F���7zn�:�	]��1�`�K��kX����)��<��hE��=uI9���:��q��UW�f��t�.`c~����#ז,��B_.+oL�0�/�L\��ʑ�Mj�jp��®!̡"C+wVA��� /Ci��gp�<T�tv`�Z�-�^u����I�ħ^>�2����[�fӐ����> -�gi�3��׶� ��h�5H}P�%��xc>����ٱ��/re/(X�W+e����}�/���,2���}�!�f��b��M̮��k�Ilw��Y��kaӢ�{kFg ��cHXU�����v��#B:k4��N�j��?ö���h���丸��r���6�R�ՉP@���?��4�!7ՠv�q �ɲ�m(�ІH�qvi
�%b:�Eo�ɞM�q�7 ���em)�ݚ�N����e)����!�q�o�M���뀆��m�(�Tey�:����M�����yd�"�D�#��kb�h:�F���Q-N���FZ1S�=пMO��M����k�RZ�Oe8$c�1C�ۺJ$��MP�#0���/�?(�����������M��lKR~�蘄�, �P������u�r��y����4���N��L�C���)��K���|���^�ލ;T������k��vG�F�l3ŪW��!�^�k6*���~��dԝ���]�WQ�	e��[np�F�x]�d9;'/�_��c�zB�;!/	׽��wL]t���A�e[����y��ElD��c�"v8�)����ёhfR�+��}�G��e�'ޛ���(, Й�.~	 Ng��)������ne c1>��:�#�-� +:_/�oCO1_�!�}�	/��1��&z����yʄ>�>�OXֳ����,�o����͕�t9���ĔQ�UE��{��$�r�m,�bi�#m��|&�Dp�CK��1����c�S�
�I�w8�N�E9�:2������Έ+�&���Gʻ�+y"�U��cϳ$IK�?�XaO�j	�ZA�r���Ǜ���[ٴ��ɩ��00��4J�d3�.9�h� ���`ݝ�?�r@��6��{�QF��Shw �}a�R{`�l)P%��9}h�!��.�z��F��#�H������J#$�������%�|
���&�LL�g�7k����#�P��-ۮ^�n:�	�qZ���n�.��E���n�I/d�f;�]�vlѵo�?���c��ś�,���硕�
�����4�%\����P��JOʹh���d���f1r�����QE� �?C�[Hm>y�g�������z{]0��M�9�I;��6��3�Q����?��[�U]A�c�4[}YM�R�zҚ��o�
D1��n����Y�7��<�,a����� �*R�]c�V�4��(w�tX�28F�ۏ�iφ���;���&���M��@�T��y��G��[W ]u*� ^��;�f��8��g��N��9�~�.$ņ���J)���oZ9�b��NMw����`y>�E����!+�<|e@�' ۶~�wt��7L����2���+Ɂ�����j�<i�����ɜ��ˆ"�i�;��]��Hn��_�|�	��=Y,�1ڬ��uTFud�Mx�Q�E��	ܡ�0��)ey�!')	�h:6"��U��W7A��_��������mP�d�S�z�3'�&�Xcb�7������#0�t�K7>]
�YVf�!�K�������U&�������?�<�&S+sQ�S&�"L��cc�sN�*P7|�4�,a
�j�ʡ�9���0�/SG �B3��vC���Y0gM�V��ܫ4�^�I���GƦ�0��ł@�vH��d�Ԯ%cɮ��Ə��ep�e��2�ـ&��ɂ���Wh�~E�ɔ,�i�7�[�Z�'�`)˽cZҮZ����3�[slT=J&�qP�g���w�#�fs(�yݔ35_�|7fp��øB7L-���2G�'c �����cW>:�&���m԰K�%닜�^��U�sn>�=�=֊���K�5��3��~~��JB�W̒�Q�D��Va��~Lԛ^*����[��Ӕ���:�$������@/V�ٛ�%�i��+�_k�RR�F�h�N�� ���߽cc+$�)��R�<�KBw��V�b�[�����0�E�`��J�~&�o�ٯN�n���l����K@���.� (Kȯ�T��E8��V��x}�).oy_�*�Ǖ9s%dٸ�~	�B��̨������t�q��:Bu� ���Ó�v��H���� ai~�ҡƍ'��q��c�� ���l��	�V�d���2@��j�H���=>��)�%�t��H�9�5�Vg��z֝γ�cM��0��Y�/(�I,/�Z��Y>ܦh,�}����"o�Y���8,-�r��e�u%S�]	�r#�#Y�^ֽ'H4}���+�v�s�`�>^���k����O����y�D�Q	��L���DX�ry7)���1&1���3��!]�2�A//-Ezw�ٕ���a:�5oQs&�<��7sم.� �5|�	�Ŧ��?�'�7Q�o
67�ndkImu�9L�'�ek��		��	����z�O��\��|>-Z��4~��:2o�s��4}�̪�a�Va��i<*g�%��-ggfCO'q�!�9d`$�
G��O�ח���_��g����|���������2&o�Phu�D�Y��o����;ؤ.��$=��| �S*zE�0B�ћ�::x �Xz�p����c���wߧ�	K��I�:Hќ����e����r��{��nI�JB p
7����mr�&��