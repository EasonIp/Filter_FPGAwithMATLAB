��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$����v�{A6�����Z\c����]�rz+����D�2G 9���'��6�iΐʞ@ϰ�35Ne�X��=�p��՞�8�c����ض�d��F1
a���]a3D��yp{ೣfq����E���B��X��ӏ6���)r����=� ��3�ft�d�Ӌ4�9�6��*������ċh8%�d�.%��7>}�oꕿ~q
Hc��e�Z�QԚ)�/*r]n;�_|Sǹդk&d�Hj��?װa�O�9;��&m�߁������"Ҳ��wٷ%]C&]��ϾR��k��ۖ�ÆYmE��J(�&8h�	ڊL���d����>c�US�CKPIi�/�������⋘FKG�5�`͏�N�|ݝ�֮�� ���ɺ�G;aEf�ʨ67wԎb�rJF�#�n�T#����EmS�L��>�c�򽜨�"�~���_�(5f���bw���`�A�����Of@'�G�.���&eT�G������`�|Nۭ4Ա��K�H�%�&�	�V�e�એ%j00���Wkx��!��NP�<�I�������hi��U�����#�Ǳs?�!��e��m�HRS��,�p����L)���a��ݎ�C"�HFE����Yz��Y���pf��~�sr-�4CH�"����:�e�n�q�;�h���W������� � ��S�/�<��)���z�8�6o^)rm�V���9�ꨘ��iį�6.kъS(2}�|�_t�fԆ��Ʃ4t♞��SH���p&��M=��*���B(����N�9,��n��F��2�٩�+<�k?!�X�����܆�ƭ-۟�1k����0;���p�x$c�� ����
ᔐǽ���(�؁α�t;�>@p[�V��� ��VF>s/Cʛ�Ы�8��Y�IS&8��==^��x?L� �8gp?�H���O>&Z�c.��-o�g��!F��'����8M��z�g��M���J^a`����G�zJ�!y����@F�C�jH8�;�7㚞ݫ��PM�O��e<��ߖj	�F��!TL��;F�;�h����ý�z� �ч�4��:_t����`NU[=A��}�6����k*�����D�9+=.�nJ�D�@�|��F]/0+�/m�س��F��� :�x9�P�|�l�ǔ�R�K���Yt�J��keE7�6�UaܲW;K�x_��B����QqI���We�Z�9�h�!_��3��ҙO)0J庢�ki
�o
t��A�L�w�71��91����l����X:�G�2�fyݕ�h�m�$3�/�8!��>D�m'��Y݆�Si��܊y1�M�1�i^3#��������&-��k���d̐!�.���8S@�T}��޺m���O�t٬�߽���Մǩ��\Q�-���K�m��"/g���A�Z} �c��D=��~G�엨��i$8�'�v�>0�Z�6t��{sљ��䪛wք�M��f�5#��9�C��qh	5{�g�z����rT
�'�.��LܖSpܾ�$F�ݷ�_ �p�*�*����T�a�""��-}NL6�Q��j��l(G�����$rxQaU/Ы��Ջna�k��fW�m�nCO��i�ȅ��ُ֮�-ls�e�v�WV��@��+��2�a�Y�oNE�yE-�����x-���2JA��!��lx5pυ3�Ś��N�`Z�ρ�޸��P6j��@�_�g��:Dc�E[x�#}%
�k�=�4+`T�܅�cx�yO���$ԙ(1�D���͠ ݫ�|��hB�9	�*��Ȟ��e�<�@�8��'���2&F�L�� �:9O�H6%�s��R��%����|��MX���
$%�U]s�{f��:g����� �]��m3���<��;�/�fC�9�4�@���W����BG���{�gv_������y7�<�����G���m�2��4����G�YiU�22��ߣ�
Қ���ZWz�(\��4ht������*l��1����%�x��͒�R��K���4����e����i�O�9�5��o���h0}��C���.K�㤊B�K�����d<L��:7Q�&�4�v��d�N�I�k	������L[DRGEI~�Lx�7� ֋���#%;��h��iA�JGԸX�~�-� ��B�jv�� `gM��j[7u;Dn�@+��.c���ː�Г��k'���F]`�`[[�ꍟ6����#���az_�*�� ��C���x��(�����mb|��[���.��Q���:��P�ӥ���1q�R�ZϹg����#y	w�������T�J	x�[����	?�J#V��F_X٭*J���#h�Y�=�� �~Dչm
�E�v��n�D���%��d���]��).����T؊�(׮�J��6���M;��x�:��h�w׍5�f�bFQP~����!�Z{� ��ݤ8�p��to���)��m���k����:��A�Jkgv�����4?pFӰ^h@�T�;�a, ��1���q*?��l��o�S6}C���s\�9Z:��XN���X��λ�r�� �R!Qz\��*�|�U�$�ʒ���s�m6!��
�hawe3��a���#�vO{	���r�V�sG�&�o�Lٳes��sYi��}�hB
��j���	뇴7�q%��#U��A�ɺ /�+�E֋��Q]\8x��f�l�^��+�2Ke	���.6$�d��	gl<o��*�%uf����;�O�yG(X��B:?�y��vS�#��g٥1�ƀ���#u�w����Ŕ��2�R3e��A�v�L�����2"'K�)&�(��:�2*��y�H�N>�`5���5�T���iQYޭ\��qw\�:O�-$��9�]L Ԑ��r�P�YOh�/������\�ڞ(��nv�*�S��B)B.n���D�$�����B_y��}S�	}b��W��[�̋�bj�]��4(�&F"��KTzr���S`�j��i���x�eB�?��Ng
��$���	�>=�,+���)5bI3���Ѵ��\j�L�p���ooBe)�`��ok�����6ـ����Ze]�n�n�$����`��5�B�DAGCn�;��C�sO5]��O��G�۪�Ѿ��
s ���5+~�.+�C{oSY`�C��w#�XՕW��,��xc��B�q��M��a�RY���{L�%r�	��Y \�^����"<2n~!��1��pg�#jY$RV�\�/]�n�&�yw/����RzY�����4�k*��"5xi�Б��ڬN��ܫ7F�xEB�.��E[�Mo��s��_���zp�����=|;x�!C�b�L�;�#�
pE ��.�e§]�^R���Ncw��U��^��0�3еh��H$c]� xA�c���QQT�36Ѿ���g��=oo��d���)8m��Ţoo�pؤcXд�VCM���㤱2j+.��P����n�VO}MK���h�?@��-R�<�9����Dn9R���,�Vs#����`������m�(a�uq�bV� /[��/�`*}�'t�O�H�ܧ'�G����'��6��-b7�FH��y���0���o��!g��� ��ɻ+��2�R���D�ӳ�s�L��/X9s�'P_h��L�,�	���i��˸aRNY��Tf�k6;�4�(���j��q�$�]>9Ѧ��)���뢎�>*H$+������8�7Dz���բB�s�Q�T������!�t����Hl4���5-�s�o�P#����MMǏ}�O�%ϛq�1��w��T���eg�d ,�1�k�=�K`Q~����EX��]�-�wF�y&.�ͨ�P��dc�s}�O���S�1tu�b� �>��5y�������_��cP�B�O���7D�9{\80gl�����^��P����ta���t��
�Dw�����Eðj��,�Fo�Tc��_�'�v5J�����ꗡ�n��	��K���GP$�*�@�/��i�Whun�wjht_6�.qrEiU��n�m�[�.I5����	�ۚ$e�"P��o6����R�"┌U�)���ǧYr�H����DB҅^fKX2�Mp����a�߳R���d&����\�p�1h>%B��8Z� "'à��)w/L_��5�<e �w��ih�x���E1\��G�{L�
��{�g�} ��ac7�L�jx܇�L�䲦b�|�iL!sf|Iw���� &��6R��pmw�/���nl�!��mz��f�A��~6�&[�(>�,��%�����k�P��esF?(b����x�k�XXj�ۛV���k����)-uht��G#�*��>�\�	a~��;�,{��֎���d���mѠ�a���v1�j��lA������C.|����n�7)�2��p�k�ܷlҠ�I!<TLQAS�t��L��^rd�����:��ż?P��F���$hZ~w��U����;�#Z8\����Pˡ�ăE�4�K�*�$�R5S$������@���=��R����L�
˘}M����ga3eA����}y�C'_��'�&!E�i��f��y�T�oX}���e���R��&1����#ؽ���]a��ت-�9����~�7�Ͼ���t�)�8=b��.��qrK��CV�o��+�#y�耛���U� ��r��t����%nuQ�V�B�����h��d��|�����J@{���6B5?-�y$�qe"^=���k*y�ac�M�:-f������Q19s���W�I=�/��.xDq�iDؼ{c��8�]W�X�8��>�"�z��Ll�mYl1�A"��jhlQ �it7��h�!h�K���V��碥R���+��D_KC�/N?���G!���x��a���xԘm�%+�ɗ�6?s��������ۛ]$7���c�j|՟S���[:�h��F��I�8��o�ff>"*�Oq��<����29a�4�*���hn�6A�2� �_��u�\B�0��5�8����Z?���Z�-�u�.�W��I��E�!��d�{���z�TQ���>4DO_�L��2�^$�P�Ae��\�N{j�l��s�h{_��&�?��)��+��;uD >�rAr��J |}�D��RTp��ۡ��K+�,��q�?Z����.�?��l��5j_�lŦ[q�����j!R0��hغ���6�j�ZlW�����o�E%K�$�i�S�|G�)�����4{;^Q�0��N����>��]Z��`�yL�H�t�)$T���c.G�~�&3@�H\L�>o�q9"��yQO�rF��2ܓXvLZ��h�8�!2R+�Lڛ�w`�s�:S�gIF���!�8`@�Z<?7)D��?/yE�m���قB햾>WU��ԉ�J��/�IE�k��z=� �v�e^/�!w��s��T��m�2V����Y>d-��R:�D�^���4����Z@��LЉ���t�^��{�1-RF����	Z��,�N���U-c3*p�)�� ���b##2�=���d���U���U��l�G	V��?��᧢<��.�6���5�"y��������*܉���X53F1�t.��ẓG'�4��[�I��B gCK�B=�`���c�1YD���F��ϓl�����c�B.�oz46/����AJ4`��kM�~JK_X(�@ =A"'��;͠�Kz'���`����W���dJ%[�yVj@ ������ݶ��p�H��3̱	l!-��F����~k=bV�P.`�	��{�{�|�������{汸�>e��L��=�IrRR_(?���_�ɮ�vh�Y4A�N;rV$B����Y���# E��.���}Kr{vk����珒���U!���^����w���G���z�QIUWBU�s%��9��`��=�����ƭ$'z�.ش�CV�W�;��w�!��)�P+�H�O�$ ���V���tVk	�C򲌽�'����FkG���^~��ɩ4�?��k
\�1���?4m>��Sf%B�sA��.1�0���h����@�xS����</ʃ<-� ���Ġk�߼���!AY���Cl�2X�f��~1��)K��3�����W:�twCJ�֩��g�k����kR��4�n��e��2Ss���}����yI�{�,۰�4�s��샖�y���?����cT�^S��ݠ�^k4���a����@&)��q��~By�E�y���t���y|_���\b����is�j�ܔ�kDa3�LGVAD�مg�㚘��G�!�|�7g<�]؍z�?Ĵ�_��Ǒ��Ѐ�&�(��L͒M������lyB��#�&?ԩP�����Zo�w�h$��RpbS��c~}����P���v3�� qT�������?�񥫬�D�%P|m�g�yٓ��!E���A=|�����6\`)��#�146�C'�tތ�{u��'�q��ﴄ��f���|��ل�4�ӛW���������R5��w�t�����-:��c��x�� U�9*�I}�f��)H��8����-!�Ze\N����뙮᭡�=��+��WT�G,��/�:��`��:�n���F�/Xބ�Q�O�~G�y� �AW�j۳	ٲ�>��W���� ��8.�a�����6ٝ�����
V*��q�|O�u����"6�
a��,{����`�P���J��)J�\��p���iTE�P���QlIOhu �;���"H,���CAYr�C<.���hʱ�GX�ۋ�%������c,^� &��8M�I�}����3b5��xʍ"ޢW�0�p0����:q�<2��tyLB�u��xh�0���e�q�HU���W��Mmė�Z�YM�,~�|��+��慡��,V���΄6	���O��c�EA����S���j�:���hM1�_
��C�U�^�ܙ�@CN�@������c���M���t�NQ�C9���2�A_t�?�;���C�֫WzAc�U��e���5�7����`i��-8?�Y��
 ��a�r����Oxf��ϛ��[Ԙ	��y��/�-˺�,m�J��-P�'
���}�*Z�d�J#b��f�F�9�F\�ĕAÕI<,�#R�na�(��� �7����8W%0=|#�����o	�h�Ϥ=63cJ�#�]�y��%��-���@���%h�V���TO2�w~7�S��f�����'9��%���):��~Fj�6�T(�[��:<J"�ɡ�@�2��_z�(�eF���Ұ�� �?��Wb'�:j��P������h�;3��*̘{\�[5�$Y���4j\.z�U�`�`c3'C��E���t�zX�_�W2�Zb~��-d@R�V�I�횚=���1�����?t��DX�n�U{`��l�kh �E�S�+��*|���g���X��&�<%�"H�9������[ut��Zoſ~"~g��`�\1�;re�߮�>�"�[��-���NC-r����^
�(D�������m�嶅y���֮�����$�7����g�up��#���a��jNZ<?�L���*侖v`�9�'	����(f�~�I���$I���)d�Ԭ��K���������P�)�# ��3�箝���
7Q���t�4~5Q��QV�R ��0�^�t�K�dI���1m�bf[���u�ՖC�ÙE	��%�~��a+=}}qKL�ފ�И�'���J}E���60m�P$�>`T�8-Z���.���2,��57Ҵ&#f�������3?��1k�42�����(V$b��w�djs�x�3���Bn��'\�-s{EζO����X+�� j���ҦFU�M��?-/boɎ�'�o�Ǘ���0*�R��[�>��w�?�=��kzΗ����4��)deu-�W}_ G�kO��Bv{�y3eIׯ���m���.É�iG0�*v�ํJ�Q�q����5XҲ82���&b�6�`Y���	6<��$��J�\9�/cr*��v����1�j��ſ�{1T��/1"�5 �;�bf+	/*?1/Ã#���uU�@O��e�	A��2�p�g�~}�̊���FBϨ����{=����FԃFM��l
V��7'�S�k����,��-�"$ȔW;6���ņ���D�N�!�V��Ńx��W�B���l���o,�ü��
�Súum�x��k�Ꭶ�������T|���Fb��
�J;2��5]<0$�2;�;0uۺ�ٝv��w�g]N���m�W���]x������*I��h-ug�su�
�E�5��x���e��L��Şp��ӕ�����a%~�2���p��J&ɳ���핥{%�G�'�Kp(E[J�.txDfdBZe ��)�rl���f��4CF��7k?	��b&dU��O�j��O�6��C�D|�g(���O2q����(�>����qhB��F �-i A��aGf�x��WY�[
3��e�B����je~��6$^�k!5�8K;Q��o�il�^�:�Y�8�#!�l �ع+��6�8��$�ɟe��p[�{� c�UOwnBƨ�G���M~�$�Y6{~j��O�d��q�v�4��A��Z1ZY[��8k�~H���i���v��q�b�B�".�h���E��Ϊ�U+��o�0���'� ���,�ɗX��֖�\<?��:Ӕ\���$I=��j܋V��y�'�H�ƿ��sN�3��H(�Xy��hni��8�����إrz�\(ӱ�'��O�9��Z&�=�1�ő�y#y���}�!+�&�:	�
�}��e]�/�Ft���ym�O+4������X�/9+�d�[zYNq}�w�S�U�5v��nfLIŷ�r퍪"4� ��_��Ec����eW�,q&ç�zl��.r�l^��w�JiŜ$��u��_{�ȃ�;S?�*Mh:�v����[��h��[�"��$Tu%�ɰ�:]c@\w�o�xPW8O iI�������2�B�̫ë�;Y�x�Z�B3��<��^^{*�Z�)�#�?{��S�8��.�{q���娍5W���!ߤ:�DsH�	�fo�c\����M�ߣ�E�6&�x��-�D�&�˝~˟�V,��}'��#��Κ�#�Ɣ%�=ab��ɻ�ݤ���E�����d�X�!bk���=�^�,���N=z��a�Ѽ�R&Mx��j�5��X�1Ⱦ�s#���
�r��A�ŏ3���B�˪Q�8���R�����<�����ͶC��B'�
u!��̎>b���N �$���E�Ց8M'���"�Ȥ����U�L	F��FN�P`�v��e��%x�%�����330;C]���&=�*�o��.��a��8!�t՚e�����5l��� �Q���{���z����������E2fnb��������b <�]��r�!$s=��AYR����h�3Qm���D�5K۳�;a�[���]̦,��� ��;k?�L�r�$�V��y�p�rbM�x�-�4sYz:�#K�q�$�D�����9�~q��r]͇j�I�0$��M�Qj�>����KR0���Ƒ>��H��.��D�����HԤ!;�:l7X�ɝk��`Zy�r�r4`�?�ڄ�c��D��G澯��Y�A� J���-�׹!"N}8��5�Q�6Ř"}|A��R�h�Lv���6�о@9�a��{��}U�Ѹi���|��-�%3��:�5���-��Sl���h2�G:7��e�vg,��PxLF��R<>л��޵L �� �.�x��j(����`��FzM�.� 2��+�?hx���s5��-��X���-�Ǫ��T��y`_)���{#�i����K�>�K�)]�7Ա�]�J��'��y8˴~"�}p�����S�k?z�$r��P�܆s����m��]�ϕLsM�^�(2��}�䊑+�s�:�N���%���ja��8�ͮ�Z���Āw�m������p�n�8�s"<���#�a ��l�XI���v|D�/*f��Pk�$��y(��T:�Ȫ`#���m��e�wܰ���o�9���|�#��h|���/�,�;�C��:w��R�#ik#H���q��_����~�ޚ��U(������Rs"�V��=Q)"B��l�e����1;�$r�{+#=��z���vۮ�I�{����T=�P�5*��O�  �/{��-�m���s�����x(o�|3t7b�	�������?TԴD�� �CS �j΋v�g��;ہ�]��=��<��?T��1�DB�FM�����m�B�aX�k�-��p6����JY��S���x3����?PL_����4`D�������{�'���}�n`SFX=�5�-�����3/�&�`����"�Σ��;$��$;����:;1X���_�&3�̻�