��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$�ʩ&6� t%F�����)Ǭ_B,����Lwj�e"s�^�Qq��kډ��X�e4��h'��_N.4��V�5�!���c�y��Ӭ���X���V�t��������0��m�CZ����F+������.�̾�Z��fW-~�-�G�OK������=9pj@�A�ni���+0`��C2E���)��n�/�������-V�NX@��~ņ�3�vl��W�g�Pz�&��t�V�"9N�R��ᗊy}o��!����__��`D��=��H�҈��>�,�g=ﲓ�Ĕ^,�t���D|	Qe���|/�P�؋J��GbO�}�1l�S)����v�(����"�)Mi���0���Ƭ
�D)&|�vǥG����ۄ{k�ɣ�I��������M�V���;�kߗxN��t��?�b�3�{?O\{�f�b��f�Eأ�P{C��2�ܸ [�x} ����1� ��O�}#�P�>h�=�A��g��l����7 ���b[�)���gG��I1&R��-d�m����-��B���[|^��.N��Ǭ-ʈT��TB�t�u���M��^)�0�ۛ��U�A���j��T����XSw��,b����ӏ}gE��Oʠ�������C�������<ٶ�JpeR�29*8���T"���<�K����T��oh�Փ���e�E�NS�'˿N94�ڽ�,T�t�p�[� 7/�h�m��!�q���~	����5�`
�3T�+80�(�G�c�B�a�Lu\�̹��k�-@A�9����>��6S�Ֆw��C����m�ɏ��]m�{�Ƕ��K����4�v����j�V�O�����M�o_qP�*�2���~�<�h2���i8�f�t#$5R����;$1-�uuD2Gf�W���-l�Bac�>�sh8��釱١���Q�����:7E��0^u??_(�,�7��wtz�Vػ(�j�-��-�e��-��S*�W9�uC��l��ŭU�ߒO��'�ф��n]�T��:��k,>�*�������a���>����|��j��W=���-�r�z)~6��eL�꬘a�E�ʩ��˝+)���;^�l[��T?��z���x�Uɟ��7�*�gz��rt�K}���lfE�N�eE=�2Pq���5b��3�/����a����Ax�%��u�	=�l+g�p�w��G۔�V���|��}G|�}Q��W��n��6o<��O��f&4Pw�����O�V�yqH�U�[+<y����Lvf
�y3����������;����i��|���eX�}'`^������@�GNs�&V����.}9�/|ui4g8!g?2mz�@��J�C�ANL�b��otjZ�xn�B^%R`z���0��s{un��7�h��uf7è��L�q�)�O�0�0z��:�M�/Ð �=��6 D4dof4|����8q�d~/ԓ�4��;���TC3��?��`���1C~qK����!2J�T}�U6^X{��C���J�Sqp�\�]���G��~r��;��!jq�Y�K딞��!Fa����p!")i��/�G�2��(/���qt|J[o�w8ʐ{?��+@`��f�]V��bxƎ�t����KsF�OQʮꃬ��b���<�cuT��~kj���@烑�^ۗ�Ås�vω��U�0��򊎍z�=7�,����)WW)�[� 4��p&R����i^�s�{�js�^X��X�gSA�O��M���$�(N�s��(�/���x w)z�V梣G?<��-�SH�4A�%��I\`��bn�����񫬜0ce�v ��$��K�`��n���H�p��f�� ��5`^Qy�Zy�S<�ZqD�;b��o�̧[	V�7 ��%2�F��CT���\�?�9-
�g2i��|�J9b���]��������?�t�HK���h��h.-�����k�>���������%9����o@ϼ��S7�%�WA�w&���1���_q�袉;�A`O��j�UW��n�q3���pN��N�t{��,�EZ�LT��I�eV�6�N��!�P.�x�R$�����*}��l�Y��׍����}"f&�פ����u%0֬�!s�`���L}�6���4�g�N2w�
���<��b��H��� ��i�!��3�x2/t�.���Q���� '�4�6y�E���Წ,�!\������7D�eD�Ҕ���͔K�,j�����ɡ?�l0�>TFl;ȚT�����_�aK������D�㴂���/;�js�b�D�J��9���!��Ə`�>{I͓��L����P�-����Ƞf�3��\��Nk�S,3iҟ)#�x��|��i�&܋����W�D:�c��	(P������Z���_ME�o�� ��!��ऊC���H�-#�*����
麡�7��$yf�	{�w�5� '����$
*�I��{ax�>���CSmϔ��	�}�<q�a���u��TK=ܹ�f��ю�z��ק��:_������ʊ$�cܦ���A�-Y��D)�^�Iȷ��;Ŝ�q�#	��H���ax�tv@�*-�j�S���|�ʌ�ҧ��rf�C���|`��6�q�)��Z�k��u#�;ZE�
9��L����s6{>@����Z�ݙ�I�� ���3���ҘO��+�I#�ռ�}Q��/%�e��hMr�n1 lu��_z�s����9� ^��c�&�`��;�e\��(�S˼�U�2[B�q�k.
�8��O�U�²������2B����8|��B����e�`�y��t�]��[�0;1�`�� ��>л��'��HrV��()
�zk��6'��N���f{�7D�{()���.�5�ƪ1�J�b4���#��b`
��L5 ��UP�"���'S� ��B%g3�f5k�(�*��%����i6�YZaC���v´Gr�=7$�ɘxn�)c� �G���9����D�ҾK᐀��Nڎ~g��N
dtA��n$8D���ix���\d�������P���K6���2��ͼ�<F�yp��v�����n���s.���m{�ƽR5-Q⧑c�XR)��A���[2(��cCͯ�-�
J��45J��R�gF�̀��#`���^p��؎�sAK��O�!9F�����t&w"i����$�̶��6�1I�(;����يݮO������y/\1�X��)��BS����$Af�>3I�"���C,��g�V��*���v�;�bz{f>�?ԑ��bK�S�j��c@׵�T٭l�9�L�#�����.��-��&�L�p7S�2��m���K�,����49��83��2�W�Ӣ\���9��3�L	�])�*wՒ�W�t�nȉB�m���0��S6Ûm1�$|(e���y����߆�#�YkA`�Y���-��gÈa�D]��L� �̚*���8�frP1ᡩ����>�ۤ��C|��ח�!�1�_�w�`�g��	S������\��Ĳ'���*ۇ��w�Bq|�9$8A	����t�Ơ�$���9?���gK����,ӚAUJ4FX
d�u�ͤ`�w�?{W{o�0��!��tGT�D
���s�L�0�%��+:���$�ݖ:�R��\��.��o>ߌbgֲ�j�R%wP9����W�m�!�,���F�x�ֵJ1;Iy� J�>��$n�2=�EGy����[��l�v{��ʻ�
��o�*�F
D�t4��"��3�x�6����٪Y���-U:�6��K1֐3F]a��TZ��l��¯.G+��t�P)0͝���b �u�i3�{�������}�r����.a�������lK������P��dq.�0�6L��k���k��d�'@}�� ��T�����FԛwX�F��Uw�ݱ~��jG�h����2W$�a�a��+f�?��'n�}������b5����؜�_/�|<��Ǯ��ǫ��+|�����3{�ż�1��j��K"��hWy���h:��lⅡ�����ٴ"��9�N��,�.�S�k�26�uB�[ڲ�O�tC�b���4�V�"���4��5��A���d
�2�y�˒��g~c^r#/�A^�B��Ҽ�"P�>��	�%��N<-]��p;V�B~y&�o3�9�}L�Pal���-��m�$������{����6��b��S#��ԑb�j=������}�:���iI�0L�Qi�	x��p�Sο�k���i��}R+���.�!6���x�r��_~i��T}���>�=�?:��r����
�6=-Ѹp}��rd��fN��:�Dd���"f��#%�sQyj��G�]3��Q�b��~?�a��Ԍﭫ��M�ӳ
&K�I$�r�<J��r���ޣ�|� ?���߿殦|�� =ȵ�r乼b�ޗR#s�OƜ-��xi0��ii��2Y]�]&�-�f��6�pO�[u�ۚ�y.Y��Q"�ʤ�h_��vK+�ߺ4�0������{�V2Os�s���$��6�`�.���`4����O������*���_��G�e�t�$w�S�F�\gK�.�ǺTy��䑗�.�3kTo�-v��,��Fz�o�u���05o b�msy D畞�<�7a�������Yx�9L����6>��'Y �y.���;�W�s�
w^�D�3%C��(��nZ��3�����П�a��딉�� ��h%H�z'qF���G�'�y�˨OOH0]�GX[Xn��H�c�-L$|k^2�=n�e��|��K������N���ܪ�o�`��`�3����٫�Z�6 ��I���Շ�wIݐ�5����EXlXz�Ε����T&�k/�^��r0�����q]�3�l1-|Cc,7�De`���!9��-Ď]4}��)@W��k���1Up��\)�'��8�e����X����Hq���1SL�Ȣ~��02-)�����JA�ڲ�oli4��[%6�����8�Ui��p�wh�۲�X��+ж��z�B��v��nY����Yɔu��u޾�L�9F�ք��_/v,�P�m�i
"�V���˺��.�'�O�����$�݉$V���EVt�I�)�����q$����s0�{���6u�vb�1����!�\,Kq$
�G�3)���p�7^]�����rM��붾鉾c1:��^��(��͈����(�:���˷MH��PFuL�'鳊�!��4�ϛ���D���k�ܿ�P?Q��.�-9T�f7L�ײ�!.*	�$C!�B�>)5��u3�?�@ �d�X���Sl���]U�ZN.��t{e/���u��j��פsej��2lśG�5�r�ػR�E�AL��x�j%�<My� cT��Hm�=0u|�9�ԇX�HឪE`������P��M�X��:G<�)����&�b�	�oR�snn��|~�"+��%�Ŭ�=F_�I[m���îĭ��W9u�i%X�O���y\:)��z���xmm��(~?}i)^\G�X������m�)��i|Zn�o��L]�.j.����ؚ�"~Ӝ,	8�N%8�����F~���a�������[�kS�ԙ�Țu[�(/�����a��6�T2�(&�Ib�p:��H�`~  �۴�=C� âU���}.b�otX`���@�I(M�J��a,�;�%K��7�T�"���x3O�Y]�ዑ-_�.Og��	[	���WF|\���{���R��̀�i���db�v|�9&ڜ��i��3�m"���`�#��U+u3G�Gq��F�
a�nw�	_!|{>=�3�7K���CY�7�z񋃿��8���֢���]<A�F���F���6\,��,]�g�X���%�"?��X����e���	o�ډ��Ŷ����̛LC�{������k�r�k�r���=xG>�D��������r;�C7���b�`�+�E]��\�_���A�H���Tlѹ`��k|�P~%z\�)Z��5���K��rś�M03c�xF�gS�'��o-�N��Mes�.���l���a�u��_� IX�f�{��iE	O�0UQ�B:��5Q�po��3,U���po���I>]�V��'���"4xMu��i��T��^SKC
�3d�@���ɬ����������L\�#NT0"�Ɇ<�A��a��ɦU��"��0��19 u|��df�
��b�����Muc�7k��\���FX����]���; ~ ��rȪ��P���nw�u�+?�?����#��J�'ny�	�����q��$Ii|��6���3ހ�j�	0�� �V�N����|Zb�Nr�ܒG<ya�6`���̪Uny�K��dؒe77���d����;n0��K��#�Px�zYw�"E�ͽ�Ħ�ﾜyz���G���OH�}{��
�j�l"QG��g׮�ʱ���^���D��n��Eo�>}סíX���i���\���f��sMP��k��"���7�v�hB��F��������lwJ<�D�bS���h~N�:��4+,ps&��~r��r>Z���Y�=�)��f�Ann�RD�"(Ǡ���7DM�HD�(���9H0gVr�R�n�I
�^�� 3���s����F�ϖ�8��ّy�	G�,6�-'�h�@pE;�8
qt%%Uiz?
��-2�$��+(���WW�?���A��pmJ��A���+�%C�j���x	��^az;�-�OOt���ڸ��J�[��Gw$���u��0e�p��?Ə<�1�?�^9]4�o쒕�㹴!�1�I9�C�k�aE�(z��Zcu���1R�!R;︍����f�]/���1��ڂn��6fٟ�p�Џ�&4��Ӳ��c�u�����:���r�����t��]_"?�� Z^b������)�.�ϵ,@���dt��SW:T�F�c%�*�h��$��������\���,��h�d㺁�J_�NF����_������2Y/m.�Z���Of���"�Hl*����pЧ�4N�{��h���胐���R�P$��o��Kr�b��ӫz�h=��7viK��L�k����;D>ߜ|���Ғ��Ĵ��mG�`�d�:�0�����}��]��`6SB�P���7 ��4�|�FwX�NV��F�,���U5I%�~O?w�aRj��햨��	�N�\��ɝ	�CVi����WC��a8),87ɑOU���1�0ҍ�����m��l�d�M�~�ɠF>��s�.�Y(r�zO�����]�mE�Oi�?�"����Ez�Y=��tx��ӃjR�����f�����F���M���<*��6^wa������g�i��O,��t_�R�'�듈�?��
O�)e�i���F;`��Ҿ6-)��y�hz������v�Ř�Z��U�L3�ک��)��[v>�%�Jz��Sm���J�}�z
Jt�@������ ~�7�d�5T%\0�M�Y��PJh�l�����@��'#��#Pg-�('��.��["��8��5�}�������^3��5��㈟B/�L*f�k�\�6rM<�k���e��rf(�0��P��E��<!g���EQ͉�P��o�;c��=�;x �t�`�Ǘ�,S*�����~$���/A�r
���#)�������	ϝ�Y%x�'���h�	��A�Fr�E`�ɑ��56#�8@4<��&�Q��@�t�Z��f���W�}p�9���"
���U�>T~�%о�t�%����pk�d\SQ�ǩ�K8aޏ����Ћ��Y3v��)9c�^���F�7O&��	��7ɭ�f^�ׂue����6��9��5�ZA���XP��itUר1&���"t4Y��[�q��=pF�@�Y�D{�+���XX�#~�U��>��@fi
�fxcn%R|�|w�K� Ǳ1�Dg$N���_1uǇ40��A>��ZX��+���LG�{vTEW4��L����x�G�W�{S�\��2נ�/w�zyf])��l�'������a�'tf-,���2��""�Y5��m3������b3fl����B]����I�d���L���ŌL � �"���t���%�ȥf5�a���L�"�i:�J\<ۖ��4F�2�a�aj�L�� ���o��+ c��U�s���\V�fL�2ƹ�����E���*�]WM���}	F�H�r�ڋ2�5���F� V���:�m�f���V�ljay�G���~ l7HKmURfR��-`�TP�Et��s��`3�;�/{b����U_�n�w�Fk��۶���G �NOag$XRL���8?Q4숔�b	=����SAYe"`�;%���N7S=�A3�l������~���Q��t��V�V�g[����8�3�][�+�
xEj��.d�+����3��w����H �[�f���yY��9s�E� �-5��5�*��B��gئF�I�ƚ�*s_�Mu�����cZ�M�j��N8�:QQ�;]p)�:�L(ev�Q�N�G6D��-\-h�ӯU���
�z!!J$iZa�4��pFq��M6��sX ^�`
��%���=>ʔp��Lw���N���T�����^4kA���B�x���贅Nye4"�F��my)<����\��_ͪg� �l���E"I��F��?t��V��T�JR�?Ri�5�A�Vq�'&sI����_H����>6���s-�ARlK��*�����h���;��3%��%mϞ�6�)l�K�n�ߑ�̩�n�wP%k�g�T! ��J��@N�޲���T�Z@����%�ŝz@�ȳK�u�;R✖�q�p�o�5X���)��ʷ>�����|
9w�7)���a~�Jv��ND�T�s��5潰��T!�&u
��'o%R��.q7�?�s�c���_Wj���$[�7j�`W{'��C�S�FK�g��{u��V���v��
\��}��O��"�t����pZ��e!�si��;4���@���A��}����F�M$U|�b a��ۏ�����W��k��"��Er$еM��?G��r�k�n��b0�>�ܡO�^�6�~�����\g�%E����$�wR˒|�|uD���ױ(L(�18��g5{i��4�H�J�j��swkj�\ª�ѧxSn�"A���݅�Q�F�~�s<���
�'�e� 3��@�$2��b��9�`� 6	սLy��q�����t?�L��ǑS�oZ*���h@+�cH�DSm�bq��A�CQ�l��iZ?t�S��V�]�qT���EiȐC���'2{����ndP��w����+2���LJ@7�4�x�2�vR���=�HS�J�v�*��JN(x�]�Ѓj�ebڱ\1|��#��y'�D��۝�8¸�&41#����;�, %͔�!��k�%��ݡTfl�!���6�{�h�l	��(��^+����ݡS�Z�ӡ��k	�����wؕ��鑨&0��%�o��|��#�yH=؍y&(�e^P,�娟i&C:��T���'����7nE]�*T�Y��WF��|1?��F�L�3iǒ�-T`2]��I�X��
Կ�_f�vY��H�a����K%�u,U�G��G<x�I4�g9�����sݦ���0^�X�e�Pٸ}��t�$�������F�\?u�{៓���-�M_ш�6(�-���b
��T^��
L�fu)��_YN��K�$.��M�/�2�b�}�/>ײ�q���w�b�*�I�n"�o�������M�ID�r橙��+'���P�j=��=q�s�u��L^+�v �:~x&[�/�(t8���y�G�#�y�aڣ�}HǛXL歨�MTv�M�@D��2i��Ce�W�m��|�6����&�b�W�ەZE#I���MK��ʄM�ď��l5#�f .&qf���$���\������u +Z�Ֆx��r�H$�>��q�n����4�8�p�̀p�o9�H%g��T�����Eϗ�8�\�[���w�Fm������T[0}0�rn^ˆ.{#��
f`v�&N
{{�Y� ���.���_�}�[hS��r��ؾ�
p=�d�юZ��%E	�"<�G��!�2Cjh�9z+\{���j���c �0�4 $���l6�)��-Ds��#3W����4}�=k���oఒ�qY�;�r��Y�4�	��z�s~�
�&��U��,�K�D3�Uj�٘��ˋ5�9O��$.U���a;ã���`�8�0�:<S�Q���x�3����- �}�Q��{;���`�\5��Q�`[0�����*��rc'@;�E���IJ�q�-���amEt�gvf�l��FHv�G�=��@L��b�㣲���OQ�)��EñHf���+��;�Q��X�ɓ�y���wG$��:b�� <��=o�p���1^q1� qo@3�[T
�Bd׸��M!��xG���^�"��?��z���a����gde�v�v��l��@^}l�>�H�2F���u� �w%�NL�N�����-�PT�D�|u�%�|b>�:s:D-���O��7��;�l���G3�W�0�)zp��
����7�/��:�,��{"�)n ��i��!�����Xǅ���z������ �tnSo�,=|���<а��.:�7x��5��3�%�HY�Y�65,���SBfh'N_���"?o��ْ.:I���F��kW��((Bs"��'���d��2���NP^	w��o�EӖ�B������� ���M�rС�uY�����8y1��S![��$������ۀ^�X#�t�~���\��MF{L����u?���b�����Z���1�pE��C<r��W�C8��^���8�����㐯�Z���A2�zl�B� �g}�)CW~�G}�9f�ru���_�'<H}mw �b�CmXEJ,W
�������4�r�"�?nW����N�'��vc�a���OaG3ѵ��~�r�M,�J��A���0�x:��LFA�V�O J�C�;���.��,#���V���ً��7i��. P�y�~R�*=�w7&.��	����0�3W5�$4��DЁ���te�~_uv�a'�|�)n="�SH�cP�|�~a�!_��X,����D�F9ǟ��~,b]po9�S/a2�D�+��+!g�q�p��Y}������������~ݤ��sn��'�?��&��Q�&���K�n%�[��Ii�rgMߛ��c� ���9�7���ꣂ+�EtVb���ơ�pb�Q����](G�zк�X��O�Fs"��=@��=x��"�,���7.�x3��[���2�o��:%44(SN0bCAȕ�v����{h-��=���)��h	�LL���V08���A ��3�!f��@*=����C�G�����ຖ�o��X�xI�U8038 G���.������Җ���.XOB 䧬�ؾw8a�B����f*���/r��}9y��k٨ȥ-#�G��S�4���,}B�����Gqpy9�Nᇳ����NR�r3P�n>O�b��Ϯ��g��*�	�V�B������NF�x�8+b�~fM�n�c��i̪�_9�۟���*�-[���YJ�T�:*6p��}�//�g�3�8�&����D�����F;�'�� �f1�;i�$�}�6�*L	yw�>=.�8 iQ�8��<�I��d-y��>��`�W� 3�@3���)"�CϘ��?	X�-�X��D,�[$�y�nr�Bq�WV���7��B|����/�3��(,O)?=8�N)��!�n�\V_,�xM�*�P���h�? ���ʹm6���u�ƣ�h���j�K��c���ɣ�XQ�9jˎˑ��uV�������c+�mF��I����V�Jl�*3*m@2S��D���p;v��YMHO�;��{�.U��#m�t��U:�B�e�_�lP3v:�4E�ZP[!ߩJZA���(��0-���ƻ�ق�^V�����������lG�a0�jѢWKr�Y%��l��"��Z����0"3a�A����]��i�տ��� D�z����5���340����v$ROM�>�oW;�����H��G&̯����L6�/Ac�(}�|MM���02ق"�?#���hE����,���oUR3?'(���MK�����J3I�!eP\D�wq���G��ʃO[�z9��e"�o�w��\Q�B�CMV�nR\[ӻ��':lC����k�A�:Ies�C�E�+�f�^
M�S�\qם3���x��i�1�ũUb�6�^�6�&�O��7����S�	B	����ل��R3\X��oe[з�v\���*X�/�X�����,	��=��?��sk˼��c)��%�^���d%h���E�&��]A2R��9��o{�1�g1A�G��!�GBn眂���h�����/h)�`�T�D�2���r��勦��ą'V�a���~.c�� ��~��cJ�����Y�����s�^�;�=N��AF,��0/�{��#[7?�v���\�rO�b��<��)�axD��#�>�d��wۯ�̪����9���r��{B����񞟀��,�;j���DB�}3Ҹ�n�uq�T��� KM�6�=)!���=e�6TӸ!�{3j[d,_�n�6�f	#�$�I/��09J�ӦM�2�R葿���8���!�Z��Y��c�7���_<�L\*Q��w���[�B9�|b��q �}R�J��}�+�̂�LՅ1ݾ(&GI��.���ݫ�hK�����d��Ճ��%!��
5����?�]Lݘ��M6jl]xy ZnE��W�ˀ�)=�7'E��u�hD�t���%�!��D�6 �$r��G�cd�K}��@�4Ɇ�� �GD� ��k�c�g#�B_�!�}
�b���?��Ͱ���΂K�[��M������5UcL䛆2u]rc�*� �d�f֐ �+ݤ�qp���5�WpE8�M����Vy�-;F{�g���j�}ߓ�.�Ũ�����kގ9���g�:C'�(���o��ϝy/���ѷ�v��>B�x���#e:�����+��ǟ�B�4P�р��6�F�P�]���+�����B�p>wT��F7m7��v^an:�2�ߓ?����|�����]N+U&�So�Tt���T�	���I�5��sZ/��&`�-FW�ȫ�@���}ɤ�O�:���A�����&��U��� Ϩ� ���S��m��~��9!�1C���;cޝ�dLNZ|�l��5�%uoB�^�D⭇�H��AJ��؄�p�|���V���h���x����͸�s[^����Rb0f���C�Z�;��2�/Q�B��;��;�n{=��P�S�/��j�aw��r��b���P�~cO���^�Y�ͫ�`��<��N����EҬS�`A���]E��7.U�
F��2 ��֒��ֺ��z:���d�sB�-6C��(�,�8`����]� 7����:�N�e�"h�B�d4i�^��Ȟ3H��C�M%&aV�O��0�ɮ�-�\O�?r�y���l|����'��R��Ⱔ���j���_-��6며��5�8Z{�L��=����)3(
����~ �7��g�p�=� ��2�ٌm3�GEXo�*B�5������M:�lq�lΰ9�E�A��*ɡ�V
D��h/�f�`hH��R���7I�ˮ��Etc���s��ǚ����h��PDU%~�=��{p������B���ZZ��T�Mnŉ�^lү(/I	���Y;�u)�����42X?dw�ݸd �"�/�(�W6#"�����K����� C���	�̉����[�G��\<�e�18S����0���0=��B�<'���7F!�%��j�v����D�ݗ~ó�@�q#�I/��l�M���P�U�rwD9�AC�"�G������K��3�ԕGڔ���.�� ���Ѓ�h޹PrkIKb�H��*ψ�q/q�i�f�@����S.^��r�����Q���>>�ۦp+k�vga�q*;iU�5�=P+)	;h@��#��`����ٗ]�*,�JI_�@1@]��-��6���c��p��?���n�k���@��1��>9�f!���n�c�m��)�Db�x�!�=?��ZP����^(�q��A�t�6�R=�SG�;�Ԃ_��b�V�u����="�KvQ��؜�r�F��F].v�en���Y'��������W�E�B��A1�F�(���Xc�+IERu��Z����}���S�t@}R����t�5�m���ޡu?:�P*8�kb�n%l���+�Zt�V���am��_��R�:��4o�n/L�\4��[��Ȣ�ٽ�%��%Z�A*��{�\8�4�� @�8��!Roj���%��q�E^Q�0��ۙ�c�i)O'��WRU˲#���^�-�ic��m��x���ud��\�E��Ч	����J��K��:́3xmC��2�\XI��r��O��7N�� ��m�sl�(�k��
q:�`~��u��6c"�틯N���B�یzCp�#�1TCK�:l�4� !뛹5�]������}"�`�4�cf�)1�V$��r+VT4Y�6&�� ��V
*l�L��WoB��ݽS�
�.h�K�m<QU�[\��=�5�4��9@�Bd����F˚��n�^n��V���	4��+��HmO��2��G�Ev�Z�9�/gLy֦%�?���$�wx�o�zT@8 
Hhg.�^}}��n+O��{�����}(�f����Q%ɔ㼋|l��y`���١n@��x��*�վ3���L�FKd�i��<�?��48t�AǷ�2D4��_;�jz|9�f���t���֦Z�����Ͼ,8g:nfl�x�3�|��.a;�X���`~T�'�_��&���B큄���x�z�����v<5V-��	3>RL��p��g�${�ڄ�i}T�5�/S�>����f�@��J �g��&"</�oY j���Ԁ�GF�$�;�v�  s�//�-X`~��J	~
"=���������"��jGh�^�X0�����Τ}~4M?,�s��XFH���xp�#�%)�C�p+]5���uG*�k9�¥�W)s�V�A� '$9Rk�_�2��w,��������^�{��F�����w��&�p6�G�䓈b�>PZIF�~�e���ܻ��?&�σW����2m����O��{�T�T�����h��s���VZ��-)$���):V�"��ל:��8}/8O�B�u\y�1 �ЈP�Yi�>���zmt��y�Zo4����J�d��2�y+a��x����`����(z����O����&�H0�&/����*�?謾�j]��7��Φ��$�"�d8�H�t��Yލ�}Υ����߀��~�C,^�iB��Td:�̽-h.�h��r��9ɣ]�����GBf\���v�U��Z�u^� aU�vo�je�F�a���w�b��s��~6o`뛜�)ƀ�Ϭ��e�3T6l|X6=�J�.�V��7��C�	\�8ۢg
\���)�H-8�*����5�3dA�4տ����p�Y�V�gN^�T��N�Ȼ�eu炖$�Tp^�_�e�]��2��SYߨ�z��	`a�ڼ7�ی����$��uG9w�BF �s-��n��DS�vm���y��V�3�m������~��k�H���>ޜu����̊����Z���*�~t����n+��]?�$$a���.�"������ަ����S��æQ���ʴ{��Tn��h䓥ͳ�>sPg�z[�D98�yp�����L`<��G�3�볢s����<d�l��6�?x���I�	z%6����]��F�)�>��ԙ��l8��^�L��z�QEf��i����F"-���&$)qF���LVg� 	�\)��-d���a�I�Ey�yJ���-��1����Q>&ȡk�Fi!$ˠ���PZ%v#��X����i��V�,Rџdܶ ��Ѝw TgB]"�gbf�H�_/�:L�� � ���4�x�-Y��h14+��]]�dz^��l�v�%�\�Zt
��z�{EW���Lh�&\�+�����Wb/��C��P�<<��N�.߳n��Y��DP�y̠��(�������*�������LG���&O�*`O�N����+�P���Wh\�n�I뒡���Y���TM���NE#����(I�����vC�(�C��)fĚ���Z܆v�f����q
`J��aiOQ��t�Nc���1X�a�������*b�U�[x=�Gsk!��*���$d���ݞ�ժ;�I�ь�����+�ij�.̱L�.H��!�9���.ڗ�\�G��+dM�6�c�%g��ϖ��#�
�~z�WP��l y�r�aN���,u��A��l���w��p�t�A.6��:���,2��
�<U��a����{�"Ţ�
EZ�o�f����!��+�H�r��y�3	�m:-y��064Q"W��։��)�9�u+�I�Ϻl_x�ξ5ü���m� p��8@֏of���2]�np����gM�����\6���Z�	'e+`�[0��	ux����s�d`"���$�P^�[��$��ز�Y�kPܫ2qt��Ϝ��>N҇Y�m�{�#�l�ͻ��E��x�xSn�������x���^�Э���!�Zֳ�
��	2Z� hhyĽ�_Ȍ�d���J0j�w�5J���f�Q��嚳5��&�
{tq<����Y����г��@Kn���	L�PO{�G����m:��?��\���;_J;C�w��ٮm�=�ڨ���j��VG �N���j�g���Б=P��&Yu��̚�zINW�J6X�����vA��^;2�����Ve����ړ�`C�c�f�]���3ARPfIj�뿇�:"��p��J)dod\�ك�r�Ͻ:�.��~Od��{�>e�[�(i�-}[_�Eu�U�'��th���h���O7�s�����9*���Zy���x��1�xP�8�n��+� 7��p��l5���Ãr'|[h�M����Eg}��5���<��Jv�>� "M�?���4@�}���iĺE�=��D�Z��jڪ�/�n��c���S��i Օ�����Ch�z�� 0���]
�W�'�(�ˋl�.G�k�%H��P����ӗ.c��=A I��?2��]�)y����Q�J)?
��E��㚴?m���4��E� a���
�?�f��Ǯ�6��`'���(���Y�:��;�y5�)!n���Q�h��p��:�:S\��-���D0v��c@:�1ϷJC�3�-7_\j2 �8���M�Bye�ә+t�/o(E�k��m�Y�|d�2F��'�ծG��bO?kʄ����1���4��Y���9\�d�ݐɎ
���#{�},j\V@����(_�12�~�0;�O�@Da� /�ơ@� �.��#߸�?�1S��2M�ni;�j�і�	��n8��eh
��|�}Je_��#�1]n�WO����ܳz�]��PZ�\t���f�J�_i��wNQC k��*!���N���9������v!��|�;GD�����ϊ4~5iٴM�B�rΊ��es�9X�4�®�W���m4k��'�Z��=��[٭�}#���ڨ�V��MP�|2�����}^�i,Y���z-�5�ޡns����k�Ǳ|���2Y� �C���~2�fڣ^�W\���#�\G��jMj�V��w�Ǝ P��v���P"^��=�~DC 	1��;��q[�F䵳�W8���VנV����Xy9���~_�a�0��Oܺ��NP�޴�N�݅Г�K�������ySb[��Ad����=X��Ӎ	�K`��-���zz�!Z��P�`��,p�w�����>d��M0A�K��#�)z���ZH�Im�!�R�P�m��-Y����L�����d�ڣL����|��*��s�`$�h�W�7�rQV�:�O�y��D@neq$݀�_������S����{�@7����GG�� �G�,^\_Q�:�q��+������#~����W	Q�S�7\�}q�% �0qڂO�P� 'jc�Z�@7�$�����C%)��1��(GupY���-r9��P����ٴb������f*��B*���Y.sE��}���z:���-5|zW�U<�~8Q{��	��gu9�=���� ��
n���H����pr)<)�ˤ�/<?��N�]l��qt@;9'?��<vw��S��]���s�u{t��F���Г��T����|��s+u=���]�]8|m��u=�z��W����Nf��r����d��J|q�5{Wsy�c�������L�0q�u�K����f.$�o0�Jp�|F�f��-`����Դ19Y�ױ�ߑB���*Ǔ;�<0�EݓY`����oY��0���xi�]3,mG[�j��q�c}0��F3`r�{�Ǳ��,ʀM>���W�B"�<���C�z�@Wt��ē_ؙ���e�[������O���G�qp�
�Κ�^c�V�85��A|��2��&0���(��Yizg�޴W'�yJE*a�%�������;����`_IR�K=1�9^��_� �Ϫ&T���� gQ/���N�n��@Ÿ{��-���x�yaeW=Y���@�<����1 >�Ɵױ���/������1�X�r�/�f�~Wފk���} �P*Ox2�
��z8��
`VV]���r�R�޷�6-�].��u+��C�S�1�w��v?[��c������|�Z���H��	i�"�˭����R}%��ea���߫��3!qQn�vE��� Z��wC�=��kk�6ɁsZ���#�ts��_1�>���Aԝ��܅�y�2Vhpr��?y���0i�sBx�ъ��� ����]��i��bd���S�㿵����g})D��$��r��K`m,I�uŚ'뛟p: o��͟|�>�(�������__�/x�Q��w��WuE���#�S�<	�_sTӺ��~5g�������wAJ�x�R�
��΢�E$�f�	/�՝o2b�QrG�(^����(0�	c�h��Λ���������t�� ��y�=ti:��'�4�"*�)+���.�>����],uK�	���IٛG΀PNi�_��G�>�U`'�+l�=5�I�0��.��g��7{3!��ї�E馺��p+E`1�ܱ@
�2t�{l�JV�{�W�~Wl�B�p��W��\fBI��H��<����ϒ {��e0j"�k%M�\}�δ��x���w�V���2�s]������es��wu^�9f�X�!*3jȤ��뒗�k���"+\�B$id�NB�P040�{"ڈtY���^����l��Z	���^�ϳ�~�x��ϪPbpygVK��dm'֢���I��'.����� #J�(��n�)��wx�#Ҁ��[�'21����9�~����h�6w�E�ν�V"c���u�S�ؙ�O�fČ?	�Ō�^J>�v4k�q��Nl<��7������Rw	=��	xj)���Di���g��y]E-f�W�a�ȼ��p�uI&O/g]�kl�������l��O�
BH$C/���BM�:�*ٟU�fy�6� �x^��-VW���\����QX`$]���hE?��6@�%E�I�=OZ��ap���Tv��z���m�� �?7�*l�C�@������$�i2�d3�C�x�O�M7�`�j�/�BJn%��������c�ܲʐ@Pk�R��녅1y8��Xc�����O4���^I/Ƙ�)��u�����xfJ��}26&��Yv�
�	$�X~�} y�_dXo�/�[M9"3����\5ǁԓ����j����7�$�"tN��D��7��Ub�UV��y��t�ێ���f�z���<g�8|�eJ���%
�P�,�cW�%��e�=}�sڴ�a�՟�E� �N���a#iB��%^.x�GjR˾%�Ѩ��y�0�>u�\Ǧ���$�KUU�ƻ���Ϸ��)�a��B�zԝ���rҳ�-9��R�O� 8��TE���� ԫ���~��
ӝB���P�;��p�&���`z�;��[JU9*ُD|�f�e5B�gT�a7�g ��R�����fd���8�� J�ǇN	�j�jQ ��#^�nW̠#�O[z��D�0�kz5k?��"W?�x����J?I�B���Z =:������$��t�B�L�[��v���h� W�@�Ȍñx`=��c���� }�G��j�՜geTV?+�1̴�L���|�wO3���$�6�ZmԼ�߆�}@�:K��+Su�D�I�1��1�N���g��C����]U }���z�dvaVk��Q�!E�[.�/5�u�e�Q�ACsSP��I�3�Te���;�a�K��Z@�&wm��!v|xO�>OR��j-3u�K�����Y"rl��O��L�+<ߴ x��'��S��x��%���8!��(��%��Y}���b"<)��d�:�%���[$_�c%X�����iu?vZ��z���+�Za�`A�+g0�Q�RH�6�ߦ�����uT%%���	T/V��D��-�/��U�M�:/v�i�Gv�������P�=��������:���K-�nN�A���H|�9�8��8�b��-�-9��8*S���6���2on�G��}U"�$��
��^��kRxe�S�xv
_�˝�/��o��.mp�	%�_��V����s*��٘tE�鷘3LР��f{�|_�Ҹ�����!�iR�[�0:�H�8I:��*#��TF�����sm�6�Lն}NH�I_i�(l�8��(by��B���0!?>T�uX�"�vRi�X�/ͭ��H�xf ���׀�o�l@��Usa*�x��t�o�Z�� � �������x �XJ������v1`g.��	�ev*�Z��f�^��|�(�_/y���j@��:e����T6�x�Z��f�jK20 7�� �p�5�G����3��$h�C�NHw$%0	�`�*�go>�$�������P� +�ɪ��!�2�n��PR����JQ �v[�3.K��P�<�	�%԰զ� oɑ��U0�
�)����Ee�
3)'V>���E+ۏc�s0�*�}NO@pl$t,<�����tt}�W�s��b�"�x��Y(%Z ���_��\�RI:�9ox�i^)���L�4�f!}��h�E��J/R�Qb�OGUXG��6bϑ�GP �$��&��r��L���ȅJ6����uCm��U��U�C�V��YЎ;�3oZQ���NԲ3;q��D&B�3r$�|!"lUB�O�B���b7��1jW7)�ȫE���)��c�Hb,nAO��%^êyc��_��Tu����HtL�|� ������}���(�%����W����n�@�1�������y��ɹ�v�4�F�g#m��c����[ܻ=�m�����NR�=vHS(�Q|����x�E:b#���D��2|�C`�w�6�o߳���m���hī#��`��P��-5�Н�}����<��ba�m��a���G[�&=��2���*����BdvL�����4�\yƢ#��O$�@��~:ɧ�Վ�\g�F�.?3F ��� �aݺ&���RR��p4��g�\3Mj��tһ�cc��nC�!�o�r��p8X^�m1��s�:��-8�<���o�<������4��Vx��9��"~;����C8��̂aG��P���ϑ �w�6V=�ݵ�h��<�����)0G�ņ_C9I4To>?Y�B"{�T������Z����Y��å5(����dz6H�X���{�Z3hDX?��*bG�	��0W�`�>��@7���]��&k��]"˝p~�&Uw�aT&h�W,iC)�^�򋇂��M�6&1�ïm�M#��}��":	6Q�����%yuf��g����!���}�fE�[��U4=g�p���,����1�>��*���s%_�>)�0!
�Ђ�D��v!M��w՗1�9g٧Zǉ�����(q��V��8t
3�ӆ��M�`U*
��s-N�kI�^��NB���+J<X���b��lR68���BW��t8���Ջ���{]�]���^���D�	�{^}��S'�(V�>��M����b��Q�d�ՎM� ӡH%�i�����r �y�b�1��հ����d��?u@�)�Y�(p��>HpEU���K� �Մ�C���OH� ���GN�V�3����t=1MJ����w]���a_^D�=�Fu�uv�D�˅ ��Y�VJ:��"g�-L����'�ǘ�f^�6��s��p�V=4=JC��\o�����E����ֽ�����T��@k�KS�r���Q�3ǰ��Mav��^�����	�B��K!dě���[��bG�?D}m��U閮���s$\�y�T6;��B�s^m:����KR�%�]J� d�F�>�p��� ��h�R� xۨ�����Y%�V���(�/�-]_bvgX��qsZSFÊJ�R�dH����y���`�6qmu�t��2�z�U�xx�cѨ�7eiQ��xY_�(�bqG�SV�R�=�2�b��;Z�q�_-{��4�tysjq�P)�x׺߹h�����%mlJ�dK�C3-dMy��f3��iLº(�P�ՈqS�uA�C�������%�*ܹ+�'�ݫ�aCg�8�F���t�����q����5Es��e�>8���}���7@�C�c;�`Կ��^���V���`�(���c��l=96#h��\��0@���e�/��)h�o�tt�����_1;]�n�HD�CM(��3�f���?�Y�i0�P돹e����E]Ěgj�A�_4<G�9���̉ �WXK��� ��9c�7��P5�l���U�\(f����Tz��7N��e���v�6XZ��#�qZʪ�&��D�=¹\�"�&ݹ��6 �÷rko�$� �_���[�$ݢ�"�%�|t��$�WH����uuC��SзM�Z̾1¤0���h�XQ����n ��d+XT�bQ��>��#<���_VZl���V�|�J���m�s�NS��%1!�њ<,�������zF�kDL"~�s�>��#�����$aѯ��N��Ō�H��3������׈)�����D.ߜ��16V�Tn���ޯ,Lf�[Jd�P��#-���m�UA�f؅����dΑC5Nа��0�s]�����ܟ��i):�G	��v�=�P���d��o��m�·�_/���{"m���1-�>���9s��|a�Q�Ox,�m�y@Ţ*��)8�,�T�X߳��?<h��W�^�_$�`��,� a�^Y��z;8*�T����L�¥�B���:�U�#	7L��չ1)A�B�WV��[����b�tp���Vch�� (]L���|�r?�W䷤"8�ԙ���o�l�������o�+\�'����=C%�ĭY�;"�+G��6w��y�}b�X0uxT��2���k�k2N�+�pP�d�pA� g�rrH�>\b�#	S�A/�Ty?�,���մ����hL�J���N���+>�`�ӝ�W�dluσ�m�ޢUi��E�[�!�o|i',Z$��WX�z"�9���J��'3�]K-����\ ##nJ�V	v����/�`f����͖`x��$V���ќ�j��9��a>��� WZLc��s�n��M\���z[3c��f@���l<qc@���ͮ�S�,�r3 PI3�P��3�"�PV�lZ)Iӿ}��>J�q����D6���B��WVy�gc��Yg؈���ȧ�e�^T��#_r�G��wD�nlȩ4�]"�l�p�w<A?����C����<��j�L�h$��m�c�ߡ�TгP�#�*�����x�N�@�FC
��#߫$J�k��D��Q`���N�єm�X�-W��� m~����	�F�<�[��G��0�#^a����޽�1���)U���s����Wf)w��Q�ќ3�� �� �t����֬�$k�l��Z�*/�7{I4�	�]��iD(�.n	B�A��������D���ɭl%i#�x�fC1�����b;�,|$��{Ĉ���/��[W��d{�o�X�?G!�{�!	�Ҵ+\�3=�+\V��烹��_ڪ��w9p�-B������8���bj:2���4��0�<j��#��U���a������WbR�Ŷ�����j�:����<{�,%��GI��
]K�Y�d����;���{�$�c���_0�����,��_�E���C`�E"��ܵU��	���$�h�6a�A���[�Z����͑}^g���8�NƊ���T*N���n��yY�gJTl߼����ꏌ5s�o8FՓ/`�4.�Y�K��|�@�evwY��Nl��KTGj,m��44?�af�ڢ?��^�{`�-ў�h2g�n"ѡ�Q��ýo ��� {W���*��f�P�u!L�GX ��*I��J�~Z���ڀ��Km���H�@s6Oq��"Z�]�H���0z�� m����K��>��':_C֤�7����h!-�*�R���X����G�H^�b���$���9c�����j|�=.$�ŧ�w'��C8@F$2ٜ�BR�qY5�B�1�&�%�'iꯤ�r�m۞��X���n%LC��1�e�����CD�C��e�V�]��x���K�����ºT�8��'��RM�Ʋ��
ZAWa�h���L�(�Mk����ܮX�!��?zZ���L��D���*��'=���G���AM���,q��V���b�v;	���8�P+N���������Š�A���� q���
���"j�2+w�������v��ǭ�[�ePz���<�-��u��3�h��b�Ǖ�����E��ޢ2���F�>�;J6��EZZ��w���n������4�����(���rx��jy�e��xn.��]x����r{���	'Mǧ.`�A��ɼ-��Bg�Klh�!��C�K�v/ӎ �*�[�2+ع� +����0��-���`�����SΙ,}!ӡy�W����������� �*k�����B�������J7�Q߅!�ow�2�0X��:�<��[ۿ�	qG?$w6}�����ӏU��%G�ẕc ���K9^.w����t��6^Ү�dJi�|��#$�FdyTSj�T!�����?|Ao�X�m5�XĠ�6a���2\h�{������M��?UcFf�a0�rG�]ܕ��3��+�<��ң��X�.���:�:� IT2H��0�����V.����H�&~%P�f� XK�횱%��E���a^��ea�_[��������uBs#V(��zvq�4)�k������1�i���$yJ�Rj;"{�w%��5�\G�Q��:�T��q��O����5]Wo��\�������6�� ��w�%�A�����u�Z���k���R�%6Ϝ�'���WV6�ϮL�/g`1�0)�n�W���*�Ƹs_	*$�%�h�E�}
�V[/E����܅��e��-�5�]��"���I9am��˸����R)�����03�Č�C�h'07�?IN0?U����n�6��~�Lts2Ց���S�.;�jA�,���{H�,��lS}�3��/���tW�6��o�u�q02�0'g��������\�����G��L6E�пJB�����������X}Eƈ��\�p�[�߅���1_wT)���>}]��_� ��Q4��QgV��ϵ瓠��k�^_��_{��������l���{M���dz��R9ĝY�v��*�,W~3o*��8�qT����W����j�^L�K����n��`�y�i=F� ��!x�.f�?��P�ցW�������/�H�pÉ
������(D��@#��;~��(E)]����g�gW(��w#�u��8f_�VX@b���B<j/~��	����%�qxIm��vz�=��lG���-����H����eeq��</���ܖD���� k'̓�����w�n�!����h0K������v��(^�Ä1��T�e��kK��������R�MV�#�*[z�ISХ|�%��\��@�=�I0��̸O�~_?Q�(�xj-�{����%��nˑ4�a�U �7�n��v�h�����n?uP�|���\Ȥ��P�Ck�޹���f�fx����嫶�s"̚�5<0�@�������t�;�fx�l�Z�0�-S%U)�ڝ'������]Ӈ�Gt�ˏ�<hh�#a�,f��x��'4Y���ZN	�$����c;�ъW���ACߗ��=�JM���75V9.U�����ژ�S�m�SVgI�ӽ�{�#�?p G2ͥ �D3!VR�>DaA1��G�W���6#J�m�8�H�և�g�VN+�y޴Zq��md�%S������̿�p�g؍\	t��q@�w����2{p?��ׇ�l㼊�RL��!Հԏ���Eh5�$��}��#CMZ�p�}�X�L�D�����f�fH��1o6c�e@�r�����qΐ"W���B-��Я��
K�M.w��>:�e��m�ҷ"�=ؼ��+3����ˬ�w�\���L�����y/��������rdM��������0��:�# �減����ɱXAh:�~`iZ:��=�i	`ZIwG��{g�G���M�O�ףIh��{s���C���ʰ�8�����lTJ�:3"���I�H�B<d�V���[�rU }1����D�>�Z�OS�� �� �J��=��AB�O6�ǐ��C�h�8(�ԭ�B]0⡴�D��ڮ<�")H��IbIض��Z�E����æ��7����A���s��H��������$��,��|����� ;��,_釦G����e�C({e�R������['N��i�=�>���- ���KV\#�jD��{EJz,�3$��q#�4@¦S����5�'�E�@��K�8x2�j�4�?�)���$��Hg�!2�Z��"C��ʊ�g�=�����Z������j�HF#Ai5a��?	b��⶯5��rp۳qd	|��X���s�	0�v":, CB&%��[�?�����=�N^fo��rh���1L��g<x1,E��5�^B�P����&"�%Q:������Ѐ�L��'>}�*� Շ���37f4$*��g<rb�㖾^w���kj/�y�!z��:��ۚT]0���q_ʗ���\��	��)�NA)����\}���c����.{PX�pF�M�R�~�3��Y�g�"J���p��Ս%��Eב��~�'� �#\4:��d��wNd�d8�4�yhbuT	��H��0#/*�nr�*4�/�QS1��=*���pC��>�Oã)K'��Yy���d��4�\ބ)���z�T����C��*�?��?��]a�[WG]>)+�ȯ���9����!��)��1�����b�_����f�-S�����^�����`2@�uk`�m�_�����g՜Q^��T`�2��X�5�!�f'�==��ڼi�.z� "��"�N߰�Rp?���0)�:��W~��n��m��
�
ոΟ&F�T��`���ر�V�z/D \aV˕	`��6Z�$��̀y��r^ؾz�:�b��:]�H��i�a�
�ϣ�d�0rucg���Dy�t����ֹ��68-yWz����������Q0W�o���Pf0OӇ�Vt,���z8�!Ϗ�W�i���*���(�5�g���#-��>��&G���62�U��Cv�����/�^|Reat�C8�g�n:��֔���>���a!��G0U�FO��S��kE���`
͡Th������+�Q�[�U�M~#D�j@x�tG5�T����n��,�ƻR��� a��[��燙��l��F3MJ��l���d��ɛ����b�K��*ꍧ3�ڿP��o3T�5~b������"y*�ն|H���!g{V�^��h�uq�{���c���z�k��G|I�:90�D���9�@Z9����MCF���@���q��􋴭��A��<��0S+�zO�9�$#o��҃���pF�q�� ��xam�� �GŊ��>����*�����V�aO$���ո	jnX���']2(��'��k��V��Z�H���$�k*<�z�O��*���fEu�~��{ѧ0� [5�"8ey���D)�vM�ٵ&U�G'�S�Z��vj	�S�R�i���gd��P�DK�of+c>��v"y��
]�MO֋8D�#n	7z$�W/?�t��L�·$?�&I������XU�����K���oe�'X�@KR�]~��{���g�L���Fn�F�b�^��Xt��yd��+tMGb[g%�VJv�SW3�����*N��t��(٦-P���6���Iw��BK��� ��r�Y�(�@�o�F�+���Ǭ�r�Z�Q�_ܹv:�_�V�v�E���E�x)�����Qr��G�N5�iS�z�^�ukJ	;2N�fE�-��߾�^��_O�֢��🵍��eS�W:H�둪p7V__}d�*�O:H!YW�3�+8������X�Q�^B#L]VST]J&�(�2�.ȱ����ѽ]���ܳ�Q�yݞ\�+�#�rF��+�� ��{]Q�+Rb�ʦ�U�Ǡ� ݙ��z�4ne fs_��r0�h�r� 	/ �����u�h� J0�oH\su��uz��O���O�`�[�b���eY7>[�$j ԇ^3�j�VS�8��);ξ$�#��e$|��?����>(q$'�Do��T�ǛF�����O�w�w�_��f��P����\�{��0Qupsbq���"S1aP2�}n?ؿ&5.e�2�67K����ö�����㌏5PG�R5���Vq(���)M^Q��P��n��8y�=<_��9ѶVgW�)�AZ8G�e���E�B� �Jq�6��7:\�X���`�s�֪��_��)�<�F(Hj��2�.���0h` �y�k��|��e����w������!D��7�/~ ����9��V�'�����=��,#sj�S�����'��_$-e�S�ҹ��2j��x9��:
�.kO��S�MޘJ�UQ���M_�
l��ܐʕtɆ���x�m�}��ܥ�Պ���\�,���+��:��v^������(g]����A��<��>���\��G��sWu���V�� ��*K���SP7��O��"����o���'�ْV�f�}�uι�u��kѽ��{���PJ��T���l��D������m�J�I��L	x�M�T̲?�}]�4W-t��m]?��O�4<ipS@�I�oi���z�ݿF��_�kJsE,����q2���"
�wL��sL:�iq���y�k�NM�T�=tH�:Z���x�2��[/��Iei����Y�s��ǒ����b��u\�i���
��&Y���y$�Zո.Q��NP�Ј�"�&S/�y��a�l�J��p�}6����]{ܫP�ִ%��)�\�D�t�;iš���r����V~�亶n~:����+J�y�3�����n2pS9��~эzB��ћ�^�� �"���NVEn�(�Wr�T'xM�v�.:�(GW ЮL�"O�q9C���8I	�ѧ����F��DЦ�;.��+1��r�I��JacBe�k7�F����&�'o�z'�OME�k���>�@�����R���|�Ǫ��Z;�c"3fJ�HZLS��b���o\F�"�U����f<F$sm�I��?I���V8O.�%��0��7h�!��=�|P������q;()N����of|������R�B�J��g�#'�'[i�?d`�#���m���������h☨�c�^�|�Y�}�#* �Q!��"��O�&�t�Lh+u����Ph�������?R��̱���g��,��qu�B?�kl�y��~��#�V�W١�'��~V�"v�ˀ�l}�A�s|��n٭�F��_��Y��rbmiȑ*�	q� �{K���2L�g�(`&J�: ޗ%*D�5��~�@��¡�\��o�*}��^A۬@xH-��M��'Z�9e|���G��:�G	�{|`���鶨�|���������I�`�d_�8G�6�8�7'^��O~p�d��5�8S$��j�h��J,d��EG���H�	�B=��;T]cb��ź^.��T�׮��)[=��̠FQ|�㡎5m�'|DNI��h���*����Ϭ�q�$k�9�;u.;pN��˟5����n./5�ft�[���S;�<��{L�`:7��/�)�Z��Dm��s6��g1����`�i#��XH9�{]�݆�o|�B�7�`l��>(�f�rz�8!�϶��6�{'�h�_�|���q��uI��|�uQIY2e����B��WQhL`�a���؀h�9^��5��n�ɀG�W�fKȵ�v�$��ȅ!pw�U��y�"=ѬX�q�g�)��I;��X�6m���k�mhw�_��	��r��>��O��吨dmIV�%檷fܲ#�;"��r�Z���Y��m�3�������{9��՚��R,�-��k�@�T�N��;0�͋�4��Ã��˽�l���0�4��IƄH��j봶V@�;Y�J���XI�D��8\�%yԳ�.��&�/*�̦�6u�w<��%X~
�Q/�0��j$Yi�="}ˆ��b�;��	KƇ� N?�oS�l�xf�i�.ؔg��v�����s"'ҳ���5���|N�^�Dօ�ѣ��a���CW/�fc��Dَ����*��c4e �b�-��㿉������5=`n��]��L�g�p�}G��ݎO��H#i\�}�5MeEU��Y�LZϳ;R�d�\߱���V�\�w�?K��I�k��%��GD��$��|��!~�=�+4��s�v$�N4$���I�hl�top$� �[.���I`��]e~ױ�+�GG�{�{{��12ulh�i��6�-7s�{�q$�#�G̩�ٯ�o8ӧo�$�X;Hq>V�U_�"�H�A
%H�w����M<�lxA5��j�� ݴ@���o������@����s�yP�1'<���{N����3����wqyM��a�n���L�I��<��h^���^2G�zUͲ���j`��9=W��W��=6.)��Z��4���-�����m]��+���O�wXr��nd�z�l�/.^!N�l��7�wn�u��F�ڜ�OT��S���z?N��Cў9��uME��rʐ�V`xs���Q�|A��WG�%TbAa�54ݤ&�ܩ)�h	4�?�kg��h��u�'��'�]�KkB��z�\I�`<=$~�z5m\�m��lTx��S(�@	��(w֓Wdx�����W�&��I/.���� �l���ɐjf�Y�3��������Ŧ�m��{|��zjY`��a�S�, �J�뚫�?�.#ٷ<��|$��Z�d���y����8��&��EDf��Ѧ��F�n	ԡ'����x�0�ۚ��a��}�#�Ӑ}����m�>4�S:j^��.^I Z�O��2p��+G,����v���_М�S(����tf񞗜��-Ϻ�ca������l�R�+u�"�ԇȞݓ4�ILMٿ��q�1�`hmn�߻��A���@s��J��r2�j���M�~'��c'�˓�j�q� ��ش�˥NP@Ϡ���j����l�5r��A��;��@,���*YC3֡���u�)�橵�����[? @\�����'~S�;K��TX�Mz3�Z���D����P�s �	��i��"�P �V�l��,���3
�y�G�9��|	Cջ�4���Ûn�[�mS�zڒ����*�����̆��^i:{|]�����͈�7\m��X���&�k�\N}N�־x�,�,����u�����d��0Q�0ɲ�W����χ	���5�i�ߋ���}�k��!?���*�_Ƒ�a�M��-�����c+xg���p/v�MfKhZ�nx�~\8[��)�����d"X�9��<�kJ��n�8��IbHLSd��9���k����dq��jڒ�5�I&�9Y����w��̇�����A} ��.�����*��׹j�?d�ak�p�lC��fr9L��F�

��^���#|��	�R��m�)���,ޙKV
�$?��F�)?� rI�m#�~PcFٶ�̼��~�~�oY�?�Od� �+�N�c1}Y�*}�e�s=�QF�>�2���r��㺘�C�O����3(�4s[BI��	h��j�����y��