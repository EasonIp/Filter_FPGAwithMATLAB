��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�η��$Y��!��+��ɗ�����6����&bq��j�#�o���ٹ'މE���QD���0@���G�wAT�ܹ x�*�'afڱ�L��+�'5P�.?�JSb-+�D����Tls���(}�Mi�x����и���T$�O�lO0_Ų&�ҷ(��@7d	{xx�E;�{���e�5�e{ZV�t���)	�1���R�3��T��Q�M;��� �Zs2`�s�^Dr��f�ۄ*�b2�G��6��.[�в�?��h��@Μg!ɋ�?	�y~~������-�s%;�z�?
I��N��W-���m�f���ڽ��M��7`Ԏ:!`��qӜe]��C��+�A����Tnd����Ve��S,iJ��d��O��s�z�_3C����B���E-���hOH��ut�x�Hw=��?�oxS�O_}�2��q�_���x��#��JS/r R��o~�f8nsVK�*��Oؖ<�m��{s�0���?TN��XV@2dR~��JE�o���?:�΅%�7��P���GJ�����oW�]�jQ��a|O��t�;�C!9����o
0Z��?�� 7%#�{��O 31v�k�;�e�'�z'�5ꦢr�V����Ǔ2ܸ�/�,�k�+�_��y5���ު�FM�9A���2z���C�8����7c�p3z�5��n3/�k<���Y+T��Ԩx��%BT�q	Kc�n1h�tj5��^�u��ߖl�a
���л&�^4�Sn����mi�Z:���"����:��V�}��(�ŘXN������@(���k�Yz�z�}Yh[^k\2Wo�����V��`Q�����N�7}��������#0��l~Qٲ6B���E����x�T�/lʬ�z���n�+�H�c�f�$1%�g�rvo�n5�&�МⷳG�oV��
-���2������t#� s��K8�"�_wY=T�����gʃ��Hv��8���-�f{��#�9����.�S;V��&';�,r��ԭ"�.�f�����G�l{��6�)�� �x�yM�9�%#k�j�9���36zOZ~V&P�֡����"�O�Sܥ[e���l�׭� �x8	���2�&��=��]_=���o�sP�o���t��6R�c�f�8S�ߚy�7�r�	�P�)�5�r��lD���'�R�%��5F�3s�N�r0�q�p����vX��
�!�<b8J�08�֋���eCr=�?p#�w�0?f���J��
[��g&��jx,��x�d� f��w}q�\?M���:D��E��o��/q�8����R�Pۀ���}{�-�r��/�)��(Nˍ��84�͹�.7�._�Ǎ�2�U7��6�O&���|N�fŴ�#�f9����׷�0��-�	e�f�T�+�Z	��>䲴<��M�yY�
�L�� r��c�F�@�3��B+S�Z����n�7{ւz�u��3��wt)��ZY��@R"�"4ħ�{U$������!Z�T�!��j2�RC49��'꣭�߹�Wq��<�X��K�=Ѹf����k�~�{�'��T�m�� =�'g�� J��V�0�c_~�x�(`��t(��ve�n�W�H����߆k�O���d�π���D�Kɐ`1����*��p���#k	���M|Qʩ�����>�C偻�a:�L�� ��M6�ےE�������X���� ޑ�o�`K�UY���܇��gY�4پ���==��C�U_�֖_��z�QTn�'�ķ��?� ��%:�/���o���A����3a{�����]hQb9�}�I T��P\��lb<���Ey[}�T�H ��!��N�gƭ�L��"۵&�S=r7a]��$����ƴY#�F?n�m0���x��s�����ʻ�-sf��JϲP�]˃�8i�zUJ�nR�fE�Qm�Ճ� �d�����J%qqtp#'_���:L?�!���L�&�濂Q���*�CMve]9* D���?�q�06�<3"��5bs�HP�t]n�n��xw��_�kf�K=OB�/+j�;B#AqFa�g�JZ�kq���P�b�9�n�������p�8����gS����k��w �G����ͷ��������-OZ>�`�cةa��~�x����ɔA�-��S��	�Kһ3��'�������D�׽W���a.:	4�⺆@�EK�d�d�J6�!�#��0�@[�(�c
9!���2ZR&f���\���O�퓒#�a)⌣��^0�����[P�!vs����"?o��</igr�Q`A��oE�Wj6��P�c�^��"7F/b ��Λ6-��-"a��>�R8P����<O�=В�'0�K����D<q �3J2�9����D�4Q=2�ׁ�۳�<#��~?"�zzR��hK�zҲ�8���ͺ+��*��1�A�j'��F��|5� V
Z�}P��������;�~��z��J�!������Gq$xbV6���s�9FE����+�1�	#�n[a:��ׁ�+:N�������]�n�/RS$zd���Ԇ���_�taz= 7{�����\�1Z��MHb���N\��@��ҿcK.�,�V�[�@���3 ����^�'OGI��`t�>�H^�d�������6���
��:����m�L�E�!���82rJ��O��J���k�@��k|�H����q�M���:��%������@��.��I��q3�7�ϨV� 6�F�"���^��+��{�Nw��?�FMr����~�l�br�f�
����������HvY�B���C�s
ڠ��+���de�}��X�y��m��n�o�J]R�.��[`�(�j���Ȏٟ���i+WsvV��=���}L��]T��F�F��&^�7�e��%��{E����u&NM�&珃�Ok��.�n|��8�?��,� T�`q�_�¥B��Ϸ���k�H妘��~��=W�R�ǰ?r��/o1W5���Fֱ�&*�i���%U�ŧ@5l�[Ek��\N�ͺ�4����gוq�$�i���*����8�������`*R��O�h�A�a��'��A�s���C�Mn�4��|�q-o�J�ۨ��Uyg�ÔCÈ�F:M�f�6;�9�g��-�)��3�l���Ճ�9��`���F��8WY�
>�&�/~����l��hz�%�ٮ�-�?�eu�
�I�QHQ�zT(��>��Ё �h��8� L��yE���.V.ݩd���/xr�_��"�����hGZ�z�o�fǋ��j*O~�$�i����&��Q���m�jK���ix1�UnV{ؒ�"�&�f�ߐx��}u�_��ʟ��A