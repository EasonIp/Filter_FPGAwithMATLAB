��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K�P
����$"uI���10;�f��� u%J�Ċ����t(�k���_�ڭ҅�q[�Y���hB�1��
c�,�'�`� @4��B2݅�0�$�;fb�l�!�Y�l����&˄���ؑW��n%����zfT�)�u|nM/�ϓ�}�K�������'ꎮ�s���L���9{I�\��w:<2z����;���	̖�X��%ȇ���-y ���vv'�(g+P�nL��p��p�ť㥲ݤp1�~��sA��l`�
oT�:�^��ic3��b��2,��7��:q���.塚�E�D�vL��gӏ�e��aJ�^}1��PR�p2���5���re�������$�I�I/nf3�r��8�x�W�́�.Jڕ5���N��X�c[[�M�#�v���I��r�q@e�you����>�[ͮSù�y�LL�I܎u�?%6��Ԑ�'�Q>������Ȱ8*�T'��:��I/�U�,�+��b���9�Lǉ����]R��MI������&�B1�=��Osv4��v�q({��䆽
*�Mݠ����ǽ���vasA��"�6N���la./�DM�=���J8&��ڱy"��D����w*�k�i��U�����]�Q列}��ˍܥ*�AP���Ӭ�QŁEe*+��ɲ�V��k���J��	XM����.���^�L��H�i��� '���9G�l�`��c���q4�L���Ϥ?8uG�u������Z<D��Gk7"(��?��:eɹ�1�lQp^
���"�v[H��Ȫ�34��R8M��W@��e�n-�4�<2��J���_�bI���#���/ǳN�xہM���^Ҫ�!�+��1L�G;��ګ[����hk!Mm⟚��Z�'F?>[9�z;ysE��I���>��w�2�'�C�v�{�+��C��\�e��q�LtI�h�>����.����U�GŊ�KZS^���wwr�R�1��̏�2������X� ���F�=��Dm.U�{/�4 ����
��:a��������(�M��/[OD9�K��k�z{���������}c9Q��h�ﵪ�s�5������r�H��6�w�����ʸ����
�ڎ�n���"P��7�]>{�� ��a�">.;���h���Um��5�sS[;��z���J�VWZ�w�"���Q��o�=�m6�P=��zɯv��S�R�Rgl�IN�Up) �$��|O��.�~�Q����J��ص�(O������;y2ZH�29���L9h�������K�+O���
�f)#��f-Mi��?ɍ�d/�#TUzV�X�s:�|7j���� UJ�V{��Q�������J4W�ښ_���A鑂�P�s�5�(cp�A$��,˔[��.���q���1g�Q4���ɟ����'����6V%��I:粼n�j�8�ߖ�Y�jݟ뾒&SsOqwN0by&�!d���Bo�j����\��rI���XɥN����ʋL���J9�x��*��FC?1�SY#e��L=VfL*�1t��A[�3�pf�#��$�*"@g��N�&]�D^Gb��r3���l�%��\��">L{>���uJ��Xg��;�e[�
�c'�����ڔ�)_��� �v�c��?X��ͮ�	�n�O�S�����~�aKm� 4+��c�_�rxزJ �J����Q�va j�RCԟ��W5�J�E�؂��7��TN�iW�+��j7oL-�ȁME3�GcS� �-��)�^[
n-q�9��◻7���*������юGїŰ��E�R�2�,�o�&�H �0�[�TF���1��b�`3������@����$>�ut�4�Е���I�
_�$�CEv��օ�'��mt��L�O"�a�/�Q>��+��C<�M�y`��	�'�!��������������Ϊ+j�����Y�}J�(µ�;��,J��Z#�.S�ͬ��!l%9J�? �enJB}CmW!K�j���Y�g0�j����߆w�5��!�W�u[�i�/�
��38�S�K�:0�Z���;�ȿ��� 2$3B��C]ff����Kl� ��+��P�{����29�=��מ��	�Wu�M�{w�	�߸Q�U�7>���q�x�5x�q�:Gk�����p�75~k�,���qYP5NǦl���Od��F�"��%o��?�_��)-�+O��ĭÝ��'��$g��Ś�H3������#>����rq`����졓L�Z5�/�0��$So����̚�R�;n���9���:8Z��7^�8-�v�x�K�r�Ln�%#�3%�Y�L6���.�r\�+8ʟ;�7N��s���˰�s�S{��}4{;A���V����;�w�FAf���5��s�Ӎ�~�Uun6n���j��1@<LT�2����EPEI�G��7�L�e�k��:��_%,�����˃��t*��pù��dJᮀ���ݡN�>,���je����.��t��(��s�jc�@��^� ����Y)NqaȀO_���=�R�'�y��|1�9�8�x�(s�YMF�}5��V��H���)0�[IQ��|�Eq�d��W��� 읕4�O�o����u�!��9d����X�Ձ�?|�vDC���:tT����X�33 fD��q��*�Y뢁,���k��u���<c\�T���VYzo�?�U��#QE2�K��oOC"7s/�*���t�v��,<x�$�h�m�7coz��b<'a 蝝E�n]Q�Y�%������hr6��������q�*��S��9x��df�_�5FV6bT}5x�}���{��A�����sމ=��G��f�����1���p,�k�+���1��s��-'�kv������i���OK�����_o�^!?��u�����υR֞����1�Zn�����'���I�w���U0%^�+��6[�A3������D�O�(m?q��3ɓ��տd>4�*�	����_��}&�G�G�iqG̮�͆0P�r;�*��
Z1c�C���Xԋ��\g�|��._p�w5&�(=�tu�A<�����:����<��X�EH6�r�&+TV)2Ofg��,˴���^p�A���y�k��=��B��=Y�	��v�t�_�����VG/����%+d�P-�p1�]:\1%��R�xv~�N�h#���柋���`*�?��n%�՟|�2�v�4)����u�VA���r!@%e,�9�\
�?��uh���'!�`xq�Ղu���{��5���>����E��5;4�ha0��s��<�LĈ>�����
T�66��6|��O%���˧�?j��L�Ai���VA��O�C���d��̘'3�7Ĕ\�
���v������,���]���/E�'y�Ms�����&����`��c'o']�P��%/�x�p<���ۭvd'�]�&�}^udz"��z���.�����A<�K�x��r'I����Ƣ����u������'�h_�P�2����z����m˺����+��-a��B2L�O#�%��(9�LB:�D�N	��Ex6�؟I����^�O; ��H���g��K]���+Ip!�W!W�5�cۺ%!E�~s�Wj��o,[M`<\b�3���i��'&O�ι���D�������v�G�^�����q�(m7^�r���U�:
us��4�j�IW)8A���2��U��P��q��=���fِm7��P4�۳�/�%�;�4�l�K��כ�s�O�S��0#�e�$o<���a_�7zⶡ>�<;���'=�T�X��ӇX����
�8CyM�8�@2�3Y].C�Y;�jI�lx�]�4�Xtz��M���;믥��Oq���ɚ>0�e�|�"{GFԿ��d����Z�-�%Ԙ_&m�_+�D/���6^��{0�e������TJ���^rm�����T�=�ȱM��@��G�k�0�20RI��QJ�9�7Ҷ%��O���8�N~�m`���B�&�#�ݒ,H�Y��<\Qr�nH�׶��'K7&�0���Y��b�WB6J�3�1;9���mh���Gos��in���k � �
�y�o�Ĕ�l,?OD��x�Ի-_~jFri�=^���/�o��������&Nz�A�����.T�ӊ��޲�BsPm@��@C&���Ԧ!��~AD�������>]R��@*V���P�&��7[�h��&���]��\[W1��)ߺu�����n#���`?M�������2�]��щt�k�KﳺW�PybE��C��t��'�b�;b�p�R[&W��f�)��H�}IG?���i�2{*�5�V��c�x�T�?%��Evvo0@a�~��&��s!�:WÝ��6�,��(s�Ȇ�aܤ�h�p9<g�9<�l��T�k����6���V\4�t����=�$Ka�:���Df��y�r��	dhܜp˂�s)��"o-���p���_��&3#��@_J��+�J_?X���|x�Zi�Aa�ǒ�� �ӹ�la��K˙[��`Cٍ�jbUFù�o����2������3��J\J�1��SP��%6�Y�r����i�r�Z\��j��6���I2"�މ4;]�W��r#d009{O�M�)z���`���;��L)`Z�Q�{��P,�ҹ����\�M�,�bج|i�%�r)��@�� U�������B���s����L$:v/yEGnA`�1���0�^�_(�����p[��yX,Ҽ��7�������zH�������|b<HCY�͢�hjAș:�S��ZQ)��$c�����GsWD�>'R�l^q�`Z!`)b�b����O}*:ǆ�s�Ю{�OB⛎�q�c��C�Eݶ�����&� p�����<��4��S�����y�sV
A�^�7�!���>iH��ቢ�U2�jL�h�ΑG�a��gu�j(��O�h%�K�2��a�p+|�	��n�������:t\��֞Z��q�@m��m�2F��;(��l������fS�k���^4϶8.�����(�w��I�m�f,�B������ m�?���#<A����)����ͮN}�5K��aIS��>��[�z8?쟂ų�b b���b'uʆ'�P��-�D'ro��Mw8(u�^�G�/���<>�aJ���~W�S�pw�.Ɓ�vv�r:;��e<�]��K����Ə>Ue|(Y�1�^Gl$�$)�-qü���\�LР\;=hdO��7�W=�_3>l������U���aI��.�2�i�>"�:���R��>���'���0�
����Kl7�CI����
��d�q�!w�|m���蚙ޞ��j�Kx�܎.�0v]p�����9���S��������"���z��5.8*���
N�<"<D��0��&nO3�.!���L����M�y�����~ti�վ�w�t��U'-8�%jqt��԰ӸO{�$�?��?h��y��o��~�`G
.wO^LXHT��HD��w_Yꪀu�b��j{���EV�vU����z��%�������K���pHq|�q��""Q8�jl0��Oa���4&���VĎ�U�!q��]wU�f��Lʻ �%O��
�̆ �YY~�6'͉dӰ�a�����nJ`.Ym�Og^H�
 ������JYH��ћRۣ����E
#��3�N���j|�W�]���R��bg*�X�M��a����t�K�I���km���r	=��9��D2�>�{_f����K�����z�M�dl���_�wk,8���3J��f��ԭ�\j��׻%�ʇ_�d�_��0��HRu<��,ǊG��2JV<*]�2�g��B���z��ML�m�q&��7�
���s�'��1#�z|OS�~�6�h/ �[�*%��DvįT�<��l�Eh$��^��Rp���2!mN/���r��vE,�L���l#�8� �u��v4�.�뇈ù��gq����D����G�d��KRP�<�;��B�U����8Q������6�:Ȱa=]�����/�@'�K�C�ZY��9�,�qvQ�D�`��������9i�(�����ے�	+�$O4�M�e[K���.��� �'�5ޜ�G�s�e[KM'�<AH�?Y��%��\Ij�5G��8�5�#B��f�����4�>�h<��d�N���$=I/w���v�o":v���Z���n6y�
�}���P��P}�Xt��8R�)��yE�mɭq`�T6JHb	��/�QZ��Ս���؎N0���l���3�����Vy徒cK: ���^���,�Z ��k��H�F��GEM�������q�1�y�mf��<�?@��
����/��@jH�r�D��
�Ho�ʀ�R�J�0Tf��5���E�!G���i�Kõ>�h���g_>틣�.��b���n7D"Z3.g윽�#"0^}H�_�G�ξt�k/V�>�ͽ�*[�gC��̈́*N�1�?^/E� ���A�O�����1�'�qη7��}Jł9�Ϊ���-i��3?��B<)���쵳��]� �'wJ�*(@M�b�t[�����7t��[A�_�D�&�&���vl���_m{�d�^#���=NF<����B�T�@7�ǬJmx��@f����!q\����#o�H�Ƥ!+̯��v�N�Ò��:�L�^�2&���^��ͅ�*!��э��\��iD�I�s��Y��Nz:3�j,���rdW�B�Q{7.�f_�d�%a� Nhj),*�o;8�BǙ�o�Lo %q��:A����3�����r�3C��� +���u��L��Rx�=��Bq�9��{ �mc=���"w�@�v(t;�Bx��ȓ�&�TA(/�^ 2k<�9xF�V����/��)H����Hx_n~^s�Ҁ�g�hg,!Z�D�SMID��/ɀ_?SǨPL��z#�� ��ò=q���7��I[� 8�jxi��g�vx?#m&����]�|�p#��tv@�*����2�^r�=qmKj�ibؼ.��i���a�7�o,+��R_N emfc�%��[��ܲ!qZi9�V����m'��~Tk��^z��0�`w�j�%�|�O�XݺG-�V�����d�0�~�ג5Ԛ ��积P�lDfSl��N���4&�@S[��Y�+��g�e�ZBِYE���&y�t���\�C[%*�@���ap����F_,H�ֽ?xոJ��)��{xͶ~��� i@��F�S���`���X��tl=�\�@!�l�(F �EzP�0q����*�\�g��`�� ɜ��hX���
,�|��##A���O�p:^
��2�2JK-�Ϳl �Tk*7�z�6��s.�.���Q� I?�Ki��m��"�z����R��u�ރA�e;ă����Ѭ�@��z]&4ʺ����]çs����ˌ��{=� ���E�$�JOA8���>|S�A���k��#�x�t:��M3��5W���y���9({��|3��k`o�'ˌ�탆�U�,/�jR�T��r,��2���(%b�n4�d���Bɵ�4w�)wKyRZ�D܆��yXR��O��86Q�@�\跴�{tфk�EU����f]����m��}��5"7%���\BY���(�V��Nnw���?D���W�#Y��vG�"�>P���/�t�vZ���='4##g!���ld�����9�Pʄ�7kx�av�Y���$������<b��ըs���L�oTDR��%��F���8Hs�5��W�OI�(�s��Z�4�c���z�`5YZ������y'Ij^�D"�Ⱥ�����B{��������NB�φ��l<��*��I���˖�d	�3����E2�Ǐ,걽S+>�U/lc%�`T��/X+{wഷ�i�At�>�b G?e_�$*���/ۙ5�Go�pB���t�����y����N~"z�h�'�\�o���{0#���RQc[%�[0>�(Z7�W|� ȣl�L��:!�r��}�k�ƽn:�.�(�� �16*��0��ۮsnJ(&<Ď�l��s��c�_�>3]G�Gғf���4o�߀/�H��� ��%D5z� ����ߝj>�䨣/8�ps�I���.�ڻl�ގ��Z��'����B���I��E)�8�]�P3�ǔE2�?���?�泑ŧ^`V(2��şԫ ����;���u��o�~8|���A6�����X%A����j�loxυo��B\t�$S����	@���Ǎ<}��:/V�Va���<	S��F���Q��&�1c�Iao���z�(�MV��g"�d�H�W^���"�$���۰x4�`�P/�õ���<~��{��B�X�S�8{?�%k����[�E��A,�ǲ.O�cK��E,+��!ފt��AȱKM�n)�)r뺶3:(p$U�T��E�en��"fܔLcXu��%J�.:<I�i�����b��P���m��g�r-MzgP��;B�}k%ڸ�H�$�չ�jhb�}��(�Lz���ޅ�#\��|�#�#�ك=o������C��
� k��g)b+�|�?����%���WZ�?���OK��U�́L�"�9�RW�&&(3�~/��Åŀ_CV�y�$���T���QK���8ŵV��+�dB�HX� 
�wMS��ۖ�o����<:� a�~�4�bHF��؏��Cl�*ߕ������a�;m�)�9T�t$/�������M�U����/�@r�J�ٿ��]�c����j6<�Rw�� V#�����U1WUTL����C���c)ߣr����s�FÌC��ӳ�ү����m-����ougH������������i4{��]k*4�ZSf!��Y���u��B{��x��شM ,��,��)��VHo/lW���)ͧ�� ����T���lr�,�U��g > ��F`�h`�	�Sk}�J��\#}��Y�4M����W�`RI5`�9l�o���*+v�iN�;�>�(��ΧG;��3�~��
/q��q�¬�Q,���X��(ŅEm�?^�s��pL~���+�6Y0�5�.��LiԶ�$�q�t/M�������A�{�;�y���*����]&�B���yBj~w�<w_a�QU;�a�M��r���u�Amĩ��_dI�j�xh�B���H�19k�f�P7��T1a�tY�I��\BqF�`"�#����bŞ(���!���j"z����J	YQ���6� �}1u%M�� Fam�a����{WװN�},�ȩI�^�nG_O����tޔ�&�:��r�#��	Q�Č���Q����N$"EC�o#$+O�����;�p1і���YU�i�p�$����E~����!O�N<��#�Q�[`dW5j�u��W<a��~0D4��H��<ɳ���� Y^ ����L�뀩]�a�b�d$�^���k�����C�8�8�o�;����,�w	��I�q�� ƣv=����Ts��	!zt��
���6T�d���SX_Vl,8ʻ�Ǚ	��'ⶲ|
�[=C��<�Z�4��@�|����b+�bCL�QT�g=3�X	�F
8?<M���	hz�}�����곴�� ��xD�dZ�3��g '8�te�>QY(M��K& �ͨ�N�%�<���NE���c��wa��NH���
L�7��&����� �@ŀ\`Jx{��d�Ɗ��͢]���e�Z�M��Υ��1R)����lH�� ���'|�#�9)�G(R*��د^�ud<��K�����>�Ю�m�X)�/	7N�E\�e��,~QŴ�6W�t�8\m��秀m��T����r�9��ٸ�g��b�S��(
�s0$�-��g���ј	�SY���1X' ��|��<� ��ڵM郦�1س�@�:w�<>�;���ܸ����]�:��~��'YB���`8 5��)�6Y�W�x�
t��lFQC�P4oO�A>�_�UڇMTvڮ]��(Fi8!���⟝����W�%�u�d;��Y���.��,x��\EF��=�������6
e��R*B�^��.���3���'��Nӕ�+(0�?�����6Xҵig�H�zJ�FH}��1!u�)�Q�i �gR�+a]<��,Y����zc����"y[��.5xq��U��b�)K��>�5I
!��YWf��Z�D��{N!z��e�Vtn!���	B*��7�Sn��ZT�>h���2���c��3�lq��v�g��`�i���D��ι��S�J���֛���.+����vm���cz�nƄG������s�
	;�=��eչ�~$�������ڜ6��M� 0l�7�v���t�������2��S��ޟGY[�A<�X{֣��h%�y�O*!���:���U����ם�:L0%K��:��=U/��G&p�E�`�o��x�%i'��Rs�km�~z��J���rz�*E ��8�!�5j.�ʜ�b�w!�Lq��5����ɺ��د�1V�Om�1�!��{��x��������9�(> �l͖�E}mTҿC`���z4���	g�8Sp��9	!�ӂWEE�/{D�k�yA	o���<E��sA��7.���g�Z&V���z�'�|���FfG�{`�C� s�%ϓ�{0�c��T�{R�na`����J���5r��������i9@62K�ꛢn����u]+�pڃ58�M��*𴍁;y�T��<ZDɈ
r��o����{{���4�zKY>z�4u�hp�W�9��rd���)�a�\�ca
$��k[�U�G@��ж�u��Uh�0{�o�m��X��-p�&r�9�R�v�7�7���Ӳ-
���:�����jO�溞���&ѽ�G��mq&Bc�p��Gb�a�3��b_�f\�N���c����jr�1�{HK�K[�K����n`��֝�K�:C����;�U
o�V������d'�tb�ڈĆ'�=���G0v�~��B3C<��(8�i����u@��`��Օ�y��[I@O�QwK�_*�͠�7���.��@jv{�8A~�rYx��G��S��&5)jD5$��t�/���#ƶ���<����RՉ�Z�dN���e��"�¡#GP���6Q��i��:vt���h8X��������׵��\p��J�(ˑ!�kw+��$R!f^��O�8��O����.>!�?�#3L`���*����n��x5#M����=�������	�ބ��16g=*Wh8���/���xv�b�*�m(��Q�̾���vZL�8��&ym�E0�/k&U�ee����������_���s��f]�[�|ƞ7w���Y/7�g�D