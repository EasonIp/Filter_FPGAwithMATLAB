��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,G��U�	�oJZ�@�z�����>�� �F9!�/_g�T@_hm/a3^��(#z�dZ�E�����v�h��|���-�>����w,.��N����9Z�S�p�ւr�p^������[�G�C-�Dʩ/�Pm��[F�9�U��G������y�嫋y^ch��,e��wٝVČ=&������Qc��4��b`��B��c��o����|�"Z�G�_g� �z��ğ������|���W����,����o��U>FZ��Փ+Jucsj�4���T�U/c\97���C�=�Ay�����JH-�|�hW��L^!}�  cU��.��q��$��ޖ�뙐'B�L�J.��- k��)��_��m���kN�hh�� ���X�͍D������ip���"hR:�!�I3�Q����~�����o(��
6�? [�U���r�H-41whȋ�i5J�ڷ����"G\�!d�� I����y
v�����hg ���JS���s��Oȓ���T�\U�	�+��?5g=�+�	o����;�����,���m��#T\+գ
��Y���U.���d���c��Lr61��d.V�=�bps�Yz�oxb.`��[��ٯ�hh�u¸kJf@a�`�U�6�����"yR#������ax��7�tL����'�T��$��ϳ���Oq�-��*�ofVJ����tLwE�'Ϊ�`Z�/���8d�bx6|�=Ds�vV��&�o��\ئ+�̼���������0�3Vjޤ%�T��@j �ٵ@-�\��IZ`K�_T%D��X��٪ >,�:�b�^?;�+��?�=~��l������1��62/xU�|����&ǐaF��!H�;��F��L��$y�k��ť�<o�q,�G�?S��и����Z)@i�E�s��K���H�/8�$�azu�*\`�8��w�Z�
�F��	���!�οZ>�tUv&0 U���&j}��Qb��>�V�"�F���8�b�Z7j��HP\��Z���j��74� M�ۥ�#�x�8�$I	S�4��Q((�������k	�,��9�t�R��u:��uo<m"������-VK��
:Z�'9F�Sߒ�!2P�3Z���h�ġ�Jk!�Kx�󖆂��oG<+Ca�H�a��p��;b��w_�Bj��%t�ݤm�@Ρ��D�}Gm�1>�{?��c�`����K�Ё�>(N<��h�g�[�p�X����Z��y�$��kW�1|=�x3�ң�M{�����2��"�v,BV������(�-+�jZn6+I�E�?�.�"������ >���}��z�3�Or���bg��#T`�Bq�s'%4���V s������n�jV�;�Z�<�3/�8�Ő#��=](ߏVGHAN���F�9�,k_Jm�ڴ��$-��éfO�,��I֣"����M��[gs��L{v��ժs*��n3���XԪG�(뻓�e��K�� dY^Lֽ9���X�V�� r<5�w��a(�~de�&]��Д�%�9R��:<yϥG��l��o�����y�����Ɉ� "���w��B'�q+N���HO7�
2ݰ�ؘ}��S�(k!�:0|V2�y�E�~a��P��	Nh@(��Ķ�(�p�l�( h�\?"«G��q-iM< �z*`�~%`�I��c�}1+H�lj��e�D׹dC��T%p77����O�E =��:�1�EaR�ALm[�X1��H�� vh��?����v�
�����^�&&��{�1��q �nK��E=F!e��(�-�#{��\�}[��TU�u�6�	�N�a\ã%O�"�X^β���t8��z�����VG[D�[`c�+n�
���!�0s�5P�:���@�'�L�}@�ՑR�8��(e���A[ҋ�L
p�d<�X0�	�'*i߉?���U�U���?��L{]R�n����f���2��%��~)���o'�|�{���44�oQ��r|~� �w��+���t�L�׎5����1߸ByY�@��KZ�\�����⽶3 �k`���Z�Ͽ3w�39�`"�L|愿[>��.��P�=�Z��@�qA�q�Z[)XBQGA�������*��uJ���ĩ*P��B��-O4�B��[J�ޡ���T�+�"m���>�~��TEhX�5�h���c-������)����6�eb��}loy�M�r/�n�bJ���V�'��c!��&:+2�O��R��`�S%}�T�	�k.�v�-�:Pӻ�x� �1�É��ɗ��0�="��x��w,=�H&!;�bd"_�&����}��R/�KR¤q�C�w�Hu����2�y_ta��_m�`�t�>��,��&����򅴁%!ۓ}�fCp.�_��C���m�/��@����'�֋���om�퍃2�)��!��.��+�� �^'��ڕ-��`4�%���s/�]_�nTh��|����*�8ﷲ���m�9k�G�Z���n|�o-!���v�w�d@`!�K��b���:�gv��in)_ؗ��X�s@�H���U��
I�}wC�8�E{���l=8>$nQ����Zp��ۉ�U�c<�=q6��n@	j��t���:������<s$�<�u����.-�������)��1P�#or�5̚8vI�\@���$���� ��~��oD���ĜE�W��]��	�^]�_Q"Q`8`gbdߺP����%GCK�����V�ԺY��Pս������*�Q\c��k�_4ճ#S���u'*�o��r���8�
��-,��[۞�ư�gЅ����z��.��h��5�#^˿��@��>��,�V$�.u�� tH	�F����iV ��,h{�1+Wc�y�_��|!��E3|���Zuа�C�r�|���*Xrz�%�b�~.���f܁h�����?]�Hj��-م	jۨ�︵�trĕ�aZ�P$eZ1>Hu9�S���#|���'�����2�,�(/)�� 8�sN�i��D�(��@X�y�̨��JD	[e߽C*�KZ�vr-}%zu���f�Ƕ�?��O�E�'^��v�ǿ�!��D�^�w�W�#:ރ#YXB�I��� ��Æx��+6���hc���H��0Efݒ�9��m$�d�x����Q����8��Z��͝P+�G`�ʮl�e@�ģ��`!K9�����V����"-J��I�-�<)�SsR����RJZ��e�{���䂰�4��ON1��޷�=�(1�N�=d����o��}^f��d� 3�0��I�O*�F�:��x�	�Fk��:���FW=Z}Sd�G�7�8ɧm����P��±	,�� ��wy�Ѝ_�h�j���YO^u��*��6�*D��:S���vq뚃�SF,�'��i����r
�x��{�F/�,�P�ds�8��A�bG�5��Γ�"՚ld����C	{$DB^z~��6�gIT|?8��{|Q�˚���qF�����������*by*J�
�\
D@��/�BR���5�=�/������"S|��%;N�HӬ��!\Ċ��wԻ����(*�;��]�6�e|$8�վ1鹧�ap�'���!�	Lg�xP3؏�#i����P���:v�����#-���B�����ޕx��^��W�͸�j�K�Q^�|	Uc���ZBu2.��v����@W�Qc��o@�bv�)��#� v��	��1we�70�Z'5-�q.(��d8�x:仳���~�y@2���u�e�	+�4!*(֫0]�˝K�)�Ѻ��� �g�>7�|g:t�g�#T�:��@�d� ���(c0�� ��'M�=����2J��0�x��|��=����h�y�KN�����@a���h�9�ך�/'��ȟh�Ns��E2~�J�y���B��F���{���F��ҽ�y>, �R��y0e�%%���
��"�!Y53,!��=�'{G�˓��f����q2��,H�	e�����	��a�O{��P5�$ܸ;�Q���������2�� �z�:Vڃ�.��ZQ}N%6>�wL7l1�CE8��a�P�Y��$�xj��)Ţ㯾�9]��I�vR�׮� ��Gތ�jV%�_L�+U��f�GW�~bQ��HPʈyd˺��
��AW| ��K�aӄNl5Q��|�u��<$�9��T!�]�6jXOT��&<2@ћn�)&Z�#�}2���T܂P}�9��w�K���$O�E���mCJJ�.�Z!�Myc���Yq�g�����o���oM/�-p	{�u�@��'��-�