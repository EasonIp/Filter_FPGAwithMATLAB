��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���2�U�z�[B`�#�� 3�����E��R�=R��1��TH�G��N�����` �۠���<q��c}�޼Y%�(�"�sڙ�AӛXG�{|��AT��x�PL(�]������r�@�h=n�O�^����	�{K�*�q�a�T�FV���:`��Q�օ�H�m�Z<A�=p�Y3������ϭ�;�jHz�#D(-������Γ�Qk��c����{p������y�q�K�Ʌ&�o՗Vy��P�N�*��}f�G��g��&�W��$�R
����a��㯅�Z^<9:�G��S�kUZ($�%��]&�A��Q_�+�\�~�4�Z�:��iI��`I���E�G�&d;���;u�A���|����"n���П�d��D��+Bӏ�}��r4:җ��	���ORG�CP���|?:�8_n!����R�Ca��V�@5���t��͹��i����MX&��;kQ4�>)���3�%Z����5y@��?��?B�y2X&2��\�{ń�;�����wܸ7����,�Ƭ�DE��6����률�
�J�\�vU����T<��A.zJ~�<��=0b��d�0�lG�=k�+i+�Ʈ
�3�DZ�������y�W)�a(�G-I���8����@��:��jX�nY��W�ݦ��d�C^�Z�g�����f��]�ҖF�"�.����&��{ñڷ��C�/?9G8���!�DMw]����e��A��$�m��mP�NT;��g��{� HI��qT%([e�^L�>�=w�B��a|0?:{C���-�_�[�X8P=Ȝ�l�� �5%n�&ƽM̊�/��it�G��Q;W)��r''�I�� �,f93�?����O["�"'?F~����CzE5K%�?e�_���&�,J�����/�oƦ�M������<:�v�q���:�R�R{2���Lm�����>&75r�Ll}+���,��L���@�����)SO$r�e*O�ƴ�S	��/*�l�慢����W��욌~]��@r=J� � Ϟ�O{��v��;���O:��S�`�^����� �ۍJ�v�3}��C-���@��iyɆL��tYm.�^�њ$���A�64!��-��-Y�*�� �گ')��rل�v�:QNaE�BI��kv�9oH�d�G/��g�&<>>�]�L���>���au�RM��3Y����I��1�2����Rp�95��xW����dqR��Ncr�L�$-�}H� Z���C���'b-a�Ԍ���J�H�󐽦��=�J�	za#��@^9akz��Bf�Hk���\�k_ڛ�-��ʷ���5��L&�D�b���v_�����6;q��,n�s=&�<�I��O�S��Y����87B��Q���;U����Cn��Z�;�O+Ŧ���)�H{����<L_#鬃���IⅠ�pg��Z��#�&�.C�f�{�W�9����=����c��|kp؊.X-��i�x����#%� U�mU�OAR��a�F�:RdX�f`w$�f� ��C��xu����[c��:�+��!�G�G�������8{M{���N��E.F��~���C��~��K����	f�҂��0�\���Ϣz~�����u����D�$��0�fPP���x`]3D(oqP��n��Nq���0�u�pm�rF^��C Wt���]��bu��r��4�X����k%�`u�iɔzD�����#q�r۵F��ʙ�PC�ҙ@����כ����`�����U�CUr���i��~�$��'�"�#������w��WG��?v�0�GI���/����")j�E�r���H3�!m��:�ܞ��L,���Dף�ba4��Ռ�5��p8�! i���dA =u�7���ھ�Y��������ӰR���*ύ7��n�^a�Č�����F�]}�R�̨�u![>���+�_��_�9��"������N<I	]]r6U�ċԔZ�et7��}P,I?����Y��P��y���:�p��*]<t݊��_�ڦ��������!
b���J;0�ɨ�·�u�i��K��O_���1�!%�i�u�7�=��\l����きO����
HBWV�E ���{�ir��o%ț��T�QH���B�!�T�'����^�B�5����?�$���S���{f�#�������c:ײ6�2���w��+S�s���LO��&�RQ�(.��E�q^��L���j��q�ȼ�&����KzΑ�U��d���"�r�#q�c@��Ǖ�F5�9&u��b��	"5�̣���o�I�\���2�:0
jX������j= a�t�j�A�Gx$�!�T�f$�w�: ��{��u]8	k�e%,������ke��MH�� ���VR���D�"0��|<��v��G����*P�{ZM��<��0� N]��F/��[!�_
���R~��
�H��#�yfs���Yd
�@VT��p-�����Ȯ��f­��
vI!�n�M$rF���_���5w!c ǎ�G�`�<�L�g���;�4W��1]Ԓ\��KO����5�������Qp�Hb������U�L'��'N
,�,�<������W�4��ǰ�p=rk����)�K�T�98�I(�D.�ǜ�b��{}������KR���� �1� ��K�;���_.����ޑ��i���R���[��7����B�=���D��9OdW^-�a6����9g�/]��H���A��'��fM��P���pC�擷='�M(��:����3boR�ȶjb��r���`Q3��NS.F8j�^�Ɣ�W%�Ñ���&y_W�������n���^u��#�A��V�1�x<@�~	b��C����Z��0)��A��s�V�2,��x�� ���_�U���Z;��m��	��N��I܌�k5XG����b#rKpxE�����%Rc���P����S�kl����G���ج��Q�� .�O�al�c���E]^�*�NE�󀝅*��p�V��A�}MP;����Pl�|p�M��'�X
�Z�&�5.�n�6Z�CH!�z|�7åP�Ug ��^eR���E�z��5��K;�4��;]�+>KxHk9���4�l6��3�tF(���ig���8K��f d�=��k}t�H��}%����8V�g��P*t���GTvxJ�(|��϶��0�ە֣<:u��H�gV5�:r&��n݊���ϼXم&휘R+�ګ�E���N�fp�
�g�����22��(�n��7:�7����� ��7�#��x�.�*��e�,	����B�����p��g� ��#".�ɣ���
�!��	��(�Fϙ�BQGu<��Ӛ���}
����B�#���S�qr=v����:����ο�W�uD����y��\��d�&j��T������"R�[��H� ���������'i��+�U4Kdx�/�|Hq.�rL�H�C�9nP���s�Y0��{:�ɥ���p%��~؆�=�3�trz��� �<���&��u� �I5�o̬�����w���C��J�8C�7�������m�Y�?��o��9*cK�0�٫H�!�&�d����<a��E"t�6$n��P�(��P/)��p��l����I��Ι?[�A<�A������&xZ�BU*��@�b����k�������ze��p�!p��v�)�N��U���H/Q��Xp?�&Y�fB�9 $�H����-0 M�E�_h��}n���	��"��)Z~]�*
Y���O�^��O���SS�� "�W�A�,�o�̀e� ��o��5T�B��̀�~}�~̒�SV�2�ck����z�]"�ˏ��,�� 1l]���1�hN�����$��Ck�����ci���b�,��$*4P(S�Hn����H�}���l�� �!������W����:���_��W�lf�=�%�*�%�%`C���%طm��7���������ء��%�H/&�䭃�L\�]��Q�J|�	=_g����V���P��� y�ѫ��qռj���.Rog�3�t�\?�����7XW�Y>�b �_�O-�?]���z��(�\E��o1r˗����A��ޔ�9xB�qb��$_{�V��2[Ķ�Eտ�H�êrZ|����c��&Q��c=�L���,��&�����K�ZS<\Uu����d�]8��RSm�t��C��G{$o�v��J�DǓm��{_zl�.��9/�d܇CQ+����wx��y����4t2��h�4�ܜ3�o���4�5}$zHt0&��?��c�")��y�h�ĭ9��.=�f;WI��4}�ގD^�FlL/E��#u��,��:%��kt����GʑA�%VY~�t�G��(N�u�C�n�U_yWJ|�@�^D5o)�Pv#$��Z�/�D��ؙ�	���
�w�6��W��׵�)�\)V7�h��,���L�,���\����M�t��K�qF �jz?i#�c��b�QP�`oD�`"Q��y~���.;��{w�7yl������mV��粫��@FD��I�t�R�@ �N��>�0�v�L��)w���̈����ar�?���8�q.Q���X��%:D�oL�� �:�34�F@� ���*���sHΚI^�e�8G�o�`�_?3Ě��09f���$�U'>]H���~yt2/�?�|�P1���F�ZM'}�$�ps�R��E�#|�E�ۇ���ﰋO�NJ�����`7A�U�Bf~id<H� �d9����M�=�>�����%�����E�k"�$-?c�{��V�!"N�o�C�������Y�.:1Ra���z�����	�ܫ@ʍR�8�;e+����(7����U\n��#�)1�}�r�|aq+l�����^��4|%�Cޠ;����4uDB��c��iq�*�e�ӥ�g���.�?��j�h�]!�l��St�7��=�U]��O��[�g_,6죾Ѻ�m[��h�v)��i�b���e��IL�-D�B���T�FAǊ5�{cϖF=µ��}e���y��0�l�����:�}3��^���5x��r�w\<$1I!Y�Z[o_���&���5��:rKx��Ԇ�Q^�Ζ}ս�!Oz���t��6d�*ř����!�{`�7EZj���~�JF���
�S2c@�z��Ba�� ���͑�x���Td���7o��f?�n7��䳒�:V�`#F[��� ���ĹK:N�g�P�ୃ���PX���*j���a�6��c�M���s�� ���߰��&� &��U~ĉ���x�	ߓ	���R��W^3!��!���1���,� �l�FF�l蝫���d���YӁ��������� `��}�w��z�B�N�������;���**����AA��q�J���\�g�H)��粮Y������r�Ѐʇ�N���Ġ�\E�ʃ�g��S.o[�o��	I0����lj� ��ܽ�
�}]�NΏў�=�hZ��OI7HRj|P>##QzB�j6PVe�s��N:���P����U�	Ҷw��.�l0˫��Gɺ�FR�����'�w`�V��>l�z����f=V���{�ޘGg���/�sy.0q�B?���j�ڽ����� jm�@�'mN�A*��ʍ��	�LQ��kL��N5�f��S�s�1lǽ�R��ǖP��Rje�Q�#Đ��Pw�.�:�}u��ʻVkZSS%B,����s���%lܖwjo��;�Z/M��L[����I�@�tILZa,��x캴�)2h	����]�~�Y�䙚�ѕG}�m[:���ɰ_���$@n��>m����,��B��"|�wΎJ�����Rz��IPx�&)��KQ��D"t&��o?�8�=T+�]Ք�`����h਀��q/Rτ=��h�����𗭖�x���}纓�rK	�_���w�����C�������`$���X��r��J�ygS��iTT��G���N�p<9ըM�
H�^!�lϐP�~��l����^�5�u%Pj�%��7�l�Yz�#��ὃ�����#g��d	�(�~-_�9|ЮD���$��ˬ�J�M��}k��pH:�N3in꼕�b�fZ��]�R(5ƃl��X�T���\�|I�����0~�f�+�GQSzK��9mS��I��щ4U�pY,���У	��j7P�����=�oJ���D�>vߕb��!��C4���{�ֽL���dn�(�=OhSf|��A����R�U4�%���&�FQ�<���"3
��@ol( �#O��r�T��@�m��R�.���/R�F[΀��k��A
��F&�Jcؕ�T+w*���s��1!;^]�U�(�s���o08��.�E�_fJ&�5p�U�ԑ���A81����	�<Tf�!,�m�RI:ǳ�4�l��,�5��ɴ���E�2���7����9)P�_[Ԗ{dc���k�cYɔ�./AV��'��׌���Ҧ9��e6�RR��~�
d�����_vh��J�}�|�S�֐CX�ϔ����O��t��tDpCy�խ$"B�{ey����(�B��\�:4̙V�RL 1pF�GG۫�}�F�p���d}A��h�����b>NT͹�Δ��+��-�g��o�Q��T/�P����~D��{b��Z���/�$�J���5�F���[;p���=Ak�<�~A����84���n$��������u���s\�X.�( b�8L
�@�\�ŋ��%!�����dD�hd����%v�?�/g���z��b�_'�j��Q��:rٶ9
�F�7>��h�g|�����^�i2��8��Z�.�8j��GK�������t��d��OJ��j�H�Z8�9~/��0´�"�=U=e7.>�j_�3*O�O�Xw��
��ar�j"Tڪ��A���=������C'&+#��w�_�`;��	mE75�%Ik���J������O��<T�o�a�i縤p�|0s��xq!���Sӟc&�5R��Wd��x1^Oz��ж���I�{�3�I����Ko�*�GjCM�<e��� �"�1��U4j���+A�H�$m$���e�H޶bWDgB�(�5Ś6���I���~1�?k�n��ܘC֥��〮Va�C���1ĺ
Y@eb���+��Y��63����ZW=_��+Q ��ŏ�A��s�U��r�����=�J[*i��(/�(.S��u3��g ��LZO����WQJ�Kt�ܳ�"��B��ى��F�(j�����j�tk=4�����/�|��^���eyqYo�C���x��J�
Ls���e\���A�Hؿ���vpy�	����\q��.WS��M��Q��\2(E!vġ����޹�n�e��A�&w��d>�T���}*�XW�r�J�+�PM�3B�,�ڒ*8�|��K]���y�<�Z��L��jʹ���hL�K�3�STH(
�o����s�N��EzǄ+��)��]�OI���>gM�Q�h9,�=b�۩�{(h�-��ZL�-zK�T,���(HܰF1Z�<�R�B|�g�<�Z�$�d)����j��e���n�#��!�$h��݇z8JaH���I~�ݾ�����`��^�x茏����:�\�´P�x�-z�˱�H1J�l�W͙�vuvh���D�� �x5�;~J�	}�F�b)��t�@��}U~��?���"r`8�ē7�^���u��3�B\t�|�n��d��E�F>~�.&��J�Ǡ�l���P��:2?�z�Z��D.'8�	Zri�3�-��Ho����-�m."�s��f���;+!�r��jQ���^��@�l�6H,���.�R0.[X�z����E��@YN1�0%~+Fs�"�^�wOyׇou#��� v�G�Ŭ*{>`Ƕ@�3K��<�J�w��`���f�w��F�6�@ߍ��L���Ӳ�0nd���
��J�K�]������ �I{h�jo�������Fn�*uc��qkJ��0�Ћ���F�1�}1~�*>H���͎=�UR���Haŗ,�J@�mF7�T?�\|^��C%F�q�I<�/-�e��3���LFT��|�:��G��) �T@ �ݝ��p��k9���}��Enu�����2{|G�+N��'%��\l䐐ڟ�J_/88ͤ��D!��'P�V��%��@���-�!Ҧ�GY�M��Bu#~B�y����GCq	��v��}�%�Ҍ�eC=�dq�~���)r�ƞB$��{�lo�)�pR�-X��-��@�ϻ#L�ۼ�W��T-W�S�Z�؋
�:�HF�&2>�ݕ���=�@d�IB�u���eNd8��0� �����Τ&��7��D616�FI68��d��+	�8P�LM~�:\g�0������4� C�4OhCނ7i�G�E
Ƽ��IUp���N6�2~����_V1#e:-�i��<_�i�kP���2��VTf���J�̼^�AR��i���ow
����Aτ����4E�B� �:?[̠�`S���7�5�C���� �x�	9z��8#ۻ����[P�ǰ����Q��y�g��J��V�Aǌ�x�R��ϣp����_�C���]�V^����Hi�����t���l~��0y�)���fȕ�DF^<��P�C��N��Qy�doy�kl��l��o���<����3��]VXs�8����=�K|�GpJB��FC6y�?�oCS�� ��)�`�:���m�ǘ��GD���������ż�1��..�|L����F�f�+l���M��f�է/:!D�0�,dB	d���o+">g�2�2	���?s2ݔp�>3s٘+���"Tfڭ���z�:�xÍ�W^��f�~�-�ߨ����Tז2�L����l�)����Y �s�rA�70X�S���k��м���'�SV��m?�>��G�{�����p3��ʪ�Jj��R��)�����|�O��v�E�Iq��̠R9��w�����z@�<*w=X��"��H���4��]��e��8�S��t�����I�7ߛ�ơp�#_���]h��t���+�/b����F�=��v�r��չ!#�����=�4�P1���50;�R2�<�	r��6��`I1�7V��S �섖6�u�"2QG��"|1��&����f����jR�=a��$�	���=9U{���g��ڕ�T�U���оN=�/�U���8�^IOi�߻� �C�7���&�EwJ��@�����ٚ�|6ī�=1d(�/����°Wp���\)��������$x�&q7��}e��3HK+(qO�z\�c�;�`6�v("�tb�*;�����og�H~�Vobd���K�n$���?�ɛ�~�ߢ��������� �nlc��̀g���z���T� ��&�N��2Iх�(�f���D����E��"&��]Ƞj�qta�Xl��W��%���������9���JT�fݤ�"⯫1����0uz���Jr�	`�,.�q���d#���E�|(�5d��Xϗ���Ía:��6 ��I	�<�2 ��u�<'��Z�~����w�ݦE�.3�1 �w�{� ���;�ŧ3��k�wDB���>�b~4�@�}F���o�6��@ɗV��T�Y� �~��`Oa�
�Z�-ji��%:�4F&��,T��Y�3�ue5z� T��f��������k[%R�;Qd�z��i��	�d��|8���w�l�M����J���j�?��4ڋ~ z���ZV��Փ��6�F�(��@�,��XW	[��N�}�a���_Nͫ��J����O�$2����P��p�o�hR#�P,�A��U6e���rk���73��|k�	?KK�N/�q���BD��T�%Δ�7e�t�Iބ`M'���pE�)`�*K��>wrq^k�����R��db"m/�
�^	"��[��k~�Z
-K�fl(4rֆ�"	3[$�)!�0^t���0ZȽ~ю?_��Av� ��]�f����*Y��5�j[ֵ�ض�O5��ND㶀�r&O�"�I�B�q�:zoO���r��EC�Q��#|Ʊy�J�`QHd��,5	Wa�R��i�%'��'s�.V3'l������>DK��e ���hwb<?%X�.��+B�V�#�
�Ch�Ǹ�U/I�{$|O�7�Jb_L�&XzԘ2��~�).-"}���m�Voj'Q�,u�c����ac�ݤ���Z���W�U֣Wk�Y��iE"��I_h�tGxj7�!0I���ͻcU-Ov�QJNQ�%M���;�O%�o��Җl0�@q����6in����,_�x�A�?����իW�*�גP��=k�6p�)Kf��d��|u���t�|	s<�h��}�f�!��1V
�\~�ޘ�{�L���-�GWnT����Q�N��"�J�T�N�,���B�jx�gw�����sU-1(s�;3h����D��rL/jZvu��_��6�T>�������.�_�f�w�p����{%������cTp =��g�g������K	�a�}a%]���˞���&pA����:��/��c����D/]G�	=���X�k&|�i�l����/�{�t�A7��7
pg���/��\�=����:�m�f�K�6��P�u�0�	6��Aμ����i�]��߫��	��p!Ǻub�d�)�8��D�Z �`WՎq;T��} f���ep����)i�� �T��t�^]��j4�\!�{�m�����gE3R��s�WI^�Z(l�U���+K�v�q�D'�[��V��֚R-�W��[���8�$'O��+3���*E�ZA�� %�����aߠ=�;=�B:=6�22�f:#r��</�5�G����@[�\ܾIztn��N�*D��s趲Z�N�Dnщ���i���4��UT�gӮ�/�3�ɗ�����X��U�����fp
�q�َ)�~j��)�ۈ��2�ZG�Y��~�.����z*/�x��nmr��G3ŵ�M�s}�Jd���61<�Q��z`���~gƧ��ʣ�Q9��'��O`��+�'����"yX�NӀ���)3_e.5$y�(C`�x�����TjÁ�W�ܢvj:+��1Q<!�9��C2kS��q�b�d8/z�]׻$k��"B.��]0��ʤ!<ra�~22��n[�r��)��:5h؅D���2T����i��9����-m��Q��*� ����E��(�9zܵf��ʢ�b2)�J!��X��\@�w�YGM�h�����t���֙�Xl"ד�e�|�h0�����O���`q�S-yT@/}��B1P��$��4�m
����i�ꖂ����F��ܪ��0�9y����7�v�L����[u:���?"�H� ̖�2�"YJ�GS�M�pIS9^}	��Rz�3&�/�\._б�������@�}Xq�k�
�"`|>Pd^Y�A�`V:�|���f���?kP�:�p���-"�`Z�?'��2>S�z0~a%��T���m��]({O�0���w�-DvYV�?J������L��`�Һa�3��39� ���ǩ���yi�7�v)������'�ں�5�b2�0١�y�y
;-�
x�&���%�Gfॆ�a��tWÌ_Έar���E�����	�۫�e�$�#<�a:�[�M`��� 2��ۜ�L��Ŗ�#s��!������y�\���]-K��T��˯{���s2�.�;}�	��3�,f����\��R��!?cɍ��K@�m��$��걣u�b?��� 0���'�|�)����X�Sc��]��>��w�s��f�~�x�$�?6��(�V��H�@쾦-����t.H�)�a�&�Q��$��{�[l�f����UŖu2�0����G�6��.Ep��/1Nؼ�M��Z4\�,U��p�(/1k��ґ0t|D���k��
n#�}��r��Iye_���ͯK�A���m���=;%��af�7��+3�2��+�-��I뒞���b��4u����s� R%��k��|�M�k\=K��^"��ؕ1cװB��g;�7�uY�gY��Q����Q;��t�5�Ɔ��Y#��X�SH�c3t\hǣ`hIx�cG �z{E�&����ӫe�\�M�̻�o�߬K\�y�0�3���]P{�o�hk֦ԛGD��+8[������?j(�Z����c��op���?�r���HQ�]E�H���)�~���e��D�t��ZM��{p�)���A,ũ%�J*4
�f)|��v��R���f!����E����01�\*�l"'������>�\m{�h~D-�IfZ��(v� ������ �[��ȒǇ^�Լ]iCcZ��X�����%�>R��'_����b �x��ߟ%@����Y���j��ߘ9V�lk���1�KuH����i��4C�� �vr�4P�E������$�1�w}jz�������L��O����0�r{@�G��;.j(�X��@���zz2�B�<��(X�Wg�Ƶ�"7�mg��'�eS�Q� g�:�a1$/Ԣ����ޡ�UG3Ed0�E+����V���C��+|Q�� ��� ���������La�&�I����`%�l&��xD�� #�e��L@�=5׷-cߺ�^N����<��b��C�r:�a�4K��}F_g���,��T	\Ԟ9m��s>w�)���h��q�T;b#�!��Գk�*�� �v�ܸ]�E��(����U�+��2��ja ����;��/ˋ$�Uv��g�O8E�z�ɴ�xm4����15����~�o�Y�d�ޡ���U/xj�� ���r�f�G$�X�i�̀���<ڨ�gc��>�#����	��IA3$�?��6)~��47m\�qς���;�)<h�T�Ω�!�Bd0	�<��RC�݀P8V��;�?�@���9ŀ��(		DdD��qİsb0o*��`H�;�Y4��Χ��Л_���䕄�d�\����=;�[2�g�0�W�:q�')����f=���ݨvq�Ë���� �Ө?-���F�]P�Q�M��F����HݭV�����u_���2��>so4"��>M4����,YP˵�cY��C�w�XIC���g�|I�d����Hԋ��dg9��$��T�o�T<�m�j(��B�����P�|Hca�'� Tg>�d�U���{�K�.���Pb�R���N�N]R�Fl b��$�����T_�r5�@�w�Q	Wrw��v��~� +P�s��$ي:!=PS��Eu�v���:}����!M\�WfX�*� �j��\�i���AZ2���������i%'�����y���ڡq.�0%}�n>���o-3���U�������� �����t�m�[��#�fT�Mf�½0�����7m
F�bG]$d�;T���OG0���0���>IPm$i� 8�=eC��b��|���'s����WcJ�G��� �${oR��+�L�zVa�"�D ��XmA�L!��b�tΣN��ίw*!W��2�K�:l���9)Aș2\�[	�"~vPj�l�ёA�)�EֲU�BOXl�UsB>=��O~fv ���׻�6	y�"�۵�"�"Y���΃��h���Ƥ{]_0��[��m�4�2��L�۶�pv�5��FT��FL)���'�<��)^��gs�\�x3�}��c��@��( $�Om~�6;6'zM���p@�Ss�7�2� EA2��i��wQu.M��@��PB���9���� zG�a��/-�t�����>���8#1�.�
]Q���hU��c���XCb��_2�X����� �֎�B��T�U������W�p�.�E��	m�<8�1��e�id��
Wg�Q��>��\��
�nCab��!�+�tr��/�?��WQ}�t�`��W�np�-Qp�ghx(f?bP���r�����XV�{aݻ�=�O��+����j�c=�9Q;�V-䖼�T#JI"�X�g��̻�و�oT� �8ۦ� {_VN.EO�6����L+�O��G�Tް��s���a����0ݓy~Ϟ�a!��O����.�X�D����M�x��.i��Ț�yw߸�%�Ƥ{�����_����3T�#���ťݒ�a6�%�$RcI~�����}T�ւ���v�%�q�@��Sn�P3%Z�gU���Z��sI�%!5�}̺��e�N��z� /���������aV�s}�9~�<�H浅��_K�:5l���.#�ل-��Y�yb�7���bTԌ�5*XY{�h�zlu�JײZz��)��`5����r��h@�	����ao�ѣ�Z�GX3�'˭�\֨�[�6:йM?��c�x`n�;��v�;A'88��tӬ���Yf�o���/x��O�<�FR$c�D���O}�Ȼ��FQi�S�L���C��1��v��n��n0T"<PV�W���{�M<~��	�@Z�d+���y���T}�*h}p&��v���L�S��J]�U@�1��uB	��^��9�|�2��2�t��A�*��mA�jg�в���o�A�F�l)iKPƼ�4b�����Q���i0�-ϭM��FkK�}pm.踠�6zX`ֺH�9�����p_?Xr��$	]���{V���=�-�2ɠVd^��r��@ ��5y�`���}�ZɯV9C~�Uk�V+n^J���>����>�J794��<U�D�0�IO��gQ3؂]8�I�E��b\]	���rWy:;ZV�RYl���Y�D��`���3R�Tf�+��%��Y�⌉�Q�S_}�*�&3د٨ı�{ϣ��%�m�b-
؄�*��k���63��P8���_R�fp7�<9E�&mb�&B+���!�<�ޅ�~�-+Sa`OI����Ǩ�z�^�D�v�nk�x�"����6i��U-�*�\���q�n�L �nVbJ�UR�3wWO�A��؁�I�#:���l��]��;���O��T�?���#�~��]T��JB ���f���/�l㼳�`w&�˴�Zl𠣟:d�'#��2wr�~,�Fꃋ�r	bg"	|Up:�R�;^�h���1 ��\h��?��Fy���k\���2��5�=ω���X���)�o���Vp�Pư
g��R���m9u�a���eTD�QP��#>ٞI���n���sJ@G��M��cr��2���:9׻��o��N��Ăj�a�ZS`p�t��4*33-c�+��-g`e��r�p��d�m�7�=�n)�	�RB�f��EV0B�Iz�*���*N;���q0���c��3#���F	�H��B����5g`
]�G�d�(��;DW\F'fdh��B���N�!Ā�
� �l-��V,��$o�
�.�(z�9�+���1OI��8[V�J�&?�y �ԭ�J��3�b�O�Xo͓)� �\�#%�J�)��2#��:��+=��?����/KP`h��x�~�<
�q�H�H��%ӄ����������&�`��̨w�� wS`1�o����U��>�����Ǿr�}���{���@���7��L��#%>���s�O�[LO����h�?�Ls�_�v_O��V2�����n:�����b~����h�,�8d��8�b��(�'��f���fI�5?%�uk~�+B�2Ɔ����ǅ���e�U��S[�D��SO�/���M��](״/s��O�ٲN "��(��:�hpvs�e"��P���狽sw��L|��-Eqǹ���ߐ)��{�QO6{���S~�Q���,���X���(r�7�ѫr��A�+9q�+:h���)9nس�g��ܙ�]P7��z*�Oc��.�K��D��]�e�Y��+s���o�ޞ�������[��M����Qj��̦D۽�ӓ��Wk�*s$�g�4� ��KK��w�j����?G�ı˘�$���!O}�.O��Ĉ�B���vv�#��b����^֒��mʧ�i��EE;<����?l�vS�C���\���:A��֎K���ܞcx������@�����h�d#��y2��r�gI������lgL���D�c|��a�8���L��H�%��2z�3@�ڷ�6+#��U�8����&�$����:�댃�<��#�� ��/T1�n��l�_�;'� ����p�QG�r�=-3yM:���vLT_v�r	ݶ�/�F$�P�t�^�C�ō����p��Y_X�����6��l��� ��|C�_���P��H##�J��I[�7k[-�O��j�|�E��HvPzN�FM|!�F?!Y����E ����Z�襜��98�7���F3J3Z�q������'Jəa�Y�����|�	n
U�����������2F��# �h�U���W::Q�𿩌�t� X�Y�:���KȱW����K�R����Z}�����,���=��R����H�=��[�)�3e@f�#,���m�y5κ_�!��I�Pn��N��ݷڲ��v_pN�1k	��s�&��e�?���];��.A2M�D�`�����Hw��9#����(�#���6x`�1��:z�/Za�9���$��.A"�q;!ٓ��=�8�B�Ʒx�7� k-OT��
�(l*���^2)ۿ��t�X*��� ����37�����n�.�>-�O�G���^�u��E[l���V�$��>y���	&O��2D1r�OY5��sD/a6���io�H��M>iob/���zQ$I,��mb��W!��,;���k`:�.���t?�әPHEkI�+늂t�0ʗ,�ˬ��7�/ ��t�7�Y!���N�MX�Z��R�{�{\��Wō�*j[�����l"j�Hgz�2T�V��~��րE�ԗ����&ۣ�ث����8�'m�0�VHq.����((���{yx&$���՗,k �&z��!�jF����Ũ�I�{;�`}��&�!�[���c	�k�Ж��@�rtJ`~�1����!
lZѐ�g�{d�@�]�)Nue�k��N܅Nҷ�����/Fy�@�1Mj�`E����B���[y� �}$ fy^P�:T�ƞ��X�58۶�ށ��� �g�C`?4%V��:��Ԛ[KTaKfC�����Q\��dé�Y �`.ht�׀ʐ�t�(i[�q�zd��^=/����p( �cȕ���_�C��c-��x��J��n��|�<���V��P �v��h�ؤe���l��V�	����8������>���(���F?��Ӄ��ID��ْf��U?��$��4���d
eS}�H��N�z�K��K3Am�)�:9YIIMlh�-~X�Z����Ko`�f�`q�,|�o��_]L�Y�Z�+��h�ک�q�i2�)7	��~$oVk�}P���mXeB��z1Є�]������(�l�J8�� D*d7ZF�b5-<���+��- {g;x���7� ���!�D?M�#��&#��'_&�<���A<4���0�_N�!�K�L����S�(�Aވ�K�015_@/�BI��@�J����i%�++�$q��p�m������/MU�,^^&�q�Y��K��zG�o��Eͳ��4F<?�n
�v��1��)dP��0�},�+ؽMa\�}�B�����X:` �o��)��[L`Q�H��E2ky�W,o�
�v���od�8捚��j�p�$9:Щ)����K�����q�����)I��������B����)�0�#V���MNӴ#�X�M��	���{(������ri�R3IN�ji�������wp7-��w�����9�2b�X�*���ܮ�*���-d�"m�j���u��%F}�D�
�k�5g*�D�8$��	5��|���$:�X��S���=~���nQ���L3�/�����=5G���W�����}��iuN��
Z�!���.i��O}��w�s�B%��?.�&l
�Dv�q��lmQ�9�-�i�Q[P�����$ �4���t�2t��Mxp?��'p������84��I�z�S-���C���Ő����l���[@������&�Cz�Y���k��E��t]����mK��cSli6dt)H���Y��y������8����іY�5w\j���Ԯ	�V=/�-����&m�T^$��"	���&bm�0Y}�<���i=����sB��t.&�u�;��dqGɓ�4�Z�ײ���%9u-CqA�6ъ���b�SZo�Õ���6<Xvu��ܤ�&�t�A�"%��=��Y:	�'�0�ӽ|Ǝ�������@��ZP穾��^+櫀"���>��CĺG2H�ɔ�;�
��.܎km#��S]��9���@'��?�� J�H���9�h�@�zH-���>/�	�l��˓�DdU�b0��uoZ�71Lg��@�C�(_X�腁o�Ov(�K?�d�
'�����E����,���-AQ���Z�{@�A5��P630?��;�*���/Ǽ��4�2OKx�A�O��	�R��O��6r�+ʹS���B����=�	��A�ἍHi�;k�UX���з`�q7Λ�I�f護�@9�?Ŏ�%8����ΎgƜ߅7�y�2`	O�-�9����@�ݫ��ނu3���fc2NeP�I����[�x�(���yVk� L$򲥠Z�S_^O�.:�]U(a  ���-n�<͎�HG�F_�CLj�;�L|lu�f��"�/@l�ř��@*
����X~닊5����	y��O��G���~�$�BŽ��ʦ6�J�`7`,4f�'Z?��F�Yb��1fg&��$���!$bE�������2�z����m}�/^��^���l�HSڜ�!G��״��|���Qe9Nv�3���ζ�b�W�8����u	& eX�S��AF 7�>gk�� � �2��8q���)tC�#"���97�MtO��D����;O2����L��`ҿ3"�{��_�1�� 4�>�R��3���Gx5���!T��K(ӠX߉��4|-�".�F�%��fho�t��(H.l[��z8pQ;U>+#�a�VN����M��Z��CxJ:IZh`ǍޡҒN8�rgM��t�#	?�)��c�?�L4������Q�����3VhU;+g�9��2�B��2XmP	����OZOU�i.E����S�<l�@�f�y���d�<&g��s�(��H�����%}�ӡ��搗Tkf�yX%�1*��^�f�
�m����J�����W������	�˅�(��C�舘;`�B!h�3��R2�|I��G�8Q�����k+CwLV*S�n���!����5`k�w�!�n9�:0�	��.o7�w+-���+1�%��$>-G/4ˠ��7��u<2����<o�^�N�!�8a�B�g��x����Mț����5l��gqtR�]���y�97�s���g���>�j�<���v:�����q\FƼ�z Ӗ�ё<�e��8M���3k2�}Љ�rlX�ϰE-q����. q�ʥ�'�6����8�^Ӻ��3\ �	�hV��5ć^E�]-�R�v��߄��f��a�,��TH�O$$�?n!~���$��AɶeG1F.�ֲH���E��e<F��6����E�����Y�p��a���(��;z�K%�j�k=p(s*�+ł��c�X�SjZ*@�7Ӱ%>�n��1�c�+�p�>c��Z�����F��0�YD��@#�g�C�L���6�ŏy"�P$�B������ �N�_Lxj���>0���]MZ�H�$�N�^#;c�K
����'�x�G�IΞ�~צy�A�'��Ih�-im�7l��� �,�k֙CGv���hx��}����vx����9� �H���Tu�婾BqqCr����K���U�C�~�^qel��3��yS0�t�T�c���8��uΈ�o����C�r�E/tlz�	z"�:7p�f�2�3���6�:A�p,��*ϻ�-O5����4�B��nxRUvu��j�GE,��D�ƨhz�v�5u�p�[��u�7Eh�|��_�'l��(���oD�|��V����@��Tӝ�~K��Ã������~@hj�:ysjJL�M޿=��b�1I��N���Z��2�X�G��)��Ǫ���dڸ+6��A�c�_����fh��#�N��q��y��yi<����hfgW��]���$�@\��=�����5��0�׭T#B	��WX:+�J�֮�
f/U�@��J6�	�1�?�|HI��.�)/�3�q8J������0f�G��l�G����Ǎ�
J$4K~�\ ��7aۤv`1�-��o*��U�}�E߯ݪVƍ.aN�+��J,W齥VZb�6������̀�y�p�a!��h��_���y�O;��Xx��v:=
܂9�y%��@�:0 �)�S`>pܢC>��9�'(3!�#t,���Ў\tS�sT�3ԍ�`���#�yИ�,�����C�ؾ��_Ի��ڴ<�%4�Awp������N�(�[�M�o��e8q���5��S�w�_�m
>!MP�W��d.г�LCW5�ꮖ�U+�J�y�fj��	LdDs^w���/7��%�I�[ؚh�`\�6vF���z�u�Na�	���7�Fs
�)�<���|H��0����̑��&4�v���
���[f�h{��@��`�>���z��l�Q���E֢���_���o=ț����~��p]j�Sf���úE�)��E/������1�B��)d�ϣrz;w�����4��.֨�C2��%������4[Z�i�cz�R��B�!ܿ殗\�܂ͱD�����F@�5͹a�ˤ������?��,Y?����d�>��fY���Ik��F$����˳k�R��>�7s��ԞS�� "742�p�"��i�U�����_�����;V�ۈݓw�el�3���,kLpqsR��hs9���_�A՟�gy�;�ד�.�G��;�����҄�D݀����#++������{�S��2�c %*D�Y3Ep�I�lDg��Q��b5Y�[3m�z)s-*�;�0Z��mZ �n�����QH"(XU�P{�xi��{#_awO[[��BdB���eqZl��I���՟N����!a���m~�1C/1�`X̊ akl`�����@`��9���l=�^7�E:n��iRI���O� �bb5��1)�K�H���.P�E(�!��X�S6�/(|���s0������q��w>��C�X����?d�W����~ǣ� s�)�
���_gPf6|�Ho���Oשּ	������S�9K"�;������\�\4�τ��"gF�3��7�E�e�,�	�������C?��¨����)�ZZ9ǟ��jA��s����@t�T��@$�G���YM
���w?�ng�:+A�EI�p����p�^�jٺ`���3b(�N18ݢ�����Qi'�������C��eQ����`�n�^CX��]}�����C��⒳/����d��#A�ȳ
@ l���6�َ}^+uqZCIÛ�`��~���u�,������r��3]�*|�%����H#>�-ku���f���N�3�3=��_����V��*a�W�.�Ї�wݺD6�2�0�������D�\�|^�d�l�tVИ?lU@O��@y+�-ȫ��`��{�6Y�a�h�C���_�V���ŞlDr`O݀�bzSt�w�;
����$����5/cr���[`9��X� 
ͱQO\��_��"�Z����u���P����2X�#N�����w2����wsq53x�?X��6XU��ʦ�AZ�o1z�҂!��n���OI��Ve<0��nk�C�١�<�(Y��R�r�,�M��2����J�X$�Μ(=%�fU��
4������H���E>h��:�^����:7S�pl�R�o��J�T �P��X+$�%V"��I�b԰��ZrHS(���btș���%F��R���>���m��
,�O���C�I��/C�Ѭ?< ')���RMp��Lq9:�c[v�40�Y�����$�;q�z�F\p�'�ug�d�A0�t7K̧\H�g \��P�>}��d#3�����-~�
H��m�Uz	���q\��C���8�12�Ù��
Z���/�t5�����~�Gw^H�*Ȯ&���6�T�8".d�?��� ������]��(�%iw	��]X���/R�=����ŭ�!V��'�m=F�[`*�7�>xpV�0���B�	���6�"��(0�������l��,RĴW���Wr\�X�cT�?�t!�JI$c���-��)�L��D�ѿ5(O,K�+=�A);P����v��)�G���^���q{���0I����u�ޤ���f!�d��TY�\����U����X��*6gD<o�����S�����._lz���Fyy}R�Oԍ@cʟ�o^�]d"���Y��}�p(h:������4q~n)�EblKT�ք*d�?z�f��if/!!�%��хBk�����MQ��?,.A��4D��9�,U�T2���;P�(w��Q��u#6>����Ɩ���]ѳ��?$���"��oH��=Z0d�%Bg�vzX:)ɲ2��uq*��O�
�}�1��T���S������$iIC�e�v"4gTیx!:��u��=N�(c��m0i�7n<��7�nʏ_�k?�HJ��.
��	Hm���!b>���i����Me�(xBm`q1B{i��@��/�B�v�m���>�mE(v���!I��}
�+�n�^슫ў�,&DD��A�7��gy���9���mt�`b�4�Ʋ=@�R��6,��_�ο�K��=ý�����XbH�mq��E��h��f�c����31E3�ó���30V4��Ų��^/��[��W�<�p�pʷ�wv�֕d:Z�96�<�t4��z�6J�S6�~Y}�<<��6�_�[�\�	�#��SN�¿����cJ\Lo��m�j�Gʥ��r�ټ�v`� 塨2~���g�i9��S��ң-�>��7�3�}�������Е�V��ӨK�=���-_F8{Һ>䐺b��c��bj�Ϊ����v|ߥ|4?�Nqଽ�_q��3�jU^҂o������Pg�s:��!ДV߬�֧3�p������e�kەQ������ۓ�ɗi�N5�g�#�(�����|!���$���?VF-((����R¸!5tsY��UY��x�J(�'���{%㆖5���:?ڑ9؊S��o���JE�&qA���/�!�t
�ޤ�YKq	�Sz�W�l�]��:�j�9�����yB#�_�5Vjee�Q�}6�3e��®��,�����I��
��y��7[�td�\�I+o[��d|Lj�|2������]0l���QWm�f`�i�n���8���*YH�j� ��25Sm�Wm��{-F���6U�l*�4t��5�b��X�=�9�pOY�]�@	�l׉T�9������.c���kc�N1���K����y�NI/1aU9Z��YWuM���Ats'�Ǽ�t�����#��3�&x�5��\�/[Ni���|�"�?ц��ġ�"x��� �e��,.@Z�.�0��n��'Y3�b�w�RG�^�R}9m7}I��yM��&��G�	�C�3�P��(*�:�>fU1�n K�9�7�ݬ47��P��(z��b@CF|�%x��"�Ƈ���S���hwɏ.�6���K��s��H#ϸ1~�:�����*�>�g��>o����Z��\%x�?����j�߮��/�q�t�����'�ؕ=���R7�2�ڞ�?_�t[�?w�s6�+d��&�j�R$���!���q!�Șau�[�_�=.p�h�d�+2]�sTɋ>ԋ�-����+��ׯxoB��E�W�3[&p^��s����ӟ��i�~��:`���,���5�K���i�O(LBM��� � z��56����<�׺;O	H[���نQ�M*
��|�����G���L%7�׏�D���L�TJ،"Ê��헥R���B:�N�%�$�>�����F�ݥ9=^���m~/+Q�f9�i�Ŗ
0/��z��
,ښ�!�ڸ��\ŬTgzÐR��vU9�2����9� ���
d�8"U�>��x�'����3Yy22�Z���+�
�%�oĉ���	��4�$<]]g>5׃�OL
�%_�+�6v��T��<s�l��Y��C���I?:O*ὕ�J�i:\u.�z��ї����P���cf���l����PD��U���)P6�_,�U�ܢv�#�:ĺ��%��q&w�o>霹-�c�<��,�a�j�ϼ����0��E��o�-Id��Oݥߋ���ID��������|�;��($s�X�K�&��n�*ڧ�$I�I�a�-��~�7��<b�Ю:2����%��E>�'43��(�~<�w��R�ff.g"]�3�;��@�^�K#���NE뭑D�v �_Wۻr!3���uO�X�a�Q���=���8�Un�F^1yb�J�T4�?��s��+�4��Ļ��	�	l6�e.H3W�V]�_�I/��DT�%�^�ap��u��0����F�
�\��J'[Z;�R���]�2���H[�/����Vߪ�rA��qdp��u�	��~z��<�i| 	�I۬P�����q�j����/P����s֯�#��u|�'��d�&��q��z
w�A�����5�L�!��8��>6�ͭ��U
���4$��5�o����(2���fO�<WT6�Te	!	$ENHap�}�a�NXˑ*��DY�H�o��2�4���z�]��ݐ���t�{��O.f�(�mwn���@v�z�������#�s��f�w�>��X^[�rE����;�4H]��lBޏމ	u�<��۔ �j��I� ��l*
��vG�w..�sF�Cn�p��h�8�1��l�8�� Q�_wM���.�-g�)��������{�}��{�d���f��m�gֵ ����}��{�I�?��*;tDO��ʸ@��h�#���G�t��P p�K��ks�Ds�6$�(�5�0J��7�/������ib�>�F�TiնhPZ���}n+�h�p��+��8�;Է��u.ckųa���kL�Y�U#��̯K�Okh�ҧ���t�O�(}b��mu�d���{J2����bҾݕc��9�ԫJ��EsQ3�-�*���8|���B�=S ���o���6�{�ßqX��(���m�_
�A+��uUv�qCCT���0]��Z��M�4��S���"gA�V{%L��q�RN��Z�{�)[H@o����������L��Ԑ�YS��l�5˟:72��Q'���!��*��b��1�U�o�#�ߢ��j�z�s����)~�6`q_6E�o��`�l�{��C���W�P�bI��/�>\/��*�ױr�Bc�Q��ED��}�0�������CA�"�2�ohHR�����^F��=]ceCK�P��}a=SW�`ϖ���2^T��s� U��y~CϽ=Ȯ�;<��I��}*��!b98i��f�g!�K1��?�鵞N5*:blw��E$p/~$䓎������ �U��$/U�_}�����S3P��d֊�D7�D�o;���}��R^�
\�-Y>�����(&�A�Y�b�pTy�� Un��75zL�K�4&�"%~����h��Z�k�*pi��;z���⡣�r��\���z����o����'^��3��gGo�x_��Y�f��H�#j�����g=0MBo_��7��AM��{+�`�7���<����]k��Ԛg/�>оX��g`1���F�\y�t����7}~9�Et�s�BVu�_$�#m�d�wu�����K])�L�j�yu%vS�s)��%3�n�ʸ��;im#n%���UU�<�Þ8ǰ��Dd���^Ҫ�w-Ls#�AA��Hھd�n��h�������`�2*b��\诲�T�c�Ӂ�7Ƿj�Ӹ�9�GuKj`���YW�(p��ҹ�Ω��T06k���˟�afT;k���y�Z��e9��Ju�8�LjXEm4�ߖ��K��>��J��K�g��FI�0��q����z-�[�V��g�W�R�Y&7��@���ƒ�QT	�O���ꦥ��
�=��+N�7P4�g��}�t�r�ϴ��!�A9SN���&y&+2�)iH�ÐoAS�2,'�� ��n`{/6�#G�����Aw
T+�� D�r��|��!���tV��pD*��>!�tNe0�])#�v�[I�_q�aP���Uሴ��u�'�Qx��TPtx;�|�����{:�S�|������@/��<6�Yj��'-�C�~��1f�s@M�*�%����s����"�Ť�9̢jn�|ͤ�����=R��DֈR+
���<s���K���~Y_�Ы�[�i�iJ�=��'����RK`Ǧ`�f�*���+��ks+�RJ�İ�w7��3W<�cj��W��� ,t�SA��{����*��2����2!C��N@����׺�s����ʖX2��Q�CaV�\��J !�_�gƮE��=���y��[��	���R��~}X�:�FV��|L�0&H��?r�u������|-�(��V����N�5E�Xf��iOy�{m�N4��*��t��v��X0$���'	_F�LW�����Z!�~\6��6�L�̲��Ӟ,+��˿��&Iz�⢸�����Eꦣb��B��
z�N0 �����QŒ��(�i �F=3��������D�h���X�:%�7&���RY���tR��:���pj�A��K^��g0B�+:��vm�ǰ2�q�b"Z�6���5<�*qO�@r#c(��Kxj����8u����;-�%�ն6~Jh%�~����U��6�8�IU��[��@�r�rqH]k�uƯt�%<���A�#��xBPg��;>Yr4m�aw>��#�O�[��S]�!��*9����]���J\��؍Ht?�C��,�������ʻp��'����(;�w�2z�i�z��1̱��?����R�K���S�|I�a��[�SmAA`[/�H�Jd
*�j�%a:C�3
α�m�ˉ�_�tV,l���m;�P��W��wp3k$X'q���r!�T���rͯ��h�+{���V8�C�P>�ߘ����u
4�0�4���V�I4H%��MDw���-=�Ґ	V�d}��V�(�<�u A�x.�	�S�Z��i hb\>Vê��~1f�H@��:A���'�@�/�	tm��.�Wv���������K+��7a~�>�
�BK�	��I&��D����L�W�QB(��2��r�a"�mܶP���~2|%�o�l���D"��/[��
�n3����B ���.�mm���H������R;���~#��rZ���!����lb�6ꢝJ�#/�C[C����h��F�D�v��/pQQ�h�u�r;?x��r7�ZpB,�>��KZ���"����
�X����WU-��1h�w�&�����
r@2>���\Ql��|�7��q_��p|�����}�pǄ�M���N,�kL�I�д�8�S�-�@�9M3~V(<5mЁ�����a"�ߌ��܋^��Q�Ŷb�����Y�gw�囡�y�y;�~m3ܺk��VN�䢒+���U���2prU�?��)�.Z�y;<��Ÿ�H�����jW�;Z���l�x��P�����v��]n\���t(K7�l�۵�븀X�A�J�J�ɑN���|;��ߵ��d��;'aS��N�uP�h����T��f��+�9�2�z,�q�4��3���Lt�&׬B�*��g�9��n(J��ۡ��SNK�ȸ�[W�'�N{�>���\ �l���絺z�� M�x�m�$A���粅׮�{e����%=Ɛw[�&��7n�O��k�\�{Q6�zg��B��樆M��8Q�̤��϶#î/�9l+q�ʾ�={3�v�C������j{>�$�kk1%"�0g��&P:3#լK���ޗ�fn�[d$-���K��	�c�UWT���b7]�e���X6�`�����i�JC��C���v��d���tS�Lu��m�sh�w U�;�(���Gs��~�͎����b�xm����-B�78i��`�3�|$1H���	�Νv*wu=W>���o']�oK����;<<������ͅo��V���{��u��֙E1�:7@]f�?Ua�h��lLZ��qH�<���tF>���!�T�Zqb��,���zW��s�j�&�	����6��}�0GX�˲��	vr-�>KTQ��ΩvBξ�