��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$��=c��7�>ݦ�G�ә�U�� ��CǓ ]�R�iCe*Ā$�����D��r�Y�:;21��*����M��*�3���|�C���ͯ��U���V-�/��0�b�t�^�D�M<�Z��c�z���ϔC��9��|�wi�ʍ�&i{t�����H	@��?~l�^j����Q`s��
��lS��IHGӰQ��@�\U�o�2+��Ik��dS{����ؿ���Բ��B5��k�� �����!��$��a����+2��ZH�|<6�7�+�}QY/8�3y9��٨w�J�T��m���&��b�ֶd���^�����@4]���cL��2���P���s�4�0��q� �zՇ�����^d[0��ᪧ��Tpƨ��|��cd.@	`� �<(�a��5`U;$%�;����?ŝ����?k�t	$�~����1z�'�Ʈ)H� ��Q1�>ڛm��0v�>L�ř.�_蒜=�=k�H&vN��hN��X���a������ui�t�P}�Nq�;u��D�+1P)��P�t�Z4\��S+,��><�"؅���
��s�Ya�c�N�4�a5[�#N�]w(�
3�|���m4�mX�����v�yݠ�� 	c��_X���m�_�c[����6={9K� ���=y����"� �3?�?h�Ft�& 4�zTA�w)����k�K|"d��c'�Z�8��|~f���kj�GQ����|Q�^Ãl���Ϥ��sb���:M���~�Iq�80୸�䧲%�}�*�᭸��r7O��������W�D��m��"`b*ʒ�2��<�����B��&�~�R�{��ѽ�N9}�DA���
��������H�Г�OӮF�ҏ���v�b�V:���ؑ�n���1o�ڂ�͖�n��S�z������(������&�s��|ȽU�5E�?�*\1������q��6����CY�G6�	����ƞ�g��禰��X'5q]@�<Iڈ7z���2��T�/��p��}&�ۍ �8`���>v��l��8��N`����q�Hq1��ԚG��}�Nߴ�1׵�k�����t�'XhA쁺#�N�.��1��9)	�{*ͽ�4FVy����z����fϙF�����v���ȼ'�����ӫΥY���.x͈�&�/Db�/jWL=ϡ0Tke���L��~ŕ��L� WK;�@�R߰��$q�Q�s���z��//zV<���LW��,
:#��:�0,��}�קf�Ҟ�7�CR��f#��nݘ���CP��T�P�֋��� 5��cH�	JO����Ò͠�Bc�d~���umt^���/�P"%���8��f�o�կ��A����N?rXm(���T*,od���	�yU��
V�+�a�\)���C޶��o�q���L˹�tY�9��&�-�zUց��w{����V��X1��[��-�����-��Q$udk�m�dF���2����#O�!�ݤ8���	k�� �笪T�SL�P���G�b��h,Vn������������ۻ�-���w,\7����$�ƺ~�4`�� /�5΍O9��� �)X_������@|@���Kd#U؂q����z��^E�s&�� �W�4N8$�d�V��x�opH��-~�@0��72�\u ���/��x0��l�]���]��U���M���p��D����z�������D�9A�l����`��6�#:'-���A�~�[r ��!�h�VЗ>�!f=�U)*�fp2���\k��7��?�Ճw,�<��9���VG�S<�����R�0��گ�ٮ<��r@��Ej�4�Q�Oi�~p��`�'Y�Ɇ�ȅ����ɠS�����C��ګ+�G�l�A2էL:wÁ�t/þ���`錅l��{=	��p����S|��6��Az0�X Y��َ��(D��D+���H�b
6���W֨/L�G-s7�y�k��|��H�c��R��<!Yc&� �fw����5�7�h�O��VD,o=�`F� WB��i)o�}�6E����l�R�k�k��˻��]���Ό����K�r�K�lA�E��
��D	��7�;���WA�/�`z�1e4����o�AT��g~���B��M�|�"��� �Q
�㭠�ELz�@\������@�Og��7��D*9�6��/mA�/�X��{8)4�(A	D���v��\"W[��7�y�΄��1T� ��ڽG�#IbS�_m(��a��`�� ����
X��1p��j!ӼX�Wd�L�� f�>\�8�٪0[�@�ǷfJ�{S�{gD��"w��d4]�uhij��v�`�4���ex;=���XL��i+jG�����)��&S��o�0��fJ	�B[��&�f�y�N䳼��q����]�G���P-&���{������׬B��Oc� �Ʋa�����&L)Լma�o�sh���D&�5
�PK/�}�^vԼ���mN�\O�0����j.j���B4��e��Ɏ�\|�f�H���]�m�T����k�3a����=����<�m��WS-�(�,�[����ݽ�1�r��:9�5KQ��}��zV1��[�hɒ�鬅�==�o�B���[�"�o�w�@6��e�g��g�0���%�i� ��1���O'I5!Oy��9JZɶ��3�י�m��=��[���uo��B��=6���q��7�z�'jLI(%����v#���h*BbM
��w�$�$�<�����ȷ���!���ˮ�DZ⎅���}����b�&Y21��*R�5�u��3��D��R�����=9�̓x���O�5��k�2�G]d��;~��fEI)�UJ�Q�yU��_�|�x-�D�SIa�~�
<q���J)肾��9n�v��ϧe���~ն\���i���j`�H�Z
#����_կ\bA|�R�q��5��g�2�B������H�?>�Y�������� ���OTR�b��r�W�bK�_����f�+��UT(C�qƳ�0�݌�5��":I�-[BX���j��m:�Ӣt!_j�r_P�䚁o���lB$����s�~�Le��\8��PB��!�Й�E���@?�L";�D>d��|��:9,�Mp/�k���F��o�fD��*f�?`H�o�ம�^�L�����ϣù PTA�����9��g�Z'�j�7�>��:��Ź�)�d �9�1��6B0�B[���f�.�����e�-@�nW!�����Y53�S
�l��ѵ�=�a��Cly�Q}��5��\v~��$��"*8��t��}4�p����Z�&���<�uY���SG��Rd
F"���$��۹��>�%~��	PD-l㜛e��/U��0��D���i�0/|R�K�{7'^�a�^imx?�v��T6$��v�Pp��y���-���cn����/�N��S�(M�L�0�詣Y�)�hgdg����@�!�[>ص��!l��\�]�(�i�_�R@�X7���Bcc����Et��Յ�;�N�Ui)�Jk:��qI��U>y��	�Z�\jMA��`p��@;p��|���,�9��%n�4D���;RBh�AHW��
du�r��U/w�"�dR����\.>#	�/��#O�C��>q��&HYM�7�kI6�h]�.�8�+W+�6�w�٬�`�{E��A�hP��*��I�+vf!��9��4���]�$�_v�W騋n9���(�Vv�iἭ�F��^���f�f������*8<Z�h��>u��B��=�-a�~�&����T~%	��V�s-�#��$ G	�#�>w�����-z&���8L�%O��olu�?��꣒�2¤��uB�a�V��F
]�R���+�Ui��Oh��t΋B�$32Q�4<�s�6�@�v5�Z k�"���4�o:�ˌ��g��+�'�A��Ô���S��FIHu2��d�H���3��N�-��F1�`���X񫡣e3{������e>:�ex�:�.8,�w!휺���®f��%D�$��ONq6����}S��{'���W�C;�� J�(E�R��6R�������ӕkQ't����R;��ӮI�^	�������p�w����6���K�w����B���K}�]��:Ј2��B��;��b��М�p�Ym��Sm�:���?:�Xtp��.�����`ͻy�8�F*�Rx�!�k��O7��S�� #㈳s��_k�Y���*n���O�o�01]��y�N�4=A|EY���1n#Y�4�=.Sk?�ȍ��!1u޷��T2���	����W�T�ߵ�u����*M���!��P���� �(�T
l��*�w�&*��^�_�BFqvkS`ƽDU@5��ӕ��j2�:���������Bkb���u�zQv8{����&nTO>EѸ�F��0Q&@�k�4uYU��Of$���K͝��M�_��ͳ����j��VL���;-��g8�O  ��%���*8C.w2�!��N#c.�<�v`�}&?���p����uu���%�8���zg�(R�I�?S6$�#���r�ٺ2/E]Aˡ�~D�ă�R}X%��at���.
���6�o�8��۾w��pC)i�䅋�	�/�{�]^�l
�q��c�Ԑ�����Q�D�t���#'wQ�V�$�}��/`�x���桓l�My���4�v@�lH)ԛ�Y�oͳX�;�`�[��O$�W���a9�(Q�U	�����l[��$�n�NX� k�78I�����E�6��%��5C�ލ~A����T0tӨ۲�'�[�H�m�/�S�G uqY,.(���ODM�Mw�˓�d�Js������|� �j�틋�H1/@``�ulR�>K������4��b{�»D�Ij��0��(��G��S[�4M�{�T�av��J�ϑ�i'M�&FP�@,�j��`��f��@-j��c���o>w�� j=z~��>3��L�4�r	�־@�:���6X��ֱ!~FPF�H%#I�s{��9@�9�`<�Q��#�R	v����NE��hJč�*��H��e)��r6$,����6��:��~|�� ki�K`�Q>����
��h�C���t_�I�]hX(١���(V]��.:^g#���0��^��~�|�\�O��-�%p
 �=�C >��S���nfBd�@��-'\;�H���(�x�n�4;��V�z���:X��xQ�wwFG&���]�<�h��M=1ȍ����b��]���r�0��6��fzT�Xx���#�|��E��]}�4�*��Qj}�^6^8�[e�������S|������Cp�(�5�$Dy�" (u��Y��R,�2���aK^�����7e�TG�3�Z_5��T찍����R�����ߏ-_KZ�]_��C��:dBέS�C����v��?��ME��
Y�́x`�y��As9��]��Gj��Ԋ!1�Ƃ`�����RM�XU��mh|�rW�AT*�Ϗ|/!|��g�i �U@�Da�F �f�v>�n]��V�+dZ�C�o9}?�Ɲ�@�,�2�w'�^i�vΰ^�\}u���s���4ٮ�8��<���rm�X�ª��H
�h|8�v�]�GǄu��wN�J�Eh�}L��A���`�+!c�6o��D
˼C�:��B�!a/���]���b�"Q4P�ᷜ�q�\���#����z%+r
��^�+(��7�z���!��-��[ �����f5�Y�/L��:K���PFKl������s����4��f�SPs�BVpM���5K���Y�~�5�P*��g�~Nbk=ך�~�S�e:��16Ӿ� �X�hA� ~j�U������^��ŲWӊ=JBn52��Şӡ���~����Z��p��p���5nտ)��[���@{�c�$ה�|P4Ļ�۰���B֜��N8�8f�mT���t�Jx�f��N�˥.4+ �vCM8�8y�	�՗ Z�l�Xe��>CG{�\�q����j[c�{��@�8U�6ao��l?/��c��t���<��)����k=V��,���$�H�Ό�:4L p��B�3nsaC�i?Aߧ�I�z�� �(f���81H����Ъu�#u��d.��9����Gz�Zq �E��wM��5������J����_iA^��m�8)xl���
2��1�Ф	&�q���9s���%u���_�˫Շ9��#CL���+tMpF=�M��0U3^��S��H�կ�\���1�9u\����n�|�v�H��U	�;R��k�5�	Q�~��/Yd��`*kz�(��\ ֳ��e�V�U2d�6w�B0�WLD��ٻˌ4���zh��E�~b������H�bta�*���j��c3�/��V�_a�ʎ��sˊ@}��T�{�ʸ������JY�@�y�^���nĭ�LE���t$8T�
��Z֗�s����#� ��#0���߶�DRp�7�L%E� x�����O�?M>���(S������K���Nː���d�-�j$�/K?P�;�`$IH�p�0�����.�dq�Ƴ�����h�K���Pu�L8����g��f龵4�F#0D��طȰ�?'����E�8�*:a��LР��X�OΟ|��$'����a�;ȶ�x;͎u~D��z����w��O�ki�UZU&Q�yp���<�R�d��w� �xp%�#?gu�G�oN\Ǳ����	S!/��Y��s��gBJa�����8��Z������R�虀f��a��ؙA�BF�g��^y�QG��W����֎�U�0��I��?�a�ϡ����d����]o�a2���4�<*��N}��R�m�M򶇜��8�����H� X���|I�ZE*ӻ��ь�K���i]~g
���5�O���o���\<�ף�E�^V��ِ�e-`$�gQ��A>��s�����neM�=Wy�^p� ϣ����˒>��~	���?��l������:=���J�$���u�_�;��a�7����Hv�%���uh�(d������E�m��r�$���v)o�4Db�$��p�3DЪCvl٠�K���%�ow>Ӟݨ���&�N�Z�ς�8�?�5Õ�En�-�P�ǁ�N�b�U����_���Sq����lrh'��9I� ��7&0��=E�u��Yq��YIQH�޵"� �
Tp�����wl�Ugx�׀/XU9�VP��r���Ѿ��e��i�AG�ŧ�k�!Zn�=b�)�����2��z���LY[kN���~aܻO��7���]H��it�%k%�eq����k����wO�FF�h���vX|�����2c'b��#����q?���mkP	� ����<��j`w����,��ԍbΠ����/[�bM��H��~����Q��3�?].��$��_F��K1��9���dS��ye���t��h�d�+2�"ko2�c��:�pբh/�1���2c����4B�N(�k��P�ݶu����Hy(h�7)ߙє^�Q���,/Kw���j}狲M��̵���g�
�.��\?�C3F�Z�{��A
�(�M=��9��?߱v|���\]��_5��8�B � ��|�Y�{�g��\����Y-���/�q�͗��I�Fy� `�Ͱc�ĵ7���8��ab�R	J�t������X�o�hn���?�V��9��ܨ;�g��N ;OA��:�:٢��J��l� �B�`��q��:T��U�����|�fuh��4���ix�g�,�O-�����T˵h9"EH�#�zwLBb\ ����6}I�_��i��C y���
� �q�L�Ƅ7��������^	��V�O
K��~�s|����D^���r��L��a�����~�97�"5���U�$Kb9+��|I��*7���Ύ������gX��c�����K�a�IZ���jK�fd�^WN��r����;.�xËxx5n�T�M?Ka��(��cX'�Y�n����Yݯq�Du��"c�S�X"bS;�
/�o����9B��fp�M��|��a�З��$s=�E�^W���W�G����Q]R�ߨ�Y�[����Ҡ��/��*.����h�X�c�:��v�H$!?�e�)��w܏�.��_� h�Kz}7p�6#)�a�΢jn�y��
�X���i��4�l�-��2�׺՚����v3�T[8=���|� Wi��9���Z�ʹ;�c5��q҅�p�������߾C��9��]�
atbs���I$�"�g�ǌ ש�X�B������(L�" ٓQ�V��Ψ��E0~��}"���2�="��-i������.;U�R^y\��-Nj)Y�yS����5���R��Um��Y��nz=�CG6	N���LG��� а�.��������!�N���E$��Y�xIc�����0kT��;��nv�\h�5��8����R�E����*ՇÕ�CZ�m�IKJ�^b�v#����w_��di�sc���q�~M�Z�$�@/���/��p[�H2�\ih̛ܶ����u��}�)������8���i�%��Ƭ٧b$J���95˚%�W�Bڞ�vtoO�!6:(QK$�c�;>��Z(�cdsu�#Xִ�Ƃ,/c���y���>���,���&��vD�p�	맦��[���`�{:QGϦ7�SJ�l l�"?�u`T��#��W�)z�7������T�3�~��VRywo�451�?��W�:Q�3i��Qr��E��s��i�}or���q�L�@+0-��s�Z����LImӓ{	}s.�8^+ޯY���V;�7:8-�/� �Zt�
��M�m�{���[����������X�#�1��B�M���W���;06����
l"�Y��RUϡw�&s�