��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQ�k��s�#��ݎ�4Jh�}������!2����s���kW�YCu��ߥ� q��j3��:��ʥ�C0�S�m�lf@q����.{�.��Wgۋ���ʓ2v��K�U�@����vF63q�^�6��\��-l��P|<��K�@j�﫞�[�dp�'iz���vAƆ�:�M��(�|[Q4w�P�k�O�RW"I����E.K�^�k������f���Y���_�#j2<�.��P.�v���dŔ���0۳v���d���_�b6���+�٢�ɐm�s�[k6vp�t;�T� ��F����cI�V���K�-�A $�X)�'�G�n��?8�������o6�ge�EI�Ȧ�ʩ��R����l���%@I�!;�0����J��L����H�S�v�H\j*:C�m��2�����U(aS��(b��9�Ǌ1�~�����_&�F��h"��b����&4^��Y��L���N����,��7p�
S���h
ADw�]�>�A��p>)8K�c�ݣK5���U�z�cJ0�b�e1R��cr'���d�4?vX��^��,��Hkg��������F(Re"��yC��\�04ئ_�]	_}���!��؍���b�?Ց���� �=�������<�`M�S�Q�Ux,�}ڧ��Ć��׿n�B-�HB#�8�HK�Rا<��s��S���Gvm�-FMV.�=�>ى �Z�$�T�flEC��Qc�ل�7������1��+��Q���-�d���S��Df~�l�bp�[�Me����k��{*���= �&��v���#)y��z�̋b��+�TY x��l�܍�N�r�R������c�a9	D�t��ÉƲ�ݥ�9��*�9�4%��HS���I��Y�5�,Ia�0��DS��H��?>�Ӹ&(�t��{��iܟ�H�֕�S�}|c�_73�XN�[�.֛�f��cd���A\�}���+b�v\y�]T+��f,���iye6؟�]��/E纼]�)%H��aL3�"9�MՈ��ay�:��&�p�5_�:#Z�6�����}V�
q�0͊�8
ɣ��}<�B@���r�K�����Ֆ28z?�,�d�ͳ��0�������aW�� gS7dL�����#կ%j5�Sz��@L�����f��)>�,+�%�Uc(����NBḾ��mM4�z็��|��"S|��gp��-��'��ߕ������U�ܲƢ���r�˅V6D�,�X?�\r�����Vc��:�,f�]�A�qp�e��,҈���K9�I=]�Z^�@����Y�߲)�."�'o<v�V��u��_)��%4��$[�Er���ݮ����l���BESʕƛ�π�e��<̢���_/����75�'?���<Z.����S�G?&���[/�K��	�i����,��B�$�)b;�92�l�Ţ�٤��o��oMj�O@k�ǭXˆA���"��iٙ����yn�O?���)Ŵh�q��6#����17A6��]�9��]�=6o��u��g��I�c��ۼ�"{�%j��f�׷�Ȯ���Fs.n��~7b+�%=���1]��ђr�t�*�� v�����ʡ���
"Tl��kϞ�;�F�Z��� Pl���D���Ϳ
~p���䈀��]���k'b#��B�)E"�N��W�Ҭ�(��W��� �N�'+����I#���k��PK������$��a�V���j��$�Բ<T�	=��� @f5��ٲ 0���s�7��İM�.�;���N����Zy�e/���m_ޯ#	D�!/��K��������4�e��ѕK�O�a#��df���x�i�����R�se4�����^D��a-T>|�J!.�.WP��D�g��A���pE��8��D
i!����ń����&�:ؔ7�ѧ�K�Q�@�g�����҉�������(b䦳�;����.��E��T	��ۧkb*�u��X9�]ҳ��w�c�h��
�K�uv���v�Bap	𫟡��0�m�-7�2�=Y�1gr5:����$+���sRA
�s���z)��D�?hM&�JЃu�D����~_:�"� t�!��n�bJ��[���*��v�7��8���2i�Ì���IO�t?��r�U�f�Q�̻��>
�a��2@@��D��ZK�����;v�?����u�R�$c�J�2˙�s���(T�{Ԭ�Aa����q$X��A��w5�oI��jQ����c�L����I��F��(�>33��
l�V��y�w"d�(���#� �Wѭ�VwD�ꓼAI%�0�CS���K@�H#��8��C��S+�WR�Qt�zGp4'���*�ô��D��]A^�Zi3}H�/����0���;}�%ܒ8��)&`W�gy$�B��WJ�r�������Y�e��P7���~�F���FW�ֈe�څ/�h/�Ă��Mt5���o� M��&( T�j�p�޳���2�®Mb%)�TPH�s	��)Bh�A��xk�,# �*j��D�şFb����/���1��ԯˏ�DP~4F��%�H�ߺC���6ãyaY�O H��8���e��o�Yb=�De@�v��_/.L��Fo�4�eu°�O<�2󓝤�^�:��G.���?m!^65^��ٷͤ�Ss@�d-�������Q�����*	���t~�Uh���`�Y�
¥��\䮌:ij�Gi�o��ʜ��?M��R3��/,˕�9��R[#)u�H�џn[�@����I�|��X�7kUn�>�q	���0��lu��gܼP���`�=^M�,ѿ�]"v4u�y_�t8:o�d��QY'����Q���-�݄d�V`L8������t�%9ИE2F�E)�0`zy��͗ix�g���ЩK�>OdR���O�/V&X
�d�Nd] ����Xn�٣�d�
��JU=:��_�C-�o
}�������J�J���%@'��~NܰL� �7��`Lc�D���Lp!>�q_@{\H�*^6��+*�ۅ�,�,���������9�Sy�E+⑦O�l��$H�ܕ��Fh,;��6�kݡ���͚(����J'���$J���}L�P$�k[8�C_�ݰf�'�B���*R]V�9+!h+�$hd�M9�1��f2���}���3N6k�����(8���_*sL�{�g/�Er6���g:�<H��?5)���$�e8�4���z����iz %���6�۪�**�=�UO�t�~σS�J"�F��!���Q%(e[���ە�,��#�
?P5YごHZ�0o|�q`���;�k�Îv�I>�#��Z5s ש\:=���J,s7��.�q
�E1my:�m^�(���*p/�ر<IZ�;�F@�:`[#Z7n2Y����m<3�0�>U�6yc����+��&f��@T��ج����$�J�?��L6r��u4��	/��5�uՈڱ��lHЬ���j����#�A��f�`����c]�}�"�|:/�8>�ڝ&���7V��7Xd��_C.���1݇'c�����Oe>���e�sgv&aQ�R���5t}���'h_J,�����y<{I���O�i*v�(��S�s�@�#&l�(���R�N�&���L��(8�!���v[�߼�~��e���%�a��Pqn[���v:bJ8���M��fB2�"R�"���sU"1�7�dBD�ƗU����$%���_�yh*=\X�RkRs=�o���.���C.��&T����B�=��)�q��{h�R_�+�{Q�$�����~7��%��> �3Ef��ZZh�R��fK��Wԍ��V�.�*��S��j/.�y�'�ߺ�zD>��l޹�מ��GIR{�4�u�k����w�����S��e��m%�9"�&��Q�ѩO;�*�ֹ�;�Y ~`������!IŤ�U�Y��KG���X���q�M&/ gcdg�Z�/�Ҡ�p�O�r�>�^F����2���	ʪX�+�����̈d�(��Pի�>�Ś�W15���]��N�_>B�DZ�s�6��Z%`���O�ƺB�6rG�c�@�V`o��D�������.FC��MZ�bFo]���=�c���p�U�(�a�o�L�Q%(��22���a6𲻪La�/̇3�G!#�<��q�z�/b�_���b1�mTv;�%�m�� 0��p{[?lm��z��(�*ʉ����d+A��?�/r���Q:ګ�6�hS��ބ��{�C!�{!��6�To�����:!�H������H����j����̚=0��YO�3�iT ME*���Ą�ۢi`	� ̦�5���1��X�FOW��4c�ƕ��/�'�XkrL.�e߃zX��hRq����t� [w�4%���W(G,B�%�a�	hN��0��"B2̪���B]`s�����Ǳn��;�_i�5��x�B.'{�Qz3F_�I��\py�����V���	�����!��ɡ�'����{\�M.t�$�N{���癇mmv zw����g��Y9ʚ�څ0Z��D?�`�V��SV�n�|��������2h�$�Oi�c��kB r��ͼ�J���r��bҵ���e����|i�zբ"���Rɴ��tex���b��c�4��¤}�,IB��Mp�©/����b�y����6L��c��*̨�Ak�]`����y�҉��A���]u��ecO����-�]2���i���wǮ�>>���f]$~�r��?��B�($&�y9W��rV�KR�q�J�~|r��tpr�S���~��{Y���߂#�Kh�>7�ۨ�[�`5N�i�Ғ�qL��MR���0�@؉���-��T|���7D��@�=��[�qʎR'����M��@_���8��P�v�?K�-�W˩Q;+�M�VLr簥�3Q��`�(C%L�!��,cm���Z�����Pa�U�N7���%�|�	/��#���D0m���\��ۉAЙ��^�S�ݣX{�oH�[H'��w�=��"s�C�����USz�l�V���+ށ0]J�Q,f�1�TA�t��_-�� WhT�p$m�DOrfoI3��rf�V��Y ӱ��J��8Q_J"P�?��3̑�(���ڍ���� �����H�tˇ?�	@�J�n|:���:<���l3�o�L�r.pof�l���NƟ�p}���a4p��ol�uO܄Z�Y<�=�Y����t5h4:�tK׶i�K��n�>�lvH���~6۲�� )���F&$�*��ɑ���m��ê�3�ZV@'C]��A�0/8����]��;�HP@����KQ�|��ư���\?����H� �?��-�|�f]KB�(n��Fc�_R}������A�& "����sQu�$ �:�����,`�E�ǪyV*m���aeT�S���(.����[���TV6׍M��].��k�&=n�Vc0`}
J*$yE� W����ݽ_���$t��*�L,?�[ξ�HG4�n]<�rw��˔̙�ⓘ���_t�Px���\�/Ρ�qkE�����fԮ��CTτ��d����Q�8�>Io ?F-X�ᣵ5��"eYp��J�Wm�+q��|\Ҟ�3{�Xl^O}���һ�w�y���l<��΄4I�jN��=�	�P �n
���a������q�w���p���j\"���n,��._�f���#��c��^�����v.H	��[��|��o����T����8^7Y��~5���Jz;ZlAN�]qx�P	����.�
.v��t��c��ˮ�Vw�.�;^��exO�Lu`����vVË䢥t��/�S �VH�?Qw������0y:`�8�T��GS��>u��Ơ�y�����6V�t��&2�,�C�F�D�B��2��u�3_6P�FQ����D�k��(:[�ARm�&�v��$u���� �/[9�_�l�p�C��PTR�'����O�y�.ev*<�4��{���@�iIs�t�c�=�� =��Mit�������v�mZ/[��� ����X@���ʁ@¤���`w#U���)�2���4����I7`�TO�$D�O�ܹ/�CS�Zs����עt��D���i�Q����FcѮH:��O�*)�-q�o#'Չ�*9�m\x�c*�mwŸ 	��A*�n����5���t��l����j�ø���ڞdQã��5dG]���PS��c�MX�,4���D�6�I����|�S�<
�FdCe�5���Gf�L�7����S�C��R�i�'��2����R��c�[�hØ,1�,���HD�J��!U>m-N%��%����{Pl�3�d�;�7BH ��V��]:��@nN��5�sB<����� �J��k&��n����!KB���*�F���"FW%&'�hER��d���?#��y�F��ё�~#��k`*Ծ�qdȆJ[�{���y|��6��V�>m�O��D7�>��T>�� T���Q��E%�� ��!�j�c�F��_M/&����\�SX��!�Ђ{q���.#�	����'�Q�U4���I�;mb�!�߳�e �-0��A��YD=�8ܸ���o��y\+ؐO���Ӿz�?��� �^w_˿��I�ܐ5�է�mhILT��%�m"f����#�!��6�󒊡�=��6/_*7���dR� I
�0q�5:A�N�uavБ3O��-~?:�����y�}�dնO��\�/}[��I?פ�s y!�8�A`8Q�[��;M*���㵋u��", �pɓ�G_���JRS�+����Ø��͏t�MK^��Z����]<��F�ŏݿ9�4�Ew��M�~��)��5]$dQ���O6��&��őԸ�<v��&w$�K�KT�2�M���G_�@�$Pdu|e�'&������� �qҥ 7Y	k��2H�F몝�`���"���z\X��ߧ�R(���sZ�� �eS:٠�@K�)
\urE�w��"�;
��	�쳆���_Q����
�|�_M��M�6fB�B+I*���T͟�
�^��j���6$�B.{~V�7�$�p���3ˋP�S��g��T�g4ν��p�h�?���D /uy�Uo�Y;n�q�eS��r̔��������U$.���-݋7�t!��4��@fjI]����Vhʂ���Ҡ�Z�������Z4d	�ӕ4I���:�f��-L�����x�5����شH���i|#+�\nsepP�6��q��O���WH;���d��F�c,e%��v�'�v��-y�I��u"��M�Z+Ka��>1��
XuYNj�g�wy'#U`�R�\e���)�-J��pv��ν�������|���=�b��(K ������8���!�P�"�DFE�nW��
 Q�sşFZ�yџ�e�t:���X�B*Ű�Xlh%�#��7&�Ԝ�j$M�ǝҚX�z7��#��3�5,5D-;�3k��@�ʨ�
��4�!�<��/}�gx��pH���/ӕd�u��-Y��Y+l)?uj�#^ŁȪ��U��Z�����y�:��D�Ƥ�� �G��-;c�w�j�v��`�>��W+��A��*�YQ% ۩��~��f��i���I|%�V��g���H)a���g!���۽�F9~�~�,F�l���MV��W	���ˍ��i��N�RT���B�H��W���6q�JP����/���l&f��(?$��z@�HP��TxF}��cܤ���g��fiDEDc��˫�X�B�п!X���4F��	p����|�e���x�}N�!p'zk믺��2z�j��!M~Q�#�YJOB5sC5�qo�@
y�)"�!T
?m���oi��$�@�����E�6Z�d~�Pl}I�r�(�8��N&� c�e5�2P4W��y�Nh�2�l%���1ډ��ц2}2q͛�4b���˨����o���dg�e�f`!qVn9U�T��N⣄	��6�����c8v=�O>"Ӧ��~��0LN����p�l�CG��Uн��.�DbkiC7)|a�g$	'?_����������w��t--g�e�rx�ݕ�D�2}az"�f�a��jL ��&��c�b!8�DD��w ��o��%]M��f$��3b�ǝ�Y�MB�;�f<�����5��e��{(����Z��`~������Xx��sR*��=9����,N�2��@}qW
/��$�y����X�@��Y��Q�X�U"~
��&�u'W�T����x	�����>��v��R<�!��S,���ǟ]�":��J
�����xM�#I�V�M���M�����H�fJ�.|s�fR�����2 wtG�� �$��9>��k!Ǩb�PV�9�G�����r��4�1S�/�m�"&�zz	t�Q���ll�_]�xk�K=��|m.&|]E3�F���[�k��4�9�T��g
��) �1w�![�F���C����q�)�W7����b� �8���O{�ߏp"��!#3T�6v���Y	zk֝�d
�K����>@}�5�������TT�;�	��uq$uI�pPVײ���6�:���"U�D��|Jv��&��u|�&�������[���U���A�A$�e��7$	�O���0�y;p�m�����o������:�P����y�z|��A�3.�5��Mj)Z�~�}�	0����֞E�:Da�ϔy�3�WØ+����Ŝ<]���y���]���;���7�`�����)�ع�x���ȸ���<g(L�Z"	��u^:�R�<�s��&����.�jN�A������5<�I0�Zi�v�r�r��9:b�ܛ9j�v����N�_z���d_�{�z�" �AB�OmR�m��?X��͒�%���xG6�@���t� jΖґ�p��H��b�m"f��q3�0
���|[���%F�m�2�G8<�s
�!
5��fv�h��B�ռ�
n]������o�ۏ�8x�}NC���}O��0P��������wz�ȷ5:��p_�D2�b���L�CaA��\z��/pr�A�t�@�
G�v�����t?X�m�����J����jQ1�Z5Eb��ܛ��(��ʘ�#�"co}�F�2�`�=�ސE�����Ab;��/��{$�#ZsZ*�Ob����Uj}�)v�?��%�ېA�7b��O��բ���gDR�T�!��2���� 2�@�(N�h�ⱚQft�R�0�1��߳dxL������ ~$6q6�ږ̂z��lV�K{*��5��+H)YW
��
�k�^[��*+�,#�:P+��V�˹���ӷ��#�N��*@�d��ب��BE�����nt2MԭΨ u��u�[���O�d��H�	�)5���KP�^����_~�����|1��!��`?y�9��<����Y�m��~D��¼��A�)�yUK�*�l���8-��!��Tf�#>Eڏ��F�p�����Q\R���v��HM�P����k�49ȁ@q�q����T:�f�ˎX�31>ͽe��"jۚ�SZ>i�zܵ��=��^��%��r�cA������<�Z���A�*��p��6���}�%�b1ǉ� $�_�H�)vߢ�������>�{8	�"�G���,? �����_$�0�*0R�B�~Yˑ&�~|[2�x�MY�	1J��M@U�P��f#t�I���Y*T��~�BY��I�~^�7���v��b5|�e�jT�8o���Dٰj����8deTTx��|�g`��0��Aṑx�d��4S��[�����_u����
g��k�/��I Z}?����)�flm�v$O���f�M� � �����+�2�S9�`��Pf�j_��>�\����Ʉh}��NI �)�����@�7L��(����l`���>�	�[�.�W�eXd�3м�<| :퍑����P��WJJ��4:�f��Œwj �%}xEz[�/��������,C4w��lB�ïV۫6��_����aưߙ[���J�1 �X/&#$8�b�e~�/��2������h�M��"[�WO��!���/�<����)"���D`�"�}��#��ү%��������w����N�t�V?˘�:�WfH\!���l2�pވ^�l���q:�| �D󾋊�a�
�Ɏ�t��o����d��Q.�"Gm��?�h���=�1.��`�,�ӉkXVh%�����q�ڡ�1�1Oxtm� ߣ�~�Aژz;�g����e|`>���ͩ__��
x
� ��D�����$�go#����������d	��k"v����:έ�U��lhKމ��wK�ȵ[�UR��FP�a9������yT��O� i�'Ӹ�h� ��+�i����ܾ��ܵ�I����3����ﾋK>� �&�ߜ�x�����A3���g�����؟ƌV>[�b ��R��R�L�ӻ�P�Z�o�*Es5����#��j��齣�!�Uz�0��|85&	��Y$�&c�P?�>����m���'N�=���;��Eb"�r��FA��m���&K\��Q^T�+}""��i�@Np*9¤�n3��!�E/�y[��Y��<l��ۜ�6�͊���ͭ;y���)�Ι��e�T��n�v�R�(9+Ь�I�R$P��__�����H��SR�\��M4��%��d�b����hj��S^k��9�J�G����F���_��(A"B8T�WI�4�� ��g	x�b/MVL`޵mT�)��,�a&HÝ&��h�GR|����M�w��w�)dn�F�� J��c�؝�TC�3!�-�{��������:�BY:d��5L���f���Dv��Nӯ�Dz8E���ts��r<3�u0�v���d\kd�W�}���pSw��Nb�x��D?.�d�΍�2�>�~A,CE��x��wU�qT���ǜ%+��m :���Ч�92�P��������
 �	e�����Աu
S��⟂�_�S=�9jR3��Vs������ޗ���f8q�P�ǙMϨ����jۇ�UbcVY+�	�l��`�
>~�gCpC������Aߐ���ǹ�,��WFǴ��G�e/`r+3k�9ӕ������e;i]�)V4�k]HA1��IO\ǧ��Z{�h^-�����-�RlO�z^��z�%��S�>���X�RS���%�Wd����4ᰡ76Ƶ�Ӏ�� �M�B���%����y�j�e��vS�6��)��y[����6�p�~�T���G9�=+���/Aw�R�]L(t��q.FjXO�t�x?b�{�Q�?-б�����V)����l���Ti�t����ы�X~'�o4AN̂��{�u��=�x#>`���X�~7;ti���4t�w[�wp��ҎsDV ��������G��
S:1�WR�F�~�$E�(����qX~�'������Z�j�w�M��\�M�xA�">�G3��CT��\\�gQf��$�$b��둾�����#+�U�R�/U ����ez04��T4̅kq���� �Q�����F���[��C(�=�;:���I�Ӫ�^/�-���4����v��y�y�e#�[V&Ȋ��$��zn�*���#�V-fac ��Lm�K�<"�g���Yşߋ�q���0��49������^��2�LiR� ì>�B���\��4=r^'z�����w.�!���jc�)?�r��9�("5�����cU�H#Ab������D�S��@_�����[����((t$Ao��,�)�o !륌 ��!}gK�>�T]�D{�<,�
؞���0�x��,�@���T���ī�X�s1W���%�!� 
;LՊ/�B�J��}��MU�{:�s�������Mn�����8�l�+�B﷗���Ӈ�6ȉ��4!tp9̖���J�h<�0�5�)�G�J$�n���s
�Q��N�z�͘��b6S�6!��H��W@�5�6O���x~Ф_
~�Yޤ�n�6�����yԡl� _�g6R��N	De|4'��~���wx�6k�p1Vj��#b��Nem�J< ��:��������`��q���l�X�Oao�`��UJ	�:��{�C���%�\Y@d��Ԑ&=a�:\�JK�����N�Uc��~x 0�y��4�p�; �H� 4%�<I|� ���t=����c��I�Oߢ�W�0���v�(jkn�(Y�z1���[�|�q�T��[���\l(����@S����̌�3�z���z���R�gq��1�ٚIU�p�\�Ze��Q��d_�;��
+�g���IK:��O��8�\�s1��:�7]8������t�X�R��SH�9��bck.#�&y� 7�?������S,2��J	 ����&�����W�,�p�����q���/�ZP��R7JؗSZu���q���仞�$R;e���5<�]�̛�J	��߼��-����"ťEa6�V��	&��L�p�p�V�G�⭘�
m��+�H�I^�:�	{�5(��Z#��X�S.*�吓$���L�7�[��ܭ��c&�!_��L�d�*',�Q"���f�r�R�Ԯ��O\�q7,�I{6�����<�D�_";��G�t�X�23f��w�}��D�-�G:�-k���X�SϾ�?%N��d�����3�ыkP��[*��8`d'G���`����f�'7��೤�,�5��g/�����ܹxWS�T�2��%�[��H��6���p'\��T�.\X�Kkx����96jw�>�����Ƭ�h����3\o�,�������Ml�)����hm���t��=�~_*؛n@i���% �vB�;��9N�8N<7���إY$ojS������t_к�z�f�4ޗ�팭,u����������6R�J�U�e���D�Ԡ�É�HP��7D�{�K�Ï�ћ��pd�|��٬*2����I�2~޹��V��.�[�.F^y�z�u��T����0'*X"8�u}�Eܬ8�fzg�ߒ���Vni?y`�-KM���ٍ��~��П���A.@���(�-uL +wdQ����]b�^O�@Ԕg��Y0`Y�C�B��;8�H^��B��	�d�ꯉ7���>;_�H[�	�s��`���_2S!�����b�B�&�|B�6�ɿ�M�[y.A�i/ϧN"�_�"D��d7�TNĥ8#|��ߩ1�um�SQ���07(⤁_�����y;W�Jm�9>�����:bBM�U���MB�*&p�:��f�6�x�j�{�M���*������=�B�S�xQ�(ic��`\t�����5y�����^��J�~V�q���=�?[��%�dL����&���O�W\w��^9剐��Ճ�i.��=V��=��Ԑ(�8nLN?7�;�-���ԧ4G��q@;KJ.��,ç!m���v�s��ϝ%�3H0��~�L������*���;�X��f�z	�W8㾘lq-4�J���#,�}&J�A`����*��eS�]Y�/a��⧁���ӡ��ړ��ui��e:���������V��[�Г$>��K�؟�>��,�3i��x����>��B1��c�r�(��0�Wφ��hk1]{؏kCy\�su��<��u�,����J�O��<K�G86{��:�(��f�!���`��n,)gN��A\�?4��)H?R�m44��ޏ�N��%�_������y��U�	,��J�+̂Ѡ�C���z�B�������lM�&��������uJ�ң�V�>ak��a���!,ΈBFV��	�!��VoҬ��W�,�X�~�L��금\[j�L���x��%m�䂠��o���
(a,6'��C��<FH�P�ڍ�� Q�c%���፴� ���x��XH�<����H�O���a�L�r��� �\t�KЀ�~Ha�y�B�Û�);m��V=�;W&W�(��[r�dВ�RTa%YT2$Ψ��bt��6���𼓢����-}�_h�v���݂@W� .��.GK:�ZK<�F�ҍX�RT+�v�����\Y�xT�Q(E=�w��#���Q�,6���� �J ��=�̵��;�s�֘w�a9��p�=�k=Z���|�JH�O���Q|L5ѧ���2i:
"�r))8���F���G<K�,��]��	Y�ڵ��X��֚��`�wä>��}�	�@���?���6�����\��vypU��`��C�P����N��?S�=���_�g��hF��ATY=��}]���.��+���� '�����J�7��i�J7k�zD�-a�~���&�3�8��k��d�S�0ʉ�4��Lh'�a����K����-�mb4,��Lnݤ���K"H�E�k���h=* v��ƚ�tr�,�Ƭ
t[��5u��%��M��e��Pw��r��!͛���9nF��At)M��ܚ�Y�2=NX?��~�q�~ȅ������@��!"�{�Sr�HUV乇�}^����wK�\�����;V\#�{��i�M{Z�=���z��5���vQ�1�-a�Ms���WR���i^���o&�DG@��������XŪzP��H�-V�k�1��|�K �{���`Eu�[���'dp*MU~�y�{'���:Iq����ª�@,�3�C�w��$�>��-�?<�����B����\z-p�������g�'#����ݮ��4�d��&Z�S�3v/��\����v� ��͖l�ʣh-0Y͑�?��_�"N�<u�%]�2ʉb�\[ƶD�AF</"\{��v#{_.�/�9�=����Z�.��C�2m� ? +�������`��r ZR��M��~I�Қ,=�ۜ?%���:e��)�$��.��<#>�]�-������c�L]�t�=h�쮅q? ��}c��Ʀ��k�B!S�!Z���=W6Ň����tX-��e�XQbJ�Ă�`�#�!�I!�䓠���b����Vx�l{�� ��FD'�5�E[�H�3�5���h��Tn|OlA��)7�j|�C+� V�{:��_8�R�6'�l�B^�V`�G�Fk�v�əS�v���ٔʹ�Io�����ֵ��}r���,l�U�1B��u+�ͣ$��=���iw�%$�R: .��R��7.\T�>y'VHP��	vS���&z u�j����oB�c�_�&m%�k�k!d�ǌ�.O*�.ۛ_Ʉ)T��0;�u��+�.<6M�ڋ���|�%#`ؐ��o�� )��Bɘ	� O��K��s.�f�8>*p:u& V�jp�#�.Z��  ��CpU���Ra�?/�����1(�0��͎�k'�9|��1�ii�$��ᡈB.�q� dY]�J�^��~3����D?c�O6Rc��Vӭ<0c�Dac~R����"�`;A��+���*`�Wy���ǒ�p� Q�"�^':=f��9%4�\?v��\�����0ȟ9��������v����7���&�?16�'�BB��;�)�Р�v<�օ�Wc���^�Q�W�xN�%rO�H9�Jr"{��-~�idӳ��l��A>�9��]��(�4%5�qk3��;7.��u<�1���=B\�spr0K��"�L���Z�<d�,�]��*BNI&�i$V�eM�V�[��!�(Ǎ�Q�-3���&1����� ��'Ha�>����2>}2*��)G|�i)��;}��,��D{�>?}�_�J�A��a
�>��N_,!k=̭�'$b{~��T�c��2�H�[#Qs8��rJ�b2wx�X�)ބ�����˅���B�hY�)��g������:U�T��Ї�3J}�qwՅ�C���P��?�ڗ+	dL	E�%�e7�c�}�.�����+g3{��xJ�Z�C��9F�o���W��p�b���=�gI��I������Oz�i�˰"Sr�ԣ�}o$C Ч�{Й�	]����v>�c���v�8���_?��ĭܺ�k�	%��Cӷ� o�RH�����=Yo�}�\꩔ـU�����y]���u�{/�+ �'1��=&>
�b��շ	e�f����mB�m�$��ب��8����z��@��CH#�J�Y8�e��h^�Y������dSd��+��艻6~�dYk�z$��gq���*	D����3��?�  ��Ԟ�V<�u6��W�@?I�mJ���}����
��x��"��R�F�ָ9#��[L0��5amSK7����I�d�N�?����P�0��zwO��`+0�~���&ӚR�V+~UT�}-��A�O�"hO��f��g��DM��Z�.�?Q�ʑ~��ƭ�I�(���,��)�Z����8�RJ�k/S���	d�$���h(m G[���dMTyz:}ڡFӤ�Ở2C͂�K+~�<������8V<�fyB"DHMc��Sc}��p"8jH�9��Y��2����A80�|Cf��7�y���߶�	��[U�1�ގ����*�3`�E5��Н��+��4��a�#��h���;ȃ�%i#��FWs���W�|K��,��P	<�nj��#��h���bG�Qa��@�L��+�6�I�M�Y�wE%ܓ�����.���%�x訁}�}�B]rY��E��$"��Vה�Y.np���_�\[��d��-���n��)��$��q%x���h�ڕx��	7��j5ʅ���Ѷ�>�Z�É�s�i	��ͯ��G�U�R��ׅK:9�7�(����W3��p��w��~I8�O�������L@+$�|8FU3������mͣ�!��w?�~�D-hll~I����&\Q6����
�A1Nx4#8�trF�PT�q�����Mg��<�*�(v�u
x`U�GJ�UX���Oۦ�r��RNÂ=�|��췑�޼�V��?���U�����,J�|:<�1�5��n�V'7�	�����O.qН�o��[���Z�;��`���~�%;�١R��۷ON G�����Ȼ�@����l
R&�Ի�,;��ԍ�~��ϟ�n<Z�AH��v�{-~��V�a�}�!mI���E��>n�Γ������X�>�����lbQ������/��h9�9!Q��?&+�X�0��M�MC�U��Z�>��c���y�  H��v�Շ �#�k<5�޶a?S�Kv�_�9P�"ىh�j,�]��~4[c��AIC
�����xF�Pw��o�٧i���F)�p�q�y�TW�m�@�M(�y�|[o��-��a�yXp��D��2Aá�zC�B�ޠ��y;��#VG���R=a�U�"��ݾ�%�]"�0I�k!��l��W�?�j���2���+c�(��@�"�"��4�'u���́p�.�L|��Y�@���m��E՗�T	\=�J��DX/_Ȇ���*����տ%	U�W�R����%�0&K�RW��wg>��!˛0��˵��V�a����F���6F���f0 ���#$An��b��]�8�4s��o[1t�'��<i �ڞ�Hؙ�����W�HO�}<0������E9b��j`�Q
[�k�J��g�J0�ZPT��b�\T(��!��ha����9��B,��Wbf�)<i�(���'75y�"Ƃ��m�
Ӵ-�.z�d��L��t��ddh����\h�/�^���c$F(�ű!0)r0t�f�$����v��_��}��/2���8��g}���ˢ|�nd3�dp�h��FWԩ}*�[��"�Z�}��%��㮖�	��a�e�<Y�����dt,���t2�v܊_�W�7W���x��n�q2����?<��-���A 2�௠
��7�2�g˳�ӧ�V�}+���A:���E�Xc�RB�*Θ�>Q��&��rWs�p#�5�#2�z�JA�_%L����*	�>R����K:�m����8�BRL!~�XO��a��*n�ܐ�	l�7t:i6z��_�(X�Ô�\�m���6^�қ�=�?�[�TN)v��O��NɁ�юb�u:��p�#��]���h�0�9�&��1�oYR�q��m�41�ȏ3+�)�2|(r�0�sd]�L\y�15�����y��~���5�C�˂~��<�҆c	����Үu/5>�z����|��u-�E�M稩�v�GJt^fM�o���+wR�bf���$,��Ρ���^���&�(~�e����C�J&�1����'C@�!r�J[/��X��y��*egWS���rn�z����X@�ߐ�N�#F�uПn�=6rh���{&�� O6�Cȍf�����a�iw�w����w��$��R��S���9'��9�����'���A����ހ��ԙڑ��liR���Ħ�/�?��7n���G��4�p�^�P��r���LQB�n�Wh���\��Q�Ӆ��oHS�w�%#v�"��F�5Z������6��R̛�{�(d��H�W�=A��,t�(_�v�
�w%U�f;F�z_�V� -Zt��	��.�adMQ���%r>�L��K��
r�?C� ����Fzx���!(��t	���=d�{��JQ�g��s.:0-6��Bj�X��(�)I �s�Ѓ'���\��=��}��@�KҊ�a�2ثZ	Ue���wi
nh7��K�{D��FN�A",��:��a@�;�΂��R4N�i<b7�&ե�j,����������d�!�zg�7ہ�cw�	f�4�*,�P]� �O���G�b{����f��4�s�ɼ���U)����:'q�L�|�r�?�:�/�yÒ�U	+�����Rb���}���\ �@X@��+��D3c���۸��T��#�S*v�{.r]|�_v���X�+?W��F+�_�5}w����jm@���R��lߋ�{���d���W��U�ȓh[��<I��|=ͨS9P={^��X*s�������8���Ę@��{
�o%vw1�r�;�n �pz8<�U�(���V*bE��9f�Ēo�.������P�dNBC���D���U���^p��{�~P�8)ٿT]p�9`U���ʑ��db5�=ݮ3��Y��8��|��s~x��q�y`~��3�L8�?/����mߏv%�R��`����0�i�����@���R!іե���X�Y���
Ο�ű�X�1�aꩈ��'�S��a��Fr>�z���ڿ!_��M�=>��]�%�*��A�=���ns��y%��G#J+r�'�O,���/��G���l1P�+�GTۖ�@P�$ht�E�$���M���ԸL�`�m;�N�WM,���Aՠ ^��D��ُ�d54�[�v���lZ�e[�q[t����\A������?�v�X�cxk������-l��ç��Lג��Y���<��+�a��Fߜcw�����%���2�{����3�-���־nN�u�6[�Opkc�-kڍ`�U�c�B�V<pI:*g�@��P��#��&�Oqy2\=?����R���/�R��S��3#����k3OT��Y�*�1*��z�"͔as�mTt)Z8<GӦ%Ԧ6����#X��"	�+�c�	)k\�f��}�ė�l<q����<���I�=�$�fޱ�6k(�q��W��y�%��x�QQ������p?_bK6d����j�&"�Z '�}�*Dɑ��(�֜���r�O�2�^��p��m��j�D&��^|��Ii# �c1fp����G��L=�����O(N����d�NȤQҡ�]K�����>���ZM\~�fx"J@lx�$��H+`���ɄQ(<:-�˞	��aM}��~o������}T|q\YW�]�9�n�33�$EFj~[譵��d��*��5'�O�HN���\��f�Wy���y�����C��}�W�uF~A
sͨ�rD������&~�@�7zL��ۋ�	t���H�7A�
��.q��@�k>�'�p���۠��D�"�{+�D6�#{4�@e/9�8I-(D�?��p"L�9]7/
�ŖKLP�[��GNt)���	߭#Qp�����"X>#�>/�����S^,��D&3�z�/q�A�������̰��Z�Q���K�N
�8�g�k��r��*��u��,WO�	�м�`.�p�Pv�[�}~�n�@(1f;��� &��]t�%ւч�߆z��(`�oY�����j(���R̅	ȩMW�?BԂ�\>��Mޮ���wy�v�p����_�3���O��i�������v ι�B���@gz��S[�����R���
��m�F���tH���W�=������R�{iܨ���h�@� ���1��js�|́S�F�y-���`,����[��,�˃J����� ,��'��(�+�#bΆ��%���o\�LXY��s3���Wl4��W�m��vR^�mU�}��F.M���v�p
�����|�0{��r12԰�n!��ى�f�4�C��êܮ\�|V�����(gs���_ʿ��h���/��b��U�@�q���k�&����E�<����s������|"�r
{�fzIuB����˙�ǋۥ�`K+�?�(\��X0mGm8���Kfu
��&{s�m��m�h)���pRfqv��D;��|��ɦd8Լ c����({� �lD3���B�p���r���y
��&��9���i� ;-`왉�Qz���|���v�Ϙ�.]��>>�	�c	G����\���H�Gz���}��� t�K7'z-t������+��c�P�"��{�W�n��vr��S)�!���_`,�dR�w��ՠ�-�+���M���Y��
0�b��n���|����z��e�S�M3	�A+*Nn�M��.6q��e�|��l����c��Y�i�[� �LW�2���QJ\I-d
T��đ���Ћz
���fc�.Ǻ�P�ۙ�#�)awfo���!k͚���h�@�b�?7C����.�2"��n�i
��~��\r�!E��1ʜ������qO?��9>Kߴk�á��d�X�	i$4��Ff�;fm������tJS'4�0q��F��KnǺm�g����	��Ã8�����ҍw��T���xy�/�������QɚC��ۀ³�Ms�y�������Lij9xLK��D�QB�B��0��׆�.�胺��1	�d=@��<�wn"�±�
Ϙ��Sz�LWk��SoD{Na/q�v�5��4H�^��,��s)���)�|���E��o/O���l��0�(%���n��9:�ˣ
�d�2�����P��f%���D8&@�ʏ���x�r~�S�Ck��=�[�y���iC��Rs�O�_���Z0�+\�7�n�!1s+8�Û@~4��Q��|��d�/>�:"����z�8�YW�+7��F)�~�JPW����KEA��ɹ�x�r�K�u��k0�R�xù�B��$�x!�8e/J��c���u�cx0�vR�K���_��=X�%rڍnԬK����|��J#��jA0��l�o���}ԍ�M�;������=�˯(n�ʠ�`WI��y^4n�6�Y�|�/���ǟ��P�d���2�ג��ǎn@�]~���l�tX���ͧ>ar7�l?��B�����c�V uE �Ψ_�!^�K�P9���������I~����i�
b�eu��Fi�p2A�#u��
uC��S�����T��#�@�
cT���t	r�NM�)U�hV���슊�;�O^�@�{S-R���o�n�&V�?�C	f�K�|���w�7|�˛�����N��S�,���AJH�=2C�U�LXN#��-՟cC�K���>;��?����i^,f�� .r���ʧ+N��؞wk��{�{\�Fcl�}��WBT�(�e}�e���r_6q�t�U�!����)�c��ʉ�K޾�Mw�$�����k8���{�39���i<�ϴ8M����#�)�8Ya�M�{��G'Տw��Y��G��ݕ��N�"B�C�1�EX��Dϼ��S~w]��3���O�����T��c�Ϧ�`bؓ>@j����I���WeL��	]��F?,�)�|��� BR�kl�3�K�������}���m}'n�������-�S;C�zR�,�ȯ</�JhW���
Z6�"l�/-@�/�Ҁ�D�II�4%-g"��Ԧ�s�tW���)>Ov��0��A�o׾��z����F���qP�s�VR�d?��f8%\���8d�@����?���j�4:�,Z@S��j�4V�('�26
��~	��^�ƂJ Epxq�@Yq�eiA����5�pc�h�]��Js����Lv��}����7��Iq���E��$�m�"U#k����.�:p���-�#���Qb�㭻Q�d�?�4�z�K?��S;+�Y�tf�̦�3K�a�,��>��ЇH�w�euNM��Z!6v��b����i��=�O�����{��!|KB��}q��jُſ�u�a�Ģ�׫�+׹�CS�<%�����ҍ<�x��%�iی�>�dZb�R���[�r�m�M��W�D����H��n!�����>���W�U������셢� ��/6=;��}�T�ȅ,%/1��V��b����U�"l�`=�"A#�7M�8ݴ�2�<#;X�#~�����s�MxDU�E;�)t��-w�cM�wԶ�_~�M�'@����Yw&��`���z����1�P��g��@rs�����IQ�I!������u��s���=���֥
SG(T��pAϠ����?�r�js�0�ĞjU���;��m�����&"&Ir����ׅ���-�Z���.�c#�6��B��� ���
�op�K7B�>�C618��hܧy�ݏ�x<�R�$|.4����/����ڻL�;6�O+ɊQ��8��y:'�:ӈv�,���)�Ő���"�K����� �6�}g��Gw|��@&��e���׋��%���h�S���&mMEӐ[l[p���M���M�}���Ÿ���#�%>�H�d)N����.��8&�=���SON-Ә�rB� ���;ff�_���SI\�C����������u<Ndc�?���D��:~����>�	�¿+��XW*�׹��L��	���+>��9���}<����U	[��[H��3k3_w�dQ�>����
����*�uT��̈́63����&�M�|�]a�ms����M)�`�ݶ_n�r�Q=�R����u�	�\]��8F���՘�m�����b-��D�9��X_��lu�T��\��,p��r�V9b`	�q)���A|,�'�Ӛ���<4O�[��nLݏ�d�a�k���Z�!USj�9 2^P��6�r�?�_��82��3N���QX��9��OZn�U��tJE� y������0�v>����*܁�2k��&�\����H��&�HL��
���J&��f /B�_�݋L(���KR���K���S[�J7����s�A�*=Ks6�����X�4��Q&jpd�77<�ݽCK7�-k%���锪T��]Ȼ��˽�Ө�{"�n���[��?-�H޺�q��X�Ad���4����*�n\����c�����+$�t��`��"�f��#ӧ`����ɋ��:r�U��L]�@!�U* ��V�L������;P�����k�QW��%��!�W*�뮬)s��]��A����.�*W�r����7ݑ��̽�R����l�K+��q��/��e��`�-�u��a��(}lۘ_���S����xƓv���]Y�oM�/P�/��u}o�#g�g�z<�f�k-����1��E���52���t�[���Al��"�hY��e��3��Jh�
5G
���]�z�d�r�3�l8"_V�F�z8�����Q�f%e�$����O����ϭܤiD#L6�+2���U��7��2�]���F�X��<��D#���V`�G�	�]���,@s��.�*���;7���r��)G���fe�Ѡc�����,0E�y��ҡ4�9�Rmr?yu������q�3�[��])o,��T�
�1>����FP"QT쳷<�-�S� ����s�M�l�ʘ;�_��������_"5
��x��?;��N����/�GιK@e���=]�X�7Gdp��ː�:�i=��#N�:;4���[��ʻ0��cZU��Jy�E��fϊ���o|�I�M�rbx����}����i�XG�7�s�}_5�QݟJ6%�,C"pa�M�j�'����@R���ք[�*�arA
I������>!�В�	qo��,j� \:_�	�VM������0����lHtB��������LPo��_Op�-�BY
_Ye�|�C��퍪H�;pn���ip�u�Ĥ!80�}����BkF@�%Hȥ��(��؊#��da�7�ˤO�A̍���%v���mT�ٰ{�A	�H��� �PH�f��E�I�E#��D>�e�c�HE)�olHԘC�������m0�}��H�f]/tShP���n�BW�k��t)�f�%��B��,a �m;�����]�I� 7��:�K�a'�D�aY��SZ^~��!�����hX��=�,�j,�dgX�B7��H޲	�S]Ԁ�k�-�1
Χ��<
&��t�G�(�H.�������?�Ÿ_"e��{2ڸQ.��s#-�QB���TZQ���_�Ya��.R�vb�y���b�C3�3���}��(�t��6x{R䙛�_�!��c����և�%Zo��f���a�%J�bČd�EkCyF��p��G/����}:l؎E&����ׂ�d�B�/�6��܋�A)/33�ʈ��5��*��3�"��B��L���ƪ��?*!�6��ّ��,�Q�i������<���/��.�	Po��R�y����KNQ!(��OL��(i�k{L�����<Y��NR��H��hn�N2�a�b>6��{l�ҽ/±SJ� u8@�%��N3���^�ljk�9��b:k��d�V��2�r�܏UE��fy.�U���rZ,O�EX��gބ���J������S(0�E⊏ z�a>�/H?�G�����S��/ IKŜ=2�j�h�NLAx	Y��+�pb��dA'Qi�%���c����0c���(3$�,������ȢƟ�`m+gS.�����z����-�wDI����*z; ��>��8q�N3r���������|P�Tsn٫H\��a��+:�iD2��.��ΆY�$����O#yk��4$���=��f�~7:[(�JF �����S��'vN�vv�.��&�P�B����{n$Ce�l�[����+ڠ���A�c��ի�E���Q���w�1�g�,���C�n�~P��i�@��
7K�C����"�s�%�7r��ӳt9Kp�WbLif��	��x࠺�X��!�v"��"��?��p�h�	�Z��������o؛AK��D��0���"*�1��Cf��0TjVЕ�f��@�np�@�F\�[m�P�=��7#�~����}��~ފ�xy�����q�pѡQ=��y����h�X�#`�G�z�3��J��!\���PX��Y}03`㋽�G��|e��,��JȬ�ӻr+�0<��I���#���uO$�4���Ճ��&G���)"������jm�IC�ۅ�wnԇF�,F\�	��.j
`��9ڃ�� of��+��<{=��/ t¶����EXA����%�At� $���]� hB��iy�e*v���D����-P�dG��B��Z$,tE����'�Bwdv�||3�|�E�G+�dRF�W�EI����zJ���c����H|L�<XO9�f��t�p��Ϳy�A�q���%f�����'6zD�Z�1R#q��M�Z��q� �����UD+S�
q��|,��R�d6o_֣�fOOĨB*"�� r<�9j�eH�c�y��c3"q7�R�ݔ�}6٘A��g����A(��u��GP������zφ������ =R�X�U���3���Ζ��*h��^T��s"����áנeW����� D���55*_h���׺`�-#�\K��{��c��2h�28$��B�Q�����vM'%���E# WA�T�����c�$�T�]��؂#WV��OS�kw\��v+�k��wp�4=�Z0#����dۭ��u�Zq�u���Q,�E�F�fm�8�v��/^����~%��"Rs����"�,�j]���I���\�e4M`�,f^�O�0/m��g��Y��T��*�����^��h|i���{�5_;�%�h�T
��?��4�;Q���kRw$�s��6�u���V$_���g�Z���	m�Z7}s�w�#���s^�ʤ+Ae��O�K9dFㇿ�	@�*G>�2���:�M�v�x��p�
&te��=��~-]O%1�g��b����H��c*��E�ӭR����h	�
��x>�,V-4bq�M�Ɣ�uZ�;�u�����hO,P����¥b�AsR3�hc�w~��+���ҷn��@��6h="�����$��[�:��9'+U��~µ�X��
�E�l@�\�y��@��4�X�)��(�!����b{��'3��9U����oR��b�ݍ��c %���,��#�K��,���ys0�A|����C'�&�:�5Q�"�>{.�E2�d�i�������M��3�i�g�*��`�S�P�uc��Zz[�r9&��2�ɗ���[�e��ym�pc%�e5ڜ�W�bm�N��Z(�/���\�B����9fè)94�h��Ni+(��pN��B���^>�a7#چ[�b�����`U�W�]ŢrO �8,�S��f�f��G]��;8��?���oT����9�D�֤.3G��-�+��id�w�Ċ���±M_���@K���C�TfV�k�#_����U,Lы�F�z!�=���y��1۠;��-lx�����T� �y�l�2ib?C!l7���b$�&�-yАk�!AZ��4��b��ʢ������۠�Z�!w�^^7=aC_��Pr5���7�V���gݡ����E;hp��rƌ�D�L�Z�/V.�����!V�`moс z߹�PtM��K"�z��i?Gk�Q5B��Sj'���)
��Ų��G��+#��v�[�!��ρ^���A�1A��Ioz����=���W����s���e$�u� �E������2������� �<�:)���-d\%�t���i�$pJ����}�����i�LՔlޏu�S5�}����)��$4A����A��Z���0ؓJ���|P��r3�h}�Kϔ��į�I�ؒ��fNP�.�F<,�`D�d��d1�#�
.l��p_�m�a� ��jR^$N��h���66�˻��{q'\)k�IWD����ɌhN��Ev{�v��zV{�`�X��X/:��:�Fa�L�3e<�|����B)�c���o��D&��Km̀g])q�.h��]�bc���i���]3��v���*�Pq#�#�d&�L0�<u��QL��^��-
F6�A����_����s�����&��	�~7_�5��e������+"*�X���ꔉ�!�Wh.> ��|O����,�ә���K(=_`�m���Ҵ0����R@�D8ӫ�D�K�렲�(���%�%%v�]q$����0��.���9}Q��@L.��)��$c@� =�wJJd��n�a}��bl��OTC~W��{Vt�5Q��tĜ[	���7����}*YJb!P�B=�����V!��YV�pM�&SH4J�~e�h����%A��R�ئf�B;��vj09^g�jg�Jn	ߔb,�����|n�0�z+0B#Lׯִ��c��E���ym΅�`�Ui�<mc����%�~<�P������n�+8Y���c쌾sS��@0^~����Z�N�u�F�\ ��,��؏k�D�@�ؾ
�� �#iG�7Y�܉-�{���T)��v]���%5�0�}�&��Z#�w�Q��馛V��%<����Ƶ�<�W���hVv�>� U#{�N�Af���R������S0�&�l��*A��ީ�4lN^�:�#�
u��PDƾ%���L�0���Xҝ�ى��U�%�KI�Tef.��oZWi �,AuW�j�މ�S.��$+�ܒ�i�5D{��f݆�Y��gC.�w��%�V���H[P��{M����5�F��%"�V-a)�i;��)���E��Pk��mfm��iF�ڒ��X�o�MU+A:�������@Ɓc�S�u�4�_�q�j;���*ʁ�R���nGH�>>�O�2����|�݆X�?#�^�S`u,g�B���`���ζ8���j|��\s��mǉ�`�K���1�IL|��*���E#�Q ���a5�8��z&>�1�k��j�A���O��z�MD	#��2��^y���`��߸�0�!��}�y�S��6�-�v^J�|��8���tE�`�@~�J���� �S"�&�O�7��a��S��Rf���us&Mi���#�Z��;Ѱ�}�)�43v����kΓپ`�s��G#D��Θ�\H_���c�Z^�D1��>���.����֋�OM���r�rg �`�jו��L���)�e�h%��~�dJuPW�Ui6�@=��L���c+���v���t�W*�y	�f�mSh8`;�[�Z�"�頔�q����^"�26�7V��y�����a
ӏ�޹���o����7t��V��fҼ�Z��6�￩��DP��j'E��%�[v�b�񼰿K�:թ\�v6y'�`�"]��ʿg����@2��>�նw�S�{����&��n���Ƕ���a�҉	ٜĄ��%��56Ln�]��Χj���syc+��Zxr8_��sÜ�84�͔8]���-�\�6��hݶ�-{�{�J��׻Jr�8�5��@�i �_?����P��� ��u!
��F'�,3&D�bAemz�qWC���%��>�|M�p�"Yk�Q�R����|���B4ͫ�G8P�&��n&�:}qT��Q�F��q�������k�4g�
U6�]"w�6�,{������N0�N�s�E%��p	�K�;9Y�_>+�4�����&����}�"5�Ds�|��E$��D�*f]1��vdA��j��������Th�T�_.3�Q��P�v�͂�-��9͘����B�k�"�0���|wmNW$9�vg�҂��g��p ����hH�jk٩��H���B�wu�s$N�0��i6�����V�"�X��t,[���qW]�(��E���	��E�([z?>��ӆ�V+x�垶X�u%S�te$:蜥I��6��Wf���	O�VQpL�L ��cb���77���%�6H-��J��V� ���weM\�+�|Y|���@�R�����E��N��p&*�e`�|�'���Ű�8��{q�ցn>إ�9��� 1����G`�픴�Zͨ�=e���'��	�A�O��c��g#KO2�ū�O�&�w�ڎ��tC�A�Y�!G�D���4�1
��U����j�����n�*CL���fݻD�T����ɪ����v�tO�SH�vz]z���:S��f�4��Np.˚E�������rZ}b���\S�����o�Gh�R�),W1�I��ʞ��Q>�p�&e�L�E� Lu�爌n)G��b�$���G�Rv4	�`>��m�$|YX%N& 3_h��ۋJwq�w��.��j�Si�q❖7���1�_H� �?����.�7��B�ܕ:^�WM2sȍ�����R�&�"&n'q�Q�Uq͹����=��Ct�b���v�0��t�-������[�6���cS)�vi�(ْ	�X���0":w���F�C��܄wd�ȝZ/þ�`���\AWcM��='��Z�=�+h�u6s����LE�����Sh8̸��C����Ov!m��H��q����>���`
|3�����vE�ݧ�b<ub�q筭�[mkS1�wy
'x̩�|bB���R�Ғ\�1b�C���z��M����K�]�F/�;P�օ�˛��������`���I|BEOd �VV��Ly�fK�$7�����zY�]#�pq/��+ȵ[v�>KT�2vY��~����d���H�EK���w�>��|.�v�z{WSi��IԐ�8�r�9���.��@j7Ӟ;�b�S��J�ԙ\��}���Ia3��8W:j�	,D����6�Y�{���B3C���y�4��p�l��iz�s�f�r�Rl��hD�*<Qj܊{S`j�A�w�$�eQa�͔+�l�u�$E�_"�����(<���w��b�Գi���)oyU���,DP-���e',�1XNQ�y'$��p�v���V9��!w0$��ģEx�Ŵ�=�z.hPw7��D�fU��\���'Q?�
E�
	���6 ?c{�"�=�;�G%�Ѝe?��c$'��.�_��6}���{�ԙ��y�9��1Y�=J�AL���n9#�I����kpʊV�n���1םf� N]��^
����-\�U����th�����k�RѸ�r�[M_SL��/���o$�y��\�.bU%�]���^g^�\�{棏��Z&�4����J`&B7�[���s c*d9ƫ��ّ��y<�b�-Ą��u;��������[�w��Ç�l�@�TgL44����l--�!���g+n�f^֭�l~
��Up��x�bX�<Dr�{�+Σ�8c&���Ѻ��F����������{Yp�ez��@�m�*��}
Ǘ1�n8����yqV_�iù c�ETL}0%"$M@PG���֨����x�l�� ;0nb�ŌK�����.�w���\?T�4!�WSw�s�����Pa��n�o�$�N�,�`�-���f���U��
Z����
9T�Z�.)�q���}D��+�´�������K����}��yR�������ú/Y��?DV�
V��M��
AB��<]���,�@��ni>wW���l9�v��Q��r��H�DL8�����A.쐻� ;��;�^Qp�����W[rq
�%ћb�A����L��G�&��FR#8ڀ{��2��1����L+dݨ�?ű�18.�s1j^�ᦣZtJ'%	4��V$|&�z�K�P���?��i�(��[����#�;�b*�^��:T��B1e<"�7*▅K�t��=�3��m�DSRQ $3ְ�	����5�5�� C��Uʠ#<-�0�����%���	�Y�5/�Yx�QPԾ�ɡ��.�	I�9c��-r�:�'y��r���ډ�2�s4sQy~�ЂqC�G���\֞�nt����k��д���:�i�0	juݕrg��vA�&��,�зh�g����4�
˽��	C�`��ϱ$b�s���u�)'��Ф�L�W+�h��`��e�m�A�6VPAA��9��S�\1��`$��nl�/�\��,��ܞW���i�#��go7&�细f�<�n�1�##Rb�5�ΐ�%B{i��^d��5wИ�\��S�7�ΐ�S_��"ۤ��"/���:g�r(	�?��J�9��8�p���ju���*6��]��G�|�މ��a"��3�)��r1�[X ��' es���Hi?/��]�9&T:�Vo�dr?�35��cWLq��Z���i�FDU_�m*,�Մ�T&��z&�9	�\�jT���3�5�0kk>pÅ��������J+��T3���g
Ѱ��Г�7�*�b�~e��<���YV ����w�J���-s��6�bvS�m��8�/�u�V�}±A�A�I�y�)	M�^��X��5��0��o����c���d0�$s�jU����}���q�Π�l0�Y�VC� ���H���D{��wc�#i_ʀS	0Ea�) �H�S��b�^~�5�����a>y��� �\��NP��"�>�4|a+�S)9�]���S�[#1�Y;���I��oe/% }�m��j0(o1C[�ƚ�}�1AG�Px|e�|��ƪ䋵�ߤY+�lo���3��n�*]���*����M�|fM�5L�����w��{ݤ�z
?�8�V9i��
��/�v.���;L���^a�8�2���[jp{z/wЊ�e�����T�]if7��e ��R����[�9'��&)�^���D���W$4�=K+�Y�w�m�q�)�@˘%�3��2�S=Nݣ�%Lt�E�R�}6WE[��;�S��Ǉ���w8L3�]H8�D�$P3�h�|Li�М?�W(PX��k�W�O�(�{\����4�9]o�P�N�чW��W'��^< �>X��r�*ר��V=O��������T@z�L�<F,r*b���h�hܛGl��kV�k�-9�6V���3��u6y���2������E�)�5D7K����d�gݷ��w�Z�#��p>j�M�b�p����!�Z��@C/�烵�f����z�#���}8�tX+%'wS��:�u�׆�l��mX����
�ֹ���H}���f� }x��}&����{<ěF4�M��WL�ǍJ���x�&������4p%����5��gH��$�2I��c���dչA\���'��̔�=��JW�n��c��8���U8H���D���\���kͯ�{���?�l&5=��emv�/0�>o��*�����Ύ9�$0I�0��.��Cr�dgR�s܅E�-�k��o*�a[�yi�I�p���l���P�?Ա�FTe�@���L�� ��<���I՚������hہ�?�0mV�ؒ�$pcE'��,����[�b�egi��I��_Xqv�*5n�>�J-נo�3�/>o�ZQ��zfn
��zNp�kU�̠UNM>P	�����Ԝ=�0ԓI��>d��I���G�,��<�!f�����D+���3
%w H[�+I�ĉ���nk��v;�l��A���!uH�wu1�m�cf?��^u�2:�p̆�)0���y������ jh��t:I-S�p.~�>�{��&30�b>o��d��nm��l�6��kDp�	�i�M�5�Y�w�NJ�F7O���i�ThE3��En-��ߢ:��`l��B���FM�io_C4^w��������.ptä 0�5S�M�Ag$�'Y�&|�-�X���j欌t~5�S�[��s�l�6C���Uu�}Av���n~&��s.�t7��U�ʴXW�D��bʝ���Y��+���z� h:7��ٔ��
0u4cFl�훿�K����^�p]In��5h�z?��_�-+���ר#_�yu�`�)���^�P\�:m��c�&�͵X,�Zy&����%�`����f�D_�) k`byb�bS%&_����g�W�܂��א9�9E6�D0�{�����S�-[�h�A����)}Z�W�s�R����D�}e�-����庻�Lܷ��aw��V���C\�%#��k(��,������G�(��:U��g�P.�n��o�p{�0�q��Ё��Z-����7�b�|���O�F+[>�~	7��
A%��h�Ն8�Ֆ�Ȋ��~�8A�^���2y�}h�����P��6d�L:�{�2e���!���L��2��~7""��i�51�<��_������h������P�g��������Bhe�d\��з!��|gF �0��C�%����ݰ$�m�>lJ�W�l-�5:�L���be�<��O(�� z�;T�+�x�ԩ̧d�3S`���>M5�:4hDw�����b��wY_�daKx]��#��>�@�}}�u�Tj���|$��TqE&wj5�N� ���j֝��1��b��|j��v�g��g�#��Z����M�!-���m&��;J��1W@yC����R(�/uy`N��z\�أ�?��mȖk�Ln�S��P���D�ئ����=�IkF~�c�j��3U�y�@���>�@W��������D��ߪ���7�!J��{d�2��H�,	�!�/���C��RV4!�x�d��J�v���f�l,Z��M�j���g(�e+^�:��p���	����x?��Zd}���h��y*�@|#|�	�U@���u���K�z�puE2ք�n4Ak9c
�������Af����⮗��
�4�y.;h-�5&�>ݲ �b��p������z�8�͏Qv5~	� �R���m�鯅���s�4�WrҊTʍ�%E��Dن'\TMp|���W��٢�c���z���SC-����Ǝ�II��
%��˻tҡa�'i�N1��*�����iVa>t1�px�D���7�reD�,zl�X#�gNO�wj���A�+��2��]I�5������ك�Y���-\C���덕��LҨKˇ���VU7$��7�L�/�3�Q�'�l�w�]�I8�U�}b@���(ݕtx�Q�B1�d���pjjJ����ƃȘ����%x�U��eg��4(6U8�t�lK����z�r��)��x��`���g~��GY���[JN�ę��ս;W���`��W!�*8�HdᩝLU�m�<O�̊��v�O�*�fry������5a�M���@`i�aee�jb�9q9��7{ z�U�S���搋F���J�yK���پ~m����Oеݧ�+�hf�&�?'���@�45�� Y�Oڢ���ndV-P3�ԛ�o�c�|�oƵO���L�+�trfl�(�;$Q���\p�i�;{��!�D�XS?)V�)$	Wm��/���v�5�f)��p�0��wiɶ�=su�����A�_��*A�g6�&}��p#E�y:'J�1`��O��Ѩne��i����5���(��Cc1Us�>]���Js�K6"���e@I �-�"�:6B�,�RRfW��L��
���c
���[3�/�m�u���Ŗ�ns������A�F7t����Ù�u��}�ƯI>�����d��©g� e�7ym�p�~=��D��Y����L?	�	Z��`
�.����\tK�Vn����\XJ)�Uo�Y@-��fd�N1�	�%��_�D���K��â�DP����ߌ�'�>�����y5@*7�~�2e�뉺�%B^��d!�wZ`�4ˡ�����+�G�3am�kK#�*�W���潼�O��?a.���u���핊4�����#�����Nж��t鋯#>T~�e^������+Hl��J5Ѯ��ⅪM���[�Ei�+2Z~0M7��7����a��*+jk��ji��T�2N6����1��th�u�&���˷�mŇ0EN�6Э,�y���|����$ gYj����W�_���i�D�:6�He��7!n:���y�w�r]��E(-�}��{.wK&s-?��TI�-�%J;�`T}��s����|����r�e!�!�ZwAKS��X F��"�����,("�)U�5�) ���T�X[;ng�YNd!��h�����cڿ�2��گ$n��q
����s���#%=���tE@iu��!����(�=�M�
�D�E�w��.��wl�����ͩB�pp�r�뉸��BUĈ����b��A��޲��j�����4gvS}���7�u��&#�X�M3�j�#�1R�|�\cϪ ���l�`�˱���M [P�{O�ɤ��w�r�\�������c��qI�S ]Ln�3���h��U���R�US���uc3 e:��AA�!�`�+��J�~9W���b�����ԯ�#F8Ex��]�}Fu�wz��V�F�ղrЧ�Q����"���qR�D�ײ;��L�uh���~�x���Q>���	���Y���U��U�����<��-�eJ�ډ]��i �#��A�:���)���6 �X#V�Q��Y�,*��X>�[x"�O#�8�63�1�|���Srq>� _�;h|�����7z�x�#]��6�=�=߫TlY��[���}O��0E���^ߖ��H �%�q��+pf��#u�@I9p�͏B����t�ER�*dKĔ���,H�v����WѬи���I1|h8xB�"s�>�5e}�P������}��w������w^t��ڇ9�[d� �k���2�[�1_|:)i�^��zU*�h��c$MJ�4!��z��d��?����XҘ���h�>�Š�o�D�J[�2�\��N���Ob��W����1�,���~G���,a�:�_ÿ�x�y�Ԇ��X�����4��@{��s�_\�3CF��X�Bܮ�PB����{]10�RoG@���*!O@F���ϳ'�n�{�m+��!�A2v���}F��Ō�z���Ej˼>�{O�����IP���Ɍ�kм�[�+��]g,<�Q�1�<B��#�E�.�G�v�==ݱ�|�P5�o�	�^��E�8��]䯂uxR��Vܠ^cwJ<����q�T�s�}g FP�����o���i�}�D�w$�Cwn��Ob���J/YP�e/[H��<������W�l�*��I�-��ËZkEb���y몧�9�R�p�`���G��"�� ��55������<��L�K�Z�?(��G{+�j.@�������9IĿ4�A�s@��OA����vD��v�9�PJc�(z����{�uXD��)�~6�ܓ�g�<�s��/�� 5z"�F���� �������韑O;Q��;�����r�=3�t�k�0�� ^�mU�c��Y=�߯�1�n��T�Vs�[���+ZL�/W��������]�k�T�ս��T�0�d�����
��tIbA�YQ<½I�Z�R�&R��2׃�uK�T����[,F�|��)<θ�Eóz�R�wگ��:�OMl3 ���7\�V�����Č��H�L����x���l�Tɫ�q��F�ť-'z�,.گ-� ��\�烸���F��b�L?�Ϫ����iH^�� �1��/����E��.�5�x��3X�n�����,�B +zq��z�5	;G Pjxc��� �rw���69MSա�ۭTfh�D��sŧA꾴�	S��b�%%2i~�ݴ0^��7�,Lw���P�"����<��^v��j��,h%N�ۣ��R����~(�O93d�6P�7Re(�L����&7�m�`ݭ�x]8�2JI�ͦ���e����W��ϸ#�16�������&M[� ��`��$��o�)¦~Z��nf��cHK��X���2���;��.>���Emd���y�.� �L9���R���w���e�}�*���	�К������~�Ko�kr����&�]�Rk
��n��)��Xۓ����V�X��K����'��ݬ�q��|����hζz�C���cx>e�h��?�?v���v�gqd�ɤf��3b0Wx��"���yʠz��i:�&���e�\HK_|ߘ2�Oи�P�}(��y/Ln=�,Ƕ�Ure,����!tU�
f
��^uQ1�5�C�z��U��	b��Rx����,��:����2L�g����ƥ��%��}�$�o���.R*��=ʙf�W-���u�g��(�
t��|�Sf͜�����/	�v�˧*'dT�fi:̆�Y���\�-�r�����jX�o`��_���;<��^u�������~�s6��n�ߌ��_1"��v��k��dx�A+u�mj�\��nl�7sۦ�Y�����X_�lj�[��b����u��<a� u1�άD#�^)m�z�k�9��hG17st�x~hѼ:H��'S���-BB0�߀�4��#�}0<�.�����L���CU�%L��gg�T�!�YO����J�tq���>�?#���	�H���n?z+=�kD�Z�)z	[Zn%�&6��6�阶��{���m�Q�H�$�#���ț���q7�%'�ZEeIt�9V˧H��s�O�z��!�f� ��돘�U_�e�Ի���F��H��絗`�Z�f�BZtu����i�m���G���o�*{(M�ߘa�%���i�ui*�]�2,!E)6�ץ�͚�r�<�q��X�Y����9��{�*�@�OkkpI~�Z�I���b�S�w-RK_>`��o	U�	��m�����t����o�^hUʔ>��Ҵ����`f�R�M �6��4>�8��?m�l���M����ͳ��B���A���p]��Q�@q�ci��X?�V�������bQi[�_�|IN���Bn�uǗJB�YW`�:��.��C������3 �>�����;ɒ�A��[5;��i�[�)��	1��R�꜕{"�������e8�WVs��'�=+ `H�Y���g�wr`�++>�c���=hD/����#'O�x��|j�>װը{�P�ϻ鑉�2�G���]Ơ֑�O�	��Um������!���7��N���V����]k�V�T�l7�K__�H����U|6~]�ުxڛ��Lk���\��}
(�.��B�:�� Fԛ�vV{43�����B�R��y��Ԭ��Z�H�j�@��x���R� M"k���9%{���h&���Ԝ���t�s0����]�!hL���m3'����Q�3h�|�b��:��'P���}��c&]Lْ{XI���w7s�<�9����j�If|,��zJ9��� �ۦ}�#�L�ԡQ9��t��x�)u��>�"���M�J��}���uE���b=��0�������xS���5�"������`��t��{(�-j�$�ਠ2���� �E�K�ǎ3k%澠�V�������q�"��ަ�{h⭾������Ⱥo�{�؊4����F��oe�W�5|����f?�	]�t$�)ڶ��	�2/�7e����X�@��7�f�Ϟ#h[����@�q�2]e�V%S�	h���Os�#����[mtLWR�L�~te܎�&���.�I�ϖXQh(�>B:����*�	��$Z�"��ΒZ���܁vL剈r�zn>�����MT�~Q��M�p,#W(�x@Q������F9�����1W��Yn�wP�J��о�I�B㢖��o���)�͏jK��ٰ�T������t���KZ�z�)�iy�F�������2�M('��T��
�Ŝ	zg���SgN�E"O)����Ap�{t�s��#(2���\�z"��0T�����[3E��	KyK� o�����P�bM�U��;"�A2R�H�������Em1�epv������
r�h�[�y�`���8�{\4����\J�����Z'���aCt �8�%Ѥh���h�h���Ζ��ئ�"u�A��U+����]�"ǝ�G�d���F��z5g��Z�BE��u�̅[Օ��6�����)� ��aW��A��������+�Ӟz��3�Xl�t9B��6�Ȓ5ް�SJ�(Q�UcU>e$�^�`�Ƀ��.\-/{Õ���]\ �� 3/�
��?�sTjv���9�x��X0PR���֎���Q����$��	�a��2I~�"�����0�䴯ǀ��!�e���轀X��E�e�y�����4řU�0Z<�碷�q[�]�ʹ�Ahc,N�\s��AY۠O\���]%a/��X57���V��Qļ-ܭ�s�fu���;���v�=s�`�5�c>ы�k&-�v�nG��:��*�$�qP���Wo@��
NO�$+���<H�ZӚ�>��)g�Ò���?.��{���ES^i�5����]��\΀��QZJ˿
gѬw*�>m�]k�q���8� ,����d�[��@��&X�1aJ�U��(%��Զ��,�0*Bb�Ϳ�$I��hd+�!J��t�U�$���� ��e�>��f���K����o"C�{\���|"�Z���D�]0���e~�����c]Wn!�K`[�j�*�	���<s8
E6ʹɲk�=�|��<�b���u̚�U;(G����o�?�⦽!�t�X���[���影�Ns:�&�K�X��c���eњD�o2`A�_�>��SM@�FAݜ+��ӈv��gѥ��Q�T@�� �H�P�����5�u~�h�OD�����d�,��=�{F��[��~ɩE̛0N.>���e��3��.GV� ϻ�C��O�b�*B��@9����(P�Ҧ��jUnp���Y[�IA#��Y��s�6���Ð����:�d�-s��jyڸ3��[��b�K�Y�3�@|
��۵������'6���VzƯP���?f���Bc��2�Oe4M�c�/�e�.)�W}�܀��[�F��9��[�Ǝ(���1�:1�G܉��1���ax�
P�� ��.��l�DXL��*l��I����d�`T��+ H�f,'�g�Ћ����s�u�����K=]^-4X^��g�G�r@��ٰQ"���^�ERn,���u��'%���z��b���{o�_��"�9���R��[����e�t�5��=Yv.AFS������:�:4�(���-�Pϕۡ?Pq�A���mϭ�^3����n]��U��	eJ5O[J������Ɛ��8���� XӁ�\�g��Hlz�(�\��x~��}�GR��&ҍ�8�&�;8w�r �m�oԇ� �����j���{d�?�+ZeR��w-,�T� 0���1 q��w��v}uq�Y������l\�X������ ^�Wg��Z��c-X��]l�bh̚�sJweԀ�|/|iz[����<ײ{i��5�b�=�.��_�5R\�p�J=׍Z�D�������3T Ř�=�p8-`_G?�*�Ⱦ�����5%��q������B9R���"uR*�x������j�|-��I
��%��()���)qK"d�Ƥg�������T������VX�
����OK������7�U=.�ܽ�LD��J��p��=3) T죏>��_���b�ӎ���CHp��v5�9H��Ϋ~�3��@t�<���Z2�N��c3(�=q�>��}��:6Pި�L�m�G�p�scW�5^gf�;��s)�;��r����ಋp $��&Ho�&�3y�ԑ.�?�lK�Q/�r����x��-Ĕ�c�`e��_M�*HD�v��}.0q�>���gr��G<��lO�SS]�(�c�P�Z���j1��˲�K>��;�bL�v���]'�K������O����a���ɓ���ʕ;�;�p�l���N�V]��?k�붭��q/���07zh/1Z�����Ń����]�����Je~hs��o3�[p��<����N�|p-��o��>�&�����IuȮ&1y�C�T���g�e�����2�_.H���Fnbi�;z����2 Ь�i��Z��A�@�ö�IƬ��-��R��)�Ό�0U���E�ͨ���J=M�B�i=�d�꜐�W�kL���P�w≮��0�ͻ)�b�φO��5AS�x�>"�s��B�6�"�h6L�N�����;:���8Q-�\�.��hEK)��&���S��6�m��h2-��[��4�1� I=~�j�7�Ի��y]:­!kx�!2���"�5���G6'��N0e�!�z��`�L)��/��c�ܾ�C�h�r߳��gJƈ0�|f�#*<d��H�'o!���^� A;q��I����񇨭�B�8Gi�>�wK��N��O�eت?������㽵�+Z����?��vDZ�q�`���DO� �O�_�P��AL�&�5�Iq�ʕ�)�{��K<+�Q��xlbh�I��T(�cSxͣX�� v�c-��>����W�C5��W�|#�CfUo{O��2��iSE�
�%C�Z[	w8�7b�D���0��6%�X�2-3pʕ_����n���u:v�V�q��x�I����9���Ѕ��U�|�����>�6��N���G�qkj�7���W��+�k���4��Kz.��{-c����|eP��ÿ9r�{�|�h}�2r�]\v�Y�j����>�<�-x+<���G�鉝M���ć�[�Ǯd���L��s�8H�8ſ�gB��,xʗ��ZKx�J�#c���5?-��>g��;L��y/���f�m����\%����jw���^-��+������A���^P#�.�d%�&��1�l����g�S G�vaX'�;:@�ֵ����L��gF�M@@P�f��w&D]��e�s��$|/)��Ip/�#*��n�q��q��{3�_��N�2�^�-"ء����z0%O6��Cd劦K���"&��VG�Zmk6��{/�e�NXR�Y�w<�A�<��>nS����8%�������=��{N6���P`�8���(���]
;����g�02�$˟Әr	��w����j�������jS��Pt��-x�$�ď�����+�b ���i\�����D�F�x�F�A�宅�ڴL��T�:���iگY��;a�y[��GᲔ&iw�$�:��T[S,/��qޯ���1�P��I@��K(809��ՆHphP�b/��6��d��_P�T�<�o5�`a/��o傅t��O�%�EIN��EY,M�!�����Ո'dB{>Ԩ]{42���?�i�>��_�Y���B;1dT��:�pg�A�
2�#��h�]Yy��iO�y���5�]� ���K�d��#�TM�ϖM�ٯ���0�r<νh{v#� W)r�)�H~�0��ݛ�ͩ>$�9@�lϖT߼��aә�LMX:�E����Ҝ����j��sL;?�0L}�q�Gٚ�P8�;�y :e"_0Y����.`���<���I���C�s=��4�F���z�Cmo����Kr�q��?��mG�A�)	�Y�s��v��1�m��m�Aޤi\��8N/�L��k����P�`0P�R��>uE&@S[���h���[�#g�����+�x�Z�ĂS�����6W�f��5��k"-gm<Ͽ;�YT�C�u���);�e���	�x��)&5l�<�X;z΢��̓;QO��If��&2��%5��/���R&f5��z:�w8����yȴ#}֋����'�1���R9�4�oc>X����^��5&G���!�-Ӗ
/G1� �͜#�r�D�e"/�	�;��c~�w8��Ul�yx��1zB�&g�N$�+
�
��u��:���+B���6����(m�@}J|��a����D���7�Jb�3[��h�J%��ۑd�=g�G�J��j�����$���ptz�Ȗ���J`7�����1��X���sٝ�y�����߬>�y�)Bi������E=(E�u�(��G�Թ���kC"���7���~�0ӀJ��	�D�m�ϼh'5��ϕ�Ņ��f0L1:|�l��ź�?�D^t�<u�$�Oa9��@�Pt᥆�t��(	Sc�����]m��m1֨6sZ�I�Ҏ�g�tϦ��e`f5� U�
�)�%Ó��՛M��հ���t�iĘdr��k��t��9��.�@����\�ޣ��>��a�_�g�nnf�M�IȻc��ɕ�E:�ǿ.@��]�MM�#�]���1e��fO���ͫP�6���wU�m\un[-�A2l��@T ����+��rMH��-`��<�d;��6�#��mQrZ`c�L(��� &��T8m�ߝ,Y�	���v��_���Bu���
}v�o�τXy�Zy�㡇���RQ*�oľ�@��"��� l,<I)PN�	k�.W3t���'�Y7���b`Voi��� ��z���諳HA�r��=g+1�ѼA��]�c��� Zf�0_�y�8�����B�����wP��T�^����'��&�:�3�N��#8�gK�<$�C�:˽��L�
�E�j��,4Zy���+FH�j=�H�2i��G�o��̯���ӹ���\Hae�	�@"P&&�@��`�nY�a>'?�ܛ�1��4�-/F���M�<L�8tǎFU��v�s[0q�a=(e�n��������d�|�	�W�˵�x=��
�k�	�P��r�EO�=�d��T޽'����������OH�����`ɨ��62�o�}� (0Z��v!�y�q�7VmdR�-��fk$����<c��G�:Z��\���|�a�{B ��}��߼�f�`�����2��%�b}�5�� ���g-zaȈ�=2�#f�b`���k�"��*�;c�e6�y!��+cSթ��*�!��sSU��� ���v��^B��wl�k�Μ�kߥ4��5߾j:��G����.~Z�����L�FW��GF�m�����x&��e:¯�D).6VX�dy�"��� �9�䊘���rWR����G�:TLP�$a���J/�c1
˱�k�l'=u��d�DC��ȹ��-U�g
���j	 �q�C���6J�!p��tn�P��dc)}��O����6C}C�?�J�N0���f�`��Cd=�BJ)��\"� 2���`��i
�1��gн02�_N�z@�/�=Ptq��,�z���i���Y�#=�L�n�,q?��7�6R�|��*YQ��ӽ��3ӵ���(���S`�7��)��x��y��t+L��������/?6p�������a�=
�AI�Q�DwІ�@���P�DI��,P��쿇��V����Y���C:�C��(�����G��2�"� ��x� ��=�!���Kt��	>�R�{��ϼ7�v-U��iV���5j�r�]�y��w�#���e�t���gȈz8h�YT��!��W�2{|�_.*�\��A��u`�rYTd��WP+�z�d���D��<�n�Ks�d*�$����LMh͕<�[
�[R�V�be	��\N����˟#���A�q^�h��1�pN�zu� �04�v���+�L���T~Um�o0 �2U
�پ��WP^+���Ha֎7X�*�J]�S�v�lU�g���{�B�k�1 ��a�#X?�����N6l���
E�	D����X��	�H�_S�c;�V݃j5�;h�>�S����Ճe�e��� ��L��l�ط��*��RJ����w}g"mڏ���n�y�]�����gO����`��A�ja�CNT��g_k�a�/��:t�,�����IILy��]\��h~�8)g��}�r:�h�-vxv	"�F(ƞqx���O����<5�����C��avj?9�A��j%:M���]�,w��"�Q��f]�y0�6�.�v�'�l�E����(�o@iv�?��5�gl̷��kJ��\���	hW(�h0�3�x4Ԋ(���H�]8[�9
DB@�b�o����_�Њ��C$�,���n��(Wp�ab����NO����-��r�������%%�#ζ��,ΤX m|�*6}yK3>8Y5�_+t����i��{/z���Ζ(J1��n<���#Œ�gG��(���B����>j�}�$}Ba4�RZ0�t%����Mvm}H"�I�z��6xU^l��aW���|pȥ-��Tg����]���»���t"Sa�A�8�������=��֚��ԨT&���4��J�q�z �ċ@�̬U[���g�Ry�[�I�?�)��%����s�c�=�O���6�=���Y0��6�E��xM��&����G*`_�^����K>�Ӻ/Aa���#��r�s%]�z*��F=����,B�HA�vsY�8Rѐ���&�~c�a���v����{�̆-M�4ؙ^��R7n��;�K{�m�E��#��h�
	Y����D6��e��1L� ~�.���>��TW�`}S/ >:���51��wHE�X�iS,3 �k_ƕչ$F�6G �ܟf��6�������H���3���- ���d���M���������=rk�$Ro��_^���Ojf��dW�[&y*1e8��Z������B��L�[vH�z�I��ߦZ�̖��݆ZO�@'��<��T�LPݦf��t������&wx~`�A�G{���v<�vڤc$����Z�f��2���ڨ���"r�f�90��9H
ޤ�lF�yc�멒\a�s35�Ȟ4��"c�[��Þ���."�oK�/���T%���Q��Ǭȃ=Μf+ؐm�*�p$�����Ib�UUS�_,6��՜Qg��#/O��0���L��	�ɪ�]N6q�Kq�~�R��W���|!8z�亹�,{(` £���z-G� �弐��d��oOQ�^�Ibo����5�Ȱ˿Qo*^�cU�]:^�]j�C�X�D2�V(�N�}9�H	hJ^4�������<l��G}�f����S1�s|��2��&�XN��Ӟc~?�_���	�z*���ߚ���A(͞�X���U�p��d��L���
F���z��m���(�$TK��s����U����=��ٸ{��~�\��7(�<�+HU����yx{��o�31E�����0~j	��(���z-���I1auA*v#P���`�Y8A�cj^��+�� ��z����s5��F��/#����Um3��i��C����<z��_""��^c�L2o!【��")��U�$n�b