��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�J��"4�=�7(�T�JѺ�ő��,\��s���ӣ�F�؏�����;���Wt�R�0�d
��nF�æN���8cs�����
r�8�6ն��8%�yU��/���@��]z�Zb�/��]�,T���<c6�
B�E�"��yk	@�� �o��b��zw��Lh����8�a?d�h��~�N�~I��c8G-"lF���M���j�_R���os+�"D��R�T��~�F𢠥c��l��3Q\�� ����pq���G4�����%������=�G�N4iF�M�}}Q>h_�rV���U�-��q��?��	�q.�z��p�<�0�X�eIH_�%&����j�	�(�(�GH����!��^�0؋;��mJ�a\}0bh�B�\C�Mȥ6譭i:q�:��%[�+��.��wm�{���Aj#¨t�]��(i�Bkhg�n���ܱ�|�a��i���ʵ��?}�&�	%p���!ۃ����Rq��G�2���}N�-ħ�8&S�)��c��!�ğy�U��^1�+�(���̉DH��=H����SƟ�8!W�M��ypm�=�m���\ J�LQ{k�|$-�0��&�6�K7�d���r��?l��(��<��̲mM4�H� �a�J�)U�+P瞭�f�L��/>P+�f���z�S�T����">
\U���j ٞ5!G�<];�x�	w���t���@�mu,bVb�F�u�w�P!d��l�4z˨�Y�>މ�?+���0)�3H�g	,�B��6V��sδg�D`0�l���B^�%?�hF �=8�e4ôo�h���>��bV8����:�̞�k���i8�.�f�r�ce�4�̏��9 �s���#������8u� 8ׁg7�a
���V%%��D���󎆀9�B{#x7m��f/�/��`C�/o�Rڜ�R��!�&�>p�s�)���?�C		�	#����?�ʧ���A��ڮ`9������U��b�#E��nMPsڥ{��w�\q���:,��k`�i�r�D9��7�Z��3g�j���g5��j���ia���Wb�A;F��KM�q����N�C�l4f���qDB��V��	:�,�����wLs03c~��/�{����Z6e�0�.(%�¯�O�0kGcs��3���#	)N������_o��`�si(�r��@��Ay�?��Μє�m~2i�z!m]8���~�6�P)�_��KY׍�2N*����aB!.*V ��?�I��;����|�j������V���_�39�;H`���\Ζ��;D�,��sh�,�W�9���-�;�x����$8o���ZM�3#�	�C:�ٞD^�Z{R�֠Z�v���Ξ'j�� ��'�4s=&��O6+pjCU��
)UJ�^���3��<�>��s��\��r�^��A r������\�,��L2K�y�j���~j����:`+;פǯ��U����KiY���ܳ��=��'�h#�{���^��g�ޱ{k�N#��Ě ��^�-`O�t �9�_�s�|Fa�����jN�FS\��䓌����H��խ�Yp���T���j,*�� �['��ٕ>mޙ��$����<t�	��G��Q�q���]����8���������2����+�)a�}n����d-�H<�ב�WW����&|���,5�1m��k���h4�����m�wޛA�X�"SNT�fҕ�2�_��+�ۅ ¼j��xE�!I�-2��0��OCE�l��ak��H����N�Ϣ����́B�G�_[g��5")oΓ ����+i�ʆ2y()�q�\@���\���FC:z�����ZZ��˧X�JHG�4�^`��3��/˘5@�&M���ӻ�ߜ�i���r�4i��h�&��Ǆ��I����<{�,o-�\��0[��V�o��"�f����.��D��,��=G1m�ֵ�x������S�%�껵=a�l ���FY ���%�i��p��*�K����>����{�~8�'H����T��?�����T� N
�IA��)n#<tc�Z�N�.���䎻��07�p�hs����V~��'��i^�5RM !�vn�H�<k���$		{�*5��'ol�}���;�ֆ�c�gR����;Xe �L%;���K��q �[Ma�R�Yɐ��a���(�'"�qV��:��Wm��D:8@��Pr؁5r�_6���} l)0���Ǭ9n���%H}�*X��jy�A`;9q�bV����2\����O߫
t$�i�&2W�����Q�u��|��Z��V�7�YOF�t{G`��mk�nO3����t�{��彨�`�KO���q=\a8�i�^����zU�DԾm�K���RÚ����Ӌ���J�{j-�~�l���R.�uJ��3Wpܚ�m�o^��\2R���qt|+���[^��3�x�O���Z�JI��u�i�z)�R�͒������fχ�T�?�ikӈ|`r�{�P�c�Ok-�Xp�y-��L���K#�X"���#�$�	ɮH��ӫ����.n�c%\��j�>#G��u6�͔=[3V��d� �ݭ%�x��%$�Q��i6�ɩ.��E�d�}�l�=U�H��RUi��K`��JYQ,r�z����j#��g�mj��)4�C�C���I����ƙMdi��Є���
���9|V�U��j�X��(����9��=���<g�^04HY� 9��|/�V�������º��n���x
���6�X���b^*Sn�1��tCdFd�"%9nY���Fx���(\��Y�A�:�;䭭�)[�]oJ�D2>Hx�A�
�ݲ�p�����sA�i����4v�9M���>�1IWq���O�i�i�MG2G��$��� �+3��:2Q�vwJN�V|�u:���՚V��t��=��w�+\ R?���t��33��r̚^@g�et�p�Q�����z TQ��qm�8I��/3Om��(Iĭ!I��UQa�6�/��Qo~�U�z����5�&W��]g��w�M^JCbX�+13K�$n�ގ�F6�Px,��#�0������n`�0�/�I��:�1ۇ�%�#Q.���c0�@��o�ؗk"Qh�ú��O��2�����1+���}�}lv��/\�b�+��xQ�<,(�w\_:��T���(g�M5�[��P���cY����H�B}_��Ƚ�����@K�0F�Jq����*�]����-�mS(z��{�Jހ)-��E*�b�+�BW�&ִ���(b@����]9�*-h�/�6ɻ�����~��A6R�e��fG�֨L���
�'�����U�KZ�=t��{��rv�~ J��c�@S��Y<�^b��n�Q���N����(Iۛ�,���I3��I�C���L|x���ql?��V}�8��Q����w��������7�:�1��ϋt��wnC��K�C?������'�����Q�u�`�Ɛ����f;#}�<���q9B������KN
91@ �H�GY��d�3dl�\IIB>��`�(*F������N,���P%��!n7�y���g~�����>��� SR6M���Y�KlF�".��'r�C��H"�cU1�9l��#Xh��Z����T�-�M�7��0� V�t�G��tuw��S���7Y2��_x(� �n���k�҃���H�k�����q+��SZ�³+�Qӯ��7��Ҩ������k���$Gal���@�5\�kBĶw��!8YS�<z���<�sPJ<N<�3�"m,��J���'%�3i�M�;�v.� "wA�(�{�N�R)
k�c�<\,�w��8V�W_[��Kl}�R�h`cQ�[�NH���~�$c6bSێ ]��x'{�
p�\,=�6�V��q�ԸD���6a�:J�Yc��R��	fS�I*
H�ƽS)[
떍r��V�u~���k�������jH�߿�|�b���s�-��}�Um�_���NPv�/]�d � �^i+���([�����/ �(� �c��nm��@���w2Wg<���&�Y�j�K#�� �w�ڛ��a�W�>8�pŏW��_�A]�[d�U�c�U�թ_{�L1m�P<D*��&�EuY��;8�_-�T��Ǵ�8�6/��OL���q�$�>P�j\	��ֽ�0ޞ��5�=V�r�9�ĥ��'B����,����Rz�J�b��k��������+ta�σQL�k�̨U��EW����P�����PCu('��GX���$6��^�g�������l�tL��"�*mv�jt�4ȶ���dNK���c0��aO3g�=�1p\҄Px8���<yy�o��3vk{�����-�	�����\Y�bx�:(A�F�}�7��q��_4�ӈ�Y��� D����&.^�bt����F�Ԏ�4簿�D=�i��Ch^:��1�C"�ٜ^p��7��6B���Y������Az�@�CS���Q�H�����x��P��]�D�x2�f�����0*�`����!`�^��6*W��;uop�Tȼۖ����{�o~_�����z��=Z
��j�K�Ug�����{�Ow��� ��M�E�z��L�M�}P:�|�;Jx����CL)�����\Bk*b�u@�J�V���1z򿇍��_0�k,��I=��$�7I�6>�a�*�e��l�紶!��q����qGf2�������.���S�]���C�́�8KvY
eF��(��|�x!��_y�i��w%��I%M��w�}�=j����\B�㕡�F0��[6B���e���z��P*���[�w�"���O��L�P�ڔ��N�3�&����B��x����~����Ґ�`�*}�wk�J��!�)m�ڙ`o�@�-�g��[���2���~��G�'���_-a�ڲ��Q쐰��n2����B# ����DhU���&�S����!������.,��V[���I�ʙ
˾<���eق�r�e>�fe���s���O�M{\�c��P�%��
L+Ѣ��%�!��6�2�Ww�\� z��,��z?�
� �uڦ˂��_��H}}o���i������gy��p�T�
�Г<զ�P���y�[l��;�R��R:�Zɓ�Oɘ���j��"3�J3�����Q��ыD�[$��|�*�|�[E�z@��9G�j��<=R�;��x��(���8[��Rx��l�M����E�>��_����u�����qK���9��~G�4�G,&��470@x>;L�m��c��>k7�zut��b���C  �O>i��
>}A���-?��0����!A�I��O��<83o`v�+�X���*�:d�EӇZR�y��2~���o��BG���T�G�y��(@���3�?=��m�6z8�O��S
?U��P��˸i(%`�˨>�g/�p���#^��K�Ə#z]~:���UWr�W��^�q�LB��|Ďd�� �<��_^��V�Di<bl�ki
�O��G�&�;Ė�,ɇ��=9�yc?�C!DR��z����o�qX�j���{�:*׶�<k���ah���X�*<q �h8�I��"���~�H��qN�$.�xφ�8�-mQ�E&��ōdiZ�lS�F� ���Q��߹�po�D����>�4��(D�0���0�ryr�r;�&v�*�9T)�(���Ҿ������?&��� �7�y���Eh�)T4�R�����M����t~��^	X���	����}%��d��ƛ���i!���g��{"�N�ι�On$Z�MJeo��I)c~�.���H �J������cLu R`R��w��b��&0����3'd�t����#��S٠�-�hQ����9��Q�/8���<��u�V4���q��Ot0����2�������}&*�#>�T[�_]#<(h<CgRxy�.ŝ{N$6����7
�[��}8��� ��o!�+ȏ1�ā��K������EZ��c��$��|VJ��]
+��6R��!�A*9��6�h
�z��PF
|�T�S���i�����wbu-{��ј�yW�!�E�-}�xemcL�DX�����k��X�n��
�j�z��R�췞g�㻋���p��U��;�D9V�lڃL��̱t�O@���_�"�ы�E� ��T��C?;��@h���p=]J�VO>k�9,�H�2��_|�|#�u��9�f:bk���(��p���p��; �)�x���%��S��6�W/�,��c.ئ�C(�(��n�͂X\�l�?�aA�st,��znmУ*h8=C8�S&�h3E�����D~բ?ɶ��{���W����̨�EF�Q�����wr�i��
c��,N���K�zJ\�Ғn�O掩�a.�'�Z�z���x��ov��o�*[�/v�I�!��g�ׅ}��V��HE+4k�K��3w�U��NL�*�J��U�T �H��C彂ϑz[a�`��H
��JWݛ�xAt���uFe��[p�	����R<;������ -GU5o�T>L:
U�s0y%�_�ۑ��6�7
�*��9����21p~%~I)�A8X�ob����I�����&�z[�}��~�����69�z���&����hu�z�
SH���wI��8ل%:�}+M����K�<q	9x��� G�<�I"j�*��fۨɌӢ$6s ;��jD��Aݨ��� w���{���#��V�7��+[������P���R���;14��`��Ay��X���Zy�� ;�o4?��q�$����_��#���W�֐���$.I�����ӳ�fޅ̥dcpñpa9q
%��ȸ�54�X���U!\�8��r�/�82�V
b�O�(xXd[6F�������1E�2%���H�]�o���H�EDͯi�����{Cc=��r��>V���e]�����N�'�]L��m�	�&����ݭ蔴�����C�FKk*��$:��2��AK*�8��h�ػt���1�L����ņ���s�p��|�W����f=r
�e܂z��&5y�Ί���ĨU���+3�Ur��旚pp�������uƜ�K>ZB�v�q�U�g���l���7�'����]C��]gl���9�<�aǆ��N�j����4��H��J���u풽��^�l3�qm�<�LM�4���Ĉ �".�aҗ�:T��.;��i�D��S�v���K�Nu:���3R����q^�cLF�5�ӽB����T	��9�ב��l"����?'��Ҕ��z�9w��?jMY���gfC/���k}�Z&a);��2v��.��o���̑Jh3����uv\]�=k�&�w؏U©� 6Ȗ ���atz�8(#�Vm���F�yBsډ#�0,���e�wϋEǊ`X]eǇ#�ds�����h��f�%k�� ���7��vV���xa�0�Q�Gd��7��x��nl�oZ�I�������F�m)��d��K��	?{]/�U���U�_~K���,�P�JWEʽr��I`��������[���yI���'�"t�q�a3�>�o?�B�x�	���ic��͘�_�E�[��F�������D��"1�2��++�e��JJc�h,py�L4Y/��[���N���[&�49X�ˠ"c5ouޟ���_>�(�[6���v���VM��"�-V�jF����v9����.v����6�6�&����>���.J(�bq�X�<q��K�.;�w~�$�s��A��Y�q��+��z4p@�\1h��e�]C�^$���" )�inY3TS\�z��<�(s궃��r��G=/�Z܀`���-�i�TД��w�ӥ�=/����A����:6��ͥ� i3��)�]&g3z����Hj�w&���W��=q.c�-�t�.���
�*�W"�#X<�U�v��\�������clŮ�6��^"]�n�j�B�#�,�qS� Ti_��֎�f��5��IP�ܓ"���`[�bNrո��aA{1��Ծ)����3�Tghݭ�m�BTo�R�=�$��m������X^��cB(�݀�ԙ�j��Oi,#��e
�qR]}<,��y��47�qjT�K5��/���.1���o)v;����E�"��w�q)�*�0����/��EBH�;�3�s�L#nu��̬�X9@��tx�@��vQ��ʀ�i�(��l��]#O��l��e����#�v��ڼ�Fo��CG�h+m����$4�S���P���N�Qh��3��'��K�ĶkW�����;�S�W܇jV�)�_P����'|V�,��^2�cTA�1۬S���Ff���Ttl���?�W&7�
��?���)�W�u�X�KKm6��_Y��^Y2��N�A��Y���R�l����%K\q��'�o��P��7�]
l��Zn�m|�(�94˦�j�"�hg��w^-�ڡ������׍�h�z����Gh�Q�s֢w8��w�����'�M�>�I����}�7���V��^0~���z	��v}�&�r��j��]����63"�A��6zw�I�dC��o�k_��aX���;s4)�'^�
���~ʜO`����÷)���0S���D�?�Y���kl惾q��}9�7+@��[�$U��A�El��$��Moַm+>�k�օV��P�Z�H=��i,ux�	ڦ���ƃ� �P]�Q�X�AIh��D�]��h����\�� ��RxР2?�B_�nV2�隳�6�&:Qq�tg� u[\�H��_b\��y=�������J��p�q�;�I%���b�$f����εu?:	]'����)���@��z�GĖ{���_�U��Λ�V��-�,ӭK�w�Su�?�����tT�B�����"9��挲�pHѤ�x��&5)&C^?>��f��_�"(�����s��%7���$�ia1��2��V����C_�Ħ��ا��y�-�G� ��xP)�[���P��UxiB�1��YCL��_�>j���(IjDo?��uRJ�U�����ϗM'?��UJ(�z�Z����s.��N>׀�8�@���NXl�e<d���84�f����D�{a1n�[F�E*�(+ �]�K.�$��\�l��|W��!��ƴ��LH��t�d���N�� �'j�����P[�p� ��Rh�
�r[�(z����Y�¨�؞�����mٿ.�GJ��f�z��A	J��N���Qܴ�B:N�+vcz��� �߻ԁ)�E�@�C�K�&�����$x����1Di�R��PzJmz�hAܠn�϶-� 'W�N�F��{�P���Z���پ��ϔ��'�3��9�Ejyv���gU�ݬZ]��z�-�k`���
��>�1ӵ}8I�����_,������R�<=��
{��h#�����6�ߊ|��G`(.���86$c�����R�QP!UК��w<��a�DM�NTx��9�����~=�D�h���m�jw��>�٦�֣�A�X� �����~�
9c4<��/����ׯ2��9�
b��}�)�NҜ�dkOi�Q�XOe�d\n�:�C�=��&VeCц`�av��0�M� L�z����O:�?��\� 1��7���߇g[�1<c[���n�o�\R��V��h#_?��]�q��"��'���̉�t�+��^��<����0�f��^���߷�v��}�j}O�T�6�<?p>��;L���;��۳ܮ	ߔ%8�м�N!�k��z�Ne����߬��P�.x���mX��$0�'�i�z"6�=�  �{H���H������p�=��ùα�&�K��a�=��r���*�����A�������2�Q��}�5��@���(��=��S�1Jk�¥V��o��_e?/�t�:a��zX#�4\�ϸ$�U阧��~%�ɓ��P�C�l�M��c���g���}`-a+&8*��v�C����x��j$Ac�ӻb��A-��I^^ ��/��폍9bQ��6x4K����ƾ�%��,Yf��K��^������g�)?gYrBu.��D�픣�=�O���H��� �T�5�����oMT�*u�F� r)!:��n耷� ]>��I�e�b/ �H52��Q3]�tl0�oo�������mL>�o-7��ի��u��܈�w���%xk�|Up�P����c>����B�pۮU���Tc�����v�x�T�E��+td95ޏ[�}��u�Y�A���1a�f��[48���#��X�Z�=���M��!�Y�B�_Z���5�Q�,�{ƨ��M}��i�g���mg�>-S�3k�&������F���E�C�5���xdW�Oix2w��-�&^�#��Z.1S�t?�o���d�gV����btWr"���0��B@�;�k��H� cYA��~��i4��P�s^6�N��5/�%qS]�б���bZDQ��2�ic��9�3��"�w3�oW�����.�t�f0I�
�
�}������p�$���B��"��]�Q��uB��D��(ހ֥��g�GVC��u�F� �d|��ut.�,f�O�dh�(~�J��ȍ���#)���J��RB.o]@�����*���^�*S� ��ľ7U�ͪ̸@�N9ބ+�>��IʊZX����o�`$�J.N���0���f�t�
��	�p��w�n�ڲ �p�F��K*l��x�;ӌ\P�wȡ�=Fv�*��c���y�x��2�y��yp
Q��}���G1�Y�Ë���<�#��fS.��]���tNلV�*�<Wd���#{�������,T���f��$��jt�2dZ�'�1�7[���*���۞h��ʴ���w%R��C� �z�����l�Hd��>,�s�\5��x��������Db��{�Oc�ỗ:�(�:�N0�$����/\��`�\��H�&O��tW�f%o����\j��9M*��;�ptLM��v�s&��vK	d�o��1"!$B�&�k�Q�\�Y�l�x>ڛ�2��9��FyT#�؉�yp[��$��:�� � �����C2>�*GG\����2��.����]΍���o*W��ғ��{��)���?c�qt5Q60�P4�> �P�5�Qa�6���
��-%��B$���(��6��3��)!'�v�j�������0O���l.56 2D���)�R��i�
�<L���犃,��C��9q�3�ԓ�\J|����s���q[4��J�y��|[�IF}+t��CX	�10{�ґ�0�(�0�uA2&�r<��j��VBɂ�;���b�����
�����C����A�гi��H��ϸr�1�y�o���ىrl�⎗ou�e�tR9�<��i%��I��:gk*���^o���ˌb�v����8 0%�a�@��@|c���;%�4�h���V�9�>��[����-T�Noh��^����Q9R��a�1��F蹋3�_��t��� ��}�/�������/���btXwl�������4Ķ�T��y��+�,�.���LV ��"H3��"5��zB�L����z��n�OS�j������c�0��F��D�Y�����KN���=��2��n�5�.�'�Uȭ-��U}�a�e���tT��� &�Q�Z��z+$�p�e�5�i2��Kc7�h����l��^�V��.����0��c����GY�b�;Oq-�����o�޻?�e�ͥ��7��\�;�x�`�= ϊ�2�z^nk}_�I�80A�ӣS�#�щ��M ����J7�58j�+o�*
f�zJ#��?���{ǣ��b'
�=��܋%dD 0��|�+���`�ܾ�!�J�����h9�W���uG��Y�'*6�a'�̾�%���҄a�߀�?h��>���*k�<�����@`��?�4:��>|�N�b�si���2�K\��#���M.EBT�O,��e~3	/�(�R�͞k�Q�U7t�6�C��n�C�2������87�(�N��M�k5i�nT�2�}��=��u���)���`F�[�,��#T�η3�z�p]8?����;h:5����4bf��49X�q��@c�uu��K���yF��!�"�-��8h
��ѯ�����x�ݯ�X �>�^��?��E�7��=
Y��N�11�F�3r;/�������g��3V�٤�K>j�d+=<tXoE)/��HS�64�I�`Xx���a<N!�W�;C P����s�E�}$r@CF�)������N)O������@�
z���(p�8F�����R�o�ii�߽6YT#0���NY��H 7e�����(��;�I�92uw����P��#�%c�5���
`�nn���aT1����eۆ�g�K��R��Ao<q�<yfЁ�|��)k>��n'OQu��SRfRY��cm.s����V]V�U�C�ێ�U�.���p����r쀔�cB�m����G{���»�&F��18"c�W�/4w\�q�[��[N(�X,%R�%�v�:��(����yو
Tw�fE�*�g(�%!S����$�`(��r+k/9�ᢃ�s���ܴd���	��S��V�9�vb�+��3M9d�������ka���@�c7u���j��A���+�z�F�(Ƨ�
��_rAr���Q��B�-���A?" ��!%2'��e?��m�9<��߸ �Bd���=Np�E&A�$*�\ e���%(�(2)AVr�U$$�5A�����t���?�����/|��S��4�f�8�I�ϟ���[F6�+�SC���UM��`<�m�)�X~R�IbKB���~+rp�&�v���B>[��LC��H���٥�7#W���t�J�,Bo��n-̨�� �JBӥ	��k����G'��!ad-���c@#�ⅻ��0K)�m@�Pґ�a��M@�Q�����[�� 0�n�e�"���Rio��#�����S��� �, ��x����[��@7�.���TS-���熹b�Wk������E@q�������w�5�{6�OO��g<�2@ކ:��XŐ5-��L�T�0At/XZ	���)�h��f{���fQeJ.YW��۠O�2�Z"E�]��@�����{� ���C����r ���.WИA��߉?XQ 
��O�b�孓Ȕ+w�+z$=Y��"}J6�9�˄�^�d�ҳW=��}9�������;�oF���k���jqr �>%��2�N	uQ�@����������SrQ���E�v�,a)9�e�$�qM�,��o�����r������u�}�"�Z�$[T:��&%��77����7�\K�	�?J��:0�<��=У������U�-il�l�ib�m[ۢ�F�2��*f�����e�A�����H��Y��j�T��5���܀z��^n�-��pO�f���F�ݸM��4�ǋm�Oؙ�K��F��]�A�l����؏��ѶpHL@�=�3-��Gt=��z�.�Q���i������О�ieNyʚ��,g/���Dfu/r&�{���t���.�!�<	�y�J\�{�5�>z��0��E�w�x����Y��8�6�8�@�>tL�����7��4��N�{�Ō�G�\F�L5>��fIH?�@u�G'�miq}٥0fk>�B�G�c��;=O4��9�o����Gm�;��6��B�v%�LcXe7J������_�����yo-2���������-�E�k���N��:V�fC�ä�O�.���'S�#u�)WZ ���Ї�^�3��Z)A�B^35\g~xn��ޣ`��ȇ���M���5�Sզ�)W��ᶁ5�3&Uު���|��Sp�Չ�1��O��j�G9�����C���G^�K[�rT?�^s	.�сIY�׸�%3���Y7��S=d�dsn�]4	�p�%�$!���j@�_��TJ�]�u�`�Ε���;*������d��g�܀�*����w����~�Z���6#gQz�)��8�b�!�8l4=Q���,�-V�}���ηjʈ۪��յ�Jm����obB�,��V�g�<�`~"F���2�����C��Y��7�a6��u��%3�/�+?9�Ϊ�{�rm�9?��曎��(k*���k�����v�=j#�!��E�n�X��[��A)��B����r���LL��=��q��w���Ud����|^�Sп�L�Ӟ���9/;�.,1��8Qr��Y^����v�S�N.ԛ��Kq ����Mp4-�1F��e��}D��*ţ��o�W���U
k#��M}�ڨ׻Y�)��d�_�4�Ja'����۷-%�<�`�W���c�W����tx���XȢe����r�{aL�|�S��*��&}�v[�0� �ȯF�����ȪO�/��Ą��We��9�_W[� CC�{�x���;:����
 �Ŷ�dn;u��c��k)�ӝ�V�3*��_	S<��+e���>@E�=Q�7~C4�*���E` �5�
8xŃ��n!r�\�&a������y�
Q�҉N��ѯ�D���<���86��
^H[��^a����u�߄zW���t�v{�L�go��]r�,ܪY��k��* ��0@����1Ƭ�!3��K�6v���yQS��+�w�൞��G\�|������->�&ftc��׋e7l*�&u�e�4�ː��@l�y��°������*����T����D���"���wJb��#ک+Ek���qy��=�(AV��!�.�'�vdJ�P{{��j����ʒ[�+;��8��u"Y�2�%��s��d9�ٍp���
����� ���nPcA`�����Me��5�,g3����Q��G�k���G:����;�� )�A����^T;�:�O
�(�ʟ��$�� Ϧ�f���87g���$nc���O~2ia���#/9�>4���JՄL�{�_��RN���G�^ˊI
ts�����k!+9&
(��K�,���b�䳳�!W@
�9l�I�U��I��\��X´�g�&������������>�����$�ѿ�+q�މ	i H��ǋ̗KFb|Ŗw�5l����Uc���u^i�!E�_�����p�v:��zg^�K�By4-ħ����� �&rw7C��,�Ǻ��B�#1c�x�����9�&�KNϰ�꫍�z��x��W�`�1����	�cy;[&@�?�p�:A����S���,͍�q*��eӨB� �)e��y��������Rq��nˉ����k�i
��5sq��e�����s,d�~lAC+�'���k�8�q�gq[!7#Q�����	S�|x(.���IET����D��ҏ�LV�F蹢rS������ĭ]�H��>nߪ�)&6�Dժ�����x��q�f�=[�{�]�vrD���ÔB6c�04�ڕ-��T�1���i]@^*��g���r��~�3x(Y��Wc��1��������%L��׫���4���m�}䅀[�c}�f�G!m��*fV���՟#��*�4n�!���y�b� Ò�����,�M`��KWt:P0�� ڸ��G%Y�N��t��?�� :$�nK���F��s�\�s|kBw)5%�)��	ʾD�@�`jm�ϴ����`@�7��P�,�{�E�l�q����V �b�N�����<��n��qrBp`|�s/��ǰs���*!�[p��.��!����S��[!�������7�ȒX�d�d���('4>��cH�fg�#��<�����д�q'9�H������Q�]�(���Z깷p��e��Ҋ��˘>C�kSz>y	�|�L}�#沑j�V���@K����5�
f�煳������`��!"2�:�ͫA1Æ�F�\/#��k��yjQ?|9��[��-M*�$�1;i�?u�L7���asO*�:ꯛ��u�v��ȍM�B1�
T,�*�D+�|�m�wU�ר	=�����br~z]�����ȓ�Q��������}.#�Ϲ-�	V�` p����+]�@�3�"���Xv=��O,x�e/�L��L��/�3ڶ�~�&}v���J�o2qyv;s�x���$2:U����Kk�q��q�����*�gS18����	�"���X�
p�=�)�g 6V�_X��5j��������	�]<>E?��hKI-!&�x&k��Pz�#]�������B8kc��y�����lR�OF
Y��ʓ�\D���6m�����܋��P�u�A[�?WTGZr�O��ef͎Ty�Lߩ���((�$���
���ޡ)�
�s�1T�C�24�)��^��f���1[�ᧉ���]PwM8�}>r��nޱ`I�B�����s�8���
J�.@���#��2��=�V�w�+��^�Ul����;*fJ��U�2�����9����}M�ή��?KY�`f���Ն��������p|��ʂ�"�7w�)-�`=s�{|��:١f��s�t�%ck*A2?�uze���#;��5*�\��\Ｙmi5�()��N?lI�D	�i���F�m�X�
��*���Q{��pVY�s�md+uJx��|HF"]�'����Xx[|_��v}� ea���\D�\��z&�g��Q���ʱ,<��s�-�vz������j�
�\!mJ��?������e���q�u-1ӱp#�5�i�t��<yP���o��`����ϧ;f�ʣ�
4����X)��� 2��-
9	��6v�5�[���(yJ�	!�
CT��i`֡zV|n��8^��0ʭ��jy��qm�����Y��\d�4��bZ2W�Ƃ�$��J��6�Z: ���9���\O�j|��'M����ӛ��=�'��&׃gU*��Fhkf�f�Z$�Ud��4|MW؆�V_ŕ�Qpv��/	�G��m4�|��y�S��PR��m�~6�4tG��q0�N�-�_���?e�Ɖ�@��F���-r��Xr��Ƈ��z�!�Q���:ܱ1\�����Xj`�!��ؤ�ٟ�;W��o��f�Ru9��"�b�ͬ���|*�����"��H����Lh��L5.QڇM2��O��ѯ��9ҵ���@�pOJ���]���=�|��-�
�4#�fY�&=�\����σ���r�L�b��T_������yˢ��?V��R����V _�.��C&��'Z��)f9r�$��{�a� `�GC�b	����#R�H(�s3����W��p;?���H�8�i�M�9�~A�9�p�8Y�l���m<�%4�f$�D�2�ka�Qe����kÛ����-�wiD销������o'%:�J��J�n/k���<��Vs�=�]=�����l�dӗ%�sW��?�m>�n^������^1�M�<&sC#l| ����v�\pL��Wl��Ο��Y
53L�Y�#�T5l��x��ߗIu��m$�WYO~�o/�R�eQӴT�3�,�%�{�r<ˎ~�.-v�C��W�;�L3�[;/%�.^_�fZg���r,�����_9��X�*��]Z�[�kV���R/��e��ׇ�X)������6��B����(z��V�P�d�R/���sA%�޼��HfӇ����X�ф��`�
��������!֙
E߯���Zyd��HQY�DV�yu$ΐ�ȣ��/���5�U�ԋ!{�ZQ��%,�1����]GEx�x&����m���2���Պ韵�7�@kk>�]�k����_1j#�x��!���!n;�oC�<3$��,T0a�$�8�:{#�y(i;�����j4�����L��U����;%ۧZ�1b��DX۫^��3 SԘ�Hބ�8�(�^���+�p��	���E��;ʌ����:r=��3��܋�i��"��Ԁj��ey~��t�>��a�$��oJ�`âk�Y�巀	�C��|#
]�fvS#y,zG6�kQ[�#��㣜~[B�>�׼��@:	m��P8[4��6;2f�@Z����H���t{~F>3#kjO�>��q1� �f��+Z]���G�*�5%�E�J��i��M�'C���(��]�&4#=�Gjm��E%�÷U��U��x���u֖���D	�ڇ�,��\�	1Q�1�:v�%Q,������o��@؇NCy�챁�ƙ��{L X+���+>������O=Sú�*	��\=�׋G^K܇��G���F��,��Uq���L:�}����{.��W��$��L�����Nq�\�+*�Z4�PE�C��#C�ۼ�`
T�ӃY�
,���|v+����@4N,�T
X��y����qWc5M����'��b��)�c*[��l���n0�g�Z&�������?�t8F����
�w~癮'�� M2�	q鵙Jf0P2\��А������\�`�f�\8Qg�M2���.��s���=>c�d?$��7zw�.�H�� ���mT8�4Ą��S�����=�Q���<�')��p���".ߗ7�g����!0:��A�ΐ��a�ҽ;�l��')��jTHT ;*W+C�!
��I��j$�yq�tU�
�[b6$R��^����{�꾏@�;��X�ey!�*,�X�ErF�:�k͇	-��T�� e\g��'���q�5W��&qh���Yr��6�H�t�l�M#��