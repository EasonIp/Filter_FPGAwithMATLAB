��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$���c���D텎��A�/��"ڂ������N-���G�i��B{�ёl�R �O���$��Kv��Y:Fy���Ur�^ٶx�k�f�-gZG�Z,+@��G�����@mz�u������1�PM���|�0	��ӞF�I����\h�7�R -x��ö���m��KQN�����	��ڥ���e�ɚWc9o�^픥��Ƚ}ŞPeO��c1��ÖѰg����[XX�G��vz�ī/�x�}�-�wx�(��$^�~-4R˯O홽�����0�%;t�;PFw&�#N/}��oF�^G�ם$�ڍ��tm)�h�.[Nz�������Ύ1)p3n�p�.[�A��Q���vY���t�]wG	�,��+�����Q���kC�>m�����F�]T۞2+�� #�^�+>�2� �`��{pjnG~��C*(��I�W�+
bh��U�����X-�L�ӽ	_�Z3�Y�r��D���Ͳ^����i�����<��o� ���c��bG��N��!�n�<1���G$������:O y�U�L\�V3V�b3ս�)�"N_]^�b�p��C��G�8�8�o9���("^���	���O�����h}��2��qp��Mb�pqHP��{X�v%�������
\A���z��ɦ� �?{���������S�\x��}��]�YfL��%^`
l �����YSѯ�Nƶ��hׇO�$R�r��qz�{8he��Wj.�%[x4�Qu�9�J�(�j2<c/�Ou������#�+�`��R�q�PLQg�	j�����^��@����N�zia���K�iu�.�l���V� &n�:űu{��Dg:	�o~� ��?�y��鸷��q���a��%�F$���	ڗo�;,��p�?�r����!Ͷ�:'��f��;n��$h���V�ד�u���'�a>���W�*����8��{@�EE,{!�MB���
23G�yF/3эϫB�V㝦��K����0 ޅ>�{��O5w%k���D���ȥ��Ƚ)n�� �LE�ऴ[�	ʔ\�M��BH��� �D(].<�V����%�z��Rh�<U!��38����NhO�ݐl�E	��"i��A#�&�i�>|���>_)�|��k����o���>D�hO��q|�w[ɀ6QĪ�Z
��M���M�Qīh��v�xJѤ������U��1�y��4��o+�r���e�2����J5��g��Ϡ
��jO�d-����@��;��K-���E�!a.k��\̌Xl�"�q��	+)��v�f;�"ctS��h�)�W���/�����-ZwG)l����ޣ
|ڽ�D~1Fٴ��j������E����A�F���0���ԂG]���C� o�g�ho���%� �<�y��n��ǭ҉�	�~��\�]�T���-w؉��q�C��������6-C>�'WfKkz�Կ���o[�c�ӧ��޹�Z��6��A�k~w��1�i�@�_�����Tk�$*Ԗ�-G���K���AJn�����Nׅ\-���y;�v��hH��ٮ4�9ۜ�ڒ#衩9��<�K���4m�:��տD8U��� �<g���z]93�����������s���CZ�-����(��R����N��l&�mp����#/��,�us�$���Ϩ#�2+�����\e��EZ��1��\�������x>��}�����"���h�� �G�h�:˵���D��P�a��>��ON����nxQ| ���e8/��Ɵ����]9��f��~�q�R��\��"��E�Əi�?RE��(K���E�b� ��0�L˔粶q��g#� �ܫ��ہ$H%%�Czw������7�E' '�� ��X(�b�u�n��ܧ��-��Õ%*+%,�o��7�������|kv�Nja�{��a���rߣ�9�$��	�CсIY�{�El�fc^���#�O��H�I��������s��Ƥ�2�0��.��x�a (���cU�$c�tm�KrUa+J�g�
p}H����2gJK��|��	N�R��NC�T�9��I��䡳U����ۇ4�7������r[�����$��򬋸�E�vdP{�٣	��S�c�
)�ĜIl���Y/���f�����ߛ�nq���iw� ��A�X����S�UK�� �Rs��1��ɽ2
SP��]��W������KY��q���O�u�B�ͬ�5<�i����$���pc�΢�����r��ɇ�u��C� @�A?��M(o�����p�{��L&U�o�R�W��`1A��$�Q.�{��V�x}�����P��x#��˪�(۱��!���L�4�2�"����m Љl®��Jҗ77_�P�P͉�Thȉ=h���m>efM�ֈ��:\��dq3�I��=9������21�j�L ,�}Ӆ_��vI�|sJc�^j�ly��XiX}c�-X0vd}���s���;/Ф��Y�mŞ���a��Т�(ݰ�:������Z����n�|�4L
�w�XnX�o��]����&_��e�x�=��lܯ�6��U�S1�Z���>p�	�`v_�F���4�?�ґI�z����t�n6����/ґ�r�芥d[(2Di��:�Q�\*����Y�����Hv���?ɛ ��8�D(}��C��=����1��qms���@yYS�x���+=i���K����FruCA����<Z��+%P�{�z�PE�qoY�1dәOT&�����s����3�Pļ��]�/�+9�5-�U]��m[@Ad�4T��eb
H�3����:��C��Q}4	�����0��(�m׹Y|��-V�H
,Q䇄Sl�U��	e���)n��ܬH(��A"�I1�}�w�V�@,�[���{���� ������@���.�d�)�hm3d�i�ɨ���6�Q�2��׋O˹�����,?-+*î���PSx��m�)ԐqB�e�;hj����Y���>�k���]|n�L�H��u��ؙ��9�=#A=��8%CÝ���VXq�>�����'�b�EC5�@3��M$�>_V�A���	�����f+��n�����
 x�����Cdg� ���<3�Ll�����;}�n��+1��΢w��͂p�v���N8$�ղ_����6В	��w<՟d+��	�o����`���R��@}
3�kw�Bj��A���i������^�qֈHԜ�U�{d�w7D5�]9�׬c�2F=��A,�#�n�(�XnH���߉e��g��X,�:2J���1q5C�r�[`�'1��x�l��_* �j"RD��Ƒ`&�8(�	�O�/����2�ǎ�����
nٮfLy�kҢHO�!�0F�GE���1�´�z�>N�hF�I�^�e�C��_��c<_�6���y��Vdd>�%4�0Nhq���s��3�f�12j�`�>PʍG�m�mZ�?�U��� Bq�i���f��[ϐHK����e��W�&���}E�X���*h�y�QN���{�~�;��c�`|��	�Yu�dZ��s�yTi������	yp]����oi��@/�<7x���`�T
�MȰ9០�f�z��h�m�ɦ�R	 R��T�[۳��
C��:��R�M�gٖ�*t@�FldM���fE0�����������)\O��<�^����J%�I�7>*���.r�GA� 	�k6ĩL���wjF��7˴��|����T9%"�R��3צ�麟���y2]�8����:� E�s�CH�4,�3JW���G�죵9�٭����?Y����%����q���_��Z[{t��$�2b!>��sj&5�U7Q���V���`���E����S[���	.R��;���4Q&Jj�:�"���,��#>��tϵXcm$�T�0�\�����l�]2UQG���r��-�g/��>��o-��#v���
� ��&�'p��?������NM�'�񜚩�&
7��s3�Ŀ����G�� �}�R��(q�Ű��3��)�=�t�m�xP|A�1�FS}n�JO�B�����t��Mi*�~� |�"o:2g����@u��P,^�FF3hD�2���x���Ox�ZƟ7;�^���!Z�O���Io	�IY� ;�f�7=�GBS 9u��򋦊gown6��_�b~rw�Bi}d����2Z�%=��l��k�q.�n+�����q�$kh�
-D����>��'��BY)�#cǩ���K���./[7�*�_�vв��
�d�v�n�b;�Q������E���h�бj Q�#-���G�8�	�y��3_����us�N�k��ꗱ�f���&�k�2�.�]�s�� 8 �&8d]���]�'R`'>��J�IAw����hc&{�-:����Q����A���1lAn��7��l��Jq.-�ѷ�j2�~D	�"�4�yPK$�֢{\�ݧ�/DҐ>����o�����||���6��!�t�q�sꔔf_< ��E��ǆ�_	�.�׭�t�e�����ϭ~z��uy�Ű�%�1�U&�~N�H�L�%��c�"X���إbcՂ*��t/�WIES�L��;��L�u*(#�ɚ�t�.�{Jc�z�z�p�Ye��Bo=C��
�ȱCΥY�����ٮ`>O�Lָ��;a�.hj�K�[�{��G��&_d�\d"^���`SQ%'���4h����I�b�~�,�E��XJ��;�oFhr��=o��
Ӑ8�T��I�3�˖���Cˊ���~O\�"���%%�;_R|~r�|$e:���&�'P^����ǝN������E(�.
�ɒ��80) ���O'�y�r������{�Se����wHRn��1>D�)z1$ ��!��/H�"K��׫hS���s�%�EL���*�����7�I�osPYF#�DP(�,d�=���{԰���E�E�W�R�V����=	G���	��"�L29JJJ�2]c������V8�NY�d����B����
s���A-�[��ܒ��&��K�jh�����F�4S�QÃE��C7����*��x�ͮc.'o,��������ǆ��?胮R�G*������t?�u����'����%׻�����������Ϝ�(@������l�&h�q0���c�[b���ցLq �e'Y�����ŋGHi]�)>�����!��*�� �^�F?>ѵ^�D�7����̂a�|��G\���	�їgh�3'�~r�ۉB�����^��$6J�@�i��_�ڇ��l�MO�����
 ͓�9���i'	�`ȁ޽�0�A+_ɥbH��O ���7Ǳ���X-i3���@��͟�1�n��3үD34VC���G�es��L�ȍ��p=�c��V%F8�n;�� Lj�6)h�P�AD/ZQg̐T'bX��`e#xX�\$�@#��X1��Ɋ�޴��C
/���eM��g�K	�9us�Ra��j��_}�(δ�D�=#r-pz0�/nj�ݓ���A��B�I��8�f�y|qZa�{�J���L�������O��s��sj���jH"ҧ�c�V;��L,�Aoth�<�ސZ�}�|�2�M���͘����nL{YOy�w��ڜț��]t =�Z�ݛ�� 3��ʋ+����G�<�%���^# DA>�Ez��c4#�N5L
�%Y8B�R��
d��ُ3��� 1��u_����\q�|k&Íl�í���|��k��I���0�����G�6Q$He�4�Π�ʪ���9*�-/O<��*���,��-��9�RH�DR���p+�yU�(�f�եe|ԝ=m�I�R!Lk��dm��1��V��Á�P���N8��J�fWU�z��&�5�!��E��Qt�<;>�5s�e����K_���$8�4���������%�f��0o�e0�$�x�_2B���;0H��&Tq��{�i���<�cHշ6�4�5o��@5�e-f��び2��8v����eN纴s�S�R�".���C��A��E�?�J�M��"�
�)UN�9:;n
���<���=�����F��l���_��Vl|�tSrRpK�v��v�+�T:Ӑ��h�J �=���)�q=�T��<!Q�|���{�A�{�A[���K�_�6�U�!d�EZp��m��-Zm����ܜ'^�t��� ��w$���
�Q��E�5GH�t�+ P���;�ܴ��Vt�)�� ��*8aGJ �h�v�_~v���<qX�;/-/��no���e���J
����<�]�6��^�B�L���46ȹK�o�?F��@I8�Q��ڷ(��#�T�׳��]���ƞ܎�7�������O,�h�H填�?8t��(X�1T���`���z��ɷ�\���p���	�F~���P��t��o��@a��$�7���g���Ś��L{�S&`�I@O��Ј�]��t�������ޕ7�i�(���~*8�;x��YF�k� #ե�ӕ��6+��V-���
�^i��ݪ����2����>%U���<����M"t��]>����=�<j&AE����F�y��W'V\��]����.��״��&`M(��2%��`�O���� �������lT��'��E�C�zBn�L�-�)`�c<&I��t��h1�E0�W���lc� .X���W� ��^�����s�!��ync#7��}��NV�$��FM��\�k�����WW���c�>4ml��>�6��73��,�|�l_L&O>k-�>2Iӫ��S��5�MȽϟ�x��0c�oH�喏4��k�\�s��	�/��W�l��!9＾O�Q:�le�0�?׌�}�"f���p�wg��4�s1T�"��D��f���������FJ�F�ڵk�ҝ$*�{��`�6d�iwnD�2<�k2�F̡	�טb꼥�$��1�ɟ�Y�?cJ?���,!�2�H�mu����/
y}��+�.К�� UM�b����尳�%��]�wK��LI�(���o�M�g4���c�x�%����1�v�%�`�W�߂Ő���SZ�{�fi�9�c���%����S�3{ƼJE�����^��_�,j6���e4^XJ{X��� �P���M�8���\`�����iD�T�x�*)MX
�x(e��}Ҽ|G$J
\��8Y�5 �v�߫��'��4H9��h	�5��28�;P"kχv��D�R�I�PQ&�d��<��a�-p~A)��a�k�6�˩�֚���8<l�\��:�f�}���ڕ�]����I�)8�&ʍ^W�b*zUe��f��Km
�-��^�:��.��x��yu7��Xز�F��;�-Pb#�S����ɇ��xC�41:��Vr9�v�[��q��ui��K��j�MĊ-�"��p�X�wT�f�EnPtvvٱ<<�䬰���Z���d��z�����`�`�r�n?B�|�((�Ԅ�pՀ<�T����q������f�&��pI��"���+\p�Į��o��N��Z�mb�x���=��(7.&����_ ���R��#���J�e��u�޺a:{Q:Ji.�q^rT#(��3{���ݣ�I$�I(�'ؠ�����k[گ�yv+̨��ҍ�R
՝���c��&�@�����BŌjw�)@`E���S�j@��CS�����u��@Yj�0�[�ۄ1�^�p�����L]-#�� ���D��~�#��'�Z=�D�7�WH6�"��D6kc�*�H�SЄz+&ƙJ��?i�8��8������p��_���Θ�B��k�ʧ�7n�S� �� �&.�(�y��6�W{��)��R����~�(S�j�{pN�3�۪?3d�Zd�|�!j>��$��M��8�Y2j+��j.&���@5&� ]����1=��Gl�"����o���;4+]������z�.�\�&;�(X�VԳ�{,S`��$휒c���hUi��El���ڎ���D/��r�2}��F>�� r���~Z�ZgNֆV�?7�j�����80����h��z�@�����*[�����N�p������q_�Z������z���O��H�qb�����^�kR���Ľ��\'#�i�1�D����.�j���v��b�eA��gW%xm6��q�D*�k��>�{�=���
�w����oˊtH|癶�l�A=�tVHR�e����{ ��L�e�l
�>u�+���?���J��� ��3�"����UѬ2�	脰�v��D�'|�
��S�0=�y;/D9sF�g����x��i*����i8���
	�L���h7����+�V�W�:Z]�9숳��x�Ŭ�IU��ub�Na���H@R�P��09��_f?������*����tP����;�y\�I=�V�`7�U A��1�c��cث�']_�㽼X��r����U4�W(�o�TT�k���4�#4ݑ�,�4r����]}:~�_-�dv�jaT�g�yG��? ����,ø��_ذ��,�����cA(큭�`�G�����q�N=��H6LWm���C4�9H*��C�OI�\��J_W+����F�����6���F��K�hx�+���譧��OS"����+�d����V,�&8Z�7���Z����;��x�:
�Ӡw�q%)����]vC��b�����Qؔ@#��t����""�����;��n�(���RƓl�w������8��9�w�a�>$��d��N�ڴ~S�$���z
w.X����C��&�ux[� �.'��U㜳<�?nL�X~x���1a�[H?t�H+y0b��i��\�ҙ���Φ��՝����3�}($��	�=f�g�Rq����"���bC��f,7���I5�l���rf�:�� 	��u�7o8!��CwECҸ#�o�&�'������S��	�^�9"՟]��$=���K�ğ�G�.�d���0����*�����!?L�)��c�)�G�<�J�Z�!vb�N��,�\�uQ����ty&��DS�0�8p�JM��/f�1W	8��ݛ����5����N�|�'���u{?X(�C%�"�F�=I���tpFŦzǢ
�U��.w��<@�T��'�?)��l�r��-��e�-�_}x#���g�U	�G�hL��E�;��kG$0��聿@��,��p|O�=�f"�5���ژ��}e5{%��j`sx�k�Ǝ*�����5l�k8�3�i��x��=��Dk��4�P5W�MaM

��~�%^gؔ�R�@�����'��1mZ�cyb�lk���F�q�wy%A���Bnhu��5������ӑ�a\���+����k|t����-���\���K!����*�����Iޑ�N��DۧiL��N�a.�A��8� Jf2���)��R	�h��}�f?�Ѹ�o��u��Hf�:����&��u�|y��Lx��D����c��]_X�xlAn�4 ScX�0iᰲ��V{=��~��>]s�zn2�?0<�t�v��M�Ԏ]{������J�{cN�ymYj��e��o=��	3�@��
��t�eև:$5��TH<�֕�w,_��CmZ��z�d��^�Sg��5�V~5�?(�B`�7�4����w8˩5�Z)�E+��*u���U���60�O!�sk�]H�yGK-=�g&+����~��@@�_�����P0U��\����w�z:�Q���h�(7�#�J2�Q}��P�|�8B��gl�"�\\�ˍ����Ey<~�p�����ű0����	�<�����o�d�4
,5>\�R���m~��k����-oG;���e�,�Z��0]���844��PP�A����%5���j�[�WG-�b}��:c�#��Ba��� �B[]9G�'%�R�V��[�Z����V[vaL��}�z��RW�����di1�x:mz՗Oۓ���Z\�*�<ȉh��}�B����3���~wJ��B��2��z�����􄿔>��@�i,�	M����L��g{��&��FP	i�d��`�!�?#i���k>*.H����L��-��^Qv��؝t.��;F��T�?c����o�X��<
&����W�/4T"X�t2���P��$�V0�@�St�께�WʤX��̳� ~CĊ<9bb����N{|xw���s�L�6��+Du\�%�3���,��!2GY b�پ�7A�,���-�U��ݍͲ?����>�����͝�0JS�A[�-��j
�똨$h/�X��K�7��M�A��Z�h5�^Z���4*���q�|2 ��Ro�4P���h���:�
�n��4p�D�A��@�=�o�4�`{�c���Y��\�u���>Q��	:��ٵt*0��-��V�U�,m����gC`��A���i�����`f�Q6����l�[�*���5�#Ls7f%���CıP#?O��.E�U�mq*!�-�9o�_�՚�׾0��R�q�C#�q�]��~WpWߒ�\w y����9�ʇ���y0m
C!�|������k����]l9���G&2VD��|2٘u,xJ�p ������0m��;Q������1D lz�Uh�)T9n��	Z�T�JKp�&��/�_$V�6�N���b�`��ǅ���G�;�x��� �^/ �/E�b,Px�f8��ؒ�139��`�e�%�38���q�����R�\�S
���AƟ)).���Z��r�D]z����=�'*��q-���c�� ����H�����K�%!��k�A5Z8f�8��3�Br�=��U��Ct)j����x~�	u�,���*P�pL��,�q��H�4�h����8ю�H�N��I�5��b��4�|�$��E� ���`e0����鄥�����ߐ�_��z=�L��I��������M��FcP�{�/�mJ"�Q��zƙ���u3�A��Y���̬�u�+��Q8i+n�3a
���+aH4s��cp�b���c�) ��.�B�¨D�ݣ�-�ThEZi!�Dː 7�� +�zڝ?���x��~Eg�����2�6^�O�6�}C��¸�I)c-'�;�	`Θ8��ևgߔ jt����ܝ�ɾ����ɞ�`�7��tY1�G��v�c�'����'ߵ:�=�>U<`�et��=�4%|?e;���S�_ʓ��6��$��:��Aڗp�N@L���vnp�c&r�akm���mJm�Q����-O��m��R��R�g)�<�}C��.����0߽Q�]��U�3dG/D��w���R��%1pb��}/��z� lN��C*�A,k-n��;#���(�~%(Q���|a�����Bs�X9�RlAΩ��)��%��O �̙6^0������[�ڛ�w��숐s���RV$��ԷEyAA)�m�Ӊf���,���;_,�%��`����g�x����8"9v%���[p:� ��ʡ��n����