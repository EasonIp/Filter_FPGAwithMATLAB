��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e�	X�Dy1V.Tٵ���E�n��i]5�h������5�xA�� �d p���h�t�?|�q����b2į| ��ע���8��:���y�HO_����T�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬��q��lv�ӥqA��I�vݼ�}m/���GޕN>�ݳ)��S����!11������䌴K������8�9;�	&`��q8Å�U��@i��`9T���_T`��:3�>�T$1+"�R�)� �=*��4W�P%��.����'�eA
�\7�4�$ʕ@a(���$r*)�b���)�v%Y���nʢ1k	�nG��y�k�nOG���?a���?�R!	�jp�V!X_���1@��!�W��~VXn^�(�B�S�2�j��c�Y��?R@���t��d��.�Z6<�+���=� *h�I�G�>�;M�-�UY��'h�)4r�a?�yɦ\��|�Ǽ,�tТn��T2��%]���6�\��i��~i�&G!f_ѯ�Y�����1�sg9*8c(`ܨow!_]݉i'�+V��T�0CS�((�������k<�Zӟ�.g���?��âE��uaD,s��f�}Ht�����=����й��u��34T�~ӺZ��ԄL6�p�#�)�
��,	]�Oduj3ʫ1,>��b��JoP�n��S�)�K�<�D	��g�p8 �sGySU�!����,Tם�,�%��IV)�q����y-�<[կ���ZT��n֘�-���,��}R��Qx0C�<;v.bp�'X�50�bG���	�H֮'H����8����\O;��MV�Oإ4�7�؅+�]����f&�3�;�CI�'*��eU��H��T%R����5:=��[�w��w/v�&/��[��If&�.1!~���S��k�q���I�6ؘ��k&��:�*�� ���H� ��w-��@f���@\�%.�N�֎A�.v%O3I�{���h�CPFt���� ɰ2���u�C��������})ԷE�}	s�I:dzW/Y��7ns�l���;/͕:Xuv�*>|S�>`�<lmШ�c9��&��&��k�Q4Q���m�=y���b'@�gLX�o3��N1-��݀f��م--t84�W#��$Xv�L�W���L���Qy�cq*��t �z?DS$��t������)�;4,Ē��,Zۃ؟��T��[� {��F(�KQ�@,
��,�s,vΰ]�Ķ�dDH�wKD�ʘ�#���?�m�:<0˨�ӛD����[.� ��;@�BCs<m�
�6\�h��,�Ɵ,��T�2r
͇��gS��~J*�SlU�>��Z�d{*�He����=��N����"a6����Aް_<�jCn���7�FH�(�� U�$���R|�`�����8��U�E���5l�����>g��n0�ݣ'[�$�*=QX7*87���p��7ۉ��ߧKX��a�����z�����I���")6KR���O�"U��2�`��ڎYݷ:���*V]z�����Cw?)S�O�(NW�v���پ���'F����F��X8Du�H�*�Lh�b��>�1�J���Ш�*�h�`"���.~�eb�>e��-m�F��)�S����݇��+��ߺ�7���N��;['�{�nY��+��/ʈ-���e^�$�8e%��<�q����>��[f�'l�w�gs�u���1T�|���YuE!�2klLee��K^U~�D��{�V!T@*������ImB[���\�x[J@{��6mܥy�v�k�n*�a��ӁS����"BI�ef\�l"��ϕ�)�{ٷٳx���00�䱵/7$N+�6(��t<�!���6��9�i!�O!f~�7�D�C��OC^�l{�ݿ����~m|�8��:�%�Lg:�pw$�s�v�Jâ:j� �t6L��-�Uqi����W�&�̑��hߺ�G�� x�u��z����0�K���y�,��*�8��j�W(��"����o��a��ͥ�b�QF��zJ�0��8bX� [�[�[J�M%^x]D�tO~����^*d��aa�����J,v�+�Ȇ�$�j"}����K��E ��Pؠ���a��4���0˅'���D�dU�Z�IH�?��}+6�oq`0�z��z�]y�J�|�L���=1��GA`�GT-��w'�4�LJRȄ�.Wۆ#��5���vrU̐Y�t�`�<��u�&��C�G2�����Zx|����P���j�~�����c�**��a��}�NN�ff��^nj$������M��w�{�Q��/��V�!���fc�4������FDڂ�w$��Q�o�¹���jl�%Nq�Bd0�oZH���C����{OZ�q�ء�b�aJF.B�I����AT}g�����:c�Y��J�~��&�axV5���J:ጛm4y���4��f���=�fX:7��iِ�	����I#j���I��bCr�� ���#�Aώ�O�
�k���%Ad�{�����h��Ea>m��{�o�)�=+*�h�TĪƂ\Cv�?mɷ����r`� 6:�Y��kfϽIU�=����Q�������!�°����VDqk]Ue愿���$S���S��d�V�"��7�:�I2$ ]+�H�^�~���5��
�R���X_�N5�IT������Ce�ß�N��HמX���WvX��}�Tr;���^�U�tmW;*\�'ƵV�]G���*��ѐ�/g��~)KG�Ǵ���w�p�w�R
={6.̼�-ͨ�;���C�|�}JN�M��1�r���{jgD<L~�k6��?+�%�!�p�9/x齨Ԍ 7��^�0�<[�����ޙI�_&����	{�{���g.��Oo��F1�Y<(�w�X_V��xcf�ƪ��g��bS�M���mݓu�
&��;�����������}���؆O�ѝ����Ф��T�	��_h�k B��y�$�E6�~�3g�CN���"5u��Q�
Zw�s�'	$c���>,gS$C����
�;_�w�*OK��\I¿���H���a���f�l
��0���' �:
�K�r�ήA!��(��[��# ��.��ɻ ⷣ�D��c�x���u�T�$^�=�.p�m]���q�ڀ)���z�������a-�b+t�(�}�+�8�����'˭���đ�;�ò�-˭��@�kۂ�ʹ����j�z����卼VRDM��I%1��\�ʍb���5�G�D�㷴&*ц�z���<_�_�6��]e�5U�S/�d-j�-���n��4ƭ�\֣;������G�p�X#a�W��Ɵ��1�gn�y�e���q�T����I���o��a�͉[ы���w� ���Ʈ}�2a߽���b��wdi�8�ZH��B�83Wݞn$�I����31>��I�(�$����d!V7����P�k���͏���������]f3��O�0���-�ބYM?��X���<��n
)����>�9q����D#c�cT��������|W�|8�_�����$_�bp>c�6!kD��H��I{�^2#�p�d~�ij��8J\	�>Q��,�K���TS�aE��ap���H��Q����^��~%[��h��m��wk�
��Je]+x�D��L���K˩��O#\��7~��A�~�w1ptc�з�Y�O�E��kж��m�ԥwm�5�\�k�F�ɧp��Ī�M�L�͋X����5���w�R{��4��:�@���8{	Ԭ�T�N]��4_�v�b���.ج]��q��K��i�����,��D��L�:�0l݃kG�������8�KA�|9~]nZ���o�LnDC�`��i:�^��B�g�S@�m_϶&M������(�4���ͅ ����]���RY�Z���K[td��Gt/�tF+�(��i]%�'�(�f�L�-)%σ���]�mC��Zoc�9�!��R����⟉�Q1Iq�*11*e��m�����]���Iەٳ�l(4��R�h�ŚÙ�vZ6'���1St+EHX��ހ��F�j�_����~&;E�fW�X�Q��l3�ɻ���^Tނb/*�Dx�`��`����lI�~~�6 9#�$������Ox2n<�`\�h��ҧu���[<�b���`$��ĺ5���G5��7	S*�o�%2���@o	�7I�L��H=U��#�����4_+ �7�b�S${�ڴ��C�������.T����yR�3�<��#��-ـ����1��Z,W{D���š�Zά�4\*�	6�S�>�s��Ir�X�/�"����U�tm\���.��MbD�H@0�*ہ�X�>�E ����;_���4��:G��Q�O%�J�N�W���Q�e��%���]�z��1��gjL;=\hW�� T7������=�'����=���	zƫ�>KB�{�?� ��<Y��	������.u�L��;�Y �D�j�Ū6'O��[�q�����ARc����!�k9TRZ�S�'�=�H�p��h� z��29^D���T}���sE�}	dc
[IV�2�-���?��|j��8o6���h.l�������$����-��'U���@�S��oN>q�n���4��2A�y�{Ԃs�l���F�:+�X��AP�9 ���Մ����������.�$ڠ��̭^��EE�ڲxd,��d�/ zD/��c~k����o�� �+Ec�YE�P6��\X�9�j��!�2�L�Ce����^UԘ��1�"�D���K�'��J���A�N/?=g�m�k[�I 
i���r<Ncv׮�YY|��t�M(�+�Ƒ�n��ۼ�H;-��D寷�8���`gt���k�0��Q��sN�(sg>8�پ)S�F��c�z���d=�{kA�e*�L?&p9��o�vqY���׵���7�j�X��;�k�b���ܡ����	[�vT �~�m�W��2�K]�b(�9��	(�hwr`�ߘ\����v�:T���I��CY�9�8�����ő���4/g����s�Z���`���u8䚗:s�D����#t�ڡv�
�Vn(�L6���G�m�+[��w���p�kET �9f�d*��J�ĸ�[�O���:yx�Z�Re}���	���3}����ׄKJ���jQC�!�����O0��8��6^�� �z;�+�^�\���'�3 w���sFy�q u�;Jz���,����`2��}��n��e��E�&��(���NTj����X�?�!pw���t��
��ǈ���j�_A�R ��%2/l���T$C(����/�@��(��)�����2��&��]	�p��[:3�$I��y�5x�hK�"�@��{	|��6���g4�Ǳ�T�k�[����%�\�]E@���]�X�I�+�(so�����	/���|������Լm�@9����e2Bh��S����@#��i	�6�P��(s���U7���{�����:��p� �?��u������f����Q�2�'�z�#*��ܤ &op&t�\�'к��,7��02/�ԅ䵁�zP]��}�)-�`n��]�o��P���#k� y�C���q�Dl�M��E���z��3�_��nN0���2k>u��AP��%ܥQY;h�.�M���������b;�V����K��D��ȟkEd=*��#ӓ���mm,��6�	_�a��oS�1�̵c	�Ņ�_�,l�c��eNZwn��}�#��;�%9W.qQR�^١��b���m<��(�̟��~��#O�8��B�G�e����|1)�մ��A���d�ܞ�)J��{�!��٧�5�)w���Mr�P*6� �H�O����땕��o��yV�_�������3�������"_L"��]�
��	U��I���\��7����g>���*N�5�1M:xgs� �Ѩ�s��ʴ"�`W��a��2*M
���."|<�$\��v"���%	�P�c�`������&0xH�/��p)>��d�s_"����IQS��%�4X��E'�����#yÆ|c��q.%u����<u��0�T+����÷L�ᯜ���Pv
�ǲ���X�M����i��z#�hD��$N[L��ξpy�U�񠯠�Ӯ�\��:3���#d��;| C�{Lf�I���<q�M�Ъ������8�q����oۮ��JI�(�J]	*E�~m�����g�5�͜��4%��%���&��
aC:/2���R�,�ٳ��q�?X����fK�O<٫�njȁM{U�:�+�q֙�9Vv.�|F"��1��u4����ށU�Q���妎��a9Su���,�+C��H�k����^χ�޹�yvS9f ڒIO��:s4R���"5���X�o��Z,�4 &�b���#�i��`C{sC���qP=]�U([P�M��F���u7�O���s0�gxTv��t\P�y�ʀ4�gښ�mh�bV�]0�jQ58�Q�� ^y24%���P'p<p�'e�u���YE��A"X�&�X'4��5�E��@Oΐ�xeHL]e���~flZL�މ�Uv`���M����&9I6ƪ�(��!�*��V�·��I�[��� ��;@�"E睞G�'��|���;=���l�����Haι�F���݉�3�lDa��Wa�C|qWf3_*<Wv���}1�~@��9Δ��+��ml������NoC�2|j���8�`�2���g������1�qX�n�E��X�H�M�gJ1���1�Ƞ�Y�BSA��9ĕ�Az@�בq{)�K�5�ԟy34��:D������?@����F0��G�yף�����d	CZ+>�@k������~���o��m���Q�}q��'�M0���ʡ��E�Ґ����3��E�i"��v��+�<_�s�2%��on����H���0������^�'τ�K�+"�;g�>L�o8�穽��/T� NH�p�ߙq������Z�R��"�F��n��ϋ�"�zJqq���Y��{-As����ި�S�D��A��|�j���zM^�A�G}�H@E&�f�ȕT���� nE�H���|�z�3C��ُ���|�
Z���fC��s0�2r�� qӒ̬�=��n��{ڦ��/B��Y>q6@�H&��� 1;�oq��Tq:J� �L�w];�u��б�U�;�Pj+��sr������
�W��1��G/ ~k9+�+Un�^΅���BH����R�����c�+HbZ%ls5�G�K��5Ʃ��f�:N�"x��
��NĬ��͛OV�T���0�$"��\�n�	�a�`_����^��6����)���љD4'��8�:�z�{�����<cd,�9��ZA�c�k�.4M7SA���0�����[��3Yud~cD�X��Yu��.`����c�c �MC�Gl	#�n~�j�����~Tͯ�szE����|Q=�,�n_;�mu>��!�����OBK�1x�}�5�i���aԏ%�ȶ���`-ٓ�6.�r�I�X,"��.)�~�!�V�i >��6/��5��Z6���2��sκc'�c���=��N��V<�<+C��<D�\]���uQ�b{j���Bس�25��7�%7����`�F��k"�}jb�T�1����/u$���>�����P���As�=����i{�`�H�^�&��m�<V�5S���۳<2�Z�<�1�dA� �{��:�=At'�?`���AA_ �m�V�ldKA�-��^��Ws�0�3��WoQ����#@�k��W"�+g�t�(�#Wf��U�XѤ�c�Ͳ����9�/t��n�2Y��'�5	>��eM��;�+O���f�(�8���1�Kч|��_0.e��+�����&�`_+��Ig��p�WaK@���M"]�wC��F���d[&[0ݟ���Ԫ%�: ��T>}Bb<��<����L�C��b��h�u�q�c�H>W�u��	�����cʀ�^n���j��N'Z�r{y9��1��z�w�D�W�߯#&�Һo9rF&�=�KJ�:��<s�1��VC�+� h�H�ZK�1r�A����53UAQG�MZ�&�~��I+@rL�#�2�f�U�/��N.�E�ȫ�|�t)|�f�Q.S.н��Z6�kΉ�a~m�^X�fc�	1ޓ��}z�%~��%��X��-���E�d��T�k]D��
����!�0aJ���.X�6�?Q��b�����\v��8H�ƃ	L�s�����i{�K�c��|&g�� ¼0ÝO�<��Q$c��A�U�oQM�=���ﻦ˳�?2��ߪ��F�V�,��u��E�j�ZsZZ�'���ք���mS?wI�)K:8����3mZ��7�ext�Մ�����GI�*�Q�>9��П�>�3N����:Z<x��L=��Y��Y&�[��}�Q�V�}r=�6_����N�%c�Z]����"�k�6�a��9�Ggȁr|��3�*��>�kC���jD�Tq�_��L�!@�R'k���әzjcٱ�7�_R�|t+�P+e�Z���{�kj��~�v%�~M�c�af�<1_�X�؟��rH�	�N��\b��~���~gX��p���vg�¯B�9�,_Jt�;�f
 Τ�ؓ E �����D=��|W{��ޒAh�O�i=I��U�,��|�,>X�6��G�]����1e������n��ns�H�k�s��R�ɲ2Gn��i�D
f8�I�2�9�����
���];F=d�QfdU�>�bl���fO�S�a����wz�e=&ux$m�m2.b3��j|�&�M��ag0�;�3F<l*cf�; �K�^���T�jm�O�дL|�o�����@�FSx��<�7y��^9����8̞P�k�Un���6�J%M'h@~�eH���0"EӠ���6�u,F�\�c�;�N�/7.Մ�7����b+$�W{sk��J�ލ�n�˫Bc m�pT�hott�hL���{��g�3�)��Ap��:4q�wQy�:�Ee��y�6Cݠ~�a�!�i�O'�Y:��17���g�z�Uv����L�T�\��c���5�#ȆЙM�E�hƕg��D9��F�����x��d�鱜�R�0�N�(ads���P��,��rR�We��9	0��-Y(O�Z�%�͙GM7L���XOe��x��ym]���t��l^Vt��'W��w� ���#k*�z�PC�����)��������r� ���<Y�!�v��󏦛�Z"\��x��3Hy��1��8f�T��4����J�<ў�������0JhEV}G0�\��Q����/�+u�z5� RlmuF'w��\�A&�-��5�������j�$3ys&��|�l�4  �����A�lA�$xN���ٗ�,.�q��u���8VgK��;�ɞ��KRKM-D���e�O����b&�yW���_썜aD]����j��)���I���4v<!Wr��!O:#�)@f��58��f�O��]��:G�&nPP��~{[�`��|��;}3��?:D��~��|��fܑjO��TjZ9��?��%�b�饆|j����4-�	K�ܐ���v4Ͼ� .��һ�q�s���j�����;2�F�%=k"�M����ڳ�y��+
���
UȬ��� M>%ﮜ�	HM$�(�K�����Ö�?��\"���g�~��Ԑ	���xr���q-��G�ڃ7ע��u6�C�P	<2��;�*=�!o��h��L�3)�&9~m���4�XS"�A7�x_ԇ@@84Ɂ������"�NE�=T@E;1-ڮ�s���ｺ��B#�GAM`��R��Xz|�}_����)\�2����	�'j��������u�ʲ�5�?���^X��>/Ы���������F��%���X�N��xc��=-ovq����FE<��J����<�y�m�`���r�[��]vj��!c�gk�����IM�W���I�3��x�wЪ�柯�2h#x�����aVS:�����+h�>��E�����{��Ƙf�D�A�>,�W�5� �Q@�®K�gW�1֜�Be��G?�Lߞ�iv����v�?��y�Z&��c?���(!��b�V���wl����tB:�@Ӧ?�4#�ӗ���@��R�6V�j�>�I��� M�$�DЂ3YF�N����4X��iE��'������&;M�^O_nc�ǐ�΍�%`��7 }=��n�1*�7IQ�[�CÛ�ÑF�kHF��.������ѓ�Nb�?C~ 9�
D-���lW+�J0�y���sT�r7�����n�P��b��0�E��~S�\�V�-B[!��v)Jҹ'js�����Q&��M)��k[0�{����zF�3�����Mя��x[M���R�aٜ��~������Js���.9u�5�	)���Hܹ�\��r"�eGh��i�7��|�Ȩ-�%��tg\�LZ�v�h�� ���=Ϳ��
.�௬E����~]~l2��� �*6��-��qD�nĉ0�[V��!K����57#���˜���H��?�7��r(i�F�+U7��]�iI�p�A2�B����Wd��f�k���ii����GL�'�-ٟڿD|Z|�:{J�c�i��>�Ҙ eo'�yE�E�A!Kw�{���V1��wh�V*�Hf̱�7jw��EU�5�pV�0P�MI��@�B��lS�k���}��H��DM}\��G�+�G<�o�k�	�����)�@IјY�>ʇÙ���^y��\��>O	��e�B�J�:�3DE���דh��|�.L�^1�=��(k�h�w�"x�(�Z���?�����]_2��K=��m+eE�3�R���`�!�}ΠA�G�췺eäIX"n�YH9j���B�����}x^?�͇ȡ���ÎAX=I����WQ$�/�A��_����ak�h���N<�S��1t�&�!V>��=4d"���|�� �L;��Y�D�ۅ#�{�rwR�� ���#��i3`���yXA��|Y�_[�D��f�(B/#�B���ݛ}^{��]l��6�������z�?�1�oَ�4��k<���g!9}�B���+8��7Vf Q�F������)9.-g+9焙t��g��0B��ke��s�1����X���6k@n�T��X�$�SI���\�-WU���|Ǯ���L����T������'c	_��DAx#Q�g���;"]�fF�q8~�J�0$�0��	C��e�,}0��'�6�/\Xr��{j5�v�]�y��bk��Q�r�"�Tw0L�޷��ȴ�'���4�K�"�(i`���A����.�H�R�X�`�_#����l��	�t^ڌ<k~-������p&��t�����q'�Q�[����l}��t�����5�P��p'����{uRZ�5b<�=����l��Eo$����hfD�C�&�>����"4[���3�l}�����!���Ŕ�3�3�o)�}�@�骻9� B���ܕ���kHpO��mY��LN������
f��҃?~�L\�����H����[ɩD�ŗ�R��k<�M�%��jZ)Ʃ�B2����t{CE��]R�1�I[���A�f2�>�9��R�"��*ݱ
CKm��1��}�Z�Jr�Ю�#�z�#����A��w�g�_nM��ics� �sB��F�s�'�a��-L;����o>O�������������b���4�*ۻ��/bb��ߖ��7g:Bx���M~3B�R�7�>)vM[�a�U�~�\� ���նQJM�Q%�)�z���\e�K���zB_ַȪ8�97.diW9=�S���sA���
�t��-�Q���f&l4�Q:ݏ��(_=506���jm�kr���}q��^e�̥�	^�����E� �Z�.�5���e8��L󿋒�HL5���~�EL�����(d��]&C�����
�O��ݓ��2S%�`�`�z�C���cU�u��GE\�r�Lx�� ݦ}��zxo�_�K/
;p������ȱ�7�!�Ҋ ���t�xƤ?����k��8����@m����ߊ��;J��%�	7���������;y\�����r�Szs
��	t��%��n�\,:�pn�Y�2:P1-�7�cr����[�K|�Tk{�E��!��h�;U4p����:��{F��f@�S���a��=��gXI�+�����կÁ՟�Ǣ�d8�:b&N�A��I�DbTA�z���� �%k�jf9>%�#��Xt����E��$ɁpV!�����ZF�4/]�`�A�G5h5�X��w{RLD++�mn �Q��ز�rW)[Qp��FbX�3C�0����+˸aӹ�Gi��T�~�8Q���ev�{6ӹ(��B�J�I�-7g����H���ui���ˬ����)��� ��M�� �@�3��!=ܤ��$�_�i�Ԗc��(���}��ь'��mk[���l� �����Ө�m���k����I��Hэ�~�,�t������ChF~$iڧ�vyM�m=��CK��I�3UԀT�{���#¡�:�������=��sy���ksoUoD������N�(�90p���/J�8d�e�&�%�Ta��^>0�W�Ɯ��%w̑��?�_$7Ӱ���l���he-_��j��d�P7�r�[xѷP;��u$(ED����V*r�(