��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�L��58b�Y��u�m����RVu���?��6X^@��&(N.t���G�]
&Δ+w�Q%H�]�j�7a  y�2���c	�a�}�"�^��k�YY�P��C�}��Rp�Í�Y(��DR�k�4�ן�ΰ�;�X=�-rj�<�.��ϱ�����P�-�9� B�0�"ۓ���H�&}���]vRT�o�"AJ��pD�?�z":X�9���(O���^Mh�o�ʢ��Dct���
K,Q뵠W6ʼ��_�w��a�ܭԃ��Ӽ��F��5B$�B�+F�W]Je|�I��`!�Mt��N�΃Ƨ^� Ќ�}���U�O�����
@��.�f��hW����q<��I2��P%��ɍP�6�ˆ�ԂU��:X��AR-�K8�u�ͧ�*�Mr�?�&B�� j���C�ģڌ�����d3�HP�`�Cq
�2��]���#��渨>�%�bQ�Ӽ�S���CSfN ����ȍ��3��z����\"�IE����J4��!��˥SC�xx�/.F�ǵ��$Y;�Q�8�$�we@;���4` �@���d��u+�/������J��~����
@>��A�-�u�ΝCpF=�[��� 7��8]�>/3�U�OA,-�j�U��֠!�/_Vn�Ս	$&���'-v��`k����B��D�&�7n��&�:�O�qJ;�£{�
 ���n3�W��Q��nI"��`KtgH̄���@�ա<$ɿ�Н��
p�C�p��K30�w�~F][uF�;,��PM���M@�@���Y��p���R��� Y�b:�/�cdA��q��΍�7رR�9&�::�u%��R#{�xЂ�6|�0�4p����	�g=��XR)��X�p�B��p���Co��3W��ܛ�oO�W��D�a�RC@{r�N�!h�%��GEcV�aT�Ŧ1''0���{�����WRT>Խ��Zx�ٜ�:��Mi�Cx\��m��}�˷�<$�qd�!9$�;Q�b͵bZǩ������UG��.)����N}����h����"�p��4�рd�<'��+L���L�
��l���� H��񨝧FOh{K�7cg_�F���C���t������X���m@�0�s�:�Ѱ���>�U��LpJ�v��[�%��+,f�e�:�ر�E;�	 em ? 	tVR����(�T��J��#�!��ڎ�����vQ�w1�����B�r���4�ڸ ����A�G�|H��;G���r^M��C?ϑ�"���"r��EѬ,2ZFaz�%��Vi.\�g�^KH
9R�?�������B.&I�T9�&�GX�D�rɱB$���	}8n2t-��E��v!պ䅼�~������a������m��D2v:�ܤ���^]>u>5��K�4��P J�=iB#��2I2�z	������t�zDϒA0�/�ϩt�A�I������n�%�0��#�P��dц��gm�mP����P���D��<,�{}|I'������ ��\�\�Jn��CV
���h���K���܇�;�	��>a�]��&5�$��e�b�8��`�]���Q�K:��!���m�s�����H9lt�3�#E*#ݶ�~�H�ʉ��JCmo�x�)353vw� ��^���5R���i[��ȪvVP	iz��QC�Hu�3ˤ�R��"��A�VVmH��L��	ϔJ'S����%�k�J׍j0�S�plm��~}�@��!>[FD_{��x�Ӷ��?�da�c�>����9H|[��##$�1E۔~樲��s�1Vo�> �S���#̯��.%�I�r���5�ĺ,���W��cɛ*d����獆$'����;��1H�x�D�!ܞ�{{��{���˹�Gk� 0��`���Z�_Z͐9p�䬍�
��c��{	���b���b�O^1���1u/�v�uHDږ^�i�Q��[3�c��r>Gh�4S�nd�Ǉ2���O�p۰�e���)��9�@C��vu<������=!狼�&�����%[eS��$�������𞺖a�V\w�1r8��Xh���b��M4͌����� `.h�(�<�~ƞXÅhs��[`�;=�H��p[�v2��D�[�]W����5�^ƈnG�"5/:4WL=�rI@����~	���E�3��r��si�*��gT�׵�W������.��mZ�W����F��(bs��ܪ~����ct���j��M��'6���������.8by��z�a���h8�d������������Q}�r���j��|�p/�CQ��hn�z�}1ݭ��JS��6v@
�Z��*r �8��5g-�%�:fI��5������m�D��z��� hJ�������>7
��1�B�F_�e��c�|��}�Ԟ�w�6��a�%�/<�0������,8	l�s�YSr�JY��b���5��^7�nɾ��5��=�o)M#�?^k�����%D���Ϻ�0�gGM�H�Ƨ�����o���v����	�i�#R(?�?V�-1��oW�Q.G�~Y��q��;򾆁�N3��yMĀ�x�EN���Ƙ��(w,�����f3Ќ}4���}��?v6$Lgӭ��f��f2����i��GzlZ����70���]�2���;7=����2�������h�\ c�i�����ΈBu�U��e�"z#��� �U�f�3]���_����DX�Ê̓W�)�|��_x�˱���b�l:#�Ee�6�߃y,B��	5���M�A�P]�e�(v��������2�C͛V�?�Ug�Q7�l`�l�(�k�g��N�
�,a�B=u[���h|�|r��U�ܠ��SO��O5U���N�J�̈����3���.��1�!��N$�t�(
��t�h j�m�Sl� ��Y[���7�@{=���V
������E��{Ûx��ޒ�m/�Z���D�?46�.'��p�J�1���W�ae�
�/��Mw_�� ����w3�R�D�,*�*?�����E�	v�������D��JA=�9����ŇڣF,�z���	}��m�h@���[��^��>�9�M��0g4�	��G���+�m�lRZ��Kpbi��w��[�nd��D�N;l]����"�vxG}�����-Pۻ�8��	�8������m'hm�?��&:vU�hr�H�s�/}ޕ}"ri�qΟ��'�1K���������.)��{O@�:9A_�q˥����P�ш�l��_?�!��G���~frr���zyx�@��R3y��*�]����C �:��XU��¢��ć�4���(�`ۊ�:�R�G#�)ݩK�� K�˱f������y%���*� ��