��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�tڐ�!��Q�����xZ�H��V�� �]d��� ��h�hQ�/���o�~�կ>?�5�z�+|��"D�[�!#��.J �SJ�Ҕ�5�Y7�0�f[秡3ڕ4�O�~�	����u�Q�Q�H��)*��V�o���}m�'_z�8�y�@� K$E�R�5^R�Ԇk2�vv�#�80����I��JI,3)e�nU���i
�R?�T�ƴBǡu�1�\����+i���j�;�*�z���o�ć�I�-|R�JZ���ڸ�$@��p��,�	tB�=�`ZY�����%���H8?�����0<���dYA�b3�
��F�i�཰�ܞ��=��X�W�K��{��eq&S�-���>�n�4�%�0�#��q�[O�'���ɲ�E?t"D>�B��T�"�;�|���q�����82!��.��@3z�ȸNb0�p_��љ��9��Z4�����3��Y&ݻ�*�O��j��b�$��ގk���>�d�K�*E�@���$qT�Ѥ$��n���t��m�Q��St����+ ?��=�W�
�;��/I�w@Qp��h��c���@���^4aٝؠ�Ғd�F�	R=�!�$�a�B��y�9t+'�`!��f=��B��o�D���B	p_?�����jmo��+����-#�i{�w֔�J:�!!"��� ,����z����ҝ�Rc;^�d�C�/O��(<C��E��D���
nc�����XJ�䪫dR�i��A�?Y�����.\k�S���"�����-
���*"��s���2K���?b�.{�>��6�_��:����s��bϫ�ʎ��1ݘ������?��P�h������_h�,�|�c�g}�C�����k���ćzG)�犵5g&E�p���A��3Y7g'��{�9��"���!=2]0�xr�$9W�[U
�Ǒ���D?{|y㕤+|y7|�t�+�ԅ\�2�f��rl!\��ՉP�9*�5ޗcL���do,�:�QZ`������wj��k���0|%c�d�h�@��)���9�W�C��k�'��-�uYe�Or��᧮���<��Z�Z�YD;��;�-@��<k��o'��Бe��y����^ֹ�.���3b�~'i�T�k�K�_H.WXt��@�>��3G2f�ȰG�wP�,���g�Kă�F�z_�Z���<�O|�z1�_�������×.��A2*g�2g��C���V� J1�YͶ��^rt�X���;agT�Wt���
�zl5�W��@�7�71���63i�\s.���
~6��OV�ex���~�i׮dAts:�lW�*9�=|rcIP{3c�2����z�E8;����H�y����1�R���e��d��M��N�rZ����0=��]���]�I��� ���������`מzuȲ���{9<�;=nGQ���ep�7�r���Τ� ��gj}������	��O�FM�
� �(�����؉�TlS�x�So����(�6�J��YXĵ��1���ZZL��T3�L�1�r����e\A����X�H(~����{�0��֤��ޜf��b��@9,o�Q�s���K8�Q�e~'t�`]�5TVodCv��K�*Zl�[ծ��N�.�$���5�)��Fz&+n�;Z����*�0 /��Չbr�+UJ��� �����%uq�GO�٫��}��;p��҄�'1Hڸb�"���l�N,�8�Ͻ`7P�G��N�|W>�O��_��)-�ʙo��j�� �ʗ��[x0R��
cq����L���p>N�O�Q�"�4j����{F�5Q�s��_dc�ΘO#EKbpz�<���jc�A,eD�Ty�L��/�s����!3�3u�fg1����E)��#���zIp�y9U d���� *��Ե��x4���k]���?L���ZD�ɕ�,��N�,2��������h��MD����J`��S�6��E8����|��knةW^v�"�D��2Ј�+m
*�Q�j�S��ܙ��g^�;nJi~��WR�*tƚ�r�����{|2M��ze)m��8��;��_�7��坳E�ߛ9�_V����i�K�:������4w�_�o?��@�_��N��@?��t^R�_�G�b�X��˚�'�_���i	d�=�4�>�n�eX'�1}�Bm}��y�Cl�E�H=�3{уx�ΐ�W)����/��N�[�s��v�V����\�66��2��w(�^����"b��MV�p��Eq��'�����GG��6)�޹6<4�p��Yݣ����p����3��q�t�3���ڻ�ݜ�=[p`�O`�ܥq��u)�o�߬>�{#�5�V/tf���px�2���%�9��\JЎ�"O4{V�Ǘr<Ѷ�!��T�R�
~���OxIb�DʬaĮ��Qo93�����a>=u�������	�8�X�U,1�rP����=i �ٜBb�@���0��L�.׈v �BZ�PɆ�&B ��E Um�T��H
�4��!��tr|"�v;Jq�x�������i� .����L ,��=����m�¾R�88>*�E�� ��\!:�8AWc����N��t�>��i���@�-`iY�@I�	��بx�_��J2��A�/��TUi�1p��
��nG���k�dM���gc*�q�8=��dhgɀ�5�����M��J�1?J