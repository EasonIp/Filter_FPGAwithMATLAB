��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$��c�\x.-�M��h�T��Ȋҵ����[�Z3gAd��d�(D�SO{�Ȍe���mKns,l�R�Myƥx0h-��6kWǔ��Fi�1���w)mUu^���9.�k�ecܷ��*����ךw����.,R+��7��fLf��IԺ�7%�0����������� t�M.�h����jɠ����&�l2���v�FZN7�N�?Uz�Y��@߃s�a����o(��� �I=)ƭ�K����)T��2I^!��M������bj+���3��qnl[�aOu*�睕)��� �Z���I�_0a�-vM�\����;��Vj��7�I�}C 4|Jv~I���r���"��%cn��H�j�5�/:��!m�u��dk=�l�e)���Ã�Ȱm]��p��U�K8d���~&-�`�݄ݣ|�a){bl����Z�~��=苀�Ӡ���;~.q�hH�?'W�ɢ�J����_[����|�TJ[s�qu\eR�˂2 k�iu��et˵vӆo���2jÑ�N�6}Aa�Zj��7*ͪ}����q~y�I�������$$���t�k������ڈ�7�$38�O��mp���5*�&xavB���Oh�iW� �Z�F�m�� ?i��L8�H(����΁M����᝷�i�#�w߱z���̳�4�Sd��8��f_�5��J½L�ћ ��43�uEs�}2􄱕�y#��i/��[-��qH�f+��>�ߏ�8/DdY�B]�zN1
��_�o�>�yVD��Z�$����:@����d�i%2���Aȣ�?P��@wU�I!�Q��Zu@�P��h��1q��ߙY�p�M��H��QJ��ggJ��>�	��� �L?��gLv���  �DU@�_��+������CO�}E3֗5��ō��Xv�p]���>�q��+^�գ�q�Tb�u�E�&��6M��f0�&��c�<W�h��t9��Jߩ�/2ѱ�� ��{v����������=эM���ύ�*{��hf��l����$⊊-{���X�D��F��$�'K�=i�&�ҏ����v��ViN� �2E7��X]�\�yį�1�����yK�"�`ُI@����^ז͎�&����Kl��fV�V�7��5�)t���~�����a�����il��G��[���b���wFJ�����������8�Bks0{����^��c��!f���W��}���B5q�>�2����j�����GX��~�=��f�O)��Q�![���6�D+�1H&�<��`B��my��B�x��v��-F�K�(��S���Uv<pR���."�h3Y��Bm�rZ�P�+�n�|?�{�Pb|�|��3�F���~jcn�dt��:�+A��qL��L�fͫ�H���-����;�����w���� �؁zNSzU�ߺ�N3@B�SE���dl{u?���Z秔������D(Qi?F�;'����Wp��w`�K��t.�� �Ө.���ƜW�Y1`��6|���n�Yy,����;O.�XK?K��|�ɠPg�ܛA �j��=qѨsI�[~�TL�5��h��EH4�C�ʼ$��)�[�2!cW�ҩ�m�9PPQ�vKR�rs��lm�/�	LYOw5d�uM�z;QH�]�zT$��.2����{�ɒ�z�Ă����C�G�ބ2�{9V�ԉ����K�����ǟҩp*v��/�xq��7��p�S+8���bN��7ݹ�I�4�y�'�bef��;�9�O)]0C�����V>�}Ťv"Gฝ�YW?w �ʽ���s{��I�������X*R�ɸ���Ȭ�ԥ`U+�~�d[/9��A�z�+��Gs{ۍ�k�w�K"����̢Y�`�w�ͭ�i=R�V���=Rv# �� ^<��c/��p^��A���~�i�����CzD�֮����PN�����D�֜�B�G�)����sOPl��i!�̦�dנX��X�L��_j�"b+S#Z'5�r�R�9���o��C0��U�'r�޳n1O�m�4Q��j$�b*'�=t>�V�?Ez��%��<'{�oq��{���j �8�n1'qFۖ<։��֣_d�UAS8�Ȳ/8��,�/6NDoz���ᇮ]	Ž�T�X)FH��3=���95q�������#fF7�A�}�R�R8~��� ;�Fs{��:AK	�M!.�5e��>��)a�uPx��U'��|� n�a���7[�HzZ3�I��أ�W���ol�\�f�k�M�K1+�:�9R�ǵ��`�I���UPQH�suD�F>�ğ�,�UnUv�B������x,��_m��f�9i�ә�J���Y���/d�Z�{��ƣ�b|���O���yɏ�v�]1���.Ɋ�D}�C|h�YY�y��{Db<L#�д�mH����Ll���j�k�=�s�i�`���y�6�%�{x���Lt��f3"�x\x-	n��o�?��![(A�M�^��ub��=�t��9��M��5%����*>�xi��p�k��xhK�a�c7u%â��A�!�?3����������_�V��z�3'���}L7�kf� z�����T
�l�[��\��6�8ޝ���=К�_�9�U4�:�r����zɘC��&�#�#�H�����\� ���#�N��kH���59n����:J'V��FL�E�m������.�Dd���+Q���F�Sk"+O-���7>���0	�؁mb�~�Ϣt�I�	�:��J�ȍ��h���HAZ�AM��XRAoِ�7K{���:�څ4���3�;.�b���]0�~m���EfS�_�g�?���R�{K�����-�_ 0��,�i��OB�б�b�ƛؕ�_��p��k�p'I"�����?��S!lǦ`]���n_(g��/�{�R�R8�+�=E��(+U�g�0�k��18k4����\���cЎM��2<2*2#��8���a�$̽��&��
SU�[e����"�^w-�jvKq���%faÉ+0Y
J��4ѱzR<"$i�d|��V�`@���<��'�d��4:�?���<D�i�s���|g0�r�F��%�a��1�"��)���{������ �j��G�L�}�{���5���m���kfk��x�z�`�C�)v�b�r���Ab�ػ.f���vH��8٩��h��`��qz��wπE\g���|��:�-�V ��r��mm����[�����@<4�#�˹��^CIЧo�V�������5�ӫhԥʎ2��iQ�� ʺf�\a��o����8���L���[*~*��q_0�Wt���[Pj��'��5��7q���i��:�\m��e�a�l&+K�л���H��qW!�k�.��Ovb`�L!#?�)a��<f���+Hx��Ҩ���!����(��e#�p�fO��	�y�w2M0Kd���%9�ѧ��^4�J�E���b9���,f��y�a��O
��B/t��F�5�jځ��>��2��r�9L�3��q�����.B��s״�W&9����`͵��؂
|��峌t Y����M� ��y���'��	�d�Qb��iH��*���%��v�1�0օ��37v����-da�;�T-�6 p��
|�P�F�n��m����v�0ũ�rn���vb/uː��<F\��lKΩD�H���Y!��/ʗ=8u��� ��$�;�'��#�l���]~A��-���6{5E��#(T�}3u��⥢���l�[��<�|�Q��Ӝ�*�*Kx=�~rh��D�f��|���@]u�����@d��������7�����8���q���'x�r��˗Jz�`r!y\�)0/J��Ӂ����*j(]>nK=T-0	�o`n�<Ke"�D�K����C`ZGb��]�F0 ��H���4C��{��=�?_������:iS�q�}\;�OJ��ch�� �-Y��U���7��/qW���.����'�+2�K`p�%ˮ��X/+-�_V��\F0��eQ�Y������p��l7����P�s��Z���ꀂ�qBsa>�v��^�{��p��RY��R0O��?6�+����c3N��c�%������2��-����Mr-���XQ���W
�3��G�A�@�j�����H:���8�e���SJ���2�\Z_ѓ��h��ڨ0�Υ�f�;�H���>Rp#B����`�6���sn�d�I�P�nvC��}-y��0=�c'��4��HU͍l��>;�"��̴�O��NO9S!-^�v^
�]Ϭ�z{��u���|��������N=�}>""�v�Z�O���.�g�x8p�&hX��h	蔪� ���4yM��mq���ޱ���[{I����9Ha]����F����ZC��vm�]֔��4��E,�Ѧ/ �~�^�U���x+D=���8��L�PQ��`2���Y�e���FmsЖ���V��l|���*e�V����.��ï�*�lRsC��a�=j�q9���#$�{�T��;mFQ)/q�HbQ`K���D�hܼ	w	��6F5� ��c/.�b�B��tRB(����`oޒ���q]��s4W�-�?U�F!7�#a���{{@�-��7�tuCVAR�i�� ��"ʼ��O�F�F��U��y�����b��+ZKHC��lT38��(�U d�>x��Lc��@᪙.|��o�Ѯ�L�����)N� pS�����)[ ��}
~�Qt��be�)������H�<���o$)]7|��a�w�KM���Z���S��ʫ��sAQ;ѳw��H�j�_�=w,�A�]]-�%	N�O ��=
Q�~<�9"�C^�:mh������M 朗�o�}.�nd�W7�h�?�/^W�ҽ��8>�-me���[)��������&�lmvAHN`�1ݜ��Li�p����ٰ�YTJ��"�m
�@���q�� C�_����4�+2a�w����ă"���F�M2�hE�`�`-��!�1��v�XUBw���#���� S@�s$���D��T0�R���Ib-�q����3��w���(���Cc&��R~H�'���i�.]��[�s�ChT�M֝�ԄC5����J������.z�j\�s�R�������]�� �)���<���>��ɣhMr��U&B�!��y�o?�fh�#����D>�����[���#��]G�+E�w���[N�~�iaPwū�_D|+6	��oc�{����Cg\ƾ�*j�� ���j�p��0]��
���3,Q�rn�p;�-@�Gb��D�2��v��n���������q�C�.��'yHgّ�4�bk'T�ZK��*^;��8��J�22[���ٳ����@�k�dC�R6~���&���Zp0)|v��՟���w����m��6NϪ)uL�&��h�T6�j���UK3�cЬ3������	gw���_ƪ
�Rr��ڇ�yx�򼎜�6vomLj��NWȠ#�S^�Nc;���ھ
�Ti]�+�&=ܹp�}(7snO�6ǖ�Y��>�ɨ�6A�ǀ���	�E��pR���{��q-ø���$��YA�Bo���Y-DSl�$�P;��7`�N�M*�~��ٕ�f����S�}+$.�H�ϑF�W={�p4:�|0wk?%�$��z8�:���}gw�a��	UR ����M���%#�=��j��%F�*r�=�F�v�)VQi���e�,�{+�<Oq��
p�ij)|�m�܄��S%cM�P������PK5Gf A�<�6�f���XUG�
��%�nI��ܴ<p��8#+GSـ��l�,�U��\���C�gy��5V�3�"�҂�~�}K��
5�뤻�ӓ�R%�p��(��H�x�`#F���cG��k���c�rzx���#P��_8���h�f�3�Тhڴ�$���9��D�+v�P�3��q9յ;Ku'x��
 �X2�'�u
�iٿ��Ւ/��3XZ�oo"�f?d��8�(�@��<i����~_��+F�x[I=��1�J�U��1����vgN~�A#��S�iՂ#��[�^���X��x��U������Y�"'�r���rb�.��ڦ����OP�a	e��he��F0'�B��u9:R�k�d��B.)"e�~��p5�8
�٨X�D�5�ыf��h�v�f-��
��W(��L��xy���ȳ��Jl�ǎ���Ғ4)���mi=,��|�an_�-�
&�F"a�dR��,��v������ϣYA���w�%�X�������z�Y�g�x�:��3�u����N�8Ie<\,�'o�V���fRnrp�̥H'<�d��P� |Fjf�>;H���7Ʃ�8�r(<�PT�F�zM�Yή�4
.�!��m4>�?B��P;�U�����dͩTt�Ƶ���\`�A%��ہqC�v:�N�6Ld^?d��zRIs�D1,~l*Wg<��j�M�F�!3l�)����(����;���,��b^Q��f��V"�3xn:0�T��p�O}�,-�w���^���\|z�� �;Z�k����q'��0���eX�JǎZ�����K�nW^g�=z$�H����'�]:k��xh
_�FxZ�)�B��U�p�~!�},�$�×�ݚ�Ɵ,)d���h���-�����\�e
A*���j���)}��¨��vu)}��������B�3Ϡg�k��:���p��k=�:��ï�P���yAV��54(��)U��Q���"�5