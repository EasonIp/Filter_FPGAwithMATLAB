��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$���B��:���_h[�y�h@��d���]0W��"��i}T=��7����Ŗ�����b�m���y��eض�d|8)O����w �����B,�������f(q�fY"p��X��V��zc�����`�=B�$�v2�A����/�}R-�%�%�|�ڝ팙���&��A�H3s�u����f�ZM=H���{��RL�C�x09�T'�ce��p�"^2���D��@�"�N�"�]dy��?�E�x�9�	�{ٲ�5Q�5>�m��?��y�&�?�2��)Ya�<�
���U!�O�.�^%?�b���NčG���<���o]I�z k\q�I�&���yF\y4�L�����$l.���s"}*Ru�k6�WO��A��՘�s"V����3xh��nvc�{�E�N�D3K.�ɤ)^z7�DZC3<�2*J9��5�Τ�74������vUnxұ��B�џ� .�	ԃd8�P�v�(���,z����,�42�1�79�c��a�e�����39�*��݈?bƈ0�����Rw�;-`��}��=z�����y(����]p����~�?Ԡ��h�2�$*H�V������H����kP���_��=�ZܵD�b�,�[ ꧰~MT���"������$a�e��:��(��?�P�"��u|��\�
�ڑ'��c��	%[�Zy7��l��T֔Gt�h�Z�#70����d�~�:Һ�N�:�U�v�*�"7�U��ئ���� �>W���d��B��D���l�{�M,�u<]����1g�;�<] �����׹օ� �hW�y{XbX!#�&�&�f�	5�pfw|o��»�8��n^k��Z`��r?T)N�b��22�_Ę�p�B+0���Zic�����G�Z��E�&��	֜j�B�"��y�}ɱ�Sy����Ԇ�m�R��/ ��*��U�;��~�������R$$�N5P[.��Їg_�g)Y�C���E���¶�=h�h���3ӿߐQJZN#ce{⠠�ʐ<� !����/�u:�(4\�}�^����
�6Ƨ�zj��M��s��+��� ��ٳ�{[N�C���9��9:6׏���4$I�I�!X��E]�]CP���-���ѯ�5i?�p�pP�|��q�R|#=�L\��1R����?k��(Bmfڬ��.K�q)Ă�]s���'�P�{��0UM5��K���hW�4���Ν2:�#8�;��̴>]����S���<�$���K� .g=Dk9���"%Udu����#�4Flq��yu�Ŕ�*P6�ǲ1u����R�`�� �14/���mw�0�AŎ�dg��癝��T��ڱ�8�x`������v,aj`m��hv�B�@�F���
b�;:�r����9:��w �>���셀)Z�����|�fdk��-d�PғvC�~������}Z��ߗ�c�*�۴�+72�����@�a2?� 1�[2�I�֏� ���}�^51���
L�p�5���򭠢ni�����o���0^s'�Ͱ|VM�Դ-Y_�01�(8�$d~�T>�ץ@�T�됅��l��yZ��^�?��u�|.b�O��V꡹������?2�ٖ�o�h��f��j.�����OģFt�"6=��-�Y�l>��w���u�%�<�L���sm�n��U �Y�R�Ӭ�A�k��n�K�Y�n��!(�������>H��rռ�����5�Ǉ���?BB4{bT��
�WJ�����2	�=.)��R<������'��;���^h��9��pT���G�F{�����Ɔ��C�2�D�D�(%ln�pZڿ��Ŭ�/!��VFӤ��{���O��ر��A�&J�{��U#���b�C�\�᡹�q��E͌��(�s�X�}�`�_��y���Ϲ�R@B"J�/2婚rr�j��*d�g�a��>�ό�(��m��ܑǰ-ϟ�!��v�����p~(NO�F��RBN&��U�m8��J~\��dC�>0�������i)��L�X�����,HH�܎�S8�R� ����K��6�Ω��"�o���х�-gY�۞Y�-�0��ݜu��Q&��e��Wݶæ,���DX�W�F�&���3ϤQFv�3���m�MI,S'4X�ǀ�q,'�$G��~}�އ��dji¬�և&��0��JN/�0	�J8���}����?�!���,�M]�!1�/�9�/~aZ����]�t.Z���^:_pٱ�x6q�J��#B�%	�|Zv�b>}��!xxn�.��ԅ�|_jdQ��G��P�߂㯱@8\���7m2^;F��ԅ��X��_�w\t`5��ez��/G�����و#��,x�C�֣^NA�a�I ���	R%H>Z�h�V��KE"�5ˇX���?:��z��g��d��p��Fs����[���MV���OB��V;Yf��Nn�c�H��;6��.�����5�[m4�4
���B�Z_�� `�;�ǣI�u��&`-���a]\�=!�
͑��:*6�*nk?�>��|!�y�#]��Z���w�����އ@W��j�/;iN�����-��&�a���?�0�	���q�<r����w��L��9���v,U�͜'i}Mb��K2\�ڒbȣjQ�����Qh!*��7u���"�H�����v:�e�o@U_I�Yk��m/X��h�6"Yǅ�h.�?_���c�/�`�
%\'�5���a��{�Eo�sp3�1|��������@�=3oX�'��턷%����dl���}��i�s��%k����v��:���J��A֥T�2q�	ȇ'W_�/�9�X4��([R4�b��2�H0 в�3��z%���:�I�ߟKEIDH�����Y���+�렞�Hbg�^��AI���Wa��epa��K2�=$9O����[$��u�ǡ��aJ��_N�"'���X��& �ْ.H�<��Cs�]C��?y�G�+������A��/03�+Hs�c巴����1RM$kk�.�H�ݥf��xތ�	��\�4�/}3bSB�K��v��v�����+��B<J��"�g7��p��G���W�;�!u4�O����vL ��
�`F��SL ����}��ѳ_��h�.�'mw���Ĵ"$��'�X�M�o����f�
]E�8��Ï��@|��R~�n@��"So��X*)�g�f���%�������L鹖J����n%�#�G�`?#S�����4�e����"�����P�˲JQ�$E���%��
�w�$V�_��^��]�a�&�]���uc��ơ���Qqh]���c��c �&��]Ku�ba����un��~�ɋK�j�&P���bj�ng�ܶ�G���S��eqn;��:0�s.��]��<�L���J5\�SmA�C��R��'���`#?���{���˃6�@���II��Px��ƪ!A�{�$#�h̦�	�����8kMe���O�������4駹���y�R�\�s��Ab	0'�G��V���$�����	��؂�5���w�C�ns�^`�(@W]9%C��}$� ʍ�,�a�Y��߰��p�����q:�g�{��87�Y�<���])f��oH�#_�fpp��'^�������9��3�b �j��J/�>F�T��X�����"�����c �\*y�^�~�H�mu�F���ʭC�,��Ǘ�v����>��Ég�[��vDp+'�����Xɯ#� ^i�H�	���m�g�9�|(!�9w�+����;3�,�=O^V�SԲ�~�� �or�����MW���qW�l���	��G��e�ʽ���T1�N'�<M(�������-q<��vmX��H�yv�x�dZ|#��*��gM��ßXj�"��7k8r
�N�C�V�2�)	�����$�M�ab�(Ɍ6a��(f@7T31D�C@�
�R�Y`����s��oKv5֣���
��ڻ\���u*C�qlmH�����I)?g����L�g���5��*�V��J�k����<�-�	��1�!�y��(;D9��b�'n�o�YR�KH��5F`K�D~I8<G?45%%��&���ޛ�i�J���3�L���ăhP�!�oگ)�y$
^?�H�U)��p��Ԫ�{χ9c�N�gS#|,�r�<Y�n���O�	��kڑ!�Wi�~P�.@��]�l;|	~����l<O|~;���Ii�k!׍4�����x�[G���l�d<@U�f,��nsQ��7�?���C�%����A�>b-f�b�DbSH�@K- _R���p��(�g���J�L�?���C�[�DH��P�����D����1������{ni���o^9`� ��i����.��F���ur`&�EyD1��<&�^������Q"�}��֞�R
6�U�֢�bg@d�����$��ʥ��,�`����n��0����'gow0ݯ���u���>:���@_�ͼ����l��_x�X��
�5�8��"�AX�1ƂV�}c�i���Cɱ��X��w�����b��q ~�Ո=6�8���:��&u�(��� h��1ah�]/+����n�����ؓ���9���e�ZSf��ҍ�w⪛ ��]�B%	#3 �e����[N-+#���{��+wM�#X���|(Ї�V�<��j�L������Wg�^,�[}��v��}�:t����.D�,�P6Z�j|%��54e[�v�����>F��� c��"t�OF?���܄�h�3�-s2�l�l0U0*}�N����X%�u|D���f����[O�1o��J˱'m��J� ����i��:�k}V����q���������`.� �v�.�:	o~�
(|̀slS�T�I�m�0ߥ����iˢP<� �L1l"����.���hK'�aK�Z-�p��s�BYX��5�㦆aߠX>����ֱ���&��̂��[M��+���m���q�H��.�WwG�L\��4*�+��s�,�J�j�8bNm�7�7mg'�ɗ����#��S��\�R�LP�;t�s�(�@QZV����� �F"ŐUF��� f�h$��4��Cu�z_O�yU!�]��d������-b���!��>���(e]N(?�˔�(IōV�r���U�	XBύw���[��Ͻki�[�~):�zp�}E8<Wyk^$����ܤ��O�Q�ޣQ�(~d2X4B��	[w23���`f��Nio{&$�>S��Қ�2�=B�c�u�Bb�� ���{#�Ge�܅�fX��n�B�%+�������'%�<�� ��R�unt�G��IJp�\����h%m2F�s�i@�k��}�Ƃ���a����?Hl&�I]Y��N]�����l��Y�8���ޑS�.<n�����;��9�"�����~(�P�0��L�ϻ:7[?u��r�U� _�!9�m�k�yqGs�ٱV�|��з�ʉ��5�^$���<1����%�l=��/������ρč�L�r�L��R��e-�,ja��G_�?I��dY$smJ� �EH1 �s�0��_��)��e�4����wy���`��\��ɣ�����\VC[o�vM�:N�^�y�$�lK���fN-�ɱt�_[��ĸ���(}�����f��u������҈,��?��F��q�o�?zҰ�*�W��$��4i�/�Z��ϫA�U�ݒ�'LD�ͻ̹Ց�0��˱�sѰ���	�I���9�N��,Hx�?����ۦP*�n!��M� ���<T�E�	)�W�2��Ha�~�k�u�2Z1	��:�5����w�qI�l����2	�h�jo�����!Q
0-�>Ti�t������%��z�fʄ�l Cm�0]�8Ʊ���C���=�o�'Pc��:أ��+uV[V�UGt��`[_�Fq�#|U� ǻ���J����4p���6Ez��s���`s*"D�ی�gޫ��TJ$I��#���~�R���"h�a<���-���=�i��6AB����j/��*��B��B���um����0:���7�3U^��~Ų�KÞn��A����1 ����WON��8#���ie�ϋC�i�ӝ�uJnaw�������ܖ���Aj&[�G�<+���,ܾ'#o!�%�ư�d��	����β徬0J��GQ�E�e�o ]���D��T a����N�bݦ�rE�,o�G���&,��Q8t�|k����]m�-��N������8�d�u\px�D�p:&9�-k8h���_e����#�qv��xZ��Š��ۖ�����7��٧)y_�ۍ}����_d���0+�vś�ޒ�g�XFo(&�
�
j� ���@K�Sbo.]#�h�����Q�B(VC��i=��g�V���Q�f�j���	�>��;h�C�pW����<D-��5Fq���u����MV�����w�#3����
ϧ��~͙b='�_;��x��&=`�"�����4�&88�n������=�7&�������4���\w}�pg�a�n�
��B��&��e%�W�l�*S�"3��vp�O@�ʟ��8�Ft;Ih��3�ȋ҇Ici*$`X��5W۬���\v�F�|A#o!��wBd��J2��*1�W*����������;Z�*|���}�d�����M��Y�~��#Y�L��M7)�y��݋E�VԷxEѡ)�~���ch����ŐYt�����A�53�*p���2������p�A�����q�NR�3���*��%5Q��qN$�e`��g���fxa�R�z�dyӮ�m�K���r�<,��S�>�^���'Hޱ��>�}�?^���5�"q�>��@�Y$�ԉk"u;x�ͣ�I��Ge�D��I@���+�M\+T���^D�T7f�z�Q�o��ܭ��˔^�>��EcS��`rG}����FX��@��VP�w����g^`e��[U���*:z�؈�LZrI(�o�U�����4;亷O$T~��|�I�v/��x�^{�AE�m�l��<���-W�Y������ó�
��<O���'�G�On���kp��5���������	+�8@^��Ұ���63�&�RpQ���U5�<Cq��=%ÿA�_8_�����_���U��<`�2�X	�,t�%�O9Z[`޿�G*�=%�,D�����!}���(F�~��EҨ�F0s�6!���O��g��J ��p�\��a��;�0�uB�T�+x;�$/����/fK�uX�e���7ї��?~�<���o�^K8��p�
��5���X�z۟��Y-35bM���e�eSm�*�F�s��_�c� J���Џiv"���W�FA��V���u{uⰐH�R���>�C������o6�ߓ���_K�2I�}��m`0�a��pN'�d
'��v�f[����I�
���ǉ�9�IA�߁�������Nl�����4{W˩Gnq	TAc���b��˃�5����]$�9�f�
�.iy����2=k8"&�[��9�D�M%������V�k��;;-ӏz�^�m�B-�����C��^yp6tC�aiCDrP�j��u"*�'��q�� p'�\�w��8wg����+4b�S��|X-�vnyyz%���l��R�ݫ�F��^�YC���b7��?/v�9j��S����++�ѷ�¯��[map%�����/߼
N�\w�b|	��G,������ pV�yjn
�z}!����0�	��y<��\�s��x�杶��w٥:g��]M7��tix��\�~n	~$Y��S��<�Jr޻�[�x%!'H��G0^�=-�����|�z�;É$���~R8�sq9 �DW����-���H���h�hՒ���4�~Dsalw)����iA-x��\���#�Xq��͡�/b�5É��C������x�OA<��w�l�T��^�)�P�.��}P�!q4�x:���7#�� �z�W�U�I˺�n�(��n�a5vI�D�@��U����wͭs~gX��tv\j,b#�n$9c���9�c�p�st�r�
��VI�}��B���]N��?�4��kZ~�K-�?0+M�o�2 ��]�Ɵ�Ku��F��hXcO��01- ֬�e�+��SSZ��n�HN��0�l<(�(�N���R�6��Տ�М1�i��P@��#Zv˻���-�d������Pv�b|��ç�'�
R���l�T��*�r��+��<9U�}
�@�U�hcH�F�&<�C};��0�+=�7�5߷�s�cͽ��n8������i>�0�+���<���Cbʮ��k�t�L��l��Z1�ҒS:_�%i��mA�*�?F�4b�+����0�[y[�� U�P�p/�,��w��g� ��e�OT#L�V�'�����z�t|�eΔ�X��W�ޫ����v`��][�ד���ǒ�G��R���R�q���H��@�/LZ��:E �x�*��u�U�Y���H�:���E��I�'��j���Oq��W��e�e7�\���	hA1)x.w위h�#��!#��'���0(���M����|T\�� ��J=���+	2�@�P�q#�7"$A'�O��6�e�N@��0�zs���� �j]$K�P����^�+j�+:J�4 ��J� h�&v���A�ݪ6|�r�X.D��1ȳ��Q4�n3q��T_��=���qH�9A��"�������<"���4��vvI#5�;~�6���s��H���](s�5�J?'E�a�Z9�PZE�h�D�`t��qH�L(]pI'=�g �d_�� ԃ����ۆ��(H�~�[��������y>�����$c|��4߬BIA����������[a���G��AdYe�7���_vUm��C6a��B`���A��?�V����gډ�,�����{�`�"ɏk��p=��4/����B�dD�U�^v �b�Ia�(�܆��$Cw�N`� ����.��5������z�����blE�O�;���A*R���h3�@����o��
�S@c��[u�c��T�A�{��AO(4�"1���`�o��zζ.7�����q9Ű�!Fw�%yE�U��x�f��;_�ڨUQ�R� ��YM��r_u�?��k!Z9K�U�z�#q�r}0������2��H4�j������资�R�(��mq���8����i��Nc���\o��ƫ�}]p��u��A�"Hb(��[��
q,0˚�f�������[���0C�m[�֏²�_:ЭI���h���Zyc�����WW�0D8;�s�/���PE�k�ӏ�*��$yWK���'��'�ȺɷA��yO�y����X�x5,]�M�n=��>�9���ų�s��_���,-�Ը&�O�s�j�-�O�t�m���Ă��B�����OW�X������bʪ�y�	Z��<]!fۂ������-��q��=x�sf{�U��W��	L�ܺD�N�]}�_D�"
�;�H:��op������3�[�.L�+��L���q�C��dwp���5����!�w���:�˻��g'��X�|��ˏW�e��,�0AL�<D?/����Up.|k`�^:.�LH��y�')�`��>�v���D��6K�E]4X���(N~�>@n�Xd��\׽$�rE�Ө�Ey �x�'��y���![vYϫ�i+����5���	FYs�Z�0Ë�l�&�+�E�5r�%���^����S�j�r8�l�Ȧ���^��$����>��t��3���p��/j]/����2r���q���!�R�z	y���#-�����0Z0�䓵�:sz��[�wm" ɥ5��%�{�0�����aP������Jˎ
Օ���{�Tx�+íOw�$�W��d�q�h�ޅ
�%�(��QxȢ��(g��ݑ{;Q�p�!Vs�*s �!����榱M%�	�G	����qԷn;5S�3�"k�x����9d�''�ܮx��:~f�:�1��5
fm�o�����	�U�,���y���I��k�x��*��yo	�43����.�cho�>�%��93�rm�G�b�~	�z�o�b���Z��<zO�-')� 	Hc����u��� �&Cة��|
�g���?;��N�W]c�
D��e��]ҕ�7��af}$C��`��OO�!�<mRF�{�jH�#�������.,�!<��*��Z��a 2��Z�L�� �T�q0q&	orx�R^��!�bb��5\��3w����)��(Dq{��[.[|�ʜ��~���� m���-��<��e��"c ���FZ�d���^.�K����/��,�&-Q��Zx���
>�����p�&.
@E�u�6�K5K?Ӣw�:`k���@��TV�|��Q��?5G�����|���&$ ��J9�S���]������ߤ�vmoF�?�֫���d�#��s&"ا�%V����������cf�$#K��P�����k`�_Flhz���Sd���W��?�.n�,+��Vh.r3����f�83�p����v��#S���S����?�K󔁔�G3���x�����K�����&�өH��s��������y$�W��̨���x�4���ųN��uߴ�b�B��:a�9�u�Yh�	I���y�du��ah2g�C�����)J%@Ы$�����+4�M�LZg]J��X$T���i@��"ʋ�?*����hrN����L��
��vF4� �����b����yҌ@�=&T AH�M�gӹ��t�i<��������=YB�ӣ
E?�������/�t��I���Si�Oқ�&���-Uu�ι(��$�#��d���D{h�f��ݍocwޭ��]A+e�V����\�[&>+/��!���z�S��լ	������@k�?���B\!5�0*�ol�A�Ng�nit
Q#��c���t K��'��(J5���D���r`����T�qrk����w��aTU�=t=8��OD������ U&������{C�Rr������\�ţ�*s�26��o�͉J�pmQ�'ޅ�4ۛ��Kn���m������3���`s��Z3<��&��N�|,��� ��ݣ؃E34�k��y�@���S�,��QfA�ʬ�&�\ywԊ�l�-��,��~X�� p*�5 <{<S8_4�^�5Uh���������i��t���C䴍��_����Y�g�Z+g�^ä�yza��b%��x�}u�Cq��c~�l
�g�����f����B�nߒ�z0'���3ז��`YLd��삜'�Ҏ���Э�!MMxX;�F�(*�h�v?f��bHi� ��?�-#������oѬXNW�(@x���D��MC'��ɞ�V��aD6{� �}���������������+� hjPZ���K�y^�3 �?+;yJB�g�E�>�� (��O�`���Y�n���EN�����@�a��K�6Æ�]�c1
ɔ���[{�)�-$� ��w�&��/VI�cm!�� s��c����b�<.J�S�Fya)�RDa5���N]��-R��dpƚ!��;��y1����5�SD7^���kL�Gw�FH�F��GK?
��{���g=8$��"�X #@��s��kB�{��_�/���k8�0�SO�d�C�Ș#Y�@��m��g]'d�\c�'q���	��k(�x�P��#�-}�dE$l~��|�xS�����ij���
q���d��`�X�������������{{��P�ţH#�h�naY�u_�=�$�4�FM����qߖ/�4���w%��fLሺ�Ԉ����h�7F�VV��Mܲ������\�7�xD�����TG� �W:�ؕF]���Ƃ�F܍p������$�c�M.�� O����Dd�bG���oR߁*s�O�2�!�y/��=>��:�ˑ��*��B.��]�^��O-�W�b4
����C�S
�*-���n�����K�l�X�*���#ճ$~A��߿�zX�⍹W���4���5.Lzs9"�oS]��� n�?\�Î�ab�g�;���_����S/]�B�B*��J�d��&�P���GN���}��lZ��dED�-G4�>鞼��4k��t��ĺr��1)�O���ء��6�ʃ��;yۑ��n�X��+���~�����`w$��7�^?)2N���x7;1������Ó����Z�bE�.&�Xo=.��7�p�l�[�*A�)X�U�(8��C��~9���А%]$�i]�E�Q�ÍH����띷�r�1����{�X�R�+ �RCƂh,ediCs-sU����'=X��d�8�H:#��Ų�ם�W�_Y��&�91쥠��)t�c�x���4{���j�~pv�F��+i�걒 jP
/ۯ�sֻ�#�5�d�����:]�F8��,�p���[ۆ�+�f��g���-q3?4�E����:�OT'�L+9��9?���a4PpFk_%yx+�q�E���\���S�A����Cn���*w�G�q|3���S�#�\"�o<3PǱ��}|����[����[BA����2s����%3�.�|0§�Rg�( ���9@�S&�5oߧ3pv�u¦>\\���N����+-W�>4+Bܭc�4�"��)B��3N��������L%���bǄ�QK�'�zҵvOn}�)�Ɯ�j8�U,��ɛr��I_��P����~/�mr�[4���X����w �J���@�.�B.��o��3~���iC��m�Ec�s�(*F �7�`��sZW�φۨd�E�H��Ԯh���0�ȸh!ގB�Y3�v�IH�����Vy[�`�(�������3���1�"��w���/�������@��`ӏ L ��/�� �E����U�ȶ ]$DZl����X\�x�n&RB`)��J���탅z�������O� �'�58��W��&��=��J!�4��4ۋt��}^���Y�XSl�TiL0�p!vj��bu�-¦������SZZ2�e���N�Ž����E����{J+;f����6^�͡:�CO+M�,�{�Lw�K��؜��@4^�ѭا]�b����m��1�R
r5��6�	ry/�]EQD`5^G�u���v�`[���[)�i�}��r��U;~��tJ@i���=2 ��	T�h�>���q����dth+�����6�K�@�e:Xă��g�P.��K�\A�)u�/YeSI��&=g�7��$��H�nn:��q��'n���E=T�|ۀJ��`��]����Q{!��Z R�No�-��̆���I#RU%N:� �����x`���s��)�m@��F` _`|��F��QT�L�#��+��m�$��+�|�ܒ�U��̄h4�c�$V~ z���\�߳��̰�z<�l�=�$W��lʽ�3{���Ute�,�t܂�;^	̢J�r[���K��֒������� ����b-L4���3|*`�3xh�_����wI����[o��S!���caV����
K�l��=��V{ҩ�N�*��ի'��@�nڀYx�!�|]0������σ�LզtL��p�[�2뚑 tWf�ϰ�w��<9n������R��r�E�|h���D������02���N��R�E@��s ��V�^�?�k�f3�,&�Г9t�衹�A�.�}��p$,�9�q��SWӱ�k�8s��#�CDI���Å�w�x��`��μNj i3o�6�lg�?�B�m��X��{=������*�R�y�/{�DO�@J$.(�I��͉u��G���t-����n��}S2e��M��#��z^}>��&�a�O
=n���	[حTj�ZO��h�M�n�㝻+����H�byj2j�3U��6�l=s�Lz�?0����|��F����Y��-�'����˞�П��/8�gӐY��ۗ�A���S(�P`8�
M,:n$0�� &�����ʲb�_�9܌���ƕӓ �23�S�=�}~������'���DG_�<_1t.��<L��5��6VP'g6���|)�J����`58�c�= (�cZէ:�r�""����N�(��3���Đ��w�`�^�uR��z��,���t�^O���
v'{-=������)J�8��Y�hI43.R)�v��2*O['���;��v�"�U��*>5��aG����pA��&lY��S��i�X���NQ�j�D7�
3Vu��g�x'W��G#�~�����OY.G����'a��!��Q䲑��1�y������)I��r���$5!\�Դ��P�u��x�9��i�R&v���aaq|^
����͗�����!Ռe��+Y� ���6e��� K��A��B�{o<�R�.6قBީ�(��HF�G�V��9ٱ�ӯ��Jy���|���b�e�:��GI��~p�! �A�qo�˘X��>6���A�3ŏ������K�E�pOà��8?�aHeG��Rs��գ�y���� @6�M;�'>:o&�.=���b���*��@BjzWc9~��m�}Ȧg�&j�e� �4��0����ǽM`�:�Uz7�PJ�byW��Zx��-e���W
y5љՍKżWZ�9;=�����C��p�ܑ���05��0��g�p�"��R��*�N]�!�3m@���i��%0q>�H�5�T3�����%�x��[��bE|�Uj��e��9�뮅;�"�q��2�;�=X�caZ���X0�/`��.t�f�)
2,�� �O����D1��Ĕ
/��"���B��3�<��[�SdOv�x\_p��F������� ����aU�o��e�\�AHF�7F���m�3���.u�p����f`I�[�V�<na�7��R���/ċ"m<uU��6�( �C�g��kb�i>>��Hy7��$X�}�;K�_(���#۬t����vyj�N�#(}�	M�X��D��XW
��&�B�B�s���Ǌ��)E��u)�賯�戛�u,��G���fL�Vt2���2B�̜����Y�l�E�{k<��f9�	�@��[��Y�%k�e7�d���3+H�M�'`�.;Sxc�X�4�<s�����Go��;]���^���v�-7����i5~m��N�c�{rǟ��(�)���Tj�h�^��6)���j�[�����5�=Z��R�Og���(�J���9�K�o3�[��5�{��<�uz�N,��el�b=w�S���W���4o�նb϶9���t�n�>=��'�Ss1�i
�mu��� �`'�3F:�g�ձU4;������`})Zٟ>a1��\��?t`+�ʰ�6�;�O:}��iPe
 \d�2�U�=�Dt��7���jˁ���CP��xv5�Zj�$7�.�_��&���Zs�O��	X/��+}=e�BeT^��x/6E4����'=*F1r�[|��& �J�P��Ԟ����Н͎RɊ�r���b���0�௾����}?�[���<���1�b�:V	
=If�l�ǅ���s�)_Q�eZ���+��;�� �U2"Q@�=gp{цy{&B���*�
��lk�"�����;
�u�C�P��8}��6�W/*1���*M�
�%]���������� �c��}uA 鷨�72���Ǐ�O��غL��]�)��1�����=ek��fo�n��Ʒ�:��;<)�_@ɗW��IE9|�6$�D���*g�Ȱ�y/$v��aޝ�ĭu��N<������x�>��H.J���Q�{�tִ����8O/fʰUtk������UZ̸-�K
7��(t��M�-zDŅ���О��
�N�sA/>WO	pl���棤��l`tI�1��QY�E"Ī��c�ףNW���aQ�8rs+��ve��k��v�xl*CK�a�JSce76ꋕ�y�����d��L��nx�xz�i{��
��B�������5:8�h6�����8~vB�"���CQ���]��|c7{�����>Hq��3#7w�ʲ�Q&�-�Q��J���n��~������_KEٸ�PR�w�n����ϒ���Ǎ��p��	�o�d7�.6C
������� Mq�d�Lxp�����[R��/�D4gcV��QZ��#l;�}�"\��>�g�Npٙ-Y�9/��a���B,uo�OwZ���~M��.�:N7�����ӂ}�v/�X� �>��z����v�r�Fzڎ�����Ӯd�.����紋2BNjA�Pmp5�2��#��t�K{����ꐔ�4~;l���Y o8WFGP�D+�u�F��	À��۴m`[K{����P�X�Y��p��-�?�V��Y�.��Z} f���Kϲ��2�����X�;�����m�ˮ��H�8���.��ߋZ}[8�|��e�I������-Bhg��۞cW��)��	��>dX��g��?.ݼPa:�_��qxޑ�7���$>C�\��Lp�YA�X6��s�7�N�KQ��Y�o�6Y@%`eǿ�tQ�MI��fF�r�2;�����yXZr*kӬ-g$�Zp��S�x�ɸ�ǉHP�C4]*�<�K�3�:A���~'_c�>��J�: �>�Kv�+�� ���w�K��[���� ��Q����SU�0G�&���	��q��O���K�Z}CV�{Zpo�5s.���B��>w�K�؊ӂ�V�E�C��/�K�+���ILV�3%ƗH0�M�<Ѹo�����5.ŔvQ.&�]���?o�<ys%���R�Es�>j�V}�� �1n�i�J�y�m�4!_&�@
�k��o���t1��47	ʕ[�V.��K���NAe�2;i�302&��md�"�Ί�z�W���O���vQӯ5��8�(�#�#���&����Q�|ǅǹ�j�g�c��f5Ҏ~ޏZ�}�a�󰵚)���}]�6��603�pC�X�y�h��1D����.�5 �%�aU�ysԖg�Pf1( D+����˄L�j�@��=G�MC�ĥv͔c t/G9$�r ��{�E�U��q�`~�WY��0xd5���=U5��H��U�}����ҹv�ZX�@L�P��*�f�3d���rk�U�W�$1Iy8�
��#c���[R)�;[Uޞܔ��D}FB�J���&���,��V1�@�ܕ����`�A�x"7B���`�B﬿{����j�3� ����e��<�t�ٴ�������K�܁^7�,؎T�����%����Y�1+J����<P
��Ծ���$ϯ��������f��)�AZX���9r�d�IP��@[N4*��� w���0m��e����ϩZ&4J������RȬ�T&�8���t�yS��_u�֖#}Y߇�~Ɠ��\�g���Sl@پ;���^��;�w�s������c'���G)���>��f�	3�=�Yw۵V����-��~��ֹW3޳6�]���t�|-R��埤�+t4���k���r�ݟ��>����M���I9��V_�G��Q�ޯK{�+nXE\^��f-R ���5g'�|�l�(J�ڒ�?�:T�Qm�:t�i�����i��D���ghTz�6��X�9�)i�&���؆�SF��k���w�cZ9�A��]���l��9}(? ��θ��3֝վ�����$������z�Qq����̢�nt�k~��z\*�7�X 7�
�:����}D�e8�+�b	ϛ�g��~�x� [�������{���|g�:�����`e;�8��G��+��ؿN�I|��p�p*i9�CB����0�y;mo4�l/Λd��	� �E]Q�t�^ _�h'f�=�c-�َy�1��ET��ej��X1(}汥�r�al6�i@?)�|C��E��x�;ԅM5$���(��|����)�,v���FL�_��L�z��ڎ$غ%��+G�d=�c�|���]��[)�.�i�6ԓ��y@s��1*��5X�p�ܑ4�p����x�	ϟ�A�!3����&J���.j+���F���)�*�����w��yص/�E��xc��f�l�`5��=p� L��Ҏ9��x9i-�m����n�T��R�f�H���e���0��&��D�=�%��1翫eZ~�?@�	��w�(���:�W�a�E�t���Bj������Y�:��Q�tly���dt�����ž�p��Hk%�Ez�##�E�b�#��8�A�f&�˶2$�I~���A]����-_�\S��X��|fO�?n�(j�Ч��-^!�E��-�X��3.?�J8�c��(t{���V^��(��*i�n6���:����z�~���>��ݽ*�M���'Z�X���-}a}��E "h_�f:�A����� t'�4�&YnÛՠ�͹���< �;j2Fa�Dw�u�]�$�fs�<��t�s}N:F�"�9ن�ˋ�	Z��N�5�e�[�pЖ.��.J��L@2�2����C߅�|MQ��j@�eK���`�*��f=[�oY˵��]pA��Lp�A�Fc�z���%y.�Z�|ra:K;��(9��?G�Ʉ��
�}�i\�"�?k����ܺ:΅�����cb��w3��(�̲�ܓ\�vb�zu]2�%��K�_���ZP��n�7�V�d4|Y�@#P��f����`�1������/�W��,A��?lBp��;���f�1�a�o�$�t����}��1(K�bv�P������^G˿w�u�� ��P�؈�P��}xb�$�bMHX��_���hM(ٻ+�s(7��f��vV��3ނ2KV��b�=""c�U���/Z1�̙~�o<�Y��>���U��1kxF^���Jh�iV�&x����z�����}����2.�#[ѩx/[�s�X�0	Ͳ~�%�7��kAL�>��#y���i�����v#柕 m�쐏*c�ރu��#H3T�@7�{?��#X)ho7Ã'��Z��M/��dK5aR���6�)������U.Ƥ� ��Ik��'2��f��Z�lM������QԢ���s�	�:�q�4�y�ϱ���Ea_h�);5�D�i�j��� �Fg̿D�iE&q�������������/z�ʜ�2�5I"4F�V�,��s������,ش|��G��P*���t�x2^�C�:�o������,��T���D@�����`e&F80���Fm��o��g�ڻ��^�s�d%��4����x.�{���5|���z59S=� ѭ��cS1�S���]*�8�'H�Q&*�og�1v.��*>7�!�Ө�,e���ITR�s�{��
ͫ�a��N��9,����_�A�V�B�)��D6{iq�_H~2\�+���)ݭ�Iy�{����f� d�]A�RV�)E����� ^�o�	�,"W!��n�>N<KO}s�L<yW��y{dv�6�����Z���J='^�L���M��5�1m犌�T�K>����f�4����	����=4��(Q���el���U�o��Y�y�c�0/�Fa�������5H���iF-J�֬|��<	���L��jV�)�:8A��T�3��k�����!��pQ�8w�r���	�m�D�${����Y
�3����V��,�?�Eٌ �ϋ|�Q�mC7���G�u4�t�	�7Ӻ�2S�Υ�
e�7��#AQ�%=��.sa_�1���MMmL�;�zQ����|�J�j�!X2����N@`/'5�ϰ�(iC�ҝ:P����!i��ԏ�:Lb4��%��А�?T D�������J���9�K�t���gts�y����U�L^#���d�`S!��~��C�U�-X�-|w=�������/����7-}�>�O�7�Cߞ�Q"[�&ڱ���\�>s��V!�z�&������fT ��]wG��!��Y^2��\����Yޭ�+Uɀ���n�Z-�f��Mx�ᲅ�B�~���U:)�-�GC/�C[�����B\5�M�� ���8���?��k��y`ŖY�����&�X����&���+6���X9�	��]��TIY�kBP�N"-�W��w���e
s1�o-���}N�Y�"Oꗡz���-����RKP}:G�G^��r��K��A3CDt��~����>i6��*냎�3�'�gAز�g��E���=�-�߫%v�;�U}�h�����s�]�y(��#^#�%��^ߌ0���~Fq�T�V�Y�;F�NS ����8;u^*���������{� q��^'hb_���n��%í��֫,�
����rJWl�o���!i�<��m4دy/t�zY{`��T��;�����be뎌�0��gV������I����VY5BŁV�0�t��@S��}��ple��<�k����ح� q�܃MlgK<{y�}�7�v�^bsP�3�Ƭ�3��}�A#m�]�k;C�M΀,����I�04}��?KǙ�4�T�c$��]�]�� i�n�0z�ɧ0ώ OdS{�;~L��d��Tȁr.�?Z����H��ݻ��r ��-���O�s�M�ю?"��b����\�49�"c�Ɲ8 � [�Y^� =�\Q�+R)'�C�@�kC���Jw9�-9 �@�\J��1����w�K�I�/m,�Z:ai� ��B���I�"�.�P�I�55I �Y��.hSb�+�A����^;�-Ls�<I���g��ͺĚ4�D�I_h�+�]�� ́8��ݍ�ҍS:�r"m�d�Ea.���)��,G������{'��v�*N�aq�\�I�!P�E�+�X�a�ڜO�������\�kPuU�?�D�)(���J����?�t��_O$�x������Zi���,�����ʎ#@o�\���q������Q��/EY���=?p������h͙�F3>�)��$(�V�u ���J ��JY5�~5��N<̨F�E�=�@��-�k3~Z�l�lV��	���s��L��}l�N���*A�K��@Ģ�zI\�z�r8O�8�z�b�ę���WA(�fS����Ś�h/��6^�>��#e�Q`�jpy� JSt��T��ѕ��M��� �\�@��C�,տ����5�F��Z�����"���Y�N��z1�ΡM�=��@�N������c:�m�d�I"L�p0 �:���}�G��y��P�Vb��_�JՂ}H�u�w�k�}[���l�.��f@����N�벆��L�5��r�C�U�����ӓk� H��/j��R��̨��ɷ��*r[U
Q{+��\�P8Zz*�4+�]���o�$���H<1�����m�m���i�����:�}�ܺ!������!�����޹2��������	8N� �٩��w����:ʰ|׆E��J)dD��F�k��d�[{��)�ԯ�A��rT���4�@��D����Å����񔵸�����[kF V}���7�[�	��m8��oL�]Lz�(��^O���֤""�u�Y姗ha�h2͵��@��kϛ|/Cv�?"fUى�� �\�L�ǋ�3C:c�L�� ���%�jc�6L�M� ���[�;T���x]#��UJ"���X�#m����P&�}ҭ���һ֘qS�N" o���E�3��a�Vx��ۺnu(-9}Q�L���#8'Gм�!39Ўq�v�K]W,�"遦+�@��H�k��Up�q��������w���i�Wr�:��BǍ��c�RV*I�NP_�<�{>俻�KP��1P|#�#�|��YN��}=p�BJU�^�|������im~�%Ѐ=���'��3����7�дY�$��* ׃��O��)դ�����x�e�U�@���oH�`mF� �mM����W�]T�I��9p��R��v�X,1-���K)��U��n.r1@.Z$}� J�f�xJ5���srٹ��?�'�;��������@�z�0�n�#����h=�eo�����a۔�����IRr	��8E��%�?+��'��b?'�Y\�,���\[}{v;��0����%>z���nds��z�7����h��Ê ��+|c9!�g���9�B+��R&u���D�\�6�ә��P\���s��0�']4�䥱���$٪.D�p�'������P�%w.{ܑ{>��`I}�	W���alx�Q}���t����k������X�˒l�$@c�&�'p,6�A�;V�3�T�m�|\����\��oqZt@�C/#T���R���+�a󧍈��5r����f�JQ|}��$�����V�9�����O��V
�:�Ĝ��$�=^�"�>�bc~ψ�F�gU%ƙ��g�f;����Q?���k�I>Z��fdG@N8��������}˘�,f*��5��b[�%�X��g�*���mQo��`�~g1��'��V��2VB������'K^8>�|iZ$��
2D��q3��7	/�m`K �k�K��^����?[���꒚�9�^��g<S����w01�!BE(rtFú�5Vw�xL�e��_.x����ʮ���g��-��pB�<��Nlu�܈��M4c��������#,3Dj��Ə�zV�uvoMm�s��v���׃��$̮0�q�M����z�-�	�1]s"���|E�D�$���?1��$Z�B���ѓ��e�²��	&�]��{��D�v�^Rz,n�I.��v��H�?�6����A<�� �<����1�}�bP8�3�j�-��h�/Z\������V;�EWrx`�5��!��������U!�Áh� �@x��>o���~�(7`��T�g#�ɶ��TY1	�=%/e�n�.�c��)����f�2��CLR�5#I�|���W�6�3DӾUw��V�U��C�
2�.n~%��s�e�������;�lAԌȈ�z��2]�k�T���� +��vD������vu+!��1ך��"M8��r�+j>�TN�*���u<���5���"H���[ޘ�r�	5�<`��#�\�e7���~Lsf��T�Y�?گ-�q`;j��'��BA@�F���҃6.���:�cԅ�Rq;�<�7
���zF�<���D�(��>���#U���n��r�Z�����6PTd���q=������|
T6������w���P�n�g$˅vI|�k.8�u��ҳ�f͚�A�9�gȞ��~��¼��	R��b����D�V�~����lw�z�	oS��ʨ�����P�|�f�G��9&�f�dn�`��um�{�$bFx�B
v��+)$���v�5�u}pS�ߖ���軅��(g0Y��*�4�nK�I>B�\A�~#�0?V�،�%˟))�!&���n��f����ܦ�ΩV-��g�2���]����O�c��p��51/W���!�Ʊ���h���6�s�&%�T�c[Yc�˱|�aV�Z���w�e�}��3�r�|d��$cЕ;���p��OX0[�����o�F�Į�]*{����)#�Jn�U6��4]���&�lz���B�����Vw�^̌uwfN����w��S�?:,�"�ʗr��K�B�/A��lcdj
�V��Ր�B���u�'s��w^�I-�����K|adʉc)�gh�g?���~�h�:(s�U���%�/�Y+�j�$N��gOƴ>�kx�$ЗJvRE^�H
��+���q��m*hd�����R��7�N�%|t���u�:ѫ*�~8c�P�`_?�|ܲ�C�Z��32�MW���z<��y��ɜ������[��v_k�d��G�=e&+�N��D���aU2�EO��
�� �h��)`dP��rM��ە�ӝ������3n��>��k��/�~��X�ouܴ=5�Lzy��ֵtY�����}9����!nH���)m����n�4�v}]���p�?J�8���ep+qY� ��-�o���O%X�iL�L�FU�$ΦE|�� ^ z������r"*�H*�c*���q��y�1���]��=ΐ�0H6F�/R� ).�D�����|�����M��89kZ�2 ����S2������o�`S�L�_���'�{�a^��U@��^�"�WFņo�"�����~?U�|U�仼��m�)J\A��E��2��,�m����s���R6��HZHds���y����=�ܯ���&&J�tC�	���46.��E?G�RPrI���f!��O盓+�]�Ng��%���>��qj"{%��Z"s�;c�e-3r���������On�^F��]%*���P2��6�Ld�o�bfE��\���ÜJ�W�"��<10��9Pڗ��8��E��,Ko��+�i�n9����5#���#U���Pô	I�;N,
p:���p����G(�H��j�{5��@��[�l��.�m����]�/*���� :�}�Ӟf��2�[�9ұ�0�O>�������q��҄����N����"�>YS��lQ�7�VNǳ_@ߊ&��ܗ���PU���~��&!M�,����	�-z� {�E�Ynf�#��gIh�k>��	�vG����EQMC iK����bӍ��t�䏐5IA�r�1�4�˟.4+�m](b���n��j8@��T��������VC/W�����q�x�GFBK
Q� Zà
�	�a��@c���5�ZDua�M��ɼ��rVؠ�YC(ə ��G$ߐ~4(;����=�jb���u��7��XJ[�
!�P<_�]�:�쪶�\,½:�IY�u� R�8C��?HSnm�㇥�D�K0l����~�}�f*�}ɜq���� 4\ʌ�D���"4�D���W��'��&�*I�۞�D%O�@�W�
��!b�/�ڻ��
?�8�?���'�V��GZ=:��+�*��K����_R���c�������9(�����"�`ip��\����m��s�6H
Cԯ̀Փ�����*�[rj3{��,�:2�R5��me�1&��G6�	�� �65 �&�FkLq�-����7U|(�"�ao�V���+�����Jw,g�F����eY�%���h����_'u��8REp�� F�vm�|�U�	�#�F01p�+�2K�GG7 廯vUQ��z��3Z@ �r�@X�(;.��q>�ۀ�Έ/1u�+d��"cW��T��`�e�M�]W�<��
YЅ�<s�:��cBi	�;'��Ĺ����7�'�S���
�2�b�	I�gѨ���
c��§M��i�8Z��Q�/�+�FE<KG�G_v޸>�yEr֯�������qT,%�7����}0�F��C����RUJI>Q���z�L����5�Re�_\ �C��=+_� �1��� ��UL�A�@,��@�j!�ޒ���/P'�aWv���౅[5+�j$�6����K��_-)�1�b0�9�hW�UnQ��2Ú�J]��A�3�c�.�{��@Ò��2��;�~��EG��2�Bli�b���:��$�[l��{��At�� ��LY�}��3��.)�y���G
5ݙ�{_W�s@���$�ws��3gg6�q#��1�6��1	�Ŗ���wk�ן�=���Mh�V�����Q�'���UE���r�t�h����C��v�� �{p#�+p�aR���3Π^[l�,��yA�.Y YfTRw�tkg�_�co�!�R�N�s��z� �X"Q'8Eb\��AA������=��p7e��UB��O�muc�����p��!���5���z3h�ԆN�]N��c�� F*x��"���z�Y��"xh�܍���N�sǢ����/��-#��K�pը��c�=c�����/�.^��-y�~J�M��8s��������������Ah��[<�����D;��Â�fq�	�Ʒ��Ԏ#��i�����[䔕�i���٠Qwkm���.��Ky���ĜL�/e�7����an#*���%��.F��U���jk5��9(����(`L��o�.᛭}%��� �'��=i�jRD�q�F0�9 �c��������]�~��C�A��-�]�s�o����$hUY�|���~wŹ��;�J9G�E}���%�����L��f񒿛����-�Q�&���g��ET�����!�A�K���9'�N/k�p���کA1n��72�O�[6���bP{4Ӗ�!1��X|6���H����?��#%Q���>�`�mǺngr]����z��B�wQM�kCo����-��OՌw�*�������j�����q�J��B����7������˸��%��sm�+���+>#�	�q<H�A�+)�-!^��`lME$���QY�iΪ�r̷�;�1%I7��|X[��Ց_y& ����$�V	��;�|[�b�ṛ�RyZ[������Q��g�]�~32oD�[ӟe�K�úgm�D�w�@+Rj�%����	�	�ʐ�� �iR��� �Μ�kAv3=U-�����wA������<?P�gڬA�9*:�%)P�4y��Aݕܕ柴�_�+stH{Gt1�ǧu3z,u��Ji����>���=]V�k��լ� ��Ł���8[~���2
P�7n���(��Sg�8�=Gv���Sf�R$�����%q�]Ǒ�.2��Ŋ�pK�.��C�w�H��O�e�єԩ�J�˙��Sv?��#|J*�t`;�u�s �~6b@���q�u���[�1��.J1)���(�l�FQ����#��-ȒtE$V/��B�h'�]_�~ԐT�t&_7W|�k]�͙�D�d]���yۓyʄ�`Z6�`�m'�Vt��ٞM��Z- ��s֘,@-Y�|M��{Ofk��/_MMw?� ҁ�[%nDoP3��@��$����%jj���j7�\��Qȭ;chb��1�޹*�yQ~�b��
���U9� ��zC+�V�f��d_TV��g4���=}�"|�3l+�ӊs�N�>}�v�<t�uDo�a:�hb��u��@jJϴ�!83m�9ڽ E�n���B��������g�y�<�}
R�0Z Y�5�K�^��u�'o�/@���Udo�A��!
�U mI�Ѹ�ܸ��v 06ߤ�~(�E�����}`�sP�P��S$�E�.2:N#슊��LZ����MQ#r���m���+�&�pfa�C�"���;�=�Nv�j���<��8a�{	���5��}onV����g_�Ǒ�R/�^+H�	O�$������}16D��bLg𿟞}z˄1'qJ���[�x���0
�|g����U^F�a�5 ��R[O]����^�b�k���rf�0/%��>��5����mv���W���`�CL~�$1��m<]ֲ�_��%.f���@ )N�k��Z�oEo��!�����]cKJ	�C���P� �h�jE�J0�y�f���'�������,v ���	�:�ռ���5�̗�Z�1�f���̲r2D�=b7�꧚V�a�H[�;���lsY���_��B�#[m�=$����npYc �����P����3\�e����b�p��י�:�ln/��o􉠛D_11�!4|�ca� (���^�������懿*�FI��Ra�cU�}���,�����Dԃ(Q)3e��+-�%�I�'/��)�PV�H<o��&yc���q'���fN�@�7�i�@��ј`9�L�^�5���ʶO�eZ�wF��u��&�O���ܝ;��㗁�(��f+���E�0)4�i�Q���>r�|����!��$ȊwY(�V&���q��qw ������D��Ո�{z���=#�޽�9�D�e�b�s��Fl��8獽�w�Rȧ^��Π�K���rqj�#r�Aw�����)����=�q�j�<%����(�U�C�\�X�z��N��Y�FE�4�G���]��ښ[��1#����xS�Y[t�r ���K��u�0�����j��ECNO��($���s�?��=̮���p��fV�G���]A�=EͪX��~!Լ�0A����f�c]c�Ԇ���NcY0�PP5%�dp4�4�|��5��Ι�̕�l�l�zJ��7��3�0����F�;I�p9�\�ݔ�a$�b�}�nQ���`N����uy�l%�1ʧwj�kn�N�օ�{O�c�m���f+�����/�Nl�-F�}TN_�I�l��[-e��0�*"y���.�-n���0䯭7!�A��x3ڥ.d[N�i2
���ȥ��G��^MjZP�a���f��\�kY����_Fd���Wb���<j�G�ћ��� �|S��H�-�2�_q���\��xeWi�9�rf̛fZ�N����ͅ;�����Y�QՂ�D�{0_d��^�W�;����\`�tW�-�@,> ��\��gڨ�݇����jtS!�܋Z=DH�fS �dO*�9�����K�Fdw��!=�#Jz��y�Q��SH����ӟ�y�;����p�K��2\�MF��;c��D(y�F�m�U��<�;x�ym��$��Bf�� "��9kN�󦼵r��\�M�G���n�ߣ�Ҥy��yM�`PF��I���N��rXq�����j��M�p]�G5�f�!Ј�o �MG��
��-v�ӹco�5��e�Ҁ��齱V7�L���齞T��u����I(,Z��4G_)�r�: �}UP �m�U��`N�$��B�5ǯ7Գ�������%}���m�����g^������
�bgeI�(�.r�e"p�l^ރ.��\���T��)�1�p���u�;K<??o�8����E�BX�pu����	���E.O�l1zUy��(��o
�73������r-)�5� �Ӕ�3g�!߈����+��.�r���p@\�ٟN�m8U����"��������g�#�@�UZ�����1A9���<�lǂZ&k�T�^�_���щR�y�H�g�^���e��5��y1�
�%T``
gK�Y4�F�X�~wO|���ˢQ���5�yn�CP���aR��[�$��I��w�"n8.[P�u�����|��8�?I͔���Pd�rm�h}�
�t�,ܺR�X+{��b��WA��)G��D�?W;o���25�u��[�VKK^�#Yw��cYЮ.��]!��h^8�aܻ&gC�����~��i�G	��s��؅u�����8� �ӊ7
�v����L�p��#n���n4 ����5�"HH�^ώ6`T� �$��~XzȫYS�e�Z}�C\����ھܺ����_T�U��lQ:�{�0J��Q�!�K�o?a�6����)8fOs@��N-���#���
�ͩ�A�]&W�z'�ܔ�0����:UG�&7W{�{8h��ʨ+�s)7sի����%v.���~���rv��a�tp�H�4 �d�A��v��`
R��4���czb���032���(�'5Wz��nh?����'�����I=N��_�Κ�E�� �0�P�U����8B��I%������Y��e� ;������X��h'Q���v�w���g�x�ٮ�Z���P��!q��Nb�̿M�gt�?a,s�4�e�+��9U6rGQn��z�ѿKߵD�(w0��3�H*�c�C�F��eF'�بN�#ڥ��`Kn4��Y��`XQ�v���YY����.�#x>k'�sVՉ{��9p�<d�Hz�9{5��{x�ܭ�jv���/kQK4Z��Ҍ6�ltŤ#'����Sz�h ���]��ؽŎ��B�	5��[�)y��#7�b�I���
����J^kӭ���<y��h�ׁ�	߼�1����ѻ�E*ӳw��oX����#��^�q:J��DD~:!�0��.���R�b����I�c����n� ؎�f8�&](<l*��j�� ����Hae��	6f�P��aG�B��t��o�ւ�`e@��6�rz|Z
}Q7�@�B�k��;���.���G��
���YJ�D�� 5�ow���x�%�G�%���ı��a� �}=�ri>���i���U����p�B�����Oc�ٌ�'ʿ����L�G%��^:C��Ie�p��S�5�����ɬ�^�:��b�+p,M�~h��J�e�$��T�NOnp� O�5!��뉞\ {��^�(*g�%�2ts�KP��׻8ab=�����-��W��2Ԙ�L��4*5e`E���.J��\�*�ԙ����LəV7� �x����� �xdhu:I\zӼ��;�+z�����wE�Y\��e�HL���S�O�<�[+�I�!���.!��@���NiE�\��1� �d�53Jj#�/8�7]�[�,�D��QIρ��)a\��d�)�*۫��>N�κD��0C�i��qń�������M� �##�cہ�0|�Ԇ�/����3�󏝪���?�Ͱʴ�'H�@Q�[�99��[����`�o&N&,�g������>z�ߓ-��y����D�A#W)~u`
7��������r���<(���7>���8`��L�/� �d+@�T{m+��
v��ڸ"�I*�ɱrh���̇��i�b���Qa��Y^�x�+1ő黜��
^��>��`���1^��{�O	 ������i�Z&��?F�\�hܶR��䦢���&�ō��2�
�jןRrs'�kI��R �ܔS��[9~񋙛��5�Q���gt,�	D��y&Չ�ç���ژ,����K��7܁@{1 'γv�#��e���B7Ȋ7�т�?ݿAi>���ʬ7�;���#P�t��;�l[�@���=+�V�O����8�ߒga��;v��M��-�o��
K��+K�֮�]`V�5�h�$��m7��d��+B的Z�Th_%\��_!�?i�>�l+��>l�	!����4 ?��n���9��p}Y	�ˎY�ը�K���w�ˡ[�K��2��؊8�a��S��L@G㇟3��0&B?2;��/+u�p�OwM[;}�L/c��v��Q��ڱ��s0�ҩDó�3�ֻ6�ߕ�Q:����Κ�J�.I6Ŭˁfֿ�6�����K2�����!޳HW�j�J.A:�g�� :�ö��vb�7�Y���~�B��;��sp����E��9r6����.^{�I`$��1%����&E�ʬ׵�ؙ��]��Ʋ]��;��J8h�T};��9�U�bN)��ڹI���o\8�!�o-^�3r�C���fDW�����>ݹІ�a�'gA$_G	��|8���+���������>���˳ՙF���Vձ*w��Ι_1B���u�u'k��+��_;��0h
4e�����YI�&R��22�~�s�����	cΖ���^0F���&�`�@����,}�?��������e7�1:�F�^�-ː(���V��;s��mϏ�������,/H=Z���ᵔ#�g�"�Z>�!��M��l���O�ޚktg���`���"|<��~۾����?�<�8Ui��\z
��'L���/�w�H�Ձ�����܍"Y�C�;��uHu�+��/���*��������-p/�&�;�ch�/��Qoic���ٳ��/�����άܻB#��N�����u���#��g-��`8�� 5m�,ba�����z�B��2�GY��4з�_�\G�"�T>�4�nA��2
ך�S�:�r�4��_S���شQ��ع�p����v�BA���:�eQS����D�T�H�V����㾡?6(��	�@��zϳ��[^�]�����&��
!��p�
,�/�J�\Z5�M����Y��P1��RHM�\_�#��^���[l�Z�0�O�x.#�+��K��׸�n
s�A�J����R�R����n�(��Qɴ)�*���Ϟ��v.k�>��:wඬK�U@x��?D1Ʊ�q�MO5�C�w��8����B���@W�4����Oȧ���%d�j等�<ŊoB������Esy#��ؼVA�`u�X����S���ϋ��;	�i!��Z���3���8���F�k�N���4�	 ��˼$���S�zW�փ�ڽ%�y�inV�Zo���VoJOc����`L��)�.#�f����e�0�U��ЊZ��Tȷ6c�~�jf���E4���g҅��zc7Vh�m�ձ-��Y��k�ar�Ŕ����.��F���b3�%R�M�z{.�8M��3�X���@mNs��j������ฑ��l�p#�$��OC�غ���֭�Ӈ1�V�>���J�RDgg�']s�ND��e΀q�n��}���񑯓iF.?�4��vv�7kt�/O3��	ɂ��yzc�5�}�8��Ii$���r2�?�����82�r�k`1���!UB�#�'�Q�����G=��f=+Лy�L5�H)C\f�3ڣ�:|�B��j9����TE�j��tP��BW?X3{�ʄA_.��lw#��Ф���cj�+z���
��L�VWP�F^��,]c����ff"W~��4}h5m����Ϣ�g9�f�ߚ���O5F���Rkv2e-*�����)�
��:�o�m��6��;sG>����S�0}i�����FlQ9z�NZ�+>��\ج���T������5��O%u����a���.�2�w �c?��4]n��ڝN�æ� 4�ž�I<��<pSګG:�G�Ƚ��C�n�mU,ޅ��炲���n]���ԃϓ���|]�b��g�B�O�(2� F4�A?�)�?D뷀9R��M2&�]�]&�p� ���t���
.v�<(	c�d��f*�L��6�@�qF�
Ч;���wX����"��6˚��n�݅��v�"����T��	���Q�'��:i�P��� bv�<"+�ҟԶ��J2�@hjK^hM %�n�	���7�۶K闟��h�e�.�M�F�������$f����Υ�Q;��[�f�PK[�'�\���^B�|�R���m�+֚�nc��@�5�FZ{��/k�Ha��P���4��#����%�����L9b�T�g�歰 dp��t"�繝�V/H�~��:�pQ����R�m�3�Yh���c�����s)�g]�	���x�ԓ��X1���D�ȓ�ҽ}\>��d!���;��&�c�dv6���)q<B�u�U1�8�j#L��Zr�I#2��6��j��d2~�1�U��"WS�	U�Z[6J���=��]jն��I%��m��Q��}9Ǽ���	�6�$.�ӿ-�ڄ���d�9G�I��'+��k.�����e6-����x�2z,6�_G�b��pQĢ�-ݟ���K�3 @�ʕ�M��JČ{ֽ�s��⿞S�:�8W�]@�{�!G��r��^䅹\_��O����i�Pf^�o�3�]�jވ���~��4��.��5N"���q��F:Ҷ�+���(+��z�8��֔O�Bo"�G�䍅N]�����Л@�6�:������5���כH~ͧ�`s��D�Q��'�@������I�g��Vgk&�/x�c��Z�ͩ���O�A�R_��{V�  ��W ���2������=W�o�㒥6�cr>I}�ީ52TV�#y���K�H�:�m�7��"�fr�F�#�����/����<H+0�w��z��ϩ��1�ݍ�f+B�#d!�����oTr��p^|Ől9�������{�ǧ��]䧊'���E��-�s���#�XVD\�eWv�1s֡;B�r{i��X�_���7�2P�W�=�vH)�;_����g��n�;�P�F-�@�*��II�˗
�Y�\�����$�%}�����5�y߰�r��ϋ]��uw������'GV��4�i.�xy.iĝ0����	��Р�<	}�{X0T�lؗ����ۉ%�R�	@��cedT��Z�6�;zp��o|*nQ���hd����hM?ӧ ,8�~��û
ޤ��DJ���Qt��s��wK��2�X�ņ��3J�2��DVi�ĈS�F�� ^���,8��g F �r��e���<�xR�/oƂܣ��2:��<E����cʨ�[��Fλl�mQ�}B�����Q�������8[/u(�
L7��]������{rR/�jD�a�2�fm
�g]$�"*�	Q�-C�5>�P-��sb/Ns�_4x��ǀ�lO������|�cL�S|*`E�aRM��tD�
�ݵ�1�n��*f����+���
�����{��5��#��勺�HK����\'nvg9�ݼЈGE7v�&�\���S�ջ��HOtR4(#�D˓~֥����=��}5�Jb���2��q�ں��Q*7��4����Nk���X��Bp3ݚ@�X���t��O�p������t�/��<�'m�����|��3�+1ͪ� �!�׵�JŝS0�-��3���wP%\D%���+��@��$�6��z�u�(���E�O���� ���Mc,�� ��$dq@�k���BH��3_:[��/�X��p�u����w�w�%��� ~`<���sHJ+�N�s>ؓb�尡H�\_��r:�OO\��?n����lJ�2%k�H��ާ'�-������'[?�a�n��F�t�ޘj�O�{��,���U�R�e���~ ��/)����dD��6�H5ɾpD���m�I���ׁ����l�UӢ д9G���>��mU�\X�o��R�5BJ�,_����q�2�{_����w�T����W'�f�ɫ�I*z�\��|�N'�-���#�C�W����[2�T��w۳(F����둪ڠ���2�/)K�L<�DX�������nﴖڣ��>�n͟/K�Ň���(q*�5<�mύ3�adu�Y�����ŪH"��4�`f�z�^�濗
[����n�;�@����0m�@]v]��L#�\�o���e3�d�Q���`k7���K��n�,�n�BӹP�i��Yi&M�=�e��;�8N�2�3��t���~f������.Y6��LJ��?���I$��3O��q��)�q�%�FT�:B������3O������uC�x�ۯ�]�2^㾎]�5�D�&�k)�`RYŃ�;)U7���'K��U�+����`4�P�"���3Π����'�~]�ͳ�d~�.H����\~�I�A"���&����X � qQb��B�xh���BMN��e��.��8D��E��t�42x�y̏&潍u@4��ֽ5�8��b>����KnR'��[��[���d����?�!��
g h�n6�Z���t0�-=� |vi�n�!&�l�)%O.��>M����r���B�`�ttI�%0\��%+Љ*ak�
�&�٤����,h�$�hI�K��Qi�{�uh�����X���!�+�v)<�!y��j������Y�1��w�m-���ĩq�Кm��
ìQ����큒�9vR�����;��{*�)�~�O�h�.�u����C�'�#����q��a3�c���b���c��)4m�78?����te>��^�b�ڄDR���dΙ���Ly���p��u�F�J�P��jHS��}��*U��~|v�B��>o��f�g!�c�m>#x�B��1�sL�ES�S�1��gm�|�l:O�=_F��\m�Ѷ|��Q
h��;����V�	xp��*�ã��̬��:U�������ml�(޽�l�n��ŏ���Xu�(������+�uf<�Eh�S�z�e۪x��-ף�f�Ji���N����� >E���K�����#Bo�9Z=������/� ƨn~��í�:�u0ڜ*"\��.jG 
	ER��;tX�+��ʤ�~���va� ����+�/벾g.�W��ú�Rj�N��*l�Ig�<,�u$x�*
[c�V�.�I���:�O���}���7l������]?-�]2��m~�u�e�/����z���f����V)
C�ʻ�%!c��=&<�I�s�܃~Ң8",����g�����IJe6���<�2��[����$�t�^�-\�v��aZH�[����Bu&*q���j�,��7R,�bVTiDb�D���RU)�CDl=`��.&�,P�W�^vq�@��A~Ԕs�9����*��^�����M��_{�@��"�$��7�fѭ�K� ���%We�0d���b,.;�nGu�S��HЄ�������W��I��9���Q�N��
�_e��!LNrtk����On���0e�N�<�j��Aw�72C���q��1x,��:D�^1}��0s�+]�j��[���f:vAxk��������.��^���hyM�EjՇRC��J�q������A/�K�KELW�3dԛ��iPm��2 (rʒ��W����&k��e��Re̙|m����w�Z�g#�7�J���h�B؋���x�q��m��98���<Ǎ�-�#�:18a��룫��/�9�I3�3�8�0�]n���vh�Z�'�(K~$��V������[�����zw��0���\���xU��}	\�A9�QY�b�̈�p;^q����Ț�9T���<��a��۞��A�t��},�~�8o�����!�6�9�4��3�AI��6�a�x�97���jM٠B:y����6�5�_ԽP۪yK��'QȂ�u��L�^i
}>��HkS��^tB�K^|`�y��W����V�.rq�֩Z֑t���֌c\�La�*A�#�e2E
�XZ�=���Q깨��o�Zؓcȓ�]�[� ݇I�T_�M�
r��.b��� &����_x���(��Q��d7�)���8�=�<���v��O�B�>L��2~��>G�������<[���zE��.ݺh���$"����u��K���:\��:�t� 
�Ͼ�qk;*)K���f��B�`C���^+̌Z���� ��uY�0�'��g+�%��y
_�i/�ͱ}>�fJ�㠈��gLJ���^��LMn���ŕ����H�8���ˎ��ܻ�%�r��}�]i���J�E�Aש����FFuV�Л�]�?~����o
Ұ�{x���W~�G�?n��DVrx���2��}�a���C�=�� ��zE�����I�oUr6��s�8z����͙gB������ZL�^������� 6�HK����ZZ+lzf�h׃T�����9���?��A~U��e³r��	 ��3<^n33K8e�bŋ�O+NI�C�-w��^W�Ͻz�A����0t�m�=w�|�	�E�#5���:~���������dE��q(���}Q�%)&,����b+��[���`�SC�#n� 
� |]%�)��R�.�g��z�j뒁�kmM��o��Ĩ��y�2�9�St���Ih���ݧ;wz@d{�j��T�lr۾�h*���3��8���l��C��₅5zG��f]�fD����A�׳�ʨI�A^�|1����w/�X@m�s<?	;����&n�L�Z;�=:��z�Y8c,�]y�C7nS�����!�Gȣ��L��5cd��Tާ�� `��9M��&g1D��>9xDۙ%#��T����)���Q6TG6�)��I�����i�/��YG&����2��LM_r������~XK㘥��oV"����O����Z���ʐ�}���*J221�߁���ZŖ�2��5ӿS3�w���
�M9�B��t�ۈA.��C��0Jy�17g�=|O�m���-/O颱���e��u�vz]��.i^/J@����b�яE,h�]q[�dd�LT8�\���3`D\B\���t=K����	���G���5B��7�f��b)����>�Na{q�t�X;�����+�z�aQ��B]��mP�vM����ǭ��,ް�~��]�m[�U�[�M���֣ _I{�� ���/ڑg2YJ��,6��Hi���W�p��ѕ��f�=$�m����8�x��Q]c�{�b���� Me��=8�*x�9
������6��j5��M(u/�,��A"�b����.�2�d!�+�cңFZn�̾�M<P˾e��e
*gsЦ��u�_�v�^v%ۙ�Fx(Xk�Q� ІH�����,�Y3�>��NN�c�@�zZQz��0����v��RvIT]i�[2ؾm܋ݰ���C�k/PLS��D�v���7L%�Q��\�
Y���r쌧�����aH�,K��u�ĉ����\���"��w��!y�]��MB�M!+G�OH������w~aK4o��N�N�TF��0~Ӆ�-��e�X�kE�>�����x]v��$]�,�Q�V<��z�h�:����	Ⱥ�L_�͒�j��Tl*g����-��qח�Ө�����������a�s������z���3P�,m� 
�k���kE��2uA�s����_b�����K�/,���ѣS1�= ӄ;��F��U8��r���_,�Z�ɖ������He
�{4�0�?�MQ"r�3�ޱ�	��q�RQ��!Q3�R�@�ߩ����	�)�,�+��v'�H�SҀܦ���ج�N͸����n�Ai1�H��5\��cћ���M3)�k�~���g}��yn�>v���N��}h����^d���H^�ͺ�r�\���mw�mR��:PQ��;�̊Q �o��0(Q����me>Cz�d��K@��'�c�z�r�_u�&X��F��1߽��QgV9@��|�����n9+�Y�1�#
�Mf�����[��N�C7�ʎd5��t5d2��(��KE�)��&���$�u�y�k�z���Td޹�#�O�b�&� 1��uL$���(t��O��Jv���jc�v����LA4
��Zj��g��F"��0�~`%�AC�8�ݿ������ɶϺq�
��>0ƃ����3T�R,AK碒PhЗ� mҏm5��"���7�����ޣ!3��̓��5hа����x���[�S�G ��i]�'5�!&����zm����f�E����Q���y����rn�B��'M�F����|ewy~�]*�ي�vb�7�0]��R�ChU�@�e� �����m�陇� ���q؛w1Q촥���̽�3Y�J�
��2�5��s�z 9ޠd	)ޝ��V�Ԏ�����97s���tE��6y���	���pT�;-�P����o��Pd(�@���Vnj�\"i� 9S���1v�4�|?U
-[� ��OLP8	�,a�GJ
B���m��rӡ P�1��(��&�{ѝ���>.�_��Eapy�2��u�$F�T�	t�4�T�R۶?w mP!e�-2@=�3m�)(�y�O�����������D}2҆�t+X���#�
Ц�8&r�um�ޯ!<�qm�FT_�?���ϝhS�h�k�b�W�u��Et댠��K��٩Y=�9_ho��-�tֶ�������r�����|J�B�I1�_�ҏqx̂T�\�����_zn�z��/���a�9V6���M�)V�<�Z�_��W���.9R�0�����B�ɣ^/������K�Y�p��%ܔ�)�_�/e&g���a���F�S�c��vE3�������Qf-���S����1��jF�z��B�ؔ�/;�䱅�2��D̆UJh�A�*�K{�K׮V��������L��-��)O�-����߱���,��tI�h��d��Zd��>�����:6!��Z�,̴ߌH-�	 Es��Q$�q.��~~��S8A��A]��|���q�!���=�!LbK���`p��btaӍ$�l�2j�ER�T� �I)1!qZ���l�e��\P�s�@��	 ��84Y���Gj>�f��`�"���*ە��6�NA1D�LRe���%��n����;Hz�j�۾�M��YA���U(|�(
M��\���WU��U��Ox����R� JL���@G���S�@�C�_�����H~�)>x�r5h#f�\ޥXצahh]�qM�u3����:I��G�0N�2��E>0W\�R��O��-;���u�6���\<JJ���ζ�a^+ź�ݓt�pW�.����t�Z�S_wbzI]1llQ �Ab�A	��މ�C�h{H?�����'S-��.kJx�o�T�ᩩ�~�{��
N���F��� Ra��w	�g#�e���:��G>��k���'�
�R�$���ҹ��	ۑ�
5��$��b�ݾ�k���̍��7	�eh�(RQv��_��l�bf�Ez�u�|^w�v´���6Ls��"]]����x^�Ǹ��=�ߢI0r�Nw.Bu��L���A*���M�DpuO�BG�O�=;�4�VW�$�)u|&Q�H�u��M怉��9����$���hv���u�T�6��~|�ߣ5-G��-t�5	jD��4�A�г�j��\Y���qkDo�Tz�r~�ݒ�Yg�]��ؿR.���[)?� ץ�v��+%_ɔ]�%����: 2Ë��%
��L��4�g{I�٭� �X�ڻ�-,�B����y���x��C?��QT�Рr��٭I?A�o]��t��#&�XRq����j���[�$��J?ˬ=G�&��3���p;�(�%q�h��$��
��[�JI>���HvvF��H�[u�Q����G1/�g��� D�"��|�3I%0���!Y����>�3�΅ֱ?B!5_\��n���9���Ђ����wH+I�O�,d6���p�������賋��I$F�8�Y7KY������piCN�����W������}�>;F�8Yļ½�KԄ8	����c_7�M�e6Zm�9�=X��ֲ��,1˝���A��s�o�mY�d:��IN]��5�:q�O��H�J �f)^eX·mm��m~ߔ�AS`����'�d{����;3�\H6�m�MO�C�ӜB=`���_���(�l�&�ǧ�ܗ5�}���
��%V��n~�FG0UFj�ȅ�5���`jo&+u�J���#,����	�"�2P���섵���c �E�1<$����x���L~2�j�Z�#�*vS�ԑ��O����z*�)�yZ�-Bc�ʊ.�����
�KXQ'$�g���%|��v�8�`�������r�*<E�E8�-?�ql�`�p�=�P>�j9%M>7	:w�����>��iH�#��E�5y�|�(�z5�u!��@Zy��d̴���._\�5	��,���E��F~�̙���-O�_�wh�,��}��iK�w��s�6|�q����\c��r�1^rAj���̬���a��)��aJ^.Ѯ4/6���BP�7�6r<��DIo��d��p1G��!�+:CEs���U4�·Ki�~���2���X�SJ��iīV�0�A��#�LM���]�N�`1��Um�����kw����F*�$�M�)$"���FP@����c����+;u�,�=3���BB_!�8�q���W�c�L�rt>�i�4���v�.=V�QM٥��䄏 ��G���]/�*_~`u����/Ih���7���(����F��	���X�L^7q6�(�o��T�b�[�w�����[=��(r��:&�^�T?�<��j��G����E�(�M��������IlyF �f���7/�s%9�l�!s���9+[���@�>�ƻ���d�$�����x��!���7����G��U;�C�EVi2m�oo4|�k�6�56L:���:��f��-�t�[q@x��t�Rn�9�u�V %+g3n����bL4�f��"P���]U��8��ʚ���}�/BF�Ɩ� %rU-��t1k$��xKz��S�7
jc&Iˎ��Y��L4��q0w�$nwlMU	~	=2U:֨B)��q�2���H"=�cJx�Fr={�LvX�2S�� ���HJ;��Q��ʠ
 �o�1���A�Ѱ	>�[<�N�u"V�V����'Y�hKX����L�X����xc.��,�L{̫ॹ@��9�u��X�����ou�Fhd�"޴�̡.�$�)���#t���+�
#�3'���3�߈�
����p���DAJ���>9���Ɓ�����g9!(3.���q�kw�dL��Ê�W�հ�-Fx~u����V�"����S������2�QFf� j�f�f�y�\n |�X���6in�iH`���a`�Xn��'�Z��K��6�\(ɺ�v��ʁ*58HM�&�.�%F�<�\�\�--���,H���<5�x��X3�_��V�H�����>(�q
i� �g�~��-<6hgC��o �񹃎:Q(��R�HSu����"�@~=�E�#�z7*w���I���)�b_yjyD�[�i�F��q e&��e��XV�~�T����fd���A/����OG�Q�42��Q�z94M�`  ����3�wG��6�x�kH
^F8��7ꔱ����m����Q�f�O*pt�4S�/���O6^���b�j�s��*���>��b��:���=f�lʕ�O��áU3>���P�~�4W>�Yd6S�|s3�:$~���Wn�\6�o�I1�o�&̡}������Z��$���o��y�����mπq#VW���c�S��;�Lz�:'�a����-����b���Å�y�ǜB���T�4W��@+���|��y�/�m���יI�:즡�t�S���=|7�F�.��⮦�Dm������;�2�+4��͸� ��=�^p��S���nl����*�]�/�����L��x)׏�����}��yE����4���hp��w�?�:�J�\䉹�E�ECӌb���'�~�^V�M�M���/n�\JY���;��`��! ;O��&8n�v�	C�:��|~ ��L2��ߞ��H/�r6�7�'�:*�fRb�SA�Gt��*�Yi.:^�R�d�U���]�n`V7i���/�*�\����m�`�k6C��C_�nש5Y�!9�B�!	��֐�T]FW��\�4�D��\J.�_�5j���sO66��wQ�B<ܑ���b�~��B5'�l�s���Ǹ�:,Ĺx��'}	�jtē�w~9B�E���]�.+1��Дf�^�*!�F|�m�(#�n Y\P���c�ź~�,Y�<��1���Csۧdj�T ���`g�f P�����]�\{iB��	J�q|�����L@N9�o&�N-�KRlI�M١��qx�CI�	9S��-6��~;u>�@�;����i���	'+���k<=WM��c�.��;"��Qf	y)9���6=Vw'�[W�$��m�s�k�9��C>/\��� �1x�ߺ�T��Л��PN��w��m���>1❳d%����x�jMD�k�Q���O/T�?7�zŁFna���X���-"U2�>�	 ~;�-(U^5"�m0��a&'O^��!};<4'��bQ���S�����Ar�ǱL�b���S��0�!<u�g�!dɒ⠰T�Q#�e+i�S�j����4E��b�r̵P+�q��]s����׹�F�ވ�u��?g�0-�g���Y�!J����pی�Ѻ��n2��j����c�J���s&�fP[��V,��df����7!l�4�i��LM��'�c��@f���I\����R��2	۔������Q�yڝ��L^w@�Pr<ޝ�c!�	�����;���!�jH���v���/����������$��*8�ש�1)C��G�Y4	�|X�ٺQ%���P݆#U�i���CXQ�"b�9�>l�3IcF���G���Z[U-��N� ��Z��i${�*�䋞�-k����'����$L��ۅA{���R|"��=c^�Ma Z�/I"z	���N)�IO��%#���М���Ӑ�������|��֯~���7Ui���k�Q4�M����:�b�T��6�/J�� $5�R����7�BP��ǅ6���M��~��� �'�yo�w}�&�fyN�
=����z�e���M����w,_�=��i�j�m�neD�}Eb��U�0G���J�&�o�,,H���Ê�:I��6@�i�(&KG{�y�_�D
i9������ݓ)N���{�.���Qt���˛��@e��$����Cȹ!s������[��Ґ�[pк.�5A;2���^�W�����h
�����a��t��mZ{��A��ݝ�"����a]�=��	�LG�
9(u�zwS4aa�5�OnH*�^ݓ�fsa�����b� |�È����Xa~m�XV���8\�횘?rIB�Q�a�N7�Gt�6å�L\���nnW��S0z*y����_��S���:��F�<T�Z���p��+(jFᱛ��P?qr�"���VZMI	��掶���X��)�������E��=��s�/��sӅ����,�
��-����(�{(֛�%ʢ}5�&.�L�W�#n�4�G6�ҷ�i˸y�X��т�H<��D��o�=￧��P���2}D՘�4���M�Ҁj�RNX�cMAP�q�ȕ��}���Xa7^<���l%�O��3ؐN�<�K't�D8/�J�S�8����F��M��-���_���{�8��?IIa�N����?��dt�1i,�p��o��}����Ёq.SF"�����Q��e������ǖ�\�[ 4��WE��卮�חj ���?�T�znm�d@�����T�|�s���lf�d�_W�Ƞ�J���A���j��}C��b�N�� �ߙ�B ,'�(�"���VE�6�osu�n�����~/�]Nf�tCDUC1h
Z�����~�TI��㻄��� �_��35H�1�?���x�1�L��=�7'6qd��=�WS����s�uhA8 �ס��c��Ɔ)��MĂx�O�^�_4��g�ѽRf�����\����u��n��Z��t���o�l��Ȯ�D}�0�30-1©���L�V�J�;qq��!�3�r�����<���3Pۃ瓸6PX 4�,�n�a�.��fU���[.j�Ę����ﷴ��1e��qAbH���V6�����]Q+��}x��X�O��~j�Uч-2RX1wu�3��|��n;�'���@�]�N���=��m��A-�h�k!�U1Ԛ��Yq�1��p_�P�M�=����������
=`C9�����}��C����N��zuo#b<s�V�� �%�� \�����q�L��	u4A�@7ejN����/��l y���_���W��A+7���H��\��x�#��r1�4L��M���?��t�jL������kJ��P_�MN蹄]�;��9�$����S:�\�4L��u����A�G޹��Q^S�N[E]���-�8�`c���/�c&�	��`{C�y�t,#f}O�c���4��N�I:X=֙�w��U�b@߷?�R�^�`��� K%�Q�0}󠕷7&(��b2ا�jQ�G�c�ۧ�3z�����P��� /�R�Rl�d[���Ę�ˌ�1&0��CH�hz�=�Zl[>߱��@y��&�$$
-�«��5�?K��ƺ� h+V�ɚ����K+��N��m2}��{���YV��0htx1+{`S�Pm{?,H9�`K!cỽ�Y�5Ak���;���z����:h�Z���0��d �06࿮�� �$ݽ�T��2Έ����B׺&����l"9A��z=��AE���r>��Fw�E%��U�����|4�W�������­���c=���բt��\x��7��j��v���p*G�N �;����fK$_	R��]���=ڶ��+Ǯ��EB�*za3���/v���Q	7��g��ED1��	H��BW�>��'�a�l�jʻ�D��Q��6>���/�UA� �z��8�t��	������fx�u�6������Ȫ�`/��r���`�	rȗ�8v̎�~SF/�e+SP�j�|���u���z�7c�72��XH��o�C�_^�@8�kZ�0�:��� 5�}I�c.L��^+�=�ޓ5�O��+�F�7�� p��Z�N�`��u��;���������y���H�/�mדڲ:�ލ�޸�*G;�Vj�4�`'�`����VV��VT���~h���>�W��1����z�(���|��C̚�Q?f�^�Q�mȢ��[r���	
��$Ȥ?!i�/� G���|�-��*��_3��7�����|d�T9���S~S�b��ֱ⦸���K��<Q����p�`Vh�8)Zl��܆�����g��Q�)�>h�C��ޭ��GkX\K;צ�O�X�3L�5�?�DEH�u/9d�ny�2^g\��[s���b�^�ɗ3I#�sX�UV���7�ӢU�rx�ٔ>�	Њ}�ׂ����a�ߞ����7�8�x^�P��YK��I<�0�)؃u�n*2>�\�����>T^�F�^S��ܸGƯ��n^�U�2�;\|u_�"���� x�%J��R��80�.nXM_�R/a� ���]A�),�8�k�g	@�k��>	��`�St�b%zÈ2���ܬ�n3;��Cc~-����[�${�����@I��K !�Ag�{��*��@�a��Z��|=9�@��֔��C��{��94[��(xK�P��\��/��lz�{�Ɋ�4�'7ҫ��>@W���A҈�Q16;qz[}�prp�*�ekꓭ"��t*���Z�@��M��%Q���xFp���z�P�����_���5�Vu���> < ��,0h�O��*�ߛ��k�ԧT\��g�T�nP�?\D>��m�`h��x%h�Ò�\�������"��/�#���*.yp��R�Ϸ�\��8侕�1�J��-�VG�~v��0�N2(>S�b���^���Dl>��f�;�K�r���,f�JB|�����*?�o��`���4���(ug���������!�U�	j#4e�p���Hg*2�8\N�^bW![q���=�5C!�Fe{�s��=\%��b��. �U����9�19J����#b���:{����#am-a�N�^nR7[e��yָ/'�>�$55�����
Z����bh�v����ٕm��f��S�I�@g	{
���D�!�c�J�U�I��nfoy[�ţ�=!�y����B=&����}pY�RrPĤ.��Î�^�U����E �[���Z|�;��z�t/�I��<cy���A�z�p���F�[�UT&+�������\L�J�����)w;?q�b!���7f�ƣF����� c����\/O8BDV6[� $	i�]�m�jc��;>`٪:P����)}`Ԯ�IK+X�Nz�hDғ��1!/��u`ڜƎ�,u�Y�;�A����,��	f@-a�
��X�{�	�0︗-t�ߕI����oF�� �)��
h
}��M(����x��� ���6��H�``%̯���>2�5�����? vH�ubݨ��Q��J��T M ۥ��E<�O�����3|>��9Sg�:�Y�uv�^��ʲ����D�g��C�MEWЅGc��Lp!q�6Wv��A��@LYS�m��UN�yG��|���k{]%��%�ߤ�|��̀a:ANu��9hLqz���+{v�ot� ]_���,��D��63��5ԥ!��ΰ�����᳈BB	�����Ѽ���S]��3�	�9��n��)ʏ�0b�c��J=2Dt� x=�c�S��Rq@�aŢg���"I�l�öʮ��)��>]�b���\'}��f����􏟴�w+[�Ԭh-�v��O�>���R "d�sC���o��!2�����a���Vm��s����}\ؓ��=³���I��e*�\k8	��D�ŵ��k<z.E.��dWr������C|M���ֹ[,a,�%��y.4�R�%�vR���.�����fv��d<D7��&�m�GcNн��������I��07�rZ��0Y�\�^�؎������#�NȚ<w~�I�Wd���%��o'�oI��	R�|��V�6Ѓ�^�Y)�����Xr4��t)/[��S�:Ä���O�M4��\���r�
�w���?E>yp��p9m2��=q�
5�$(���=R*@��5�_I������Ӿ��-V;�ϩ �7հL\k֭q�E[m������S`�a:V߰~5aPƃ����h�$�[�E�ĪR=W��ٗ*�i�E%a��0�>�S��!�����J*�8>e�
��7��Zч`�۟����M}`�T��Vߚ�oY7���z���^���j�Q9p��w��ιR"�4��-������讼NZ{���%����z��R���/:�@d�{]�Z<�D��h����)L5��_���l��Lg���jeR��y���Hh�ɕ;:BƧheE0���Z��Yҋ8���^q��𢽘���E)s��-��Q����ȹ��������Z��{�&������!� !K	hx�=wCY���6�+*�&ҾJm@u�Ëy�W�ɲ
A�Yڿl��8ܛ��s���@������g�����>�ǰ)���n�m��K�S3�ռ� ��ra��`�굋<��)t#�9��-�z=I�*?�N1��Oq��a3��D���#�"��ES	9=��nh�R��4��o!d؛�?�����%V�:�DW �>�ƣԤ;�Y�t�<W+f.
��~s<HT��ϩ�㾃���;w.�+�� �@y��dϜ�!������7�����3����>�/X��2�\~��@�@)�iTI��4��
mڣ{H�8#+�� �*Q}�^А��=�X��]+��H˙�Qr�j����^����6��/�z �[FVAR���B^���9�������x���읓��\�O�;$"�`֑H�� #X{Ǩ�-�5m�Y���}��������0:2�-�67T?��n���ۏ���]^�	�6�G�j��n�QLC� �!/�-ГO�BYp�c�h�$���1�����m�"�:��
f��Py8�.����A�ks���"����.Ia�������=�3��_���3D�yܼ�U'�p�%iK'�Za�����8'�B��U�5�J���*P��K5(��H�=]�|'����T"d.��Q��*!���뫦�����ҩOXi����-�C�?�7��p�n�ŏ2�'wR)8y����u�����}T���?�|��Q4�g�V��q��Ae�솧��_���L|�t^@Z&I�����]M��@|v�ǜ) sG]�V�V1Les�,���:3ֽ��;m<p��X���ҏ�;�ɋ}�e
l�a����o��qOP�*��ű!����C�+�M�=�"8u~,�ẗ́�����1��M�7��v���o�ՊF�y���%L�a�!U!���2�`��1i����Pr�uuEƚ���;����^E���3ըX����VYr�w��0�w���iE���Fc�	5[�IL.���#j��x,9)޻��$�^?m��F�΢P�0V�*38Ԃ��Gfr\���mQY�%�#�_���CN˒�kB�q��/{����]L/���ӱĤS"կhG���le�:ʨL�!˾�z[G[OtzV|��M�=��졸��ff�j���X���I�6h���-���p������Z��@�T�ɘ<�HkD(L4����o�a��Cǃ6Z*8���q�k&��͞��$hB��J��cO�A�J9�����*k6T��oc�T@�K�]:�G�+�2/�Ď��^W�X\�����G��1��B�"cLw!8"E��O�1��B�5��]�۳qlX�n����SD��tu�˂�#�s�rx����w�U��ؙ��pd��I]��)�R�&���y�[o�R�o���@�����������U-n��:�΋6�'��`ԁ�&QCsM�)5[�ax\3�'�	ެ �c_v��.������@�#V��L�Ey�>B����H��}T�',�L�a'���=?��y�E7O�U�p��n�g�Q�o
�ѵi!ػ*h�5���z[�T<�B��+�P��&�C���p-��|H��Gs��p�e� ~�o�I>�Lp����d��%�jPK�9{�"�|h�{���y1k�}9�0,e����ı�Fp�ЁH��=���0�"u�]��S+J��@_�z�r+�����𶣑�EW�.�f˅�o��U�S��Wsxkɿ%A�E��6R�9��2�M�1Ȇ�{&��gB�AP�������ę�K~M6���d����9���}���1W��܊���	�I�b��/�=Y�S삭 "{�f�Ş�C���X�y��B��f?(z���t�])��m0�9��y�.;���C{`*l��rW��K1zo,��}�vp�*�N�Jܣ���D�d+�w�ff�W��]����uO�̍�G�'O�&�{�"?2�lي�4ڶ)j�xl�DT�y��_z����Σ��Y�<*Qz������!�&�Y�0[ �B�� �p���\��F��1	J{@v�lL�S�t}��¿|�
�݉�<~�M�ʿNe��p{2�.V��3��06w?�+ ���8I>��kI<���N���A���lѮ� ]n��Ȫ��F������<��9S	��n�L��-�;}�=���N��m����y�|��F���>?��|�k,:-f��Ne$�|K���^��o�%b�FnԘ�PTZT^r��B��K0*��^k�>�4�˦Ȟ��L���k~7 r�ݭ�AQ�.�Zl-��r��5��ۆ�6��ӾR��ag��i����&����-�����5��WB%D�:�X�<��[j�%� �Vjk�AD���k��W����L
Ç�(��D;kl#t�I����4��}S��v� �rَ~
��0�f� 3���s�B[%f���F8�A�щ]j����cT<���q��9�&G�g��'�|�שݺ�JR�r��T�UN���@�~N�+v��\�8�'g��`��SL)M@�P���j��4�a�'k%���'������mk� ���]^�Crr��?����'u����������E*S����(�t�z����e����&ߦׂ	l�v��|���WP���#ӫp�(��8�F$�q����Z�N�r��5��~����]�p��d��§}#7��թq�n{�r*���.��V�d��N5�7пv  ��¤�Ѝ�8N����ЈUėEpA�Ek97H$�]s��y,��E�h�I"~�����̀��9��Ά��B̆�{�fa���ظ�w�^��*d��cj-��1�le���W6��ii�KKF��[j���OV�g�ͺ"�Dws�,�y�0b;Q�#�c��30]�Z�S�}� ��bH=�����Y|����S��U�$���S�p����EJ�[�P�^�Q9�X:A���Eg(l���+�X�z��í��cA)�����)0 ��^�!M��'=�8RE=�Ŷ��	�/%dC�q4�3��hxq\�\*@���'S���� ���j _�6N�T�-�X)��ws��6%5
����g�D}e�ܷ������f�(��Z��H|+��c>��{Qqf�e�����I�)�O��
D?$��x�V��,3���{�<�D�I��9Nc�2:�}І��I��ML^�E�X�>,�!��ȸ����ߙ��&������ϊi#��L�C����k�Yg>G��B*f�@�K���2�H��2pI?ůz@H�$h�J/�X�������#r�Gk12V�H+�5IkTV0�c�sؙ<���2='ң�5{�X�b,�X��������jv�����S.ط�����j��ǌ4n�ol$�8��gH	���[M���\f��N��d'����%ι2:�*��~x4��@+躦Ҍwہj{�����:������Ͽ^};�V~�ƽ�P�\蚚�x�0;`c3!F5x=���ɓ�Bf��~jf*#�N̜�!�WV慀j!��!Aj��`=�����5�6�<6�W�Y��'�2��� ���%�R�fbT��'a�?C��%q�����ǜϟ��E���f@�?�X~8� ؇�(D�`q�M�~��G���g�%�c6��`��0#�6����&��;J��)Η����+�Eb�p���1]24�ͳ����E��L�~�P�XI>����H��'еT�#����!�F�ó���j������s�Q�S���_������t�c �O�?JVbl�û�����+0��i�y|�],��`B��,��r��d^�z�8�^��Oh����lic�>%K�m�ޜ=�-H�s�B{M^������Pg��;�D�2�	��JȮ����ïi�b֜;9��G�E�&�jm�kF�FB�������Q9��';_���uQ��_��UL����h� *��@�Q[�x�wr����h��Yq4?.
J��%��1h�[pA��UF":���V���Mu߃7���L�]�\d0����d<g�v-^w|�a�|76Ҵ�(�8���B!}�"�)ad�U�FYq�}n@{�'>OG��}����÷��eV�~X�^��V�k���Nmg�ѯŃ3ẃH��2��s��9�k9�l��];m�"�ǲU��r�� ���q��C�{@���͏�����xU�h���w��7�סW�Y�z���u�{��:U֜�����#eu��Fǹ5��;� 0'{;G����<�W�i�G$7:�9�����n~��߫���1��'k{��<N�G�Iv��>A?^wF|�/�A&\8�����0e�X��g j��_��Dv||ԓ��� /��E��H�;B����ŝx��E߻� `~�bP~m�d`���hd9�5� W�����"^�ޅ}ŋ��֝�փ��x	o�`�S����/�����j�b���e
n��t([�<EǾ�3���G����.gWH[[-��Ӕ�R�uŌ[svI�:�Ҏwm���{J/���S�{�( R��@e3�,���g�M�����`���#w2�ı��jY{�N����D�W����W6L��۷O���,�1�Og�-b	JK{,�n�3���I%w����܎ ���t7�<9"�ݾ�(�7���%�͌g��Y���W�R������]z���6P���6i
�) �+�p���
W��ABuY��я��u�	�(���7a�sh����[�CP���fnkoj��>Y�1A|���g�N>��3J��Hz�+vî�j��wt�w��q��sk�y�:��`ή�5��� ��[���Z��T���{E8Z�*�Я�9��f�����VX������R̡�q7�T�]�5^�������`V�Y@Lޤ�p3�@R,P@���S^�ǖ0��8��<�d�z�^}�����i��H`�E��J�R��xr ��(�=����Ve��ԟa�8���D�We9���8���r?C�I��A9�.��R���M�pJ����;e������(���;;��2���f_[����}:�N������		(�>�z���ۣv>�RQ ]S�Y|��8�g]X��.�A6%F�l��7��Lfd~�J�u�D����_6���zLe�&*�j�hi�ه���q�Ԩ
F�C?�w����3_֖I �vI�43U�I��ME2�n^�N�H�rB��
��,�50?r���ÿa��Xf��[�K᤿͈��@�-�u̻�X�7J�y�EDtN�>!I{��H�>�o�p���Ak�@���!j.V�t����N������(x�����������8��C5 �{N��Z�H��������O��۟+�)�����T_,�G&|��E �s-]�ݚ�"p�i�Fү���|��wfkP{gYi?M��l̜����h��fG�ȷ
5�����ׅ���@,>sg�ᐒ�ea1�����i��Õ7�n[`�t�B�%�OZ�.ZI�<u�`�a)��X�v����QS������V�hs�����5�A'r����P^��w���{�ȽK���,��X�K�^��6�N�Ht����x�� '`V��1��V�i����ĺ��å�X£/�7ڲ��#�g,L�y,KD�o�  ���:M��_.�QGt�*�
�@�X`�|	���E�X+�������	ef���v9K%M?E�J�8GxJ�s�A�"���O�B��-��&p�"���ng7	Ra�=?XX����`�F�����7) ;�mi�q���d�[|I��^�A��(��^Df�+�JLɚ!X%��X�e��d�����8��5/��{�y2D�I� ���jg,i�#�w��,W�l#�'5�0�25�Vq5��A���I�J�!P���U�F�鞔�eШ�����{���ş�;.-�}��w�u�K���B?���*��3�}��1����|8��߶�#[�'Cf8�,\U�����=�z�qt|�`S�f�{�+��X��c��AL��Lvjd ȹ��C��h&pU�QZ�i̾��|�م�|�p������Ļ�&?��4���bP/TY���[X�S3������aq\=5ʁ�;��g�G��0�C+���o�e����ǯ�-C�z�yp%���Ĕoh�74���,=>ټJ�C�w����Q��PT�%I��)jM��PB��i���f�}v�pXgx�Ob��S�84���т��6�K�m�Z'E_��p��^V=��
L=�s��>1% O�y�d��{Wí
;�t�Zv_����d�sg���#d��V�R�����G����WUO@�5��#J �x��^g�3S!Ă
���VtѭP��fU�H��\B[(� U��῞�6�sU� Ͱ�������U��J�;�V��$�i�^�O�WIgq�p��І��Wq��I(�J�q����<SV��Ϸ�^�E�Rk��\<�����/d�Y?��w���ˁ�R{�Iy��M��6���m�h*w4��?��q�W��������ė���(R�q�v��S�Uh��v)�IVߑ?�\�U�D�7��󴨣rp��[g�b�,������蓒��N��YU�@�z���TZ�m>_(����0��{2�Gx�VW"�t9_z���ˠ�6Ǻ7Ԟ�.h�mܷ�i�U1�?����NY�R}o���"��k��a��k�6d'��E������Gm���ô|��4IX�̘4L�&�;Bp@Qa&X�}gN�A(�UQah���v�=ٯ�~v՗����$2�+oW^E5R�V۟�^���u��p����7����qiK�}�Ճ��=o�i�F:��Ut
y��9XO+��?|A3��Ĵ|�]7���z�S�D$��Aj{3���dtm|����� ��p���4�I4vo�"	o�0i꿾h�J��)~@���A����]��y7�"���sf(c悱_�Y��xH4EF�����OX-�*�x��yL��5jq5�	�?�`��n�we�#�������+���onY��y��#?:~,��dOpZ� ����Y��o�e�5mG'5G�Q��Z���,�b��e杨#=�ۖ�{�R	7�x�|֯�`�~��n��6��dR"��*t��a�lra�]��7(���ZH�q9*����"��L8~�.��Y{�b��Go#�L�W	��J�4R��U����f���j�иl�K���:�,l��GSw�[�It�|	(ү�t�^zʀ;�9 �Å�c��]E�%�US�xu<I�k).Qė-����ڹ7սz�r��vm��e�{/���aw��(q�q&2�Й��u��7�N��k�dib�oowS)��B�)��8�R6�{�~+�����ۥPj�Uy�sDiS�+c�fy����6q���E��㔛�%��@�&�|�x�-Y�4fi޳zQ��.���)�9E�y���=�;�	�_�4l��c\��$�r4�j��l�M�p�i����Պ 7��^?��8P����R����#f�ˮ��]}&� ®���< b����S��/zѕ4�N��~W�d|�����5�I����R���n�?����X,�^�>���.�O���J��0r���P��+�Fj���#�$��!U}�0]SwK������C�G���������qk
³�D����Z�H���Υkw� }g{�ّ��Pc"�+(^HWD�W[�L �Rۮ�\Rj�JL�Y"Yw�̡����]T���hoD��gΉ������4|g4���op$Nqfy`x����t#O�C���Ǯ$�{�R
��l9�2���Y�D8�Z5����Qs�&��FR��nnI�k�29(K~V��{G��%M�im�D�6?�4���+U�!�p)����y/�U0(T6(�y+_��En�$��=�v����Sr[���E��N�?ԩ������h�H�U���c&{^:�.&�G��R����U�/tq{�O?Byyȫ��^��.��c��")
?����9sPPrM��F�[�Nĭ;%�c��_+h� 5����7�>�nZ�F7㋝����4��c�&�tT��$`8��D�Z����1HS����W���4U�Z��0W��J(��S��q`z4vOV^���� ����x��a(Or��1Z&����~V� VOç%��x_�5�l��UC�d�rNūt"i2Qw�����0���i!�FA$M)K'�&�{�������0�����b'�%�cS�ޕ�V	Z^���pm��2���c5�w�t;v[p�6|y`�M�����Е;B��r���{q�gH+��'<Ղ/����gf���� ��lsՏs���LIbja�V����P.:�_��B1��8Z��Y��R4 ��'e)��Px8�P�bn�r.�-*�%�l�r[�0���<m��ѥ��,+�#�F�.\���Jw�M���o��%c�4fX.$������?D�u��\�[�������w��\�0�DKDL��t$,(���kuH��C8�5��m\�u]�C��K�C/���f-4T�ܘ��p�&9�pjn}HP���&d'т�"��
�gHw�R��3wCS�D�,3l<t�k����%�����)(��p7
#V����*l�I��K�Gd4�����Z�/U����L!d!�Cpq
ZkH�d>�␪���&�rSO5m�؅���Q�O���e<= �]X�%���b�mtYߜ��n9���ϟ�|��# Y�Jsk�i��s�^(�=��5�
m����va����B�Qh�v*�Эм��k�Ưd���3eLcId�5Գ�aw�1"r��|����#A{S�{`��.V}Mp@��݂�P��%HN�x�t���Gr�8X�-'�^G��ؓVF/�%v�Z|@�ʀ��cęS=܇���<��/��^fv2o�DC�.��w��$�� ����x�#�[�$5� �Tˏs�z��sWy\p^��<���P9Ve@^3�Զ��XљM��8?��K���߭�k[������>\B�mlS�%��K85�&^�2�X�(�hB�A���`���M�a�B�~����4�0n� u����@t�dF����s��M+��k�b����6��XR���S�	|^B_�� |JkCz�J"-��U�2�sq�� �t��Ƒ�u �b7��w���͆��܋�t?�}�cm�983�a�9�ϖɌJ>S0���¬�<a���B�_���P�;I����QMމޓ#{f��;�O��j��ê�~�2&��a��F�����?�b��1�����}��������A��p&�bT�;ػ_n�e%��m�#�}��f�9ܲ�u�.�.Vq�H�͌Ɛfj����b�:�1�zg�Z�\+�@��:���FX�k���x�ek!�p�	�����PC��%�
:�|;~A��t>�l��|�p�����͊�ϒ$'-N������`#�w��1W���s�[��؎�}��(К�$� �9_�X�)"�4J��~���\?��6b���6٬��۞�I;��
\W���I�����T�]T���v�Re��K�#6�2���~`�C@ή�4/�, S~[�N����)�n�Z5|��FN��a�V�8Ĳq�J轗7�v��a�=!.+�`U�����Bk��Z��Eth\+�n�q'Φ6�=&�{.q$�٦���4��6m��:���T	�z�Thc�[Z�#E�l���PTfLR����b�4c�'uV{z��8u����[�����d����[�]�x����nQ�r�/1u���_�š�A�7����:エ�Q6ʜi��.h2]�n��󄤹o)�#��p�֙���u��L���S��R�<���=֝PN��n�V#Tm�UEA���)��j���o�[%_������@Ѯ�᩶I���aN@�1�-���P����w�Q��b�Ng��6�eZwن>������^�M���܈Jvq��%�����;�4��s?�2	�-���a���_C*���-�*�ą>�{�.�:nC<j[�ne�oF-��5��v�#D(��'Ηf@���?3���)������Ր#l��Ic�C��ۨߪ��	e�t�̛�vf2�
�VH�ܩKjW��B���i�-�}��4} ��nR.ОR$y������@EA��C���̶$D�l%�� rT&�1�����/A�+>�8'�2���<�&�t�N����,��非�'��Iz5_>Z� �BS���51]G�Ӭ\B��0W���x��$.�!�4��ܗ��3R�=H|l1�#}KH��捫Ǝ��g�� �Tֳj���.��5�*!~<�
�ߋ8	�G�!�9�/� uB�0	��/ȱ�B��9X�Cz*���L,��V��3n���5����s�타�vφT��&[V�Iq�����:s��zb��6��]jz]YČ�^�.y�@u���8v��3��"�����`��Θ6F�D�]�`�����؃���J�C7ɍ�)yqJ��U\�,�&hDf�z+���+@Bua�����-���1��+d��L:��쾷nU�v��=��R~7��d�N.���|�����Ϻ��~�즍.�SF�,:]�g�,�&i���c"�����a���`L��+I;ʫgK0���]��R =�E����"���^S�����շs�隦���`���ø�F"������k�e5���հ����k�n��;���S�l$���D:��[͇�~�*&���$����e�q�k��L���i�OS�H��a�N�3Ԟ�1�k��	��1:9��(1c�	�Sf*
��,�����I����a�|i��CL��fs?�Z��EU�p��>�e�L�Wښ�k�{���PC�M����i�.�*�4_y�]����isimS�>�ؒ���Èg�Y����\e/�`-!2�[�����<�O�~�(��A��lvG��?: �T� ���H_�ۇ���(��`E�[�ɷg����ʖ6�;�� ���*��ˊ�3�e�a��4�����԰���<5⩛
�e�Y���_�6?��@�K.�w�r�O��ñ�o� x��@<S�����dA�ܗ<�@��i��t��2���`��6�8��	�q��&}^�O!}%�w�� ��P�Z��L�)���h���EoZ3x@�JIX���1�s�J�4C�V��^p���W�D lj���d��5έ�n�*6I'�ׇ�g1>E��FLk�����Rl�/I�<���F�ݢ)�z&'\�gd<�]�P�x���vō�A?��,��H�F1��2�������я����V8�C�yC��i�	�����b�R�	��FTr�oJ��U#ϥ�cz{�����nY��YԱ����������8jg�z��"r^nD�e"��Z�y�H�rTʂU�!�$�R�K��g������Mo�B�AE��3��c��s�I��	D)E��Z�j�䇙ύ3��
F�,G��0���/�Y3�M<R�����-���&��HPי��Kr0�s��H:���$��Az me���cήA�P�r,`�<����=��z��0VŦT�>���i61���h���p>ZK�� Z�#��9�I}��]Eկ~��J�3����T����&V2Ǧ:����&m�ۄ��X_���(6��]+�9[��LP�*�;#��h�J���;Τ�"%la$�v��0�]�v���u���TQ��ۃE��P9j�^cß%1̯�ވ3�x�;�0h�7��IKړ�:�k܄`ȓ��Y�'Y?Lc��#A4�u�y�����{�M�zAY��=��X}���0�b�o�t~*%��R���@XZ�'O�}k�;d�=�����Y]�@}/�:��؞ ��^�ڞt�l��Z�9Y��E)6��yKn�##f�qn&p}� �������=�{'8�<'�Y@�؅s�=oe���k5����p'�.��D��:��z֛�W[���JR�����c��!�nO3�Q}���J��t��=�:uMD/+FqUx��P��Ld�8`���n��
7�#�r�pN[�W�O��bj:�.Y���h�kɐ�-g�l�q���\�R%�`�|d-~���M}��ݱl���KS�9���E�fk6�;x�D���h���$vZ��͜W<�S�op��:��F`��U^A3W-d,�4~V�l�ܱ�W��VR��8_�,�tr
dկonj�ߖ�oꗊ��K���ZI�O�H��ʡ�^�_!�K"]�5�C��Uc����B�3���-t��61������/.}��;���~��@�����^ 	������������Zt�#z�4E�7��m��A��J�Oo
ºف�^>=r0��7�����%���& j�����߯X�9�:�0��1q�N�i������D�4�����D��/+��݀)��r���k�h�k������k?q����C���2Q �%�X�����H�� ���wFa�I����4H�t�)M`��g�l\3�x��&1��m����ɉv
�hK�D�{��)΄�g��L��S��%�)l�)K/N�6�a0瑰�Δla�)����v|mo�2���␬�<�� =S���{�8����^X㢫�E�+��p0��7�^�(L�sK}��6f,V���\�!�ܔ�_�\�:2`���@ni��K,�@č�CE}�D~��d%]W���O.5J��U�2��"��sL�(�+|ԟ�����,*�;�ڀ�B�]�l/��z�z��T5���p=�KG��۲Y(ʯ�"��:#�lz�}����e��C��v<2�?��3��A�����uc'p-�zvv#I��f��
�)PC��=�;���$,��~�*f78� +����qe�k�	L;�m��Dw0��;��h�d�%�]�f3��Q�+��'"y��2�������7%q��u�
i�?�P ����R��}n��	è z�_�	�[�]"Q����R�� �K��k�^�s#�Hm��]��/3�p�rx��l�H�K�\�����z�)k��C�!";C���!v �|� l��c&��̀�$���[WQ�� ,]�������6J�Q��b��)�M��`�?v�"5 �$ť!>��g�s�a4��p���8�d���y�r�Jہ� V��o���8�%yC��g�7�Bh4����4~�;;�Mb�8�݉$ëW ��'@�4���MB ur�����y.���kӤ�a�@j�e�ĖP���,A�p�w!��b;E�GyU��j[p�q��jW`�6`�?La�<Κ8�V������=O1��>`]^�H�P���'w���Ak�RD�j^����F(xո��K�fl��l�3�������s�V����],�}į�����T�&/BT���Gu�P��5(06�à�
�R��M���&U��V��b7�>`�]*��~>:�|b�䵭'��I̎U� O�S�?�5�vy�F���S6����<��	%��S"��b.{6���/脲�5�Ab[��n�6��y���An�}x-;����Dw~�&�����fS��P}�-[ΐ�,!���q����T�~�L5�Ih�F�kR������8�3"�`z�*���C0�v�=��.Ns|��+/��.H�+w�ѕ:��t��Wʵ��U;�:�c��� %�w�DJ�,���D���SDMP��Fv�0Ո}7)���9>*�_㛴YWD�����'K�~�H\ �!V@���	f��ѕo�\�W-��q-is��q�g�� Uzk���k���S���qb��<b�U{N[�^���[�4�Lz%�W���3�?�h6�_Dy�ˠv���>�Za֓VT�T7M���ĸv�@��E:�7�SD��5��.'�m2BS��J�@~c!%�K��Y�3��c�r*(�ȼ<��ɀx����\)�7��Y�B��n�'#�T-�Up�G��I�����Q�Xz�eZUe�f(��7�g�V)��,*����^�ȸ���7#�a�����-��UG���dw�L��;�$�y��´e����0c�V����XH�^�wC	9H��6�6L��V*5���	 zg;<	�O���'R�����B����C~����6ɠgB̥�FQ(�[�Xb��XޟnL�j|�3�-���7���B�K@�i�:���e��"���}��#-�.s����Ѧ�E���Ĕ-(��"�	�k�r̹<P m
�=�{���!0��W�忝�;@F9(ֿn	���e�Ә�5���ܜ��a�z���o�=,�[�\i���%��bZY6����s�c�֗.W�3�7���يb?9ۭ^��TD�fLc��<�:�L��U�ܺ<�]<L���Pv.9�=����x���K��g9^(�R��7eXb���K��lj���~C�;l�{P|0�!,g�����)QK����&���$�J!Z,@"��M���b��p�n3�+���Vq��6Qù\�������ڼ��幓�nh+8��F�������[���{5��kP�@X|s�23躎E3~�� ڥ|�\��Ʌ�
>@[?f��U!j�둛G�T�.;�� ��Ġݞp�p��i�/��a<�Բ�}�L0*��,�:��.��w�:��ţ߇"E�*6��j���Y�\�R�.�G�9쎚Vz]��v:߶g4>�B����ߙ'1�Y� z�J��_��^8���ʋ�]p�
7$����V/��	4ؔ�)ΰ��I�Gﲿ�i�#@"br.���r�ﻫ��rgT�AW�s�����[�->S�@˜L����q��sǃ����>A����]G:�(K�S�Q���Ĕ�`l\541���Q�]v�k@}k ��N��>Eu�~�~�F��ݧA6pdz���ڏZ�����[�/,��u�*ssi���� �Ō����()g����Y"��_c״�l�,��Z����&�h:��B?�nh���.5�%�	g�/5���ޠJ��c3����BYJA���cӚ�7�B<f����g�v �Q�]o�xY�V�A�嘨ҋ4
?���D�+ɷ�J�:�F��<���jg+Y�[�riW���\$G�B<`Pg����{�Ӏo᪱�'gК�1B�:@�`z�!I^JMH���a��{����c��{p�ۖ�l�C�������/��2����l�p��#���Y����3�;�����}"p�0�د�������V�B��������>\�9E YmzL�\����>�P"c�|�E�4Hx?��,-*�8Bn�Z�B��B�g����+���$%>�N��p�9$�9�٫X������"�,��w���}�y�
����W޾B��chcSϏ,9f=cqD��TU���"�F��a$f����	Fe��O���pS�gUw�ÿgd�%5��7Zyq�0W��;6m����>&��	�9[�Ѧ$)�
��-Hk��q���i�:''$��1�ߵFYK����@o�u��枝�y�3��UP9��f�S)�i"D�5��Tr(-HNP8Q���jQ��pe�cK�"1Q$�����5߈�pq���m��8��o�/�V�a��P�1�/�v�z�'8�(�XAp�y2�e�1�^K��K�T/ĩ�κ[�B`\�^��KOm$�����;:r�R���y�[H���O?�&8&.`R �{@W:N(���y�b�<郬R����3O���k�%V�@�������g�dP�Ӌ;�����g�*�S�5�D�Ս�"��L�6�5�ܱ��ˑ����\��j�����fp �+��wpw�G�����*�r����txs��q�8��P\�f.X������Y����D }��%�$��x���b��9<�2o�R�AP��%��b�-v`�h��l� S.�g���fy{m:g,eۓ�D�����U�+��c���N=%�&� SN_��w�3��5Z��w��e�1�>l�C�+H}��_�&�J�>h\I'xϞՑK���11����v%��E���XФ:Z�N�˼�r�B%�r�N�[����B�V��;��38t%���X^�b*\��%ZŻ�Bo7M���L�n���V���7�=L#<&n�h:��4��J��[bd�&>�������7��X,�����Y��bm���o�L���Z�g��۸%��>���7}ފTD��;�����q*Oi�)ǸN̡ ��[�TJ�	ǫ������,��B��__���И����M�G������?zL��t�s�j�]Y6TmqKR��]��#�� cx�P
�g�"��#,�81EE�A��8�:��P'6��h��P����؁�e�2��p��pGg�|JV
�t������2�Ď�I�H�<O<�ݑ�x$���c�����y�O	�Rz�.p}�W�vB5Rd���w�Q�;K>V #.ە��W7*������P�|�r�wV�Ŕ�Pm��%#���������h�����E1Xad��V�Fƛ�mw�]��Wb*~q��w��z�YAr�r�99�CNq�[����$���R�/��sk@��:��9�_b��_���i�LF�9`�'�\�`\!ТJ.�IJ7���fl$�=�LT5�;�[:��^6�?~���f�p��K����9p�?��lc#����һ3 E�zc�'��a��?�nBXؽG��$��S�$lsx��-��a��·����B�$���+�wh�#P����n���kSE�PM�	�|�W�,��Fp�6؅iE��M �p���#yZ�r�� џԠ�إN�q ^����-:ڸ;��X��� �2���6Ƿ���p�� ��K�z�O�%s��FoF��y%o�^h~BPΏ���i�mª픙���y�c5kBCP��yw�OX-k�݃��#��d0 5~F�Eh�f�A�V���9�ϒ��s& �"�Ou�����2�s/C�5�*��!�&c�xn"W���?'�˓!N#S[3g��\��HnI:�Yg�* ݬ�^l�E��@(k�����k�lS3������X�|�;jr���>���՞��Lj������f��V(T6�#���'N��+]g�)�� �( ��썥�%��hbL�o�I"i�~�v�-l��_�Z�-�r"�~qD���ɚ{���%´$��쿝r��@U�Ц`	�?V��zGq���ۣ�Ѵ!Ï�?��+7�8ȉ܁»Ӻ����H���[|>W0���辬.h
=��u@�	1d�G^ǆV�� ��� �G���G1�e�2W��\�
Q��5bB�N�QMK�#kj���hV���p|�̕'�J��~ä{7A��u���긢wc�,�u4!�$+�����\A�r��r��|e��P����r�"�*�8m��L�s@��2w��S��)��2"1�H�z�k�	(��z�kU+֚9�f���'^�(�G{<e����B�����P�������QX�,E��}< ���nAy��'��ՙ��)A�?}�1f��[x����X1SD9o -��r[ͮUQ�k�ڃ�TV�U�Ϣ�	I������Jc.��.`�F:^kK��q�th]�3G�2P��>p����]��<^k���˽��S�$[�5��j	�z��9��b���I��1RO�)6����s�+`�u�E{��)��nu�C+��wy�{�DF餍����쟴_�G[a��Fj!�B-�p@�ψ�l� ���Y�y�񈬙�HX�����>��^�6<^vF���	�F��`�L��qe:}hy��5v#�}	�*��;�~��/Y��?K�n�c	�7X�Sq�|=;п j�mG�my��g��M�c�������I]��6{`����Hw����t?Y_7{�/-�g6�m(X�K�D���Eɣ�1�[��Rp��8g!�3��CL;���]�J2~gt�����K�������p�m3�6�}�b`׊6�ld���k�e��\8��J����\!��T*4�]�\_��nK>0�3x)gp��V��,I��~��}LƁ�#��9(��I�Z�C��p�Y�������,��o;���?��_Q�s��ӭ�y��bu��E�X����ʹt������Lp���ɽ4�y>_����Вje�/�z'�]�p@DfO�J5դ�Y9�IkV��q�� P�\���8�Z`g�4�'B�CaGHߴ���a(��0�|�ӸY�D!�8����D�R߇�E̱�t�?�1=S����%9[��T�}_�������M���}�\x3����I�Չ��S:��9_�'C��x.la���y�i� �/n�V+K��܇Κӣ-�W	�����hV�?B	��>�`�1�O{�+���ޑh;u��d�h�z^�^'L׊�����!%�,�_����֦�D4wAD�X�kΗ#ͅ�u<���g�� -pIv������cٜH2�] ��
��3�a����^n�6�����̳N]�=2�fa,:���9����m�I�-��6^�L:�o2�`+|���/Ъ�7Xh/�`��Z+�z](��7��Ee1�����~V�{�H4G<�s��|ڇ����aItKz�7̸������:�[W���||���D)���������ǯ�۲0g�������L���FX�DG��օ1��ԑ\R�(�O{o�.tU`�	����7	�Rkb�R�y17ҀB�����1� ��_�<���7�^l�mő���D���$�G�f��M��������,\.�̃R,"���]����Of�L�\3��qY�W#E/�n�4U�Y���_��=�~�FӋٹ��@�M����Z�MKVā��KY�h
���A0� ��/�ۛWd:��\���\�y佛�3BM�&;a��B`
x�ML�Lv1u>�||�kv��V	�ݵ<pX1咽���ٖ\��-D��9.u� ���'e���j��(@�L�
cݔ��N���l ���ep��o�(�_��z�\����B���~�\��~��rh�X����~�7�L<�5���Դ��aK��w�м�B2
��Ja���ZL\�"�;ɼ���m������P���'�˩a��l%_c�ة���`���7��lUC�����_�����$�B��Z��FK��A��|�2d��v�N;����-��o���3u����Z���h�zAPi�_]����Q�o�u��Ju�w+�0W�����kέߝRXo=��P�	H819���3�.���h�o%" ����Cy�;�1�k��3�b��u)��d�8�)
n� ��Q�Z�x����;�zg�>#�F�.��׈SŶ�AC��MXCB��M}���R��oL+��ޣ����utNG�u���z�Z-Y�����y7��
�p���Ǿ�x�Z�`W�[�|�QЦzgc���EVɆi�J<�ƛt�:>��yB��C��|���Bg׳�V��?���7�c6�`�-d(�U�b�{ �Z]7/#4��"�^��'�0 C���1ڙ�yH,J]`�� z��^jo �q~�Z���R�	�*2��o�u".�v�F�!��+�*M�)t,�BD�S�<]n���~i(&�;d�8�T��ev��0�n���/�@��|�l	�M�A��U�O��y�n������
%�IV�֋�seq%R����0S���Y���a���LX���%L����<r�?3h���7.O,���������y�1�^�`�dy�R�V�N}�]�,��;�H3����8�3�[��+�h�Uo���N������<���H*d����mR�
՘�.��@�ݶJ�t���WC3�Z;�J�˶�*��?���m-#�*^�='���!�E��Fxݢ�+ay0�T/b�L|��I�rZ
B,�l崷�;�y?������������t�ZL���Xryݕ�)>[��9��rD�XY�4#ˋ����L��� �*�7~ EFnY� �c����N�����|8��<B*����Ζ�t�M�g�`GWJI�:�.�gb��K��|�`����e�eE�%�Ds�
�~tã���J�jw�r�Ed[k@�U�:� �%�@����Ѣ	~�āY��n2���n�ֆ�1aL���B�F�h�vC����4�2�Ů�Z�
����I�?vT��\���]HC/��˰�C�E$�wJ����_�h�6�q~�q���"̱�M!�TZ��^^J�e>�G,2I��X������ �șU�n�r�7�ԯT��pwTM���v��R%��Ⴢ��r�_��y{�D���g�����[�K�7 �0�jm��Zm�u}͹vn�s�������%���v:����L�����/����w<�k%P~���v�_����z(o06�������t_zG�^sa��:,6K��S�$����{�G���%�|?�I������\)܅��U�ˏz���O����ِ�GYvP����%3�-�v57GD,�@5����ېT�DV��@ F��$��#@��4�4��o狭��Z�3P�d���Nn� �_�Du�1�_��_,�Wgʳ`���6��׹{Z����ƶ^`^Ct�9��Os��ٓ�^ў��5��x�p�)��cZQg�b඗7ۇ�D�;�FZ�X���9L��Q�҇���f	�G_)A	�H�U��>^*r$SfM+/s�����}�F+<�|~NI�U5���Jc  T;%sꃴl����$T�ۆ�L��<��U�/��hg�T3<�������+����6�'?/C�<��� ��t`�b�\װ�� q;f�ُ'���Ғ�J�S�X�[���u^�����(L�&9j�,�´�b�vF.�]]��G?X��b�U_�POQ����?�p4��QB�L�M1�h��4�7ޟ���A��6�u�a��B�?֬��h�N��Ϟ%t�2�9�A#BN�`�j)��>$ ���@=l@�L�י�����б�D|f��~�����'�[��?��}�fQ�P"��5kC|��Xb�-Ԕ��[�	��hj�@{��l�bX���BBڿ��!�*�rl��j>[a�&0�����5����ti?��-O:�q��?�Rl���CAdP�6�Lv')�H1	���
���k�u�W	ήu�l�pU��3.8�06$���-�n��U��qy� �pE���Z��7XI��H�rԑ@���Q�	�mY7�"��l�ڸ��y�=�"܏{ؑ�"
�2�vK������ۑo�� ��TZ������y��MΙ��
D��!�>��M�Y�;ؼ|�A��� ��۔��ۅR�:�I58H,�����QH����n�xY�0�WB��9:.!�u����M��3Q�!�h׏�ߞ�o
���p)�8��i��Ӭ��5�Wc��ǎ�� �9S��]��Q�����9�u3���tiǔbU��}'�v�w��Y�t���ʊ��ћ�_��2��4�@�h�{���ݿeCH��vW
7~��g*o��^��H8�rI�ݬ����%�!`p�P>��Y�OJQL�,�o��K�#���\Ig��8��r0���=�xr'\[YH�#!���D�y6c)��S��y}��2m�]�RZ�����=V��N�\�(^h��振||3��bn��t/��f ��Lᔄ+�+�~��>o�u��q9��),��SB��&%cbfaw������U7T�$zH���8-j��xZC�������L1]'��'��J�
�F���ΛU��*W�>�[���u�К|tR�P�nSI��<R2�̿����s���� u�u���k|jV!k�/
*��P��R+��KH, V�%-�z��6x�76���{_�h+�)���C=��D��瓆��>264��;��d��[��\u�A��}��fĴ��cܾ2Ռ���Ѹ����
�
U�_ l�.�ڽ�s�?���A��%B
`�;D
Ϝҭ��H��x%﯆�uJ���N���v���w>��Q%�<��M�;���L�?�ᱪY��xo���}�MR_���".9/�w+M�bĊG?
{���&�6�U	3%Cx�F-d7�8fE/R�L:s��>t�2��6'�,e�ب�+��#�̻n�u��|����}�
UG��Q>�z������j�DZ�3N��%w�Ʊ�F4�g�:��/��g��p9�,Cm��ݛ;�ɦ�̯q�#�z!��ctlQ�kx� �b<z� � �T3�X֍Ue�)Kܷ0�.�i��{�Q��w��*x9�ܴ@I�4�՝���*�$�z�ȸְ�@��.�mnP�Q�Ȯ���-(�	��#w�LZ�+q�DU�y?�z��f��K�"��]�ԏ����>�r9�����U8��=�dc2���SZt�8_��� ����=�u���\�Oޛ��Ej����0�
=�/�Ut�/T/�,�G�k�R0�Ъ����������!ƒ|������|۟_�-�J`(�ZUTG�53��-�d�z�]�W4��j��<����u!�MK���gTTìf+S^E>wW�1� 
����>���G�� ��P�VV��̡T�Q�SF�R|1�Yp ����b�}�_&��^�������!��)�*��i�6�b{�dws�j�V��y��E��$�ԨCl}�+Vb�OAB!%-��W�
6����Ft�� �^S�4����Xxܼ����Nb+E��,j� lc��ui�p�o_���$jxö�J��5�}�{�}����q��̿�Ȭ�F��K+Jo�fs���6�?)���{��nfF���r
�Y��Ӹ�U��5$�V�aT4�*��n�HӁc��{H� r��A�s �_,����R�b�.�۽4B$�{�����M�7�Jj�Yl� �ђp��kieU��xw�D%�JI{�?A���<Yw��<�[�Yd_��[�����uTܝ��ɹ�Ӊ������lҚt�x��86��K���� }����)Y�m;�U{��C���z@I��xW��F
lN�d/b�i_�̉��Z�I�����%Α�w�/Y����Uk��oy��aGL�TOܰl��T�£EŔ(�m�W����Yy�&��ŋ�R3��.�'3�3/��e�LL�����(�R��c��k�7$9ݡ_H�]��%��ä2o��'��4%U��J��v�%��m�W��c"���6ȁ�GN���W�0X�w�FIߪ'��3'�'80 ]s�ƞYi�k*v����t+�K(�?�(�t��ֿ�w?&ͧݞ��������9�(���� :ޘ߫<z�]�勍�&���֭dTG0�b)��p��ɲ�Q `��FeX�����Sz�w�l��9&FP���t���l_*	��%��zV��!�,]��E�/��8]��tz��?� M�?�8X��)�9m���V�0o��z��a`Uܫ1�6���0Ņz]���=s;F��``ʝy��I��0S�������
��2��x��0�b65������C��w9[�19�_Y��":"����e�O�>�k���t��RK�Jw/�G׬�D�7g��%�5-�1��N|&�|J�3��%�f(S�ȱ�d���ܱ��H�%�ᴲ3��Z�9T�����? �v��Ll�Y���^h}V��*��W��q�T"�jZ�D0�$ȥ́�t���S .88��S��<t��=��&׼C�N��YNg�PG��X�2���$a�8�X�E؎���?xm��C9
O�p�@�7fX&{J�9G0���usL�D3ƀ�_k�b�em�c�\�ˢ/�X��ˈ�'<�Z���1�����/�Jy���&p*�����Ci�n�/����SOzI9� ���U	��24�������3s/-�N��RT���b�f�ֶ�P��vy;���bu1�C��L�^�UzE�h4��d�x�a\�I3�u7 %^V�/��'i�f�9��?���!e[Gn\��0d_����:�E0NU�c#��	�S����k�w���i=4	� !��I)�l���&�yZr&��I���)u�1��T���xeh�j#%]�4��9�؜�
I5�I�l�e5��4_�Rb��<����c��!S�a����Lw�_�2lH��<��Q���P�MR~n��L�P�~�o\���X������{%������Rr>�3~Z9r՚ѕ}��(?v�}lI�Y䅍N�#U!��hRSNL5A�����r6D���"Y��[XMU�I �Y�5{Q�N{T}Z��׃����5�?�	5L�#o���Ǉ��wf�v�I$�$XV��@�G���?:��ø�0gI[c�F��ϸ�ַm:yf݌f��i��n�i�2��EmΧ�n�K�t��9���3O��p��wM�p�B��A8z � Ե�aa9d�;iN���,�ؘkfs�m�rg�b/���c<���7أz�֯�#�0�k&���k������n��`]Cِte@VB�i��6\|�ߖ%_����!.pG~=�����r����������c{v�_�0������+[<���32���.���?��R�R//������k��q^��ℙ>��;J�ޭ����!L�O��55xQ}�c�ӛ,{jI<������@�n�v潥����D�e�O|��E�܏.�w�nG؋�P�O��E�[�Wx壕���U�H8���~5i�@���\K��ōm]j$���6��E�0I��7<��P��o�֭�c:$2@l�\���]�@o�l��M�V��H�D-��?�g�=�;��E�*��a��d	���( q4�E+�/*A��blC�J{�aa?x!K�����Q�l�p@�G���â�'}狉Amf�	N�$WM~?��^'����\��p*��E�cz8�U�C��|�n�OH|u:R�������j�]��UL�#����nowFJ��,�Q~�M�P���#ёk܀��4�cv�A���#^Ha���*�9��+�ݲ3z�^��n^vZp[�\����J���aP �D�^?��s���mp���jl��fMD�a�%9.kݸ!B�G���N=�b³�:�o�lwCh���2q�t�;GZH[���jS��:��H����oh1���|LIN�v������ ��d��WuP�כ��nŎ�[0~��־�s~��@�Z� W!�?�A-���^��a�&7�g�?3�7^��$[��X�i�2�Z��x@���!���d�λ,z���M��.�D��?�gb����1��sٚXN���܄N��0��	�#�.�A�%�`,��vU��k��32°�fa��+ ��ĎÇs\y�ct-�Vԙ���!�l�"(r i,�N���7Π��@���qe~UB��@1
9���ב������m��DB�n@�P ��� JB�k9�5C���y��h����>�ag$���+������hu ���:���EFkʲq��SI� N2��e%�놧�=d���\U�����z��I�7`m�����b�>�8��dF�nN�7~NW Δi���A���w�$G6����Чg8��K��n�l>�1`w_t�ں�1��A�
�|��H� �Y��p(�h/yG�F�� 8�-�$���[#�,0�>���T�*���o���||)D�B�zK�Dp��l���G.��?)�v���\�?�� �>S�&C Au������"+.�V�#X�{����T����U�y���T�)��|�;�Ag�3*�EU�jIN0,5�	��52䵝	�q�Z��3;/�����'4J
`NOI��F[��)���:�/�JHM*�lChp�m�:O_ӳ��,���7����T i-GF�+k�d	-OJ�y̖w[��ҔT�M�4	�P�����,)`�»���EX۩���E:
�G��	���'��p�D�����W�+���Dv��R�n뢂a��ψ@0�s-�N[g�˻f�$˳��؍sE�����$���j�1�]�&�k�E�Z�is3{ib�fuB>��|��R��#n�{����REW�A`t�7Ը#�g�V�e��S�4!V��9P�r.=Fp�2�k�}/4L,l��M^��J �"dd��*FX���[(H�i9��O~y�4��"�w��3[�ؕ����H@[��{T�WaJݰ��r�L�J�N�,L�N��V��&�+��I�̡��n�&����C�w�V%����r���([�GIxa�<�&X���n�(X_g��@��[�\.4���q�y��̥��/mo�I����[َ�,��.wc�z��Σ�\��'��_?k�C="�Iɏ3!�w�:�h��q�w@x`M)d��E<�W�໻�������
�8˿�"ū)ۓ��]7�5ܟL	&@��hiZ�C����#\J������g^�M&�4]��m�v�� �6y����e��>_����`��bK9�0�p�2���KM�c[�����%{��b���X��0*)T�9�ʯ�#;ChwO*4$U�K�Rz���t�q!&*Y&�|EB�79J^y��|$����5��3H@UNv���_�>@쎁Jk���:	d���%oG��]ߕ�|�YV��j�[5�O��+��4:�\P�aM+>�w�y��>���c]v�+����>ǺY:�4m�%Y	��i��9⍛�c=��F�����Ew��0S��#0�s�d�}���� ^Z� �j��#�`uU�����i��\m�1$v���"-��	e�hd )m�̾NT�k����|>���eX���L�@f��3شEN�`��h�� \Q����ej8��B[�8ߤ,�y���}��L|`Hm*��W,8����|
�j9�Ѱ+�Fh�۪��	-H�:Hu��"_�x���)�>�R�;8	�tb�X�� �$��$�U�xw]>+.(�I�1�=�b������29�Kv8�v~C���Bt���{���%�<��̍����\��,��#x�>�6��W<�� G��ݟ/�/'M��:�ᶙ!۩#�\���E)�s�Ԑ�n�+������v-V��� ����Mb����}��D�a��'|�Q�8m��HfI�p��*���XX �B�H��@����@C*R�H�b�#�	��� )��I���q��	�P�)�����:�4V�uW�~`}���q�q�+��z������Ǧ��������V{}z��� ^�e��!m�:.>X�����	Q�7�g��6X&Χ˟K���f�?��oR�t�Ż~f�f�z^�	s�ӫ�]��E���+���ԯE�v:���g��&4��������v��'�8yb�E)QP�8E�T�)��qr����g7n/`\e����UR�Ww�8�:GC�#�eu��{��[�>�'�g�w�=����ˌAp��h�U"���ƃ��9]A�h2E;T����q'[�n(ȢU�D�I�r�!3�V�.��m�[o��]����m��F2E5���&y�t�Үt�e�'�2c��o��g*F� d"$��q�W����~�g�x�ǵ3����C�V���m-��W�.2ڍ9!������³��u1v�c_��.��g+߷s��2w��¢}Q��=��mb1�nL)� �_]�T���k8.\X�-`��w­ez዁�c��;bZR��C�l��õ����y�P���d�s��%��~v�� �8�{鿢�%2���Hm[�ɐ�]��hR�B�G��g�~��?x$�|&%�R��ڽ�Ec[��^NJ�:�V��xv�-+Ƌۢ� �A{�WZ���;fݘ&f����g刏2
"�k]�q��eVݳUfX�;Y8�Ŋ�'�>w�2E6%�G*�*�)�l�Ş���ȜM3,w%�|md^�������V�q���3!Fr ,#־����x���>��"�T�֋��	����NI(��oe>B{w�=�6�C!%f
 u�4����U�5�\�^I6�ex�V�p�W�d݃�z�f�;�C.Z6Eڨ���G!���XF���di�q����pYکΠf�t��wd�^a�����W��XMaN������ �6#j�FQ�/Iۑ�D�Ҁ=��ˌ\y�����yq�����۠�zK�+G�S��1���m�q���j���0C�B�(�?{�{����Z��GWvvGO�"�o,��5�(��}B���y0_.��Ål�Ɛ#��q��V�M6IW0��.�@Z{�9T�r=�<ꣃ�ODLA�L+t�y�7G��'�3w��t�!:MSD�_�b��.t�c��P���.o��a(�
ʠ�a�kBYV|�r�����z�H]���X�f�^&����&��AK�נ~��f��G#!�}�����e�5���g�E}�q%��ULW�����̳4���:M�Ւ�s�"9�U�B�4�w��f�l1�|�t@�C��d�2x��9�fM�_.?�I�(`dI�f7