��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv {d��ށW�\���k�(8Ȍ_"D� ��x��k!��E�$��Ho5h.ԋ�Tt�"z�	�˃ ����2a�)������C���V$��#�`�R�V��"y͆����;�3��e߫�3���Oz�|3i(��=��l�H�5��5�Y�Bi��@�\Pδ錼Mst�F#K-y�`��i{��o�HkZ��?�#ŒW.�[9��	�7N~�c�­.�b������u��L(N�	�� 2����<oc��(��7����Tc����M�QA��KT��'�i�a���)@b�yΘH�eY-؈6ךv.�L�?��$��k�d���zz��9�N��V�U��#�C���p��{B����P��ֲ�
#����r"?&O��v�ԟj��$<iA�V�3X�Y�p�}^��٩��#�Iezx�VB{��*v��#OB�`�Į0#dYbI�����8F5�	�nF;L��1�U|�ʪN�k�s��]ޤw��u��u�2�J�T���1�vఝ�>�<l�����_� ���?w�Y�i���c�IR �Ä|�~�?1�$`�
 0bx���GFeG�hBI�Ot�j�P��������|)��I��o�s�jb�X=�aL�|U&��\�7Uʜ�<�l�ǆq�V������ΡC94"��Pm�.j�>��X56	���{\A��jh
m�A< �[�9tf�{�du�	Q��� G�|�A$�I�*��GB��)���a�U���9�.��M���]�(L �_�yO(d՝�۰YW��E;o'�`�7	;-<t�0{�7'z�l�>��k�ԑϱ��(�{Ďa=h�_�P�ѳ��^��l(��Ĳ��8�76�ľ�:..���d��K�E�Ъ�ѱ��ꄓˎ����,��ԥk��Ba߇h�`!|��wYz���v&?1�B]o2���߶�.m6G�H�Z%k8�'����H�8��N�C)"���w�f�����H������8�[�����c�;K��6ǥY5�G����lE޴�SP�4�9�����R`��JrMfp�ITL���l��E��M)�mpJ;���2b�n�,i�y��P���~�lB ���=����.�Y^�X�s���)��}j�������.�"��s"������!��PNH��(w����B��a+(�?����"'�BCB��.K���=��)�JC�	���W��~��H�C|�+L���x<BZn���D��Y52�]m�����N�H/J�ٚ����	 ��H����R�O]�
��c��lX��]��4)f�p�1�<���(��D-� c�29&<��%
*�g�������i���G8g��אPO<����ҍ��-.+����%����=6��Cw���TEC�lx�����L"��}�4�߆��X E�Ukq^ط�6"��p��M�#����*l��9�'.43�h��'���ժ���4R7imH�B��NA��|�=��[ƌ��W��[7�f!�ÌUv�As*CG̑�7;m巩��n�m���.�%4+ګL��)t�A#<$�����c�E~�q�x�4�����"<+5ec�U�E��NԳq���k��f��݀Z�"�%�|���m�/�H�<�6�M�9�쩅��$y,�*�4�s�("T�ɺI�Y�J#�#����>h{�XҸ�����d����/� ����}� t���	|iB(�����%w'(3�� ƴ'�� d���ʜN,V,��1ڿ
�;�a��l��}Πz�aS��ЛA���Y%�V`w�,MWU�Eb����1=�oɢ]�y�&������N�f�gU[X��\�\I�~��A��(�gTx���r��˦T1���YW���p=B��8T�qمJf�G*���*��l�5�s�L9�tq	�@xu�"�#���i�����*_��ӱ	��#�b�����D�c_�_  <�]R%�˝|�A�Dյh͢�X��� �iC u�9֕�z����q�a�4��&	y��SD�20�391�m �fu��U�s>4]��:�������\�ȭ�]�c�o�Ŗf`}�)F�����B9c�a������x�a$�=@�N��4A���QQL�G�e�bs���1мg �7��$��S)�+�G'AВS�D(���3�8��(���1ȷy5�5	���q��mv�fTM��q�Y��M��U:}5N�}��������XivS�v-��z+�?K]�:A�oH��X<\lG�K���n����&#���c2h``���a����/4���o�6d��]	=-�i�]��M������U��c*���pf�&`.����<�C��ԟ�����@��e�O0�RX��#��nT3�����~p�t��7��6q����V�P���ؕ`kҠ�XB���m�}o^2T���3�!��������%�wr��d��g`�Xo�U|��-;�Y1	��j��|#��խ���oo�3�E/ /h�5��z~n�#��$�x�톐n�`��2}$�{d��J�X?E(����qdG�`�&����"I��
�u�R������q��'�(�v����)�m���y�	s�� W�� �F�؈�q6�7��6��n� ��v&Q&��ąp���j#ӌjo�+	�W[-�85�r��.���jHH[�Vt>L���F��k�6ăp.���s��]��<���%J�Ɍ-�7�!aĝ�����vq�<@'��l���,x�5�:L@M0�/�Q�5N��`}l!n��D^� Z��K�oQ\�iK!���@Z�6�m��	�s׭����$ul�½��I���Q��|`��Nh��X��/7bG�����iC&\�  ϨB�̈կ�ϣm$�" �u�z�B0�?(�5([���1q1�wVU�)�յ��클���z�[�"�y�m�Iº�}���O��i3���Y�ZL�F��~��n�͙<�'�#+}���6�?�;�ޱY���wF�U[UjEl�W�)6�V��Ƙ������@�Fy ���aC�'Vx�+̠Ļ;G�Gw�F�~�����_i�2�}&7�B��>yp7�_=Z��Z�*r��၎��S����\S�ߕ��I�nPu	��R
tVt}��jM��b�Z�W8z�t{y�%,��G����P�ǅ�<,d��qm����)���ޥ��d��Y�$�TȬ`��hTod(����P�}�����yq��'��(�0KZWNYJ.�t�@g}!�Ԛ����LT0��K�m�D�^�v.;'z#Pu�U�*{G(6_:�z��I'F'�"�1Bl����"�*�yQdwKBs�^.�c���'\3�oM��d�}�ўl�}y�=���9G�X���_d�'1�/�C�a+-M�iF��<Վ��}2�@�<�%�<��̇�d�����
�@t޻�;(�3ǡ�k-Y�JG]�{#���X��`e5�Գ��njx�sm��j���tY��)�@!i��A�\�ot���kv>ۺ�.ړ�.ɽ�ri���a��D�T(>�+�`a^!ė�8�b��Uk���1�1���c�(U=Y=ߋ�X��ۣ�|�C����-�@�̊�U�#�E���'���*���G�BM��'	YfC�F��(�Q���z��FJőK�~���3��I��7S�3�h��ruH�8�:Zw���[�u%_#���N���k>�ZUwvl�:��f���n��w�mR��kk����0�%��{U����\茯���R�F�d��%M}�i�v,9��V��T������y�<ι��C�=a�H�� ��F� =�Z ��o1����:�j���}!�s�z���ۡ�Àd� �7�Î�z!�IK�e5�d �1Y)�X3�U�vӔs�AG]���~�*R��d>;���������.^i6�HY?9����8���*-�د��G�O�1�/W���d�
�L��}���#����r ^��NԴ粼����s�?�Z̀�t!|lz_l�x`�8�C^�nE+�|A_!A��HI�&�o�g��f�s�P���;��U�2 W?��/�A U���j~�BY[l^�`)�q�sD�=+�<�vΫ�q{G�c����w�5y���mi8϶�CH�c��4��37�@���$��]D۾���^Lz���n��2wɿ%�^y��K&��柀O$��d��kA��'�����S�}{_]/ o�_
ސp♚4D$ZU����ݰ��͵ގ�{��5��� �CD�Ղ���-74ȭ:L˛Y.p�S/N�Ts#)���D��O5��gwxa��>��W*�-g���w� �=�kb��C�6��9�qk��S��6؊�e�x�*�F�䜅�.]�#�jLI�#Ԅ�}�Ur�k�Fx���88Y4��pw�@}=��\�y�D�h�୆�x�� `��q�3'3NF��<����i�6Csv��lT,�'g�-��:L�,�R�~y	�Z���wyL^A�I���� 'f����#��4���HRC��v��Wغd9��,+�*?�?�4\��[���W������Q}[|�Vl��t�f	dq
����/��=��>�@Ɔ!=+�5�������e�
�͔�C⷟��
q�Im��@����qGB�~n�,6�O��%k9� �;�@u���@J�(��(�x�.�4���}*�;��^��I��q��T��i����Iȉ�u�� ��;%N�a�hS�#;�y�!�-��+W�)g�o�8N姷:������s�f��)�����+8k�ڼ�����i��߼c�[M����L]�ms�.W{�?6����Ʒ�1��TJ�/�^��ÁB*֭�O��]�:�۟�nry�H�=%j)K�,��t��������r?�3�`$(ѐ��?@�#�}ʰ���?Rn܀ZR�l���D	ܡIp��i��Q`���D}������{uU%_�p���q��#�8��Z�:�)CG�:pёt���U�@Z�g��t�;o�
�h#d_����1��|$�U�@�>���u�ۉ��Y���륎wSv'�H��8�-����S�l�X�ti�梤M:�)��p)�����dP3[d���-�n`��:���~�N��M��'�QKaGf���z�Q���C�9�v�?�>˓�Eز�]Ջ��?�<��&.���s�8ͬ$jF�Ɇ��%����ͪ�g%�2��!X��D Wey��[s!w�h5���aJ���bm�#���Ҏ̻��.p�gi�n���bl��ؽ{5�Ц;��3b���\��}�9~� E���8�.�y�[�q澪���7&��kA���=�� ��t晳1SѬ�k�5�l�z$썗�߶E�"V0�\���,I|�w�j0��M=�a���l͋.4��J�7�����p��Ĝ��dl!�{�����B�m�u`�cɽ�� � �?_��A�2柣f�Ĭ�^����U+��PěD��y0��7j��E�p+?!���j���!\P�ts}�ц}mđ��e�"�Q��:/���6�a$����31�=�ݣ� ��ᵁ3\A[=�L�!��+6��k�B<�N2�?�7�_��%��"f����I�w0,KO��~(��)�F��+�St0�\8U�n����OQ�Y��yχM&	�闒UQ�N!��^wcz ��C��iV�����r�C�E��D�U��w&5���4�'�R�ĳo	��*��]D�Ty��k�`t�j�iÂ̱��<��aZm���CW���4�r�潠��q�Ʒ�f�>ѭ���(&8P�W���3�$5q�컏Xd���O������1��v����7� �{�� ����`�fH�z��1[E�����lO��Ɓ�!�IapY���̴�*�ytv��Z1��|R3���5+�S-��� �����[hP�����,�E��9��I�tp��pd���1�pj��b>p�6��E�z�C�����2�͌����জ�����y�8��M�kW��id�~>b�}X�Z�7gG���7H�ie��o��_[)}� ��hЄ�x]��w�+�.���=�ޘ���m�U�����(F��8��}*"��\W�S�m�ڔ̔\� �ʙ#�{������Y2#!j]3�K��`렗U���~��\-l�	�@@��+e����\ ��vS>�/�1�J�J,<�IL+\]��>�]eI����Fm���QOoE��9[(^��ӹ��-�x��J(�#���g��c���I�Q2�r.{e4�e8�>a~�>�Fa�}�CE�9�D���QRn�Y��%�'���`�:#u)a�Q�����< �9$s\��,O%G�4)&��`�q�\���ߠ�G��"t���
p�g���kX�s~�{%�n&���V�����'�VqF2�e�[Z/+�!���'�އ@��]���c�Mz�w���EJ�ꖲ�?�2�fX�,����e���w ��!C吣v���R�{��Ʋ@%�.���	[�R��]�l��di�ZjĈ!��'.]�!��.!Xf>�c����#
���!��O�K�����2�]F�X�0�─w��
��0����US�lY�$�����j�T3�jQ�g3aż:d@������z�s�a�3Y����]k����P@Wh���7��DZv����>oڮ�Z_?~:�7�2+��t��u��[4>������x�7`U�K�yL���G������;���-toUK����Kㄞu��\Z��p�!��ĘN�u�6omc?;�����P�<�G����كt�g\�����t[����7�.���`�����������ڶ�<�4����QҶ�!~·O1�����]��tz�����0��RaĉA&����9�b%���yI���v�\����G,/�L.�8l=P���I�O����� ��;$����%���Wu�bVr��B\��2[ņ��T)��<���@����y��
VY����� �PYw���W8���Px��k(�<|�.x%��<�j��p='�e�A$��F[�d�R����.�P���np$P
K�, 5�Z�����6��z�M@���kꡝA��`�>��Ewԏ䝨Vyӷ/*E��n��}}U�~�?M8q����p+P��[�c��ɶ��l�����B�&2���d�7KE�+i�$#=� :U�]Z�qcjP��E��9��*�Yy&��6,F�2�1h���<�O@c�} �e���^<�~RK3��0֚�Y���-�`z~x�&�!����9.�;���7��yfh3#��/�B�F֚��I�l�
T;<uW�?k�I2�t���ʻy�_�����i��C~&��I���.8��@��	?4
}�|��~���.���Ot�э����%�+ q����Z{(k���x�Ym�,��{&����6]�-���y �}<�+�G�4|	Z;r1��摇
���I�h����5�epB[ܠ�]�إ8yc�cul�h��pXH��7�a [%��A�W���W�?�ژ����d7�|���6[�'fBI��p8�(��:���LG���i��$�m�"!�ee}���N�"�0$Ǆ2����<���R�CEE��	��D�';����/�*����\�rNM�W���=�8ga1�B����m`��[�,��C��b��a�-:u����77��B a�G��[-�(q�'ň��EdR�������li����G�X��	�CН��`-M�-��f�ira�tp��jup^dՙ� Re���e4}�����>!���is
 E����N�k�f���B���}}�p�[��	;u�1z1i����d���r"�S�Y!욜K���x>㧐5|�̱�@(�,�p��m��f�K~�}f�B^�X}>F����(�\�dʊ�2�E8#I�-��Q��U9��J��}f�B�h-�OT��]\�5� q��!��˝�[Cw(�,lH��5���[+[��D��vEM�/�w��"���\�ڑTˈ���ԡ$#���VaU^M� Ԕ�n)��?��dg���?C6�j���t�jXv?,��E�����
���5��.tԥ�X�MU����;o��p�ݠd�?�/q5oI�)=k�萆m���J�`�e����NL�6��j�B�{k���}5��S��2��[���#�.G�����ZP�Ɉ�s��@L˺��*���=K�RV�fBq���%3b�L���1��Jy7�Z����P���3��eN8��0_��<��e�����W����+0BШ�����Ϥz������Su���"��e�L}Ns��~"E����/�	%��Q�\�ꋝX;��6z��2b����K��(E@e@�E�dt����)����:W�#�����}19&ō��9Ա�1��/��;c]��=����!�`�Fٯ�L�1S�/�_�z��y����e4���d�3� _�z�T����@כӏ�23m����I�w:�тwcHO��Jn�q���,,_h��D�lԾE�tT�ݓa����y��c2h�B�������ZJ;<|�����MТG5Ma�dE L��M��8*k�k�rU8�K(�?��x��2M݂���
P�ia�b�]��ǥ�UUF����Q�=�~db�i<q�P��]jÕ@�1������k!J��(d-��苂(�E<Kȑc\͖Rw������;�#q�j����\T���T��R�qR>.6��xj,B���D�� �:@q��i��^�}V�^�6a��rp�y]�;�N�S9L�VUMJ]"��E�l�L�'�ɘ|N�7OF�澵�n!��T�;H�R�:fy	JM
�2N��>�22s���|������<ͷ`��JW<�K�;1p��>�t�ζh��.?�ҧ�sT�w>d��?h$⃘~C����ե.*�xps޼�f���-��%d}_[A�=��Rgѩ�2��2<���E����o�6c�����ұW}x��3�v��5��g]��&f���T�<:�A"d���0�89�k;���@�H^�\/T{��͕��[x��Y/]�;�U.�5��f�h�g���-&?;?��s��f���gN5��i�1R�dq]�"[>�K���Z�91��;w�}�5�\�z�6���	r�I)�$�R��Df�ʬ�n4A������c�~���c��ȑF �FrvII��7=L��t�@*d<qU��o�X�+�'h�ޘ2��C��V��@U2�VkW��h9V����X��.fO�]�;p7���B�e	,|��Z0D�N����N�P�,�]��vi�Ç�{��h�h�*��C��/a��.g����Y���䶊�<U�s�_��Ʉ���[��_��p�Dv����5�tW�f�¸���9k���/(��93�a���Ю��4��FG�Y>�@�*}��[�3<��U]�R]��CG�4��q��<����[Tg#$��45��Ҏ6�p���T�������������BT��q~|(9��|J'z	��Z�m�ðN2���Nt��/�> k��-�L���Բ��ﷴU���7��Y�I�=�{�}'1\1`Rx�4 ��nu��O��a�Q���r�H1@QGV�k�sҾ�ϳA[��	>MKq4��3���������-��&(	|F+M0/$�]��1�"v�)�A�L�?��}z���%���u~�>��{����u�����dy�:(c%:*hu�z4z/~�b��
�7W�\0����!��$�YJ>�{�?U�O��C�`I����ٕU�wA�t7��$�Yc%�	����v�?I.aja�Yq3�Vo�⛝��}�vO�����UR.1����u��,��C;^�BP�g)��g��vlV���N98\�C����?��
��9��FzL��C���j�
�ut� "����ux����x7e���_��۩�����ݹ �
1�2�VU�4��hKz�(+�a���0���`�˟y���k,��ޡ��9|A����$-�B�@E� ���XR���,ʠy��!�y��ᗟ�u U`��(�Q�ʼy�"����'ե�#Q��!u�4��`���-��MC�{�!�$ѩ(q�m�?#s���f��Q�K�z�v���h��[�@�7��
��IH'���� ���Ur���A��g^v�0\�mOJ�	jA��|�h]���l�%3��� ;��U@UY�X%�����O�e��#N!��;�s��6˅�|aXč�B��l:)^����P/��$�{
�M��WD���o�h�AO�����h;�p�j=���!�<�-l�&?K�I`�ckQ��ʓ�%���,�D�~C��w�uPӟJB�0j����v����>���Z�&��Vϵ��v����z��j�ǒ;[�Iy��b��$������oIƂ�3"㯮b���a�+��%S���>�>}^a�X�F������u?n���Y���HE��@���� ÜU�"���spS���W�� CdC܄USuq��iw����yo�&�B�ԉ$�1���k)��^zĩ�{�Dz��o|+��p�V�����C�S�@ٌ�u]bk4�j^�BT;h;$��t0�ɨ�I��/܃.N&�����O܅�Ţ��#�u8����C���W�^F��kr\	;�UA\�ƊM�1:Jg�<�C���`6`;>��Z�-q��U�"��r���7^a[��K�3Ā׫���D�M�_������ad8f�<�h@���}�������DxO��A/��0�i�W����{�8HC�g@�P��� �cB��t�#��w�̧�|�� ��-ib�CTx�x�Ձ[P� ��/ޯ(:�؀�^X$�R��[_,Dԕ�� -"�*�g�:���w3q��3����P���:޲�1��7�b<�c�}l��������I�t�$��Pw��7�>�,��45�
9`'�):2Ř��_��,��[<�0��6]���R�n�N�������g:���x���t�6Vk�Tݛ�'a�j���E(�UT�Y����Zƣ��T?�#b��:˞���2b�%�L����K}sxT�&p镕��������Q������&E�]�{� ^��~긔�g����zjs���-�rk��j)s?OLA�ь�/F"6�T�<MK)z��ny�=���A��t���ønN��lq-���|E�E��+K��2�.�>�`���5�D��:^��[����Bh�Mpq�.���c�(3�x"���C���	g()��Ǭ[�;�����<���Ȫ}��/c=%���7��i���kPw<B�z)�?���":�S���O�ɖ��G�b���"� ��"��`��X��Ku��m�yz�r\z9�)/ .t��R�.��ζ�pժQ4y��eē)98�;�U�̣V ��ZK!���\�Գ��]�/�Z8
��r���A�M]m��O󐫢T�9-|�L��t��d5˪(B<�R�7#�?�/���P�`x9*�
8�ejԳ;!v���s8AS0t��
��9���RA������SQ� ��(80����c%mg2���q�U�2s�K�ĻQ��ߠ��j�g��] ����2�P���-zn3��b3�f���/v�)3��J!��R�!���/�`d֩��21\�`��$�XR�7@���0Z�$/�^D��qt�oO6���G�8ʑ�� ����`�^�0xKQ �Ikv�b6����� r�㽘��Ҭ'�7;�jڇQ��13���,�e6���ؖ�0���ָi���l8Bx�,Uc{Ј�A���mqU7���M�#�p���kй�Ѩ�Y3>�a	��l�O�������!�n�9d$�a'o{`"��kN,~���Ƚ�֨�ik.���U��~ǋT����d2���n�����}?�(7QK��_gO����ט���5B@�/. 8�Qu�S�5R> 9�M�o7�b4�G^�w,��u�j仃q"9E����s2ҡĢ�>�C;=,�Gb֝��p�Gz/�2��d�tzԡ����ǫ]{����ϫ@�2q���5F��V�|��/(��Cנis��1nb�B��Zg�	kQ���v�C�5�x�d4�G�����0���o)��+P��D�Q	D𪢻�)�2&�`��\���)�|�[Ux�����~��y��)�0v�κ���0�lG���r{{�L�W�O�6��W�!��Յ$<�P[g�J�~���#o���s��@���\����z�����Zc{�_���Xrw8��*����
�Q�����!���pj�e-�]c�ytB��66���a4\��h�\���}@:��� ��2j�A�)��Y�<��(��y�?�l���Sg5�8�6Q��IIi�!�^�#3��Ô�-V�\8���	 ^�jֻ3��~���R^�C�<�\��܏�lm%}�P2L�X�,'���g��eKL�Ch7�6M[���^?I��BY=/�6��<���\�]��F\����V�.���ID��7e����cT`d!�G���?b�:0�f�&��������i�k�����wZ���PMLV۴��4X�������P,�|��۞z�\ȁ�'�1�Є:<6y�$)'pz;�����_G��q0�F�R4Zx�d �6�42y�T�����cW�|e&$<Y�n�h�7'u]W���Q�TՍ.2�	E��7�� .�ւ�V\�ޥK�`{��5��ԫ72�١B�8�����K��):'�a	�������p���v&{-8�ou���0��]k�>��C}kMs����7����.��b����~�^�0ʄ,Py7V��Z���=JQz�A�̠1`�ޕj���;�a�$hU���L^�gW��'�d�I������Q"5٪����7/�y9�I��b��P�;��l�3d¨$kw�A��|rD�HQ�x��5ʱ7��1#G^|.i��
����o�Co��j�pK����l~Bl�ֲ�^�J�z�#,�8B(����nX�_+S��M��^��Q?����@]q�ї�Wܭ(Z�����k�3�8˯�E!�!j���ЀR�01��צ�4�$zpC��@R��F%@��K.u�W��An���w�*��SKҧ��$)|.�b�w<�-4N��կ;#�컼y�����ߏ���[�Sڃ�G=egKZ«��a�l��5}#�wu��5r��p�lwP��Ԅl1i�|�^�N�a�=�d�;eh:�]V΃��zɍy�/�f��,���^G�3���@�Fj�,:�I8y^(C�W��.�}��3�Xf4v 3���|(��0�&�
ݔ��h��~jʋm� ��w��0M#��S��nVi�C�ȩ:_%��\��6�J�v�G���SOOÝP�U�9_������ �9��=8�Ql@�S�%�.;��\w��w�*,�</		�y�q,��}As)p���h�*���V����_�P�W)HQ-�.X���s�eY(����!������H�Q|�M���52D�"}8�B�R+:�������y�@�rM}�Qϧ[��\�u�T\j��!��X�MG��gu8ss-F.*ʂ���Mxs�C��ƁOh���	"���U6��^丹�\Z�q���</�Zwȸ�n�\�D���ly�U��|+Y��w������.g��4���+V��e� *ˍd���Ņx�"a[[ua�jYxɴBlç����� �C�8�k��J<:�\U�4pP��S㜃��:�&�g}�[�
�� Nހ,n��E��+���������m��h*Ac�,���d���I��%!�Lž8פ���Ja��X[�&�	��<���vxƿ�=%EֻC�'��:j1=Gu��=����d)ug�b̉x)�L��Z�~�r<�-��m�R�����72n�Da���N�>{Ъ�����R�.G�On��S@qjp�:
�H�v�}�T7�B�~������G�tG�;Y$P.�+�=�a���+��R�ޡ�B��a���q钱c���t�Y|����>I�k��X�����E�V:��9���W��֣�U���1aB����;��ys{�m���4�~��n��X������82���a��xL�vh��G���~��az�S�3������"DO�&f�j�\��0�JP{ۡ����)t��EZ�'���@BS��i��2��)��͛�{h��W^{�>�G�9%�X8�5�E(ς'b(z!oD�G��1O>��R{�N~Z۰t�]U
��X��=���s֌L��&�V�w�M�B�{"Cuy2����֋���#KO��F�*۠��|���IV=m�j,�j�-`����+vI�i�¼�)LB��7-�5B�t��g�6��<n�C�%40�4]��y���7D
��«:L�|��U�jA���2��L*c+ ~��#]~d��pik��s�m�����l�M$LY�Wvq�7��i����&W>v�|�ƾ�K��H3�V��c��-�`;��H8���FM��Y�� ��y�gR��T�aו{�:o�����WǖQn::��4�"4�^>?����J`��T��_{�A�	"?������R�n��%a~f�����ȃ.����d=�v�c��QKb��`��@581�S~�cDK3;�7vi%9�P�I"��[�Ȍ�F$br��%F�?@��uj�+g	V�P�`���d_ɌU�z\�<�;��g��4���@�������a<��@.[]T
~2�FVQS�g�a^��
�C�Y�z���+�,���v�	�$Κ�� u���0.� �Q��]J����~ͷ$&�}��z�[;;�G7�c�W�k�Ȅ՛�V�!fo��tD�)$���bw�����;Xۄ���]Y�g�n ��c|0n~0�KH:�0è��i�Uo8�2��R�N@�wJ�H����6��rPPX#�Bqj�\����E�:�+��]����'���$±;��N��F��o�f�1p2��To,���0z��ڰ�`.L�B�9�
�+��ߞ@֝�jz��P�֒�l��
�� �a��E�������e���P�q�����	�3��u�E����.��mh[�s�e�}DS�l4=�hN������!��sWM˃��`�'ǅ�_�GqI�%��#:��Y�e9�p�j�m�P5GjH����V�9��E��C��;1�"��h=�8,�=6��K�x�t5b���`	��Wɤ �2�����?��F͊��Z��+�դ�So��+��K���N�e*3��=�<c:KE�̮
�g�sd� Xm`�t�x㿃N<X�xIa�7����iB�Ȇ9��~����ʅУ�݉�:��D��?���uͪ�u�-��~Ry۰?�:K@�(1O��Z��ꀼ|^�l���\��Ģ�e�{��OR��rI"�G,w��nd�\�B�^�?���3��k!.�U��i�P�Y��#��Uo�B�xb͐�]܅oh5+^�إ˧�U�8J��g�?�ݤ�XD9/[�����#�xkZ��8l�2�
�8i�������m�Й�#�]�K��t?R��ɔe�q.R�~Q� \_/�u��SU)Ggw����LD�`��~o�`1Dk�{����p�[in�7�7���u�x����젫�������o�s*A��TKK��D.5�é�¶cFsb\��;E��X�����M��|F��g���_�Dd�|�D�Z�[=8�9�
��kڛ{�?\ ���Mb�J晻I��q.��q�4a����?�hȵ�ҵ��}äY�G�5� ��T����hףO߱��ք��!-j�\�eo�96el|����D��5�#���X�d����ǙϷ��&v l���Ш���Y7"6�)?��ĝ��9.��B1� 0��&��J*�s��kn�^]��=���;�l>ԁ�|K���I_�ްK?��&��AAo9)�6!��*��SW{C���w�C\I�C��W�j��s���r���<r����咋t��[}v�>	�**!�"���X������t�05�.G��Ta'ߒ�*0Zo:�<BW*N�$�즩8�'�y+q���+��xH��b��0�x�������z������5�Л�? ��][��o�PI��	�&bj�Q6"5p�]h�:쐔��ѥ�*�H�?T6�]�k��M�*����u�*i�s��,%�VٻDt�\Ŕ~&VF>_;K��=�i�� 6ɿ#�����=���3�H��$(ȾB�z7��Q��D��=	�.RI~P
�>c�0b|��7�8N��6��8��o#�V��F�)V�P�E�̍��ɒ(O���<��z�e�7YcX��]���t:�r׋��k����B��
&��8�;���.��Hn�]����D�o7�-�5X��y����2��FR�E�$��2[\5jΤ���a-ŜP�#��5'�%G�X�\�*KBf0���W1W���L�Nf�	���ЎY�O\��=T�m���c��?�"{ܾ#��t\����d�8��r�y���w�7�T�aDA�=�)�N��>�:�`tJG,��L�t@��~�$_f���1M���ǥ�F���c:���;������Bv]���Rk�8�~o:,�׺� 
���8�����EfWB�f���k���jF�=K�/~���ꁭ������(ĭxu��2e{l��r�꧅qѻ��Y�Ɩ�n0����}���3J�6|��S�w�-�?'iI	��4ң�9[��e(�_u%�����Gβ'��Vo�V���	G����U����X�4cŒ1�CD�X8_^��N�Ok�m'���,�Q�ǖ��W�5m�h�P�j�B��]nIUH7$���w澹��%Њ�6?��ةB:���Q����t�������"���da�D��$¹��݇/�kAE���Bd?D毙�`�����y�h��dA�����u�L�I��]���|�HP\�w:�J�pe�p��i�� �v�4rJ�����@h�-��PA=���� {���I��S~����'��yd�J�u��I�a�-ް��Hr<�\����Nc��ZJ4���D}��)ҚE�D�i��M$K
��C�H�y�f
����l����(.�o���§v�, ���:�,Ԙ��aKou�b9�G�מ��:!}��"dtk��Z@�X�J�LcZ&��A޽�J�"�
�D9������VXp�ꁼfl�.�'���2/�l��@^X�XŠ��Jj-4K&���]\%�`�v��(�����̩T`0ٽ��~*��Q㩫��j�n��Rs�U��
`CV��6��E � �LR�.A}���ƈh��$���7��r���gN"�3e�ĕ�jɈmo���g]K��C�U��:8v"�d/b��&��v���D�G�b�Aim`9�{��I|�ᜮ� �]�'&�	��q4g��'Ҥ��_H#W�[��#�g�)��S���ksV]�㕞�N�F9�?'CI ��c<q������h��W#�^����$:�7^Z�v;q��h`:�N��Rn�z�����rΡ�Qn�R�g#/��|����Q���F��Y��t�Y�i����M@�N(h���º/t�d����3m�Nm�$�:�E_�/.��`��J��uK���f,�E���.����DpM��z�~?��$��g�0���0�.��/�	��/^��]1͑�M�>'q�����د�K��AT�c�8`t���n��/5�'���} {C�Ɩň//���,S���@J+$Um̓���H��L^H��V����4[��{�,�T����4n�=:�o�ɭ��94f�BQ��r�28�Hh��2�,Amz&>��*�>o�u͡1-r����1 �c�Cr*d���2L��`�=/�4���ߴ6���(�8��6;X�VT. ��:�~G�)��&�?�b��S}ݛ՛SX׉l��Y��v�u����eV"��n �s��3uB���g����0�t�#F���"EU���+�y���c���{���y{@��;�Y��խ���Ū�DƎ�E�(nh�T�R��
y=E����s�O�����[�t%S�`�����
������zS['��W*l3�Q v�|ΐ��<�@5J������w~�eq�U���myd��-��?�h����E�4����+m���a��]�d3F&���u ���I���p-����Gb[oE{�HC�&r*�2ΰ��o�|s�mIO4�K/��V�2D6���.��X����(��a�}��彼��Tl�D9V�� �,��u�Q��p��/�͆ Bﱔ�Gq
/W���Nƀ���驔�6Ō��AVe'���6�bH�?aX��C �q��%����]>i�f��|�MY.{sņ�]��w�X����Cr�s�r���󣴯ň�/�]g��Y��ׅNmrF�?�S5�]Cܐ���P�D����'tT��!�1^_�a�ȑ�����~��SwH�}vW�`'��2x`����I�h�?zn�������1k+�0�Jt9��s[g��Ɔ܏8e�"��,�y���W��k����f'��z�h��p�����p���oiJ�rM�b�]K�0��k�ĎRB�!Gd���|�+6�5�Dů����"��V��F�7��$���؂���i�첚����s��Y��G7���af�����ۗ��,�+_�诤�
�y:W
6g�|�qS]����/}�q�3P�1@^P6�k	4�&�\���'�����J͞�~�F�ϔv�f��o	�fE��iї����R�D�~
?�8���9��<��9�İ�'	�B�V���b�zX���Xd���g}%ԃ�AzΔGȗ�/���g�bm$�z�(�<�z�y͸m�+zqC�G�`{k���j�|=K
� &�ݨJ}K�)0�఍�H9�F��L�^���I��q[b�~ +�
;�M���p���X�b�h[���fb�#��м?+�,�ʃ5)/Y�0֓�� Z��7rׇ�i�P�P`P;H�vʖ�Ҙ-}�6#�����+���O�9�2��Q8�����G�z⚙E٭lsE��5�bA�%d��J����W�37�P5�O>4�.4Q-�3`��|�Qg����V�����S�$0�-�`j�e1zs"��!�w�I�թ{�e�0r���.�n����%*+p�_s���#���X�*V��%S�7ôU�+h8<��1�U����*���n�MHZՊO7H��0���x��?�c��e:���]g#��`�o���$ܜ9�>���.��$�a6�I�ͣ��*���),ó�m&��2���ґ�`*��6��qz7P�O�(����-kܺ�'#�	1�Z�8;�gJ{8��BD��~���\��W�`:y�`VR$��p�҆���סZ����7���|���4_\��ʣ��V4���$�L�B�p�@}��n�\���$�&&a�є7雞?:m�2�2�A����@e�14W��x����zjE���f�#�%:a�
`�8j�Z?b��byKx�ڔ�+�/H<�'��*u�Z1�]��Ľ��{GBW*�����(�Җ#�*mTH
s�l��x�Y |m�����YoO"�c�k60W��01���fi3h��ҝɻH���sy�g�������"�U�=:�t�.~�q ^e���s��@S��Z��{/��S�+��Ϛ}�S<]��Q�Ę���������$�9��U��Y�FϷF�&�S��Хu�#�N��>�9T�}��������1v�U&�A$�
��2|Ή��?Q���_��5pN,�[i�=�(�7�j�/��<Mɍ~rYP�r�|B��^���d����v���绱>Ҏ�7bM��2��gU�%d�6�:mHB:S=�g�,�����.8�+�5V(7O��s[���>�$���x���q�s���D]8s.�e��n�,�O5�"�ː�r��´�2�>�sQ�q˂��R�e_�����A)����4���F]|fO�� �L�yb�4~YGdm'"+��M��%��a\<��\���kjI���u�zd g�^�Y�Y(?Tٸ@�J�ޑ�fS�2'J�����1����!�\��yL棅�P6�a@���#�H^�=��B�g�뚞6���<n��t�kuMufg��,'
k�T����ٔjyM�+����[� ��h( L��k�Drk�N���W������(����h&�4�ნ�l�
�ab�_"�f�#p��">�kp����x�]�0�h�̴��3��V%�i�bY�t	Hee8st�Q{��2�*9�������F��b;�z
y�}���9('*�W�Z����������n������/��g���h-�(�7+xxcAUi�it�le~�'|�<��UT_U3+<^�d�� ��g�hQ݆v�
�1��0�~�/����m���xu`����]o�`1����Ւ��ZO�v�Yhϡ�")Yػi �M��Pᜉ�j�Ẓߌ��!�~[a+*��\�	�_ ud�a i�^����֕��:�����H�5���i@b`���Ҭ�N���#�++����w�cG��~>�4�t7�lpº��d����i�B��!��'˧n�bȝ�F��z7�O� �c�Ց���-�(
m���.ֶ�e�zE���,(�4{fn���֚�h����~t���!��O�XN��f0�����ؽ���9B5���RJ��5�S��'��n�4��U`n�^�ռə�@�6i��;�7)���!��_������g_m2�p���(�{�Z��`s��)��Ǣ;k�a[_r�;ݽT{�pf�_@߸dv��TA��[��bczW�ʢ���[�2�UXC\Q�<��>N�m����<��n;��:D30������%i#o�h�ϾȜ�fg3���g���(!�7�#�mR�ҧ��SB%��������9��D��[�z�Ni-h�11Ie��f7�A�b�\44)fI:RAenK��C�X}��n:&#�H�J�ߚV��m�bI���/����5�e�Rp�������/�:�����_��ac
�?`�/�ڥ�­Q|���o�F��&'z�(�~h�T�fe
�2m�ZR$*���;��wB�*X�ߠB� >&s8�o����~߯72j�X%���u͏�Hno�q���l�q�ݙc��5.��̈ɺ�z� t�~�4�n�F��u��mW�-X{$��ll2�	t7]��F�ٮ�[�o�P�Fz#��?wm�F��V�`A�ܴ��)DoЍHr����&�,���i��I|��[��V�S3��B�h�K�0���!�Xh��i{eh�X?��M@�~��iՙ��O�(�o*ƏV��Miġ�Z*���w�04����p�.8R��b�m�-����elM����ʕ%1��!��x�@��Ұ�A!�E@���a�q���b`�41��]���u ;�f@j��h��6u��+3���!�)c�HS2�O�=�О��);����J�X���X�bRLfk;x���I�hb{4p���g�<A6=*�q+Z�$O��� ��n=���Ёݧj��
��!�C ��#0�Y~J��o��>ݙ����\o���Fq��#W�(�2�o�s�
��đ��|-�H?}� �ٯ����Ć�mk�qr��3���Bk�%��tm�OP��9��M��`�`�����e�_N���>�UN��JӮ��>���C�8E��y�w�^���]RO#�H{�>B�����	�q�K�p���w'cYQԵy��|!]D�C�N2�R_���
m����b����I�a#��I'Ň!%�H�4�V�VԊ=���@��"�e�/���Gwm��h���%1oxa���E�>��q���L��{�X�.�/y�P�&ך���EU���f�J��P�t�ޔ�}�V�?\��P�,�}�9���V�>�|����"����y+��?�S�|�≄@E��{R2�����TN�"���$i�}�KJ�{�t͚�'�C���K]3�v�{Eɤ�:����P��r�1b"1��G�zt�u]���7�����.h@Wܼfk�<�n�b�B���5�DB�k�����=����%8 ��(9(���W�F�������g}��mN�U���H
����cǏ$]/j��*��b�tTB��CwOI����̲]"hx���0H�Q�^(�.	�f���8������զ�%��2l��W�����+�������7��R�����4��\?�*�F�e8D�{6��3��JzNǪ� �g��*�C[���	Z�a�\�o�Q��-��s��@ݴ�&���[-�`�@��4�iY�(��ng�A�l�:�����E�ʿL�!9�P���h�!�2��uO���hI�7bfT��d���D#�-�cY���ؗ�tŒ�4u6o<d�ؖ