��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$����T�(zذw���b��6��"���k������`��f�)���y��\���|���2�� l�C~�*�hZ��\��&p(���M~�x���'������0�m��tvwԏ�Fg^�]�6���Z��]�(�}������0�Q?�p�I�n���V��dDe������l����G����g��ķ�gA�ˇT������Vi��j�(�L��,"�����{-��o��m;B���u��h���-[@tEƅ��+�Us4�;dپ�uk�ǹGj8zUe��r�?�{R�� �,��S;��n��&*�O
T"(Oh+:F���HP�����Õ1F�yy�D��%���̩��W��g���ʢn����$$Q-	.K�wd�j!�)?�cR���HM�*���*]-b�8����Q|0Z�$1���ў�����\~$��[}�a��A�P/��Tܳ��
�ãT2KTl�ۉ)I��ĥ΂�������Ȗ]#��U#=��C�݁!�HG[�@>��+���M�p=�t�|g�94j��+@��YHFO�Gx�;�ě�
k"�|,ct��V�|�݆�7���ʳ�ѣ_�1��Z�e/#^K+���J1d���̉i?��)�8��0�Ƃ6�61E��?J ��w�I�ء�ܲwRY��
nW�)J�[���K�-k<�X���4?Ec�Cx5����SY7S@䂍R��Bū<Ƽ?��hq����t���G'��\[��p?8�Nt��<h�"_���`x+�k+R�S0g�j�r��:�P~k��&$9 $���������ݎ2�\��7����H�/�艿�����n�J��xj��&C�n�(蓼I^g��M�q�aD��|��qL#	a����TVXy�H�i)4<������)j��Lؔ����/i�tn>O0�F�/�:T��p���#��*]�L�r�Oh��|���1�Ws^�خI�b�v�K];:��<��ǆ�Du�Uh�8�d�{�^{q[C�޳��E�M�c,�%���Ě_����!�W擖�ho�M��i���0A��9š�*fr1erq�=�̘�����d�
}�_���+�<$����rB|R�rC�1E�i��yT7h����Kl�ӯ��>߁����D�r6��E%�4��N��f�d+{�+:lM�~�wp+sj���8>��8Ȑ%�.�
̗�7|3:Ma�xue�@�
k��Ԡ���0&1b�^����7��2S,��'���� ���i�Յ��-)o��5����
6G�c!�Nu��δ���qD�^	���l���O��uM*x�$%`�3*3�*l՟Pd�͎q��J`���1�w���mFp���0�[�N�}5��`������?��Ͻr&�������d��<��щ;	x�����v���'�����Ȯ�sӭ���\��N��2� �w��3P9�œ8���90�g��P��,J��9�"�ҋ�Y
[�;5���=W WA��Z�J҆�F/{os���Ȟ!$	�xǉB�
�����+z褝5�"�˻3���&�7F��uD!�5�%��Ũe�eΆQ?(c��N��
�AC�˃�z�����|��I�o�����Gr���G�y�J��MP[��S<�{��f*?+5f���� d�i�"�!���
�&��2���t��z���#��t�"���Q|�3�յ)�.O{�r����5'��u�� h�ۆ	�l���u�P���8�X�h�H��0Gi���O�d]��6��W�%�����u1�r>+20ȏ�E|�dl"���H�b�˱��*�$�*'K���	_���%�2�g�����J7�;83j�e�W�_DE�G�T��	�E,� ��./\3t�1��%�yw�x�C���[��ཟ�p0�m�yw���
������̪��VN-""m*�
�ZqS���k�]�);o��~��XK�;^x����t�3?�����=�qQb4^=ޏ	�E%x�!q:��_6�`�ϱ��,n>��:��X�F���z�щ��r�B�i��N�#Z�.�0�x(>�����H��]7��d�Dn:Ә�U�?�(197�5~+�{�#f���ʀq�B�rB?}c�5�>����ֲU8A0ѢfPa�ò�L}�!E ��!�e �N��U����C]o���hʿ�����p�h���!a��B(e,�BT��Zh�y��*M?,�@�O�Sð�ou���7"���B���GnE+޺'hGn��ex�,Cʑc����$� �A���~/�1�ͣ��#bbc�4s��M���&��ۻt�^����w篁k�m���kص))%5� ޅ�nf%��,oJޕ�(�%e��>�#���ɲH�����^pkE
(`�M�x�:��*���I^���'����3(EЇ��D����	kPX/�P�!,40�;�~؃��r[�m�KL�&�PB�� i$�Qƕ�d�,�"7�[6�W�n�ƹ﷭y6s_݇��V�/gD����R)��9i~J�ʚdgy�T�]��iN~{컿��%Ф��b�ai��I�pδ���7B����u�/��R�	h}6m9�b�8ڥ��0ҖY�y���q���!�/�C߄�D��EA%���O 0+��")�x^#��%c�L%�OI��F���*�!���n�525�9���Ho{�3!�a�
U$�����9�X�n-���G�a�2nSRW�Pc�@�^�-�f���>��*x��U%3�K����df5�Ϟ|���%9�Ș�ҿ�qъ�8I��+����]U`۵zF�H	��l���ŞmU�b�[�6:�\�ap�Lc;�����~�#(S������J	�����$es�B�m��?}��N%DJ%�n2�K�'��h�!�"{.[��P��7��p�;�-c|6�I=�:��JQ�B0ߎA\�8�fB�f��x�:ߴ���E7/����sy�t^(=<Orz֘d�P]�8:�Ve3'WY�Զ������,��&ᮚ����Iz����L�!KP�}2F����@�Vxr��y��p���2A���̏o=܍��4���LkNŏu�������3��|�A��B�h��L:��Z��FA�T���k*A�� b5^a>T�A��:�b���!)�������!q�@\9L3��y�YPP%A>wf���/:#���lk��ɳR�����N,W`�t2pѩuB��(�"}Z�����&a����s�^���9)x��[�l^��;���$�#Ē�+��I�RC��]�Ň��J� �Emhq0T�SvQ�	�p`K�N�5�:�9ۯܨa��k{o�-�i#��ǵ��Iw�(b��լ!�u[���G�O�������]�]�]��1�0Som~�,�dJR�I�Y,�;s��fŁ��,��_��f�`ߐ�҄;/ /�Дb��Mz������CV�}I� j48l�p����G\�Wײ_IS��"`^�w��-�����I��}����>=P�����BW��"�G���U����6��(�rGt����O�AG�\0G�BG��I��>��oY[I�ߺ�wO������SK�-Ǧ���<2l�X����P!���fb�3C�� 4���%�^�?�߰�3K��mW����z?��n�[L9����ެPIH�;gޞ���t��N+S����D^`H�%����tZ�[ͤ����QTPD���ip
���iV��vr5���؟L�4h3��Ӟza�~�(:��Q��X%�Ķ��{.&mdp^LhT�{`\j���z�T���C^Ў|�p�n�) ��ha��̬�t�0��q�jJgvg�Z��,^�y,�ӟ�m�՚���y���=o��-�i����!����fu�����6�!��]���U|wE3���j�������qY��䳒,���U����Y~U<��g��l�[2r'l����B~��N��6�̻`���4^�ɓ�#�SDD�S5�Wʹb����D�8mZg,�Į7��z�^���K�T����p;��yL#r2h���qPf�<�ɞKۭ_�xM�YPs@����Qr���5i���W
9\�N�ۣ���\<��;�ȍ��6dU�&�:bI �Yx�/ƽ�k�D�0������:�0>�^�R:
�G��*��z�	����d�6T�t	y�\�l���5��˹��{у��!�y����.��� M+
��+���Ĵ�*�%W��J��Xţ���-
�y#6$0��zeg)�1Z�����iH�3~�׷��YA�.���bL��Mډ��9�V�M>xN�K��7!I
�b�,����o������_2��:��!�ǙV]1�:~r$�d���&�d����(��A|�w�:)Te�
���6��}ۉ��>��G�i�K:R���	��ߤ�u��h���G����A�z�\x���Ivs��K��8.�;�����ωY�0�Ϛ�Y=ͥͯ�B�����"`S����ܟ���� �\	9�=I{�ץ]�D���m;�>#�1	0�/�j��M�K� �5~R-i��Lb:�{7�Xq0�6I>]lvv'm�����'���1C;j�q�W��I�{9q_�[-+��TfOs� �;$�i��*I`��(?E'��al�>��j��Rg����FJ�Wh������+;l�6����ٛ���kJ[�Ӡ�ξyM�HOAq������M�~�dc)�|��>�mk�1����O%�]M�a��f�ȵ���80�;� ���K+R�a��V��J�(w��ĈĤ�FP*����+鏣��ʟQ
�tjo�A���<��I�FJ�Z��`=ڳ��U[����v��)(�fĳ�m�2uǯv�X�ͺ.u�ItDE�Y��Q0Ag,цy�����&�f�<��B%x�;���k_�S�F�,k�&�{� ����/�/c7�o�r"Ź�1ɨliwz8�������I����$��" FH�a�C;$O�9�L��=�����i ��+B�
���ӣ���Գ�?�E�F�NYW��̐���@�D��)`�%�ݱ�?���u�ć=Q�6�9G�i/�G9a1������L	���F�,u�v���z�u�CڛAM���htI��������N[���d�����>'����Js���
ܞV���	�K-/�yY�;�6�8�@�s��L�-K���ݳŨl~�g���Ԧ���l<��YO�l�)Kl�O�Y�+B�BV2O�����H+�+���������祥�����6��p����Vk����_
�����D�7����9;���of��^w�L0�dj�a�0�_��M3FJKT�u���B��^�&[��c��Uv
oγ�dT�7����d�W��>*aڗ=v����4�@Z�S�e�Y���CcZ�l��%�*�֗vI8��_#�ޯ��#�$R 3�8�f\o��-�S�T�=��,�.):���ᙐݹg(Ua})��c�]�@2l����0�T(軔)��R���IS��`X��b��n�`�6�X�ox��J\�8R��ԷG1 �ށR�;9�Q~�ѣ[�j��Ao��������P[���}�[_Z�y֘&���hK*v�]�Ғ*(n��xG���ZH5�
���:����r6$[
�|W$Ǐ~�pבuَ1y��P3*���v��h��Z`��̽�2�C�pF'ơ:��~�k��,������0#�l��;�����f�����0ie���/���i`!{�6}���q�ƕ�����E�}� �����X�(PtW)��JG�U'����#�$�����W�S5{/�]��志�>,2Qv���cM�û�kV�@���D[�S8�-���h�m�MRb� >G5ᙪ9Ǜ�Y�%�������X��e�l?�,��0|&���ņ�gQS���ܥ��S��ބON�F