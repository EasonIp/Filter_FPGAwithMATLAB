��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5j jQ+���t��-�/����u��̩�Xc��R>G��$b�xA�Fn�z�F�X�Ӊ��q	U�z�qG��f;���,-vl��� 'J:>�V�	��0�7"�%�˝էo%���7J(]�7(MGw�rL�R���<c{��y�y$+{���k��6J?����ye�@��\��q3�!6���J�9�I�ʋ����K�e��t�f(��oǎqz':ݶ32/�.��.N�
s)��9�<�2�B�	>?�����V���c�Kz6]��0;YTHܧp��VS���J�0�L���<�0�q�j��`��Ѕn��-޾�Q7�z��׿�<SP_b�
teuϋ$y}�U��4h!���'N����F*9� z�[�����B�'6$���111��>x/�mD����_�X�5"���B��h�`�I"+F�8 3��R�f����<+:�5����]�-T̖�ߒ"���|�S����'l��]{�`!�к���7��*֨h��3��9v�w�'F��	�;����=6E�EfW"�UB�t ����Å��KKY��Q�&�5�c�Dv��7X��񋕲	+y��h�< a�D��Y?/��Mio��dX��vz��{[�BJ��?qq�:۟�hF���X<�:��/��|�5�9�_�'��0H#��丯����Ҭ���@z��JwHy���F ;��ʻ��ÛV���Q���>��{y5H����z;���Ǳ-�a��!��m�V��Q�J:p% ��[}���*�ֵr�P��ݯD�/�Q���>���ʜąïI�MH��V�"�HMf��$�o��c�AUl��K^�!�p96;�����Y"���p���_�a^!�M-'W�[�r���pU�w�i�)G��mr���l�����Ə�?��X8a�o$�P��L���'���_�H�4�>p���-�ޛ����Xyw'�(�ha���7��j�4��<W\���dJ�����غX��X��,a�����IIh��w��x�{(�	/����,�+g9���a�G��kp�"�
E�)�v�<�e�7T=gA+���i;��@`�҈�f>Iپ�I�'
6�b~�hj��0���g�l��eD�lX�M�n���g�*�@> �c��0�e��C���k
�8���ZW^A�?�)寜M�?���^�[\�*��ţH�ShL�`��w��ե�=�}�B��T�K�XDr����й���9JS$a��J~���e7��&��}��|,Uc �rP���H�Uo����ֈ�T�����x΢�����;�-����yJ�R[AĳɊl�8�Z(�������k��*E���9ܸ�]�W3X�N�H�ӠA���
����۽]>��V����;�Β�\)��U�nyiZ�t�����.Y��/�����k����罇nИ����p���5^|6�����#9���ͨ>�g.'��Ghgh��o���\���"��Dp��*>�w�(���h<��M'=۞k,�\D;+��?к��Q�A5�Y�
��ޯOx&�����Oi����.<�T���E��t��]��e����;+�T�ù��^�r|�G^�g�-�x���]Cͩ"�*4$�C0���y�(HXL�M��W�S��ȉ������
��s�����ȹ0��Nn[J�Q�Eg��kT?�@�^c�oz�N�� ��{��UC(N���7Z�}<L������D��L|��!�즸=��Z���
\���ی����j�SE��&������s�b޻�gHi��T7�.N1�|+*rW� �s=af��s�#0�K�?�Ovvy�zI�.���ϜC�o��]A�i�š��2���GH��-��c(r���[�zB�
�QK��wd}�>��I2�  ���y���xuB�t�ܢS��	�]O4�f��Ŝ}�V���X�D�m�$��aSf���,3l����� ��;�pJ��T��H�GuR%@(���X,ZM��Xl��ls�#���񝩚XМ�� ��g�]�w�]����t�f�r�ZG�A�D(]���j�6M%G�9_���BϪ4��g[$�Е�Qq1��^-�x�Ԛ�����Ay;�ޮ�ǆ)I�C@P�f{�fs��5{>I*��gq�WTE=)MSv��J��}�`���i{u4Rﾑ�?���k:t�+�@<7[���dp
��lv���i����Ӕ@b½�m=�]����	���r�p��&��2NZ]��g��i�2�|nP��oF-d��0���:��X\_�b<A����-�*۵v�� Z��!����4��ca^� �q�#�`
<2�ٮݬ��-Ͼ�3��~�協���r��f������������O���R���0eL���A�)��041��4��/��g^{ ��[�S���u�烯�;(N�"�m�-y_.��_cl����Q��0cz�c�3s�-�dK�y��K�#���Ax�A�Qi(��$�r��qц���oY�TΫ�	l�HN*��e6�XF)u��H.V�g}��̀�^&D�� B�Je8Dmՙ@�����2���;�쇊gy��<v��@���/���=)x2��o�
I�΀ r?s]�Tmt���Ӎ�B�?�EnЁ[~~ل �B�Ju���L3����1L�A|��O�EA��Ɩg���$ݍ��֝��n"��n�g)ܘ��)\Y� |�'����ۄ�m<<�\z]���#���͡@�v3��ȟ?@<��C�9(�	>P�<�T����)����&X
��ᚍOM$����&2��5�y:J
TgrwEA�˻.��p�T�nT�s�Ge
U�9���-�y[%�6�S�^PZv����悼t���a��-N֗�R�!C8�y��G�r��8��lӪJ�����J��1A�>���*>�\�E���Z#��,_1Vre��֟���R�WE��0�`{T��D�ק�7��,ޯ���5m^�~R���������F�%�s�Y�����]ctyab\WX����2tu�ɬK!='��[�����;9X-W�o��C��-4	c�΍��r	��į�|q3Z��h�د�%D@M����.�*���}�`�歟�F����?�����*'�zŖ�
�י���J	+�R����Q��(���ZJA�9Y�����υ�xoW��������q�����*�D���]�ш�]�����80L'�}�+���Bn�©1�`��KR��#��]Y�ƀ�+l���;��&[{���X����țԥ3��6��n/~et:�w�6#]�B"i���^MaMl����`��&F��gƄ����b�����ٽ�er��g?�6�n
��\�8���SA�����ַ����q���#��/6A�ap�l�*݆z\ȭ���Yn-��"�\����Rk8��*�k����RT �Ij�\VQ�e�f�e��ɑ���b
�~P/k���C������n:�}�H�S�Ȕ$шh���@f�{S+��2������5j�So��%�	W�Q�`bL����6}�Z��$Rr�R�����аn�o�:�ޯ��؜>O\~�u}W<�dE���p�g���So֊���~�PZ��Gp�{r��e��܂��w�-g��rd����i�i��8_f������T+�@��doKf��i���G�ȻJ2�\��������/�p�&�b!U���Ȓ���7��ډ�aW����cM{\���Oso�V�-�����{x-���k�˾��B��Û�4���P>��������f�Us�6�i��f9թ̳��9i�ɭ�n�4'���-��̱�g�`]�d22S�fۤp�#��wN�cڥtk���e��A�-"���0�:��
m�L�ǃY](��G�%���ߨ��v�%:�HT6:�4����ض��y��>�(��� �>Y�*Ln�o�W��/fn��%���,,�{��X�(�����9]��@5��#��z����k�p>���	�ǊkS}����(no|b�¶"QM"�XOD��6�,��Q;�hK��¬�����)�j��.�]c�[��~��ƺz������!����G�c���U���������"x�֦k�(�zU������'��_H}oX?]�|��K��-o	�L�(�V�{RI�ҧl�l�����ʂz޾Y^Z��
~��
�������=�l�[�s