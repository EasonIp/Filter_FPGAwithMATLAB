��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$���v.�Zd>b������81Е�ߋ1[�x."��F�cܻ���9��X�P�v�>���,��'30�b���E��ٞU�n�MV�5|�fH�}

x�ĸѝU�k@l)�$w��˔�N:���,����;�������J~��^+r���ߐ_��;�ؒ<3�� K���ϹHs�K���m��R�"���ۮ/{���|���ݯ�j\,���Υ�Mn�T7��M��Z tB-mΟ8���T+=�<.�|6���-��Ik��٬�Tي��R>�M�z�9�d��u��Z����#���ŤB[|�U�ϓ�Hw�lQ�F�u���i�{��Q��ߚ�j�Q��os�"ᆛ�m����>��Q�_���~��^�����T.��Tg�4�����R���ۀ,����S޺�"������iIY�������9.;�ś��Q�3���jKb�S�l-n��b+����kEz�d�OM��SNF��X���/�;��R^��)��>��<�;^�3�Ү���$�d�{0�Z����+'!9G�WLk��"��.����w&�k��*�'�����5`���!�1A���Ǩ��n��}�)���e��U�C�x�N� ��f��䰋�9�T3hP�&T	ψ��2�X���⒥�/����_�j7X]�ݽ?��(N��u����*>h�����!����1�,���g���K�� k����#i��9"\�ƆE!	�β���DD���?h�d�Uܫ��T��n�x�����bJ��vz�M����J�|_��9��ǥ��ݎ���?��f�?M�r�����בy;MҾ���2|�u/}ԶM�#���ދg��⾄S�i�c�n�
�GB��������a��sI�xZ5RtΔ�D���Y�а{b�!#b븿��ktT~2N�1���E����	6�]��)S�aW��!�ȓ��G׵�V���n�).�+Ъ̄ą���r�V���d��G�v��zix<s6]�/p:�j�/��lޛ�X��ʥ�ke��w�/���"y�� � �~*k���G�%&�m��b��*��O�9��~р��� �l<��WU��7�w�j��TO��0������$����;��)�K�"L�"Sn��M���p�$��m��k����_m�N`@o"m&D^�ʷ���2�~*a���~�'-}�4�?�%���Ꞻߪ�5��r� u()PP
!������������l�$$:j�|d3�@������!+9g�ST`�z��&��
�:~����LQ�w�/�X�W��'�� �8.Kk&�b�e<���`�Q����t�C�즱Kq�[�y~ Ḻz���K|Ŷ�[� �B��i�}ܖpKѬ?Q�0 ��qօku�w��Y֌vVY���4����I	Z���(g�C���.�De��(���?G��C�D��xގr5IR�Ƙ?.��'H�J�p��)s��sV�U��?X��#zsyS�%�e�-�I�݃LH��`��)"N'f�D5�I��c63Swm���R�(��~3ĹĂ'q�IE��P.4���U(_:wd�zZ\r-:0��z�=�jF�N��Z
�����kO��̵؍Ѵ�]���wl�4���M7M��� P{y�u����`� i��K�H�Jγ$)��xV�)i]��u9ץ�A-k}+��`7�z�ߦ�M��ظ��Ͱ�m=�zwY�n������6�ņ�������_�]]�6?I�bM���e+������&���59��P=P����움t��b�6�����#�����4v�N��)�?ap�{%�5p����a�e�p�mq|����c�(�+�E�`)�?���_E"+���g٪)��%Tȕ-y����(�h�0�ZW��%> ���QFԛ�=�$g��d̅�N%^/����Q���g�يk%ό$t�٪FXV��c���ȱP!?����]F��.�-��Q �d:�Ʈ�y��3������7�)�$����]���]$�A�)_	���]�"�חR'�-�s��_����b9��t!�P��풞���<̧�P���Hk��BEӢ,���/\��B�\ҍT���(�l���y)��(Z�>����w`Q~k���@-��V�{��φ�ߨ�n0v*��Y|1��h�u_*�}U�"]r-%�V��ћ�S{�i,�o�O	���Oz)��ޔ޽z<%8��f�c�8q��]����Uy.g`na�����\%pD.sD32i	�mR�6D����}�T�݅��*�M�]��O	s������.p�O�y��f��ȵꂏ
X�9�gӆe
x�T5g
�_ն�l �c��%+��Q�k��$2��"��[YiJ����`̂� q\�{�B��7Л�r����؎�֔��*q���rfi~�n���4�9�˸�E�`�%|����v��d�,�d��o�� �4���yH�L)��8x���8!*�Ϻ6�-�G�2�4S�W��i�g�}�M�1fO"�*��ũi��OT}NuJ�e�[� �
A�1�1>��]�������)l��h;i冿����^u�e�g-��ȯ����%aA��1Y����@����/�y4��@<�!��w�,~�о�l�|�l���U�][>�T��dğ�{u�e�3���6�p`q�;�����jV���H|����l�G�@|2�8L�����RJ2͕���0ػB���J�Qqr�i�%	���߲x�k�j#���O��J��a=vK���2��c�*���(3�!}vP����W��f���-~���쓬�S4��g5�'�'hCA񛐡ӌ���1$z���?&'��-��sA��]��+��5���6��-|�S��v�.��y��+}#�� �������qG�5�û��˰�y/ne.�^H7�7�����=�t�.Ii�#a)���$b>���KjÇY˨��T�*#^d^��)0������
a)��,Jy��1pXq���2Lؔ6���@U�3j4}Հ����4�%d�EH�̚��*8�?�z/�J�ື����H��V���h���|r@p�E���j������Ú&����M����������Q�m҇�~�]�뜩���? b�7N�lgk��/�v�faG��7ޤ�>�E��'�Mw����G9��� cc�a X�wn�-s,w�fC�T!h�ܩ�	MO=g��%0
j5�Sv�_/X}�R���L� �Z�Š��{>��./-�1�;!aN8��8�h�0JaX���X$����Pȱb�h#+�B���b4y�K�&^�Vm!��T@��6x/_v��\u����Mn^�PIc�	!�D���͇v��q�xK�!ug�ݐ����o��@Z�G��'\PEFF��Np7�-`��zqc�$��Z@τN���v:�4B���<��y����<p
y��G�4o	�{Og6�-y� ���U�u���?� ��׆-�LB�A�+��Nޝ��-� '�
Ǿ�v�%7$�QJ��� ��t��A����[�n��^X/��Y�
�I.9������B?܊Wֺ�N��+�|WA�dEAdxn�>r:t-��m*���e�}��"O�����*LB�s�}�jǋ=���q�A'*��A+���MK�3 �K��L&�J@{�A<$%+�pp�;N���1K v/_57C�e�{��XC�~By�_ڸ7+Ģ�޻)�(��T*�&sG���4�}�{^Q��2��_��O�!��1�C�L(��8'ԓ����<�7f��=����E�#�7�>�}�X)�����G�ed���(���tT�z��2����^��_����C�׫��=E��Ec���E�l����P*a�{1�E6=��m�k)xpE�4n��h�7g�(���d�	��y�T��ݿ�A�@U��"��ʮ��E["䏔궑����C�0�h��S��HW� N�g��0N;5y�m���l1�K��t�Az�]Ŀ�P0�|�6#�e78�]룶6w�V��1�Pj�)�H�����]dY3˔�N��[A^��Jn^��v�-zԅä��7M=�ϯȭo�y�:.�5%Voa���'d.v��2�Դ��d;�q��%��)�)c�f¤]�- ������;<0�i�y�3��0��P�� cY��$}x������|cvA�S�a��bd;b�����+ա�����Z�F(����T���@�hm�ͽ�r�?1�x��O�=�j��S}9CzDR<^�ـ��sCy��?�!~�/�ӂy�PE��~>^6�9`����h�d��ę�K���/�Qs�EC+T̵ 5��6̔α�I}p�
ĕ��ƫD�6�Y���O��p,���Kh���8�ou+p	R9�:�d	;�Z+׼b���6;�q`*G��m�J���M^қi��yB%Od`V�ٔR����H�wvp?ȃ��p�%��S�B�Gу�Pp`Y�߄�Q�����~Sh��́����ֺe��4��(��h���4SKx� �\)?߱A8���#�9c9�Yt���*��.h�F�X�8 �(��f^~�6�Ȧ�������h�uP�
aɇhe����S&Ym�r�/6A(`���-f=6��#~&�MPg6֡���P���k�d�{�3~�����ҎF8�?N�EC��c��l������6E��F�d�M���M����{��)�3�;fv����lv��pD��h��j܍h�o�-@�ج�5�	���yY%��[l�܏�� ��Ą�izp�ݏ~�+�O�u���Qb)�Ŋ�}b�N��m�!fYj��D��H@�o��fG�n����W�8� ��\O���G�5~qj��my�����2s<w���{vv]|�ڵ���xs�7�H�SY/0���\�-��ǹ���[L���ʁJ��7SEP�kd#�N�꫟�êD1����B�/�,�����Or�����gp���4�CyhP��$je��C8�M��7��0�^Wu�G��.��I�";3"8k򗹿��R�v�~�g�����+��a�٠+x��:S�HV����f�,"˫��`����Þ��-p"4e/Hx�Ȟ!~�
�|����MgP�Zq�i.��̝�9�_Y�D�'��%ǔu�bڪYF����/�4���-���,�CtaO�����}��5_��;k��Cau��fG3�4�zQ���yo�#�_?;����8^�e��.�{n2*�5N�����l���J�D�3�71et���V��J¯�lzW�"���t��~U��Է�Cq^Ol��q�Ρ����}�kM�\m��a#7��c���cyL�R�$m�!���(�ƅ��o�Wg�2��˥�~�\�^�t<P�1��k�Υ+d��Ʈ��1�-l����
��`� 9X�̍ۗ�?�,b�����c���X�l�u���]8��j~�u�^���斃�O��B�������\������o+�����:S�qC�Ժ>��`3��S�P\�RĖ#��N֩�@�����a�r��q��LFbcZPkh��Ӝ��G��М[�����.O�'�h��i(}��o[�a_�!��'�֏��R�$�|��9�nH�/.!�[ס�g�f�)�3+�YR��P*+������g@!�B먛�����MtJ)9p'���+ʑ��G��0�j_P�N�;���2�S�ς��P���0'u�
bppdl^m��z�����7�
=���"vMԩ������-w�����M���$l<�(��7��E��i��ZZ�a&��`��"]k�L�JwO3�*'!ܭ]�M6�N����
��rR��d?ѩ�����+q>�:(�-b���s"e�3
�y�t�����c}�c�O����$��$��?�R��[`�ee[�wn}B9nt�g��}<����hs�����?�2rb���$E�B�Rw<���_ �����!봚w��͓�ߦ���Rg�o�)��k4�̵�Z[�<E9Z��8��(�dU,0�h) �{��G�e��p(?&~jL�%"�c��4��Y���Xʁ�B���|v�3y_�X�ʪT�v��&���E�BY�b�}��\�ڣ��[o0�֯�1�릙�_��/];r��Cp{�zcE����U�$c[)p�vR4$�HXl�gG;�:��-��.O|4N\��T��Z�7>��t� %�E�#�^4A�v�����~]�L4O��)7��D���9>MTUL¤i蒚ǛB�M�@�k*E%a|*�������1k���$/�/�]FѠ´��c���0��̓���QF�\l�x�0�-l�%��m6	�W�"6&����A܈)�S�6��h�d_����a�)�َ��))Qm���c��Y,�E��}��s5��6��A��3�3s�3^vt\?0.q�,��{�Z_�wF�vJ�'�C2s�l���b8��L����vW��-*��	r�ػ�9��Q�9���T�������}W��/�T�.�PU�f	tW�ۭ��iV�Z�톯��v�����;���Y��#����u<hn82��������w֟�`�cpe4�3����'x�4}���k��ql0AXM�f���ٻ�jj��\񁒁GI����������QɃ�����a��}��˙%�8̷+F{��ǭ��	q8���}�]@�hVS��v�H�gI�]�V�-�p��Cb�����d8����~$���^�eQT�
X�^�:�0�P,]q��{�)v�_��K�<E��@X��-MĤ3��&�ו �n��;�e��\~ه�s��O���9�.�P, �Ń���z��2�M7�qL+�z�1���7��`��ǿ��,���s7b3MC�q�v!V��$�@ϒ�+\р�