��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4d�#尭�ǕmpC��՘���z����m�0��X�fծ�+oa���}˗!i�v�:¢#��������<#}>!�K֎[�y�����,�]�glfs��y'Myh�ܧN>r�|j����'n�XZ/-<P?�Ah!LQ�ս�����]�aI�aM*�zZb-���o#��̀PZ�|P�	����ŏ�G'׼�<�-�w�.y���R�$Ei~�t�8�ix�98Oe��E���A�?�o��5cxq"XOw�at�"b?�Ԍ��'��nh"����&̆�h���q��2
�6ε��|����	ƌ�(M�ۼ���T���L�������E/�����?n!m�ʁx�A�#�̫ '�U��}պf0�=���K��y�0]�?Q% �~�ڬ+4��h�;���W��$X�Z��Q�Y�cp�V��2��7{\��u�.�,8E�s�iŋev��0]LY�3��yض3��&�Ա=5�<�����&�#vȁ�Q�,8�f�|n������m�,)�An��g�,�)s����=��PW�k-�z���b�� ����x�LsW�]���S|}x�-T{�����Li�v9������m�h��\`�+Gnx&����D���OA��9�@?�P��ߏuE�.��� �� �iP�mJ�8]�K���tf���s��iϭ�\�7a/����rz�N��U�$����%��z�Z:ǅ\�đ��ݡpx�0g�8�6�f���
�����Cq+%А����O���taqPD_���V��>_��"�`?��<$�#z���1�Y"�4���X�ݞ�OB�9����m�l�o�r��Dbp�g<֫ݳ��.�4b��;���Wxi�����0:��+�� G5�x����!X�E���I$DP+�?�u=<�3#�ۅ�tt����i�9������"<��cٳ�oR0�`s��B7?�X���X��X�oE%�_��K~d��l@���(�y{������
�,L c�T����G}T��h�XYVR���|3�7��ߺ�� ��o%w��|;*�Z�9k��t�Ʒ�'�8ӗ~�R_�"8	:`���q�^NDH0{�=�-V"���38ޚ�'��Cݳ4+*��Į;�'�Lc�gkz���VB2la2�di�.�|=��~�/t�uk����$ �D;���:cOz ���ٔ�+���$��v��	|��J6�o�ʳ��� &�:�>�J��,n���xCf�b����*��֩���_��y��[5j��v�"�׬j�,?&��C���|<l�A�������0��l��
?K\�M�E�w�0�`��*mӣ�Gv���N���%~�qH��t�8�=��!t��]����w��oBoh�f�R!'L2�3�e�(�a��m~Ab6
)Z�ٿãI2	4��:����-w�|as�9�TTTN��1��vT�;�㡺�ۥ9Y()�I���7��;邴�RܱsJl���vb��'4�/�֖-L���8
 �/3��Ӽm�4�8z{��i�h(��f�i@8l���������3w>�ΡF�^�W;%���eq����{���*[XV�|:�[�A/��aL�����5b%�m�X�q;[Պ�*׎���K��4|׆�z�ٟA�$���E���9�� ������͎��j`�'�5����%�!��dr5���,8�>�.\նE���C�[&��2&P�B�3�aFRM��
x�.Wys�b��a�BUg������BuW�lc�G�Ȑ���6�O�]�A����:�#��v��@���q��^�xQF\̧[Y��jC0�I����d�_Ã��<\�VbL(Gͭ��.�΁���#1�FR�nTRQ/�����s��(��>$Q�_��X[;#��v��`(`�7)X��W̫�h��S�N���9G�زg�f���J!1�e���i�həJ���d��@��%t1�)I�k�7�i�A�ls�v=aF7Ma�9�"��l5K�����W��u���CL�7f� �s=QI�����Mg��Øx�0k#ģ�Vb�$�o��ed��r��x�3Y8�����R�G'�O�,�ce��Fd����IE\Yn0ݬG�CVҝ�2dW.�qD�xЭQ�fi=gw������Q���Tl�	�!�� ��^�ъ����v^����D�tB4�k�GZ*����J}Z�Fm4"��6�)
��=Ē�@���4н׉�}#O;�~c�_ӎ ���d���H�AFd(����e9�&}U2}�6�om(Iɍ�뱷/����q�?��4qᛚ ߳Hx�4Y��a�k�������E𜅑��w~(�F��������4~�*�R\��	�m��%�=��J[�����7�!����Ө3b7JB�3�n��-���4�T���CER��74"2�O]j�e'�CVi8�)�����~7�d�k���O`�����ы��8�AD���*{v$!�6�߬�g��,EV��~`�cl�h�]1~�2�
�6K�`
�[�+{�K��)d�����'U/.F�,�'Ҋ���4+<$d=�b<��S�AL:�P������<.U6.��wS5�X����������te@�p�[�4�׽6����6b^���Gq�|�a���<�}4�9�`�8=���zn�4^���A�H���B���V0���&���&3����؋���@���4����ޗXS�'�z-�����\���U���w�w��D�v�6�]�b�:��z��&~�ɣ���%����|�.��~ʷt�ή��ø���mk+��)y#u)����A|n�f}+&6[2��C.��ѲR"�]��Ჟ:V������Ľ�~�Vj�7)`���'k������uc?U�����BI�j���yH�
��)��j픯�����V $��!y,�E~o�g�s�������	3@�4�=B�l�?�Y2��K�7�b�G#Z�����ir_`E��%�Ջ���j��e�m���U&�
�	�)<����W�OasI�D����
�Σ����2���c��G�唇 �B��r{�S��	!!��n?�̰��q��o�R���V>}�~tD�OU�g3Ҏ�J���?~����̛I��sD�Y%�3w��:�f"�;��X��lF+���9W|��V�6�MKp!=�d�|YW�^�����:�u�l���{gK☻�y�k9B��y-������I�Q��VF��tr��k������Ty�Z�h�<t�ysys<�ݞ��~�������N�@�4k���sSws7��@���%��A�Ƨ�.]lṑ4x)�eOԺ�\n(��=y�ϧ�ڕe8C�e�R7�V��A��/�͢	�xj�#�����sH�[;@���A�7.M�Yx� ʃ��2!B�,�U����D����O��gR*.��:2
�y�4�<�
��۸MD�mÍj�FYE>;0�*��xk6pd�j��8����b��J����@$��u<Ng��z�~uH�n�x����{��?��W�mί�2,��zK����4����d��$d�F�5^�aV�V+�`U�B�tݥ;*��|�.6�n��y����0� �C{��1���~/[K�?+?J�,�D������;]!���m��_h��H��sU�f���}qz�dy��l��'#Eݺ�P}�[�tp��������6(���ïݎ����Ca���N�
�v��3A��h7�W�k�G��D�o�J\�������ͧ��;��6��kE-���&#����V����`�(˽ÂB���!!O*pE��:�ٌic�� �@��{g��rm����p�Ⱦj1"$N-*3f^�%��bУ[�.˗�k�W�xg����2��v�φ��UY�1���� v�lt�鐨����W��Mr��y��?M��{�%zp=?d	,\��K�a8��z>��IQ��"��^o� �9��gwi�T�����L#�Fӟ��fpP��u#[���H}��'8�J�v�@s>����!�������9q$�&L�F�C�.�cG;����Iit��Hv�V�8.���N	��r>��tޫbO�?CE�(��o�O[fE��»o4���X$���,�g55���Y�?���=pǼ�>H��c�����6Q�߽d�F��T@��`�,��@��I��8���"X��D��X�^�{��&;l�޴7xY$����8M�G=��<?K/ ��eV{�1q]/Q����_�\ڜE���1~��������2?��u(��q�R�������9�K0��We �[&WK�NH8��"dC')i1�H�#�7�=i�YeiI�WPR�w�����#ũtp�)�i��,�s�X���:|�Uݘ4/�����٠���t�=�L�&�̨�i�qr��xL�y�%W��R�"
}��?�#���©���<{?q�D�h�U���'�m���'�OD��lR
��� ���ɆtQe"Hc7@�_�yQ�5�t�rbJ㓜�V���/|o ߹[���Hy!�n��oCw-h2Iu��'R��������Td{[��ǫ�Ƚ�4y5.o����()S7#�:��)Y��p�� F�wN]�Z�E���(�C$"@1C�	��q9e$P�}&�	_YO_���B;�����m�ő������F(�����	?}%���h���&��P䂶R�G��M����'��)��=�}�	�ۗ��Ѝ��o�� �
H��$�مU�B��y:q��k��+U�����Wgz�bh�e6˯�;���`4@����|��b�
�m�%�Hf�&���\U��(�E?�
�W�[�)w��ŝcTSzC������Yc��χ���`t����wrx�t�Zv��e�������F@3��N�?S'�GE�ؗ�igP��=c���U,�+�s��%4�y�Q9��$Q�����]=(�Io����z�k8�^��7�(����R�Ů�����)�zI��йO�)��4�Qr��~���c,���t2Ԯ�`y��K��<��\/&��ثV��w,��/�f2܃�ktww�nc}�o��`aD 0j��Pg���^?ȕ���^&�8�
)\o��?����	�+>4�]��������/�����nŴ�IOO V��e���$�Y9L��%Ԙ���~AO}(X�6����^�P{(M�7��S@#6И0:\���:�#hNV�L*�4g��<j"���򏫔C,��-����X��
���ܬ?��ͮ�1�o��XЛЅq��n�A@Ɵ��S|7���Dh�ɗL�W�wz`�:�e��ys�������n4��n��}��Je"3d4Ywv�u�xE��X���1!A����?��N�m��x�eCq����/fX)ѻ੸~�ӌ��,�C�(X�L�ٓ�Ǩ~�o>�C��r��ؗ�r�.�35�E�D�i����W��H$�ao�#�U��͚|pj/��vS��bU��n�B�C/*\�[�݌j���B$K\�|���8�_?w��f���Hoq�g�S�4���yU" ˈ�~���-l��h��'j�U�s5�҂:�]�k��9�7�dx,L��"@"�eW�X�Қ����Lޔ�!���S{��Z�c�A��I���/��&
�)6�+LhЉ�S�d�C�q������a=��C�_��i䛥ɋ�4w=я �Y��o+ًFdC�?²,/sƀ4��?#��/���X��s��ׇ�=P ��E�]�]�z=�ڦ��9��('t @�<	xri�U��sy˙���;��3Y��N����@F� �*�/2�{�\����)B&oV���.hn1Y?B����3�Ҳ�a3ƕ�	%��n����Y�o"��e+2�6�/f7b�<d�t�cz���x����hi݌ꂖ
ZJ����z�����]�� ����,���|Yv(��<�]�m���6C���w�$#
�S��j�B� H������JP�������iA�̶Y�a�H�O������۞&�E;��������LL#����\�\\p-y�"s�=�	g�\<���|]>㬦�H�A�k{�D7d�3.wۻz�ib�1v7�w\G��^���Dsٶ�ƈ�=��i�f~�ra���Q��a�1׹%^݈����6�
�Q�d�;!W�I��KV8L�A��;$��a,u�հ����taJa&�����3ڥP�ȧd����1Y��0L�f��XB��]�%?�̀~,g;�EV�,ߌ9�M�u���&�A\Qg�8����Ll����n��K�Cw�p;��e��e�u��*�j�#�G�F���Gv���z_�����ihE��|b�&d�0�U;�jcfK"���
� )o����o�i%`��P�,Z/�$��j6j��wFJKљ�q���<����gۨ��a��i�峺s������b��Q��|��k����d���F�$6��Lyg�\�? ��Е�?u2s�P�\�6R��@[H`D`,T��X���$�-6!�q�V�7	����J�R�����=�� ���|WmG��1�3w�A��y����aiƏ!.R��V���M��/�m[�uf|���k�P�� ���W
�m�)1`|�����r��=Ҧ���m(�eQs ;���|�S��$8��@�͹���|��l�_4��V�X��v�{��EY+1O��Ƈ>?��C%ߐ��b��kکݺTh5B'C1&<�C�`�/���1V�߯�<(&�>*�/-z7O�t�~�@�q�"J�Ie��2���"�Ozg�8ĥU��FK�SR YC(w����Щ-&�Z��"	;Fċ�nΥ�V1�WY��":էhJN<�U��x�p���;4�:��?dF(0�[6a����>�leZvJR�DDģ�&�*�z&+�Emnl��Q���H��g��
Co~���H��,ݽ�� a�ƕ�j�	�B:��8�Dt��J��p8g�M}� �ת����q�!��Վc���s=��_C��8�t$�2�^Z��O�Q$"�p��4�?��:��`'�:�l��#��@E�������2YI??�L��`��2���X�R��s}�Ad�䑍p6'ES���u�z�c)ˡC'��7�M����CU�?uي��2m�[��\~p7o��|��#w�MAVWD��X�	B��v���=��	���k�g��sW�]c����ɚ�{��RzD��uAL(��1m���^���j����ѭ:�SO�����f��#;JDrRk����ά�>�[�d����:��N?�Hp�p�);F�c��&�5z��N���B�Ӱr��5+[�t����?��(�Y ���<GtgO#ӆ_kp8ouj;�{sy0"lh��D�dG��5���� e�#�a�C��m��D3�@�v�[�,���O��h_I�$)П����Uۀ+��识�3K����Sr�)�ޯ��_��\q!�X���2q����4{�얢�OH_1#S� Oʼ�BL0�pC���jZ#R��R��Y��}���v;�\PE���ߍ�CHށ�#�Ǉ��Lʆ"n�<�p�O����9�qA��J�J�71�0˝۬�8#\�J]3�WU67���MF�������c���q2�������Q:�C����WJ[����-�J�e�⋪�JU�^�I�)��x�fi�uԬ!ޢ��	���\����,��G�u�a�=�V�S�x���3�E=��r��4�,,��b5^���2	���؜H+��r־䣱�=o�Ө��ҿ�k3�$��ޫ;�؝����?j��J��3�K���\G��2!��}����9����㚆��g���vZ��f���=sʔ2�M��[mLƥ=���n�SV�~�0Zn�z�aP����-��%����K���n;M -F�[M�������R��k�Luџp�����6���� �f�777铱���[0,�[1�h[�˭�Gj�P�����@�ƽ���˴LE��ٚc�e�ϊ�$�@\yEi�p�1ܦ2�bf2n�	M2��@�Vg.�AsNQe�(j������y/�>hO
�#V>��CV�e�1��)4��ϵ���=