��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$�ʫK�/�N�NٶU�L�Q�\�B���{P�Z�|��ħ%�JV�t0g�t�����e��k�2�hL�'�:=�����&]�aD+����{DT��A���f�%+�	*,N�~޴��vA	�(h1�0Ϟ���N<|������%�kd���y������s�5���c��-mn��]������V�B�S��[����ϛL`��.O��X�_3;��_A�W��pdDK4��"���&c���z���D;���x���+˺|.�S;�۳b������.aò�)1"����T����&����p6���aM�Qս���.��W�"�s�kj�����;��UW&"e�2��jҴh0x�8�����}UԅnƷl��������;��-��"?* H��}�ޚ�JH.�s\F
d�g�١=i�	.��(�֚�7㱫�i���r�� ��j�8�k�i0(X~rR�̿�:p�vu��pŅM�|Q��9F?���$���v��a"),R�&�C��(/�K�n�T(�J�[i�HÃ-{[.��ŉ��TM"�,![���g�b��jir��Ոs�;O��_�e�76ӳ�J��1]*�t�e�*�h�µ.'^S����.8v4�:�8e�	�!^P&�����t3�^�Gl�|;>�˪���PF@�1��C�ɟ����R��W�s�O�_��Y�+a��u�Z^#�pQ��%�>w��	�kG���\o�Ur+��p�K�JJW�/i��Ϝ�|�l�]�o�֭Ix/�bb��Oo���}Bx�)� ��9�.��a&1M�嫒& �0�l�����5��Q
�|H��Z�Zl�E|a ����=:�<�M<[ڌkT�S����ຘ�T��(�����+O�4(Z��t��	�����C���1"�^T�V��j����	�3-)=6���'le�~I�E�4��NI+�q��F���*s��h<�C��<�x����j�PV��,�����A�#ou��d��'�Pu�d6��f�YFR�_Ŷ撯U( P�<Q��cg�lݲ7��޴S붉���1c���O�������s�aj_�d'o���0DmK��FHfQ��řEF��2�4�+�
4�eP���d@ ������Ld�(s#Ht�`���&w��Y�>�#6ǕA����i*�����c�d]s~ F��4���곕!�ђ��E,D�&$7�����MP/̄�xHl}�X�fu�Ba��>�dֳ��.GX�����$����e�U�n9R؎�+�q��/}͋NSX(+W�k�u=:�[3�ѵ6�}ky�(�t�q^%���`���b:���NJ��ˋ��$��F�ئ������s���8��Ar6�KY��Ow s�����L����Ԝ���}���;g���O�:5��;�\�,f׍�swN?�g�i�蜓4�����C�vj�x�q�������=gޔ�����Lx�o���@��'Gjz��a�䴿-�D���$I~#�$|X���c��.���Fӕ*��;]�K��O��(@cm�*s��ź�H0\d�\Dj����E`и꽣�RI0�H�
����r�10���Q)w-hs����Y� S����L��%Z:�0*�"�
��m�ů�M�.!(�K�\Ї�r��Fm���<	�h�1��A�GF��7Y�A��d��)�Z-��*�)n�l���|��S�-c�a�HF�S�Y�KsØ�$a�g,�ї�U����� 4$ c�}p׉��g�@\�(I?k�/ӱ&��R����y�(��ƴuF��5p`�����f��|�.���{r+�>�|`k���6z�_�����Z �F�,L�i��3�ٌ�9��@�ݻ��MG�;$q�٭?��#1�_?�\"=��w��q�q�ã����>ڻ�0�l��z@�O�lG�c�a9��%V�iBC�1��PdA�����\xJ��@#	1.��R��w���|��7Mx�Ԕ����L{T �R ��HՆX��I(�Cyq��o�,�lDB�P�<�,!#>�u�:�(P��_n.�B�w8���4�4��n?k��D3�?:�yJ� �x�Q��v��d}�^{�qT|<f�Z��N+�W����F2K)ϧh��d�>Ue|}�� )ANZ6r��]4/���	B�Y`8'mL���e��P{i����*A �i�1�]�<����P�����:ʉ����V*ksn����6�2�L�)*�%e�X�<��F�J�U�d�lzDY���?��0���s�+�̬:�b������g$�����/tq2���:�Q���-����5)3.Cu+؂g®*a�w�x֍O�V:����/*�V-@�X�V���S���)m l���.^����QHC?���z�������+8�u�.��
��_Q�#��u�D�J$B#�B�x$8�#Y�����K��$t�
�]�f���4�s�|�D۽�[��\ETd
��2�=�~���<���"{�d�hr^��QjQ�a��`����WN�ε���}T#�3{���"���f�fS@kњ-�i_���ݷ�e�U�\��'�yY��<%�����u�@����==�+�<p�Y���zv��㌴�����/Hh1��~xi�.�z0٘s�}��Fd���G%�U��9�fM����Μ;����,��0baI��2��9��G8���@�<>�Q�B���x-p@��������=GS.[Z�׀��5��m���Va��x>��+��$�}�1׍<��cBѲ�,���5H(�9�bܤ#O;�S(Z��Jn�� �%���/�3"k�c�{\�.
�d�
���]N���Ft�)Yo�xֿ0M�٣x���A�D8�r��ʿ�W���r�kZ�����5��c���Vv4$�R�+�h�Wڧ�?�����%�������W't)���c��_��].�M���LH=L*���v�J���R��3�4�z��d��|��QN�̱�~�8� ��Z�3����C�=M%��m�RI�R��i�Y=��Y�,��9Ɯ\L2�v!42
�E��=��ģ����E���pok"�0�@ɬ���^T���m�~5���m���OM�>�S[��\<��qI�lZx�N�$w���zWD~����;�f�a��o޶��6��0��wV��\�l�x�J�"k�5����'��!T؋�_�����X��N�[
�+f�����5R��@��i���-\!�����&�OLH&�<o�ˁ�kT�������j����D�yT��)F�!�g�s��˃�@�q�F���F�����Yn��H��H��DA��Ԛׯ�.;��z�g!�S�)���&�����^�]��$�˩��
Rͭ�e��~$y�i#�M��45TW/o[J!O���)Q_:8Cq9�����SV��ˏH�t�:���{J�4�V�d^e< ���<pq4f]ƄJE�i猊�?Wa�.D��|�$k�e�	_��B�$;o��X�q ٲ���7[�'T;-O���mj� �����L�����q�����%h��%�4c�KY�:eh2u�GB�LU@�+�o�.�@�XgY�`6k��sG���8>�I(��� ��i���Ip.'z���47C�A�ڙ���HE��*�3[z�U}m�'����岻Q蝟�<����颔SN��X_]-��KqWV�S��rv��Lg��D]��u��w��w!�V@�$���y��7+��-;m�8v3�4~��Ļd�X����y~�V�|���5X��B˩���V�֝�/f���9�'�/yz��I��N�;2;[fs���@�1�^���E<yh¨�i����:Ү���a��)��jz�2�&�>�J���N�h���bQ���(3iL�a*��q�-�N*g]q���s��� L�Pj�O����%-���:G\
���)h��27Ws0w��6�Z)�+�f�2ֽ�t�v�a?-0X�kȦ���Y�V�q륢��x(�o5��6 Z��L�5�;���G齺���0�)p��t:R�E�2D�ι̂::�/2�/r�uAt�@�9�}��vW�b٤�BD;����t���O�ȈZz����=L5��(C�>ԧ��+@`�.u?Kqu���=c�m�K[�𛃏1�ل�y3T���+|y�.�\i?�w��?�������X.����4~X��m+3QMP�i{W�%�����d���,̡�9��P��pԎ�sx2a�7�B���t�n
d��x/�k��i-��:�1xL��E?�����M����$] B�����E�r�?�d2����a۞:�����s�*��W'uʠy��� @�Ϫ��e�٘�lf�e��{��H�؟h�Mȿtୃlǚ��+���6�R�O��Vm S��q���rV���M����k���`4
w��p4�������N֔��m�3b_V7��Gb9pZ|�c���jd�f�����OZ%� �$�*�zk�#�J�.�,RlO��>��c��M���zt2M�A]�,Z'2[S�X�������V�.}�Ā)���G�����n�6�l<Q��nc�P��E)'�L�B	U=Sl�tX �Pa,�(R�N8�YQV�o5i�w�BS���,����h2��W����NG��&�T�46�u���罸�9�Ҩ�gGХe�=$���3У���d����h^������F���4Ұ���T��S��oSCxwDV���_`׼��{���>��]Z���yG�qo\4b���=p	��(\���֜�`�f�U���=9'�-R���eZ����CooR"�P�(��vi�
 ��Z�wg�1�o�Kf�7'P&��+m��n=�ȱ'�4�����ʽYY����G�7_�iSw�>?܌TKR�z߰@	��?��sa�޻I8�1�d7��W��u�ŇXcċ� �b3�-�	~Q���+�#�¹��}>,���tB��x��5�=S�����3�"Ԟ0R�g�]�����0<C.��*�'vG�0&3�1t4%=�4I��h�%x���K���cM�>��ƃ.j�}xZs�h\��PC�������!2���G�]Ħ�l��iv8! O����m_�A�7�k��s���b���u�Q��K�ℵ��X��j�K���L�)շ�A�2��S!�:I�u���U���	���3�Q�(4��4M��B��(���^��>ƪ��Aaǡ��>w�GډQ�#0k����Z��������r��懯����ﶳ�YpÍK�	./=9+W����>����s=�>#H���ԭ�������[3+�ɡ�JE,�#Yd<Se��p�G`4]��̜����Z+�%Ŋw2<��Q1�[��T��s���u@e�5ʵ��˙�_�4�4�[�S��:���=��+��D:jѪ�w}x�²�� �<ęH��#@�~�'���#׌����P��^�6)�'Z �l��Nے���ۮ�"�6�>u�w��R�3�����"�wP�堣S��j� ފ͌�F���5e�
��N���r��V�n�[8,�����+`�$��&v�=o�7]UHY:�иY'�P����Z(�ֻ����Y��jv�-��%oq�t�D��|8�Э�_�F��&��iq�.�����y)z��7��>�ۚ+�� ���&W�
5���N����Ɵ1�����1�h�î�O�fy"�[a�G �*Ȱ��-�Q��C ��S���:�	ֺ�=rzg�g"���SQh�A���2p5��|�6V%f�:w�Z�5�K����/,78,,�
-.��mZ���K(�����f�r�S2��|:�k�`�vV��B��2_���U>բ���}�1Y^�u���K3�wv�}0\\��%#���{�ex.����q�283�E��s�T�mI�G423v���c�o�C�p'�Q��+��agt�kApy?I]��AI����|��­�@�ȜSЙ�ڂV^�� ն6�p�Ϯ�f����3?�'��}]�Hgj�m�]��Z��m;�?�=�Hodf�?6` ����!m/i`N���<�/X@�yJ�#6ce�$��k�0Y|P����vd���rmre0����ݐ����y>=��Q˲�Q�!�
P/�:}߾\N�Fp�%��+��Ir���C<�q��k�f���1	;��Z��h�����A���d��>#��N�������a�������A"Q}CϽ8h�Ֆ���b�� �Z�Q;nB�����1��X��ִ1ǑS�@5�*r>z0"��Y��_� ����!l�-��a��Lj�1�oA�SE|�HUD���{�ٜC���Cv���2Gk�U �9V��
�m�I��p��������2B�yȎy^�H��o���@�7+��*�RI��,81�U�Q�Go�x�ݓR�� &q{��+��{3,�w�ɦ�$*�aN�VO	}(vBd����F#���NV�HöG'�>@btI�"I^���\��cC�ժ��8s�R�p�(���lk|yq���F��;ƹs�N���T����2L	��0�&k�U67���9]����L�!�Ś4��[D�c�ɕ��_k-z#�+%�]��:+Q8����ħ�}Ч��+��oK��x����$_DN�l}w��0�W�<r[��Cc(�;�����=AbH���W V��S}���Vlh�'~�O2��j����t�n<�aA�4��2�Q<��t8�f�a���cyR�(��Qh�$F����*��}��̝	�+����5�wm����KE)��$
=����Ck~��I$���(V�GJ#�k&ȟ���FX��|`�o�6F�%�g�Є1B����2I㐊o�{9�Zc&pI`���{�����l@��N[�9�M?	{���D��fl�������� �U��v�q�v٠�VT���8�Ӭo�"��ʉ4���)�>��Y��J��� 	���4LL!>�8"��Jt�RjB��r�彈m���Q8oX!��q���B��!�*_� �����u�u���y����֢;�y�Ҭ�bX<��(�4l�H��C�	/%Жxq�ɣl;���l~�N��>���*p+Scy��.����?wS
L������m�<�o��@���X���qm�Δ.�L�oi���z��+�-��ˎr�h�n4��?U��f��vc��_b�Cѭ�"�oۓp�xm�9IEh����<��2����A��
���w��l�0SM����`��	%�!���ܵ�Y��d;Y��gz�����~e�/��C2����)#s��mNTW��t���R_Xs���MX�a��"��u�0Du��I>�
)�nn)h�ǡY���;�ۀ࿺ۅ�q��Z��^�i�4���gP� �&��ro�A�<?TWK6ڔ��i���~� L빡׾�&�n�&����
�К>)g�d�v�w�����=�D��W�0�����Fqx"wl�8��Oل��ua����	*.`��}�Զ��⸿a��8vi�����*�^�15莢Bfdw�M�$սhEK{��c),���-��:=ۉ�*��.����z()�}<RK��1T�V�����nJx�d=��o��\��b���9Ѝ��5SK�'�0*Y3�	��9��G�S����H	��oTb�V�=FD�L^2��/5 ړ�Ya���"�6lsdvڑ3��^��sdw�ٺ�k���)��q?���}|ES��K�U��5���n��>W��؉�JչV��͏=<%�+�I�I��e�)�v&1�"��c-���[�F���?�r**��e�1v1��SC������2̪��xc
��� 2�2p�n�7�^�/a/Na�\����l��"l��h�K#�*������'5;yP7?G\-q��L$��Y�J��_�\5�}و�����lN���$49D#�tDa�Œ�����P�1�R(G�c�ǖ�7;�<,���C���͔?���^oŢ�������F������N�w� �f�Jc.�rœ;��N����c�^o�P�`I��=6�}%�ԛ��.l��GR��5���y��JRep��W��@��D���I��q���j�xU۾�((�FԺ��Ug�>Yy�t�Ճ��+jo)��L�e�3}�N����5�<< ���k/I�ܚ�\�n���U$M�(��r$��v��ĺ��������\�k�E���eDq���I8�~���̐fo�K]�i��أ6�K�t���i��i=���U==؀��$�̷B������7�u��I`P^y'v��_�$}�;�)}�d&\�
3KXW�݀�d��@<z#pˉ�d��K�9!�d\��m������S���Y�F�C|&��fp"���搳5�nL�9훑J�Qb��\;�]9fօOn�\�sX�^#
~8����+J�n�$�L���Pѵ��_P��m1�U}*)��8X�L+�J;�@)�vTa�K��2��N�{�Iv�H�@/����~1�/�n��j*įƾ�׺f٪�xńmp�O�d�$�\S�s]�Y�[��Y �iN1t���T�mZ+�iδ�Z0�r�(t��E�]�)�.�ȭ���N�ѱfH�}Ti�L2su���3��&�/cgu����q�	�A�5O�y�oS����5ʋ%�W�{�%A�#.�c2q����~B�X1j�_��ssþ�+G
�tĢ^C��Ԧ8vz��x/G6�Ȅ�:\p&��(���ë�g�����Q*�s��r1E¶����I� _6D�mĤ�PLlXc�Iw�9۶�� �@�o�q�h�d�Z@��%.d�g�xAK!�O�&o�i�>F h9�*�#����H��m����wuh����|&w�E~�Pǀ�XH:��������/M�'j±)c3����\&�t�q֊�i/� J��c�����ê���m��3Z�ƚӶ.Br֡✞�4�����(P����f�{16ob�1M�֚a�'�Z3�#�lz��Nr��0����Q��*di  ��Ԝ�z^��*�֡�CUM���^Ӣ���.�Tn���j�����\'atÚ�%���{��o���ꇇ���L�P� �Ig��5x�C�G��?��S�e�V�:�P���7%cn�~�)��fKkPɞ��H���w�[+yU�������&��9���zt
�f�P}hf��@�P��T�7X�.s��;��G�l��C�8xvR���rZ1Zε�S���LMʪq�ڿ�5;��~u~Tb��M���M*�$r��D`4�š�Υ���,~�2 rM'\I����sw_�"�ES<nH�}EiBҖ�wʘB�'5�� ��G�� yXC@#.}�v��D���=E�@G}r箬cu���lM�.qV�/�K�L���pC0k�Q�w���?�_q�n����x=��^1�w^K��`�sx,��:%ͧ��t�R]8ۡ��ngۿ:P� L��ʷ!�)��Q�9�Al�>
�͇Cٚm+nh���wC���*������͘kX.t�Іx���<� 1�QfO{n�^q����
1�V�&���[�Q�o�E�d�MM�&U'��͵��P!+�i�'z�K}��4z]�Z��,�(����m�y���l�8��P]��M�A��	���؜4$��e,��cow?���ܝ���H�w�����2����.�䴨8��(� c.G9f%���Yv����x�F��p�5�����4���&,�KC���QK���*/��vQ_:ӬFz�שB�!4�����u�4��`J������+�>A:��_��
�<ij���4�Z�F�_��d=�9f�_�,�XA%S#�����#� C��X�����r��xbˡ�N�������s�U��e;ݓ���ښ��m>0#*����
^�E��;u&Da�R��KŶi,N.�U�,%�5Ö'�.�sKz^ô6v?�` �t=Dd�.�R���-�d�*Gs'�	M�.w��Ig"j6�q��
>1q����¸^�T.y����XAX��ۄ� �Ir�R�L�~�3}���vߖg���qhĐ��H�l�h�{:�(�y��Zf���7)��.��<�>x����}�����}(�j lZ0$��1��|b�_1�T����B�r,�d>�b�tk��V�d���#