��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K�P��9z�7a�U,?�y�"{�Rm�6�¼�L��H�Wl:�j��.����u@X�����b]7u��~V������[Kv�@ъ4gB�䩯ڴO����LHvUmw��[ї:�⻛`CC��;�����@L46�M�p!��ߝu�Mw�{����{���z�԰�;��^m���z
jis)"V�x����}$�W/�\ʜ�t�|��AF��`Dq%w�hTPxXH?VL�8�:�PY_��9��O�;@���0�L�]�D�U�[���P;Y�����K��	� <�k�v�l+��v��j��Ar��R�i�D�v+2�K���`�
`Y��ʝ+���u~2~k���_�?��Z����%��$�`Z,BHz��KiV�=�s�����T9F�,�JL�}�!R��!��W߳2�Z�5���\5>̲��Q1��}*:2����#&�}����XU�ߡ�8@��P�2�������Qz},�Kz�5�WW����v>� {@�Y|�Y�;b��c&7�_�oKwq_OA�����oR�k�8^DEci�#V���Dk�d��Ń�9�k�N�~�8��"�-#����Nˑn�-YPHcb������V��)�[��o��"8`H�_�@܌r8.��_|�;������>�t�b���0�2-�,�-��Ju�A)������n`��4��9l�\�S�8"�w����CR7��نG��������Տ��ѠP?쏅%���g��{� �L���I���+͖�a��.��f���:���_~ �ˬ�+/ӣ@qq������^���RD�FM{3�t}v�vZK��A�,�\����OF�C��ӝ�yc�B���~���}G�G��[��G,�x�Ҡ�8�a>w�cak��&:Dk�<�F��e�J��/b�E�:&��� �A����9-���v�2`�!6�sD�7��Cm|Z�|�Ia$�����%�撻�^��_N~���4#oQ�e��Ɏo�qx-]6i���*��r������v��^y)S"{���S�= c(1�7�n�ֱ�6q��Ra�8��Z��>��G@���y��O��`�4�/j��	�a@�C�!M�����^0��R����X������P�����Id8��zC��dZ�̼bEfC8�Rܔ;C��*Ƶ��I<���j�����!���lHj��H�X
�O9����n��{���g�d�b��W���"+�s�B)�T��fSm1z��j]%�1�>��Ek��� �P!�6�ayD���;sH���l+:q�po����+�`ҬWap��u�uH��|��.I��M��C��N�
�i�X�'�97�~�:7/�(z����ޓ�U�6�rg��(��
Kl{����y����a�@��y�@����|�f���Lj���)�G�I62�q��d��S>u��'fa�=¤�8�B!@�\�T��7 
�`zf�d�7T.���J���3p�4��;i��yc���W�ɐ�������:|��jc���"��Akg�{�a��t�z��K���E�NRq���y�7]D�p���,�sR�~"����ߺ�Z�J4���Y�L����LpG����tH7VOG��� IЊ%����&bC���VX	�Ek�b�~^a�FJ͉�n;���N>o�(�s��exҲںmU|�K�n�����MT�F�?K�?bAI����bM�5,Ƈ	�7��`i}��WĹR��c�h��$�.)(;I�ل޸j�@\����&�� �.#��'Pb ��(�|cmkF�?�&ƅq{��
��}��ĖS//j���g>������?��|q�j�����s�����@�3Z�5�v�kS0���e��Ml�>)y"�:Ah�YV�T�%*��v�JG���0r���m�;��0Ax�)�lV�BK$e��a�T���Z���f�PU�8��*�VU&뮧�~����I���nP����r%)�R����mI����,+��#>/�y;�h�/&j�/���Xl�&���A�Đx_8��`,BL����KtS�=�Jj?�Ëc�!�S��]�y�+�)��r��͞�B�Q"|H8V0r���x� >ZB��NJ��8�?�熵VhM8��uf7K�A�>D�,����oj�zPA�a���X�Tm|1�����b{濆V����T�"v��k+����c*�؍�wk�'���d�5l��	sln"��S�-�;9�(�E���H-���B6R�R}ӄMn���x�}���f�䜩����l��}= P��S����sB���c��{1|�/�G�ĔZJ����W�Ц���s�u*"[Kw])��̝��#���DYt_�1�/^�%�"�>��|*%��5O����R���a�5Ÿs�ڞ��,>��-B1�Yv��.��WU�Jn��\\[�i)
�������[oQ3tk"'�ϗu�!9�)���UT�Mm����U�mih�?�D���籔bO������:�����6Qj�����X!H���f7UW������OO��O����C��q}��Ǽ��ް�C&Wj�c�;��O�?·$4�6�(4axPk�|;r��l2 V�zE���b� ~�O��<����^�乣�[�m���H��2Dн��ѫ*��IMw���ݥ��mr�T��t��9��B���z�m�~�)W�ߵ��~GR44�%�'�Q�U�?��w^+w_
��L̘`ż�3S�c:RGiiw�
�;L�%d�Ӓh�O�����m����	�"�2��~���2�.�̻�͐�ݯ�Ue>�	�L��#�[;ձe��G�.���b<H1�����R�T �����o3��rG�5#"��VE�a��%L]M����ꮚN�hn}=1��q+}��,���P�Z�=����s`[�ƃ��G΢���R�Q�l��39� ݎ�����2�G%(+����Q�X�4˦���,,@S �>���C��)˾v���%��]�cQ�ch���f�<m	0�����7 
IJ�F/z�6��U�7w�b."�W3_,���՞�j^����zy�G�a��J����s	�u�Y���; �g������#�!wՇ�G���r��n~˞�P�����'(��s�!G-W2;�ο�+"�?Nڅ��
�y{|DG'~w�ܜ���T^����K���Hz��ۣ5��Ib�r��_�Ům�[��D�֐H�-��w�̩g!�b���3�AL�6���ځ��Y"�Ѥ�Z,� s�-�%�k�#<G����*;"V��{h� ]��܄7������>���G��
|���5���j���)s��i��[��a��I��S����x��L,,��>�[l)��*���R�5N����y�2��κ�����M�N|!D�L�j6��mW�X��b1�\'����U�	�9����x��"[���5�ղw�\L�����'���������������%�*<!
jS�mZ���żXR���N�k�xv�f�Y��9����˵��A�*�s
�.o[3˙�g�L�?���*���d��U;�����f�شv��Z��gU'R[�7��. ���e	ۦg�b� *��l&_i*�u�X����F6{�-M��ץC�d�%7X_x=8~]6����^��'�Z��Z�	�<z[�3+E�����'���������H-JԇE�R���D�6���;��:�n��cA�0.ǹ��n�G��w��I�+�&��xx1:=�0�ZŎ�k���ō��bņ�oDD�����_�N�85��ꕈGf��S�Z���J*�c۪o�Zr��e��D\@)=Y?��Y��z���Bɚ�5�|��>����^Z`��>�h��)��H[|����	s�Ȗ ����&�X�U�!�%1`�Fg�ߐ���M�����Q���'�I쬻"��<��Qr�1�����BiJ;��T�.�r+ ��$�E�L�V���xW��֍oZ��$���+�ր�G��c�zN�AA!�����P�Y�&��U�e�T<�t��4IQb�Ro8�2�svn�	cWU�=I��'+W��cos���;��a����f�B'���Ĺ��Z�"2��.L�@��ԉ{�l���T�7F�+�Ck��_�����Q���+#��J�02ż�$�Hc�@�Sb�(`��֔ZRif2`��+���8�b<`H1�}��먙��./nQ��ZAbV�md
kί1�C����0�`V��S�
=j�.���ap�dD�9-���d����?.����V���˗S+��P�?�cVt�/K �#Ԛ�	QF��o6�碢T�<����ӡ�VȦ��f�-=]�5�Ӧ�ӆT�ͩ\�[�S�x��+
Okݩ�ȥ|~�W��`~�4���������gaqf�6t�Ȫ{���LJ��;�f��B���sC�/�?`u��i7!gn�')��5s�����g(�[9�-��;|�ζ�o�+��f�L}���:�F3'>��e�e����y� �}�N��Z��Z��D��{��[���ɺ� \��� �"�6#�E�р�L@ݺ�P���k��e�aj;�6�j~�b�x�`㤝�іE�N��>⑟�G4G����ɘ�ˋ���VMd2�����!�m�¢��B���f�8j�1�ɕs�6���{l��%5��BCmV
��;ep|�>6���_z8p)/�L�(d�L�sP����y����J,e����(�y<h^
��)ug>���d4�ֽ���HY�"D��8��ٹ�����0�i���
�uP#N-)*=�G�'��U� �&+�P���s@j�p?q���АX��7KLw����!q� ��h��u�VN�uiʕ��tb�X� .e�Y�S�B�|�Cm5���`KѴ������u6>��P�F����v��B'�i������⡨c:� Bo�����V
���*>���%��of��'�̂"���\�u�hn��C���(�M?�W�m���Ɯ{<�c6�l�k�.]����ħ=f�E�QIx�U�����S=��*iD��52+o&��qj�;	�YRȓ�-�fY}|�J��l��C&��Q1���xd�4e"�@��o+d��и�[tm��fgr&K�)����ÁH��s���[��QV�Ä�ǰ;ؙ�D_���+ .Q�H����G���UJ��3�u�;�,`nPVG��	54%3H�j@y�}�e$jȿ��:��O�{�!\�r�l�mT��{�Ve�,����D�J��ߠ&�����'�T)������t���Ws���=�>� ���j�����}�"-l8�0�p����@[c0�E@"q�=͍$�^��^���f"�W�z�q�'�%{�Qg�h6O2���^b��՝6����r�Y���>J(,�wD�+�\��c����DI�m]�[ڹ���U����B�Aa�-a�q��Tԧδ��~	1a���dތ�S����#d A������'������u�����D�i�K �)�l$��x^���3uF�"#�p��[��C}�%�"��-���߱B��ܳ��t�"�g��R���)�;�v;���Z}-�*�_]�=Դ[-�Ȥ���e9΋��N���X�'�x�oO�~�yGؼ���3�(��/|�t2ÇI���)��ı��Ey2=j����x۝���\Ο/�mW���{0����lֺ��-�@�l{r*Uf��r/��X��=��,�C��:M[:�c�s�yR��ly;O�9�%c��ҟİ��=l���$��Ӥ|%G��r��5�*�D�[UkU0��H�?����*����/�����.��>xq$��h	E�Br��?�6_��+}�/�[�턷�bҽ����f�M���ބ�~r�a�rHU��8��z����K7>���������fYΙ�Z�Ӻo�C�Hh���nf8��Y�sgV�(�=��N�ve�3�TQ�ٻ0�8#�>t��ە���j0�2/������im�t>��d��O�����5L (!X��L�i��r�;X�\K�3�>LaT'$�����>,ǛaX��Fڠ�x��%�	X���zf�����i����EJ\�Ԛ�=� T�?)bǲ.�?#M�A[�$�?�S�2����웜���A�t���#��y�%�(�|�g���&T~��Jk�t�0�M���w)_4�"ɣ.3\�n�6�es�Td��Fw"�Lw� U�����9]����d8q�`݈�rt�K�V��?�O���R�P�RJ��+����yKӾE�,�sZ�7�d[��a?�{}�����q&h��
D�&�*��z�c-6f�=k��|�D��l,M^2	��(rp&�Ā-��d7�E�I�����l���Gc��i��7���mH-���V�	nvj%�*�$.p�ȑ-���u�8���� ��(�G�����pľA���`@m j���x��N9�ŵP�H_-I����(�s�OGVw��rI����-&<���Q�0xeX��w����o�J'f�P��diY\Cspqt.KJߺ��J2Iδ�q)����,'��R�f,��f�9l���B�b5&����Sr��FKb-x^��"����O�=�=�()b0��N�(�{�EJ�g��jK.��u��f�:�gH�P�ȝ��w�P>��R߭p��T�����g¢:h�zk>v<����ESy����lֿ8�h��э��i��#���$j[!���yS��w�-"�`��l�V���ï���?������Z��ՉfDKT�t:�ώ��d9eyY�r�m�#��4d� ���E72�4M'���IUt�ǣN�� jK,mg�Do��ױZ\{�f�P�U[�"�l�ۯ-�(�P���1j���� �/���dP�������� }�vF��@���r$P.�g!� 17�Me��`i���nm]Ʋ>X|�||S��p@��^��ѐ�# Zb�Ss��3�&����DP���m)����3 2M��C�K�qO�c�؍Y���U�8�U�N�z�&�P���+�`{�-ӧ���RӚp����L��C:�G��K�@��U}6eO�T��� �KgVD�M��9x�L��S�8���ZC��G)wA9��@j����P�[���`dOH�A>�
��ÒJ���St�$�W����(��P�=0?�%���뙀,�D�s��E�i!�ʍ��Q�em��M%��/>0�2���uf�����7���3�C�L�E���`X�u��U�+GY�����S�Hc�l�]bw�l6�@��*r�������Z:>��H�'i�Q���DJ��a�Ϋ����%\R5#������Y�!�a	�#�n�0m`����*&P���
~���y-*�F�=X�oyA��6!0���2��� 8��>��]�_%ߨ)��;�+ي~�~3D����@-2�w���z+��x�X����e��޼��M�y3]�v�t�a�����%����}N�*����l��w���k�R���V�]YB:p���b/G�+3��|�7��eaZ�Xvx��!`���K�P�H*?��#-S�ֳ�O(B�k�#̴�^��@p�pEN�~�c@����1g��{H����u-	�T1�z�2l�*%�Ter��m���iL`���5�VA��-�/5�q�K�p(�=S�tU�U��כ���c��7
�Ah՜E��R~��`\FH�An|Q��{�}ݥ!+K��R���r*�s��c��^��X�M��˚����"�>p��J$����ܾ�h�#�"��ϳ�gMMd$V���x��+�����Q�VA��i�(j��S*�49p�����H�}��1Z*L��F�La�!jP3�҉���Q׃��9DJ��NA�]�,^i�+!�A��z��C�E�H	�Q���gk����K�!��8�l_�`�q�	/��i"J��e^zT�U��}6:2���*e���>.��'�úԗY���¢��++__������XA}Ѽ>����p6����K��/���Ӿ�Q����;k��7�!%����`e,�,���d��!y��V�X_Iu�(Yml�Gю5Xx�c|�,�i)��)^����T����x�mĲ���R!l�_�2�v��c�|�Rp��ʀ5;V�}�~d	o������K�A"b��4��>$��Ӟ�����N�u�B� +{i��C!���X%&�W�೾$+�>���l8�l��r]�g����kɒ�����/;X����(����w�Y�
;�%ef���p��#
L��{:3����&,;M('7\D���y�8��dv�D:T-M�@?����;Hk�A����H���{T�
m|���8���"T?�1�=��nfd�Z�)���a����rU2�.e��.c���J�I��p�����%�)ϊ��䥐fR}���T?Ɣj;�j�↰�!O�h�P�<k'�S������fu��:���P�T誖�S��X��hiv�Ef�`�d���Z��t�,8����%3�g�OkX��3�Gr;̈́�R�*jc�A]����m��a���)��5�v���岦�\���X�%�	������Lx@A��:�\���~�V���^ }�Z��̤���^$��h����.�ZQ<�"2�D�����K�<��fLj��)��G(N{y�O��	�N1%t^X^�gT�rR�m �=|��ڠ#}������,�߲�O\��!n0�����^\�͘��#Ɔ:|��0�H��;3u��iq�+���үn��Uϑ���,Ko��ڗ�x��*������R¡W��u����@�)9֪k��2������XvԒ�A��޺�����t��2|�큹|��z�I3Ȝ=��S��+h�:|fЫ�7�D�֥Pmϲݖd˸��6\�8�{�z]3�L�r�Sqg]>�A|�+�����E>X�q�>�z�\�X>���%b��7�v�:!�uŎS?|�(n8�0��D�H��w��g�����)0�D�d��7���Y�bD��l��bv���Z0�9�X�(de&P�u����� "Ztb�{�d>AY��u�D�:p>�^��f���|��WY4ʵ� �%���c���Wr�ja�D����k�L{��������pT0�y
u�בֿ��6͒���($��g�DVC_v�t(v+N�ʏ�2��Q���-!2ˣd:)��9�9F���,��ts�:>硻�!�ɕo<A�,�d]FiX�M�(�)o�)�v�_P���z�/��Y�4l��	�&��-[���UR��x$.K���ʿr��/�U,�X'1��,���\N��zֆ�=�uh���+B7��[�I {�2|z2�-�Mk�e]d:�ԁ�>TP��M��+2��Ly@!+�5��ԲO�8�& �΂q�d�Wru��L)>ߺ|M�;��L�"�r���W�U8N�/����Q(��p���ŏ���f��ۀ��F d5��F�dϕ�[��hFz��Dn&Y����;_����At�=�7\
њ�]�w9$��H�sy�*���W�Ã���;�u!z��m�����6G�t���7����z$��=���3C��˵+?���o��>�Z�v[ژ�!����������-�)��3� ��{1]:
8�0�`E�H~^{���3�	}����{���t�>�yF�jl�b�
m���:`[����u[�B�Wd)# ��;e�����:���"m�M3�ې�l[ �N&Y�i�������b�A+PFs��e���x"9���KP�<���Q���6V?�����ph�۴a}Hv�y�p���ڳ�ܒ�P��Qs�Vt�x#�hGb�N�S���.&̯QE�g�u�<׈u�vd�^L��$Va�r��BV���#�h�]!��V�g��
rUe��Z�(��ך	���]���ֈ�䀺$1��4���[J�$�D$�<�&��i+�8�(�&��W���}��\%��4D�}W��N?��Yv�iG��u�	��HY�g�2WQ߱$���� �K1`>�f�Fc��
�6	� W�-�V��C	�3�bX,��0Y.��9�F���_�� �Q�@�ؗ��xÜ����X���G���v�8a���EݯHc1�iψ�$��ťQe����~B@d������������_e��Rx�?2��=��xɕ����sX4;�5Ԓ��qw�p3�#d[��~	n.a�b)��@qaB�x�@��8hiulP�x��
��W	_��TG8y\���@p�Y��W(�^L�Y���7(.����g;:�k[K�"�ޭ�r�g���K��òbgv�������ճWq�_�x�[�@F"qT`'K�(���ǻln�<�ޅ�j� #�qm����,R��Cٯ*$6����㷗�C<�Y�JFӅ>�(ή J�s**�sbe�K&B9��$��L}�R:�rS���O>P'�j;'�1@ʖ��S2�y��&�׃ eš�.��[���CU�@[�2K�fZ�	�q�>A��H� �I�?̻@/��\Q#�CԘq�L��k�n��m�J���D��1z���Ͳ9�
�=0��[�?)!Z��C�������}˳Ez]"�����HK��Yq-�,�=�'�^0�8����T�{�[���k��0h�Q��Qa7�oO�<�!`۞+HCgY�B�JnK'A�/;�3>�ZӋB���� }�;_bA#�����f�Y8������q��~��	>������^E��'��0�2��j��A.D�1�%w����<��)�Ix��G�_~��EC�m�R���on�$�@C�ZB�^�SL!Ո�|�I��\!YH��]��d8@�<�K�T�?��>�G�+s��P�`����K��g��� lMm�SX���C���M|���4A�Ϣ��;?mѩK��6�6 B�m0��ӆ������p�;Eן��ޠ @X݂�u_��=�EʩES�ΒV:��.g�E+OEw�laށ�K��Ei�ΗM�'��IA��,���M�1�)ade����/�mvcD_l�M���]}�͸�W�Xz�����'n{]�qe��o"�rW�y�Gt�2���\M�T�G��Z��[����\�bǠܼ�K�/��R�C���@����G��n��<vfx��~�'9���گ�������h���M��b|��[h�w�7�E�^�ri��|jJ��ᬋ�Fu��P�0��p�v��R���pώi	����Ɛ��s����r�|��~��>��	�"4�/�k,_G���j�
ۼsőHqy�m�dm�btv�f{�WX�\�a��[��%br����(b��4�����]p��M��
Әs�� u�$���ۑ�6�������H