��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$�ʵG�_2��:!�Bz���}��f������Qn����l��YɆ�Fw��ڹ�[��>�2��o�w
��p�S��<�&8x�'�i�LZ:	�����������R������!�L�r�Cs�noOtF~�*P@�v_-�#�q�㯨�n��_�wL�7�p�>Z�X放��*������b����y4fD+o�
�9Una괐Q5;$����`��j�+F1���'�p⌮p���E�sA� íf�ol�s�#f�qa�e�Гw��iA��>����ݘ;��q��?�:oj����)���J��d�:�b��T%&?�*�.a�
���&FTz!L�ؕ��c��L!T�uRde�!XS�;L&o: D.�lVb�i����\����,D�Pe�o�;&/}�7_k��+I�Hp��ڻ{\8<9n�����No�������ۧ�)�@d�!�X��%H�1�u�
+�0�v6i���%Z��!:��7�RI�}��y�<�A�I��K� uz��tI�U����'sg�s�?���V�.��F�G�1��6ɜ(W�BN�\��)5g2i�K��J#�0�BJ�e�>#������&:𨄤R����+	���@�3�����h�2H@�,�}�H�o_?b���*�i�D�볇�2�2y�'��C��:؇F���$%�+��50��d�d��q���a'Ĉ�DH �}��oL&'\Kܽd�a�UIu
�+c'M�,��S�^�աI����P�BC$�VC����"|49���.7�
wi���ڐ/+�!u*�8��9�Y?�K������ȷ�e��y������N�}�R
#)��)���7_�\�>h4��Smr�Wiv{y3����z�2����
�7lW���9��Q��f���"�@��B:�u��vЪ�ih.�2x��z���L����L?Ҹ�d}�G�-h��+��F ���5c��V��u�o�2��̲n����:p�G�Bz$��!�5	 ���g���;Z�(f*.fU6:mNy�5sIv>d3�9�E\�5
^Uy���V�+#:�o�
%��]`Bo�Zi5�K'�I�]D����x�r���<:K+��(#��M�'9��S%]	���]���ϒ��W�p�"�G͂��Z;��S2nN�F-Л�������߄���,e��U�� �Vf�%GT���dhq#M�L�W~��}������v)P�R�a�0^������2��V���������u6~�N/J##!�:�����q� ���Ըw���ډ3B4Y]DH_�K�>�f4�K�����+JF N��x�홅|���(^ɉ<���4mW�
�q�'YW�aO/���;y��8����*��%i���k~d�F_Zz_��ծ+��	%_�]�Ui�TD�`])D�=��v�=�qSv�"c��M���p��FBnλ`��پA3�z�`ߝ�'�+�|���_aZPG�f�h{ܝ�Z?�8���:3ןޘ���d&��