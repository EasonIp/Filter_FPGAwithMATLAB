��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_ �c��2)�}ma�dظ��v}�b"@@�c�
l�bx���,���M�4A<�r���w�$�S߇��`w���~p�lV8���
��%�4�0Q�Hj������8�Wnwx�5|%�B4|y��<���C�bA��T�N���Ζ�:U���J�::��;��B��O����k�q��Q'�O"�h$ZrgtI���IB�Q��s��P=�=�F��Q�4d�mM���v�#��D����)0 G<��^� �_�\�y(����¬.��	�y�* ���Ob$�}h��@y��y���ѫ��A�".R�]�hڳ��2��}Έ:�g�wQ� ��)��E�w��V9w{cJ�d��(�	0b�9k�X�� mKٺf�רZ�[4D��<0p?���T�4)G��L[7[�4�l+-
X�tv{Z����N�8O��B�埑{�	"�=%����Q�FF��bi@7��J�5V��n��fo��; ���Cn��m�s`%s�*�+u+��p�m�|:��d�%Oʴg�6�A� i��8��tK�K@k�W��'��X�@�0���K?n{ץ4Ej����=��l�=
q̤��+'<�-AOU^uO�����h��E�!A�M�]������w�l��C�h�a+�����?���{��}e��_����9�O�н1���8����J����j�H�R��T��f��ڛ�.}��դe��;rJz~ل!���̽v�Q(����O�i:
I>{��d��Q��r�D~;�������wB� �����AP��rB`�\$�Bg�E��Xzy#0-IA~2���A�K6Q,��z������JX��	�����%ӟ�ݙL�?��f"S���s��w0�#�����;s����m��ܺ'EY[����/�qR���@&�FUdL�m��ֻh5�33��dc���/�\���v~`�}(G���#{�
��@/4�F� ,���{;��e,m>�!4�ⷤRL0OS<ޏH\v��Ů�i�4֜ˊ*�Ӣ<����[����"�@��Z���T�a� ���\�nQ����w�sߐS0 2�k|+Y��ǒ-��v\䪀�%�֍if��kwTh��p�=^��f�*��_z� WA^0-�5��4O:�����i��!,Q"{�#�K��h^n|ہ1|�s�$R����@%g6g-���@�-lFu@�v�pY�j��=��Q0�����\
����r_������D.j)��c%�}HʏLg����!�����DݎD7a˱�g(V�Imb��!&���7_#���U� �3G:���U��BRxp��	:q
*n�W�_� �F��xS�T��r��R�� �LH�e>���G�U�`z��'�.@��ý� �.��i��}�U)`�ŜqP&�(��7轕>�f�0��a[I��]�7ᅑG��s�g{&0	tf�H�GY[i���R=�0;�e��i+ڷW���^���u2d�8Kls��[1/�� ����AM��7 TuEv���G �e�|�|}&�"�Y�����}ݹ��c-��i�-_�2P�Yї�#43NJP�Ͽz&�#ޅ����H@x-�j�Z �+����j�,�?�F�r��ĤTM�%+�y��j@���zs���(iz60[��eìI1�Db�x���g �����kA6���^n��mI���u'<ӧBӎ�-�O�7�~t�lì�
��xL��! ,�]�mvy�L R���x�iMBZ���ԓ�,�R_�L������)�Dޥw������σ'J{<Ow)�5+�
J�� ��6��Z��5p�nuM��^���卜�
\�J4V�%q%���+�w�y��Y�P.+M.��2M~%�_����Dy8�DJ��sݢ�D�ӝ�1��o�Ry��5f�B�S���f��b��M:m?3%3��si}c%Z37;Jg/�����vf��T5�:��Ny=nSӥ�M<Vp�
ϭ�7
���H2 ړY�u�h?C;T�b/��Yo�8��=�K(��b�z7���� Ve�g�^�4��Zp�c�`���D�H����O��d��<�=e"!��&Q�[K���ɟwA�#��,߽�"<H4���j��<f#��l���Io�� S�N\+&���x�z]�鏕Y��AGݱ�0���|�et�lad�6����	Ppl�W�'����(2s����, t6����:��{^�K�(U�h�;.4S��$���l�� ����.[�UT�g��2�|ϻ4@j�����NER͆�,Yo
��7wwt��"���\�|����j�BF�>�:	YW﯌���ҹ)�m?��U-��JSI��DhYE�wS�9[v�hx��\1���J*�S�VA�U�<��#��ƣ��G~<��Ed��$x�b$���5ck¢�BI��l����1�e@u�{���F߉�@/ݙ��.����7���ȃA1Ee��V�g>��yz�'c��8��<��u�9���j����	I���/Dz8"�4R�^(�����j0�#)�YC��._��HM:<�Y����.;����SO"-^s̍��\�.�z`
/����[�Y�Y�_
�C�u^�[�'�c(ΪDs9���ԇ(�����`$�ݒD�;�Q��fu�ɨ<r�%DD�U��zaÆ91/���Ͻx;6�1��|z�����Ī)���L����i��J��n#� �l3v8T�D��t��_�r�Ĩ��g`	�0$��m2'g+S
J�{弗�ͨ�LK[Ӧ��&�bb�i�3�6�2i� #���⻁_�un���}���f���+|����	�&N�Xߜ��ޜn��V-^7/�h���[֣�\����#~����[��f�#�rG�N�F�&����mc��U�e	��c�?���qc0�D��%K�p�ҕ���Z,Ap����o�tY�h��y	�-9L�
>Q������Qt�xL�o���}�m4ݜi=?�5�^�6!�vZ�NL82幾j�d�/�W�EZxZ��.(������:�<�B:uMMr����&%4!�a�V'K`��=7�+�f-[�Ϙ)���2���YA���TǏ�<�u�`���MqT8xj�ym��4M��z�m���|�,��^��Zs���f͡�����"~����m_��uI2iX&AA�B��tz��>x�Dv�Bg��5��F���%��'3�p��Rzj�iH����O��١��p����K��d�A�V��k�Ľ!O��Я&�����VˌV��F3�Uh>T�7&�vl��{z����b��׵�{fS�6���Į5��{�1��Y=�n؈3`"�����U�]�rA�,G���0ɋCB�䗁�������
�@]���@Z)���G����.���ǂL��Q0�Du^>]ӟ�O�+5�6$������&H�2��h��}�4
\���3R�@���&+�N$i�Ca�hb���GGl'��A����#\Ml�8��d��t"���^�;�P#�\�x��q�sۺ����j�7�����^��2 �y�h�z�+���vQubp{ �>_��Q�K^}=�S��'�9f櫡=�B���
�̐�o�3&���n<���pǶ �W�[�Щ;}$�Ӿz�u�p�E�Tu���M�fW���.\���~�Z��N��e0�>�Pg�i��I���Jf������Q���7�����}�u�^nṙ�5�H)Ĳ���e9����%�]f؄�x�G��c/��Q�r��?�h
4�J$�P��v�^(����enxko>1��CS��p�vl���{���a�{�<H@�����~�CӘ�z��U��W6�^\}$Z���*�v��Ң�8�6�K�}�����^Z�$'�a���s�������c`9�۲����0���ŒD��Pi� 8��^�����r���(�I���J @�}l����D�5�!��8IG��Q�>l���]��?̈1>Is���O����WP�pċ|��t��D;�Zf����h�͖2�8��&��
��(���