��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��5K�z��!��[��S}Σ{$Gx^����c��ƀPfƆ����[��s�x�rQ+�, �i��7Ҏ�D�'�@U�(ve��}ڸ<���,~`�v�x
��G�2��S{	f����*����r��zʀF�S���p�h�n��9�<�yS1�m���GO�y?�xT��E��n�}?ռ-xW��U2�z�L�o�[ �6�@����<�L�>�i�I�♸��kI�X[�{��%�s��\�x8]w�����Rm��j.YZ���_*��bo�#~/�Vr
�yچ\v�!��ee4��h�}%��h���8��M:ڂ�^/<�b�T����W�9��MŊ����8wX!�w�/���xO4J3�z���큎K�����'b�X%��\���g�	w���T�{B&�ģ�oz�k���Lyth����t�ȦU~t�%��/4\�pɾM�آ<M�O�������3��xO�,dN��N�f��6��t���C���#�岎k�Zw(~PG\U���(�u��$�Srd=�Χ̨�Twв�$k���ն�~�:��V��@��!�v���}biX������j��.��$^�k��U},Z�4�Ԩ0�68p�(=��a)��`�'j�<i���"rV�
QsD��&�x���A�cO�a
�060�pV˄AXFz�l��R�&�Xv�}�^���#�cs�Ӑw��@p�.��a��N*��.%��FILT��r>O���z-�~F\+�>W�.�},�� ���1l٣y��;��!^��	�Nfg������%?;���Ĺ��O\�Ă�b�_t
N����K�AU�|�S�x�H�tc�,�	 �S�����	�	����U6�\��H�/���C��S��{m�v��0�b�r��M7���TE�K
���.e�f�1�ҡ�����_x��V�,5�]��]1�ʊ�,�!6�	SL�lA8�}�O�C9��V�D@0o�?��!�[�dZ�.x$Rn�\��ua���˓����v��.���q�U�VIg';j��`�O �Cς����7��)a;��ab�>����"z��K�Q�X`���Q�c6=����h>�'!����4�ꋵ���Igh��?a�Q����_��1��H��V0�����fQ�ܯ�r�H��3	PS�!�?�$Ӻ�Mg
���j�S�ګ��Gx��d ��m�fj�2�Z�e�9��1�_�&:�|c;�E���s�L�i�4��o|Ծ�i���k$��B 0�*4ؓm�uP�y��k���dND� �� �j(�6������q$�4s	���^ҌIɾ��Ny�'�ip-i�����a�,�G�Pt��n��G6�T�`�����ݬ-_c77����J��XO�8O��L��^Z��2z��QD'���H���丩ua���I���MB?4L�&|����8!K	�6'��8i�T�FE�V�j�֐�S�����k)2�/��t��3���G�Q�-���`���&j�<$�:�c�,�.G4c��J�{����T�r*r|f�w��˾�R�<���3c�B[26���K�ˮ2kg�衱}sd;�$����Z�r3P�E\�1�nʥ������BT9\�A�h�ʟ����Y�^g?u_���x�^��<QI�'J*D�3Ժ |?�;�ȇV���t�U�F�;�3�z�����{|[ǭ¦~|n�l���=�y�q��3�����߀1�W�Gj-�/�:LoG��ŗ���삫�&r��hc>�qP+�����hK�	q�P�t=���"�����N��=t��#$��+:��`���Tv�`%	Ę��X�����"�r�S�������!`_Ɯ���F��Dvh��i��+N�
�#	�~���G�P�B���wЫ��.�#-�72xSx���>z��ｦNU�@F�B�,��	8h��V�}@Ѝe*ۘ�RW�G���"�P��l1J�w��)�y��,�����$���l%w3�C��U��}&޳�ab0vv��x�*�7f����2��(�<�@���ܕ����S��n�"y��k��M�����ጅ�v��v�1OG�<4t�7��Ҝ�s�g��8����u�^i�s�p聽���¼Ĭ�}�Z�W-ݷ83d���|���F>��s��<{v��gg�&!B�H%�\d,���~u[��4	��F�K��������*N�2�"�]�
��('EpA��Q�L��� Ñ�����P�2�6������nqOn�I��+�0oZ�x���]%���Ïn@h=�_�m����1��GEѠm�h^����n�W#���ۦ�����E+_lK,�8l>ibLE�������.���~����*�[08`.���Y`줽G���-7b��9��_�v�?v}@��6j�i����U\m���,�s��W:���������&�%éyc��V^�B�O!̀�����:$N�y	@y{�{�xy���8�c���>��x����(b9A0%�@\�?�D��p��=f
� I9s��-.n	(�*^�/
$FW�t3 X���=�D�P�(��ƙ)�FG����B�'F����qy�A���><lY�G������2�~RD#��D7,�8w��&C�Eȧ�DG=q-��^��
�+�$�H(F��^���<,�M[�y1��D]z�]�&�e�vv3�t�C���NJ?u�Ў+���.5 j���O����ӈ�,?!w�mp��	��WMm�/��udO�h$r$�3�.t�v�n��Ȋc��,t�g��Z.��E��ha�z�Hb��������*�:����O.˩6"�Uˊ��j�z��PA��q�p�n��e��V�߻"'�i͞#���6HI�Uc�qm��of'��SɌR_�m7Dp�gl�}��El�-#89