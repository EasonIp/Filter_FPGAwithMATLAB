��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>	��l_����b�-Vx�X�w���<��l�~�s,�ǟ.HIpd"q��o=�JQpk�e�A�:�G�bV�Q�O �R������U~g<3���%����Z.���a��L��$�E>#�V��1u�Aѽ��)�G��*��jfMـNk�=�]�Grd��o)ł�ܸd$�>L[���`�/���a��8�K�r�'~2aUO���^]w �BpPA��;˃�0?6���PDK�����!��z�<ኍ��QɩM �TM�����@%�'��Sm�;�Sgh&�F ���i��<�䨋�0 5��!(A�Z��r���P!��op��.Z�%v�G�?���?@�Dy��3��6YV�X�VB��>�y���섟��\�ߙ���2��m;#r�
�́����� ��<"��8��|�?D\g��~m��aK;�u���U���|��|�_�>����c������	�w�)��Ϭ!����͡���➕�Q�E��F���*֋Ց��I�X��E�$�S�d��R�8J@��:��&�A�oh���ή�\x��k
�O�W��ld:͎�I��S��V)������	Ƿϳs�t�����'/Q6�8RU��۹�y6�yph=�I���2Y :�-�n�|��ًQ�8�h���\�s'����.\�"��q-nOux ��v�m�1s��f� ��Lҍ�wLw�y�� N3v�p��e�~�Ve�I8�U��U~� an��At�D�B/<�PXe�+����0}�����p�ۥ�҆Y�3���;S\�D`��M�ː�)zg�RUR	�r���t"�����+���W�_Ƙ����UI�t�L�@��A�z���K��z����=
�'���؊ddC{�e�����&�R.�ǔ���j��AG�)�~��9��迡Fܯ��ЪU��x���M��-���S���Y琱� %Wv��e��Īۂڎ�?uF��٘��M��gQ�����;%{�Z:���p�b���}{W�Q��y����7/&�ܥz^H�k��d 2��Cz��N9�����#5qR��l���Y]��)� &��x�_����5����u�zJ!��J��y��ń��\1d<�"'{��|�����$8��C������hrHg��c�O��c�V�{�&ءYH/���
}�Y=���B*�Es$Hht�@���_~�ip�`�2ϵ>�1�UP�ɮ٩�G���(�Z�㸒K�.�h�b=�dw�u4�@�-�dB�'��Z� � ��`�c���)��[t[N={2�R�ƹ�����*������ �0�q����1�գ�rSq�� ��P��47}�f�Y��:H�-��,m�K�ʋh�%�# ��%�rM��В�ZG�����8�P���5-��Y=�vdnHΗ��ʵ^��������kr��5͢㞍����}��=4W�j�i���7uy�������^�͠�f�&^�'�4.��g�n�|lO�p�5�*o]��XCW�s.�S B��[G�_(�u���Z�x�A�e:6vBQ@}O##�6�Y>�-�7�_f *e��:"Ty�T�#�K���� ��.�J��H[ǡe#�ܭP7Nt�\#D4��@����)[�c"*��V[s��Er�B����@V�.��`�@��}A�����.`��/E�]Q{9M�����g����*/,ӝ8L�BE0�*Wob���y%����$�r�z�ܡ-*K��؁�X5[�����t���Ѻ�ރ'���e̜�~}�q�`,R�K�u����� �F�$�qM�G&��<f�Ԍw�U��:� wmQ2S�nŉ��0���)�9���~U,-�HΧ�/�|�/���)5�TĎ3�>N2���+"�j�5OL$|��vΝ"Z���R����aq׵�|���Nh�����~>(������T'Բ�����kk!��)��8Mn�g2�9"��m��'��Ʉ��1�.F@���uM2+
�"$�\�4�|a,�2KV�j��k{4�CH�T���S����5w&�yf�����+>��iS��L��L�]M���9��\�J����)�yd��`eКi�wh5]5���s�b��1��η�`ӫ�.Z������c��7�.�
�&�|�L`hx�p�k�| ������1}��w,KQ�\��8�8H����>4MѰwGu�N4�..�W���Re��O� �0���_�yB�A~��b;� ��`_��a�U:�'N�=.�$w���D�Z���ٌm	��c*d����V�F{}IT�Jc�������X���?���O:��9�a�`�Ej�%�k�8��>�y�ո�;W�=�*�X��U���ʲ�Z�ro$	�M���PO�
���+I�o�А�_	1X����m�c`�'1҉��Y)�}$Ɉ�!�:��6I�̽�9����r���x��&���[�X!�KG�1����f&��0�!qT��$B�:��v]>?��#)_b�}hm,�����l<(^�绵g�#��|y�>��i&�=)� R�&A��	�>��ll���f�z��kf+�'L���� �>���1.l��|Ɵ�T#�7h�կC\\��SR*'����D����[�͏r�;�W^�Lb�HfA96ڭ����0.�.�.¾]����@�3�����n�p���\9���?��W����v�2w�Z�Eӿ�'=�ÕSxq���ck!��o�'�Ry��z��4��X�c���s�R P`���]hѥɂ$ez�ʥ#����f����/�6jo���@�gDUp�Uds���'�RTs@����:/Et�S�"�;��%��8H�H�,��T�~pU���Z�]��������ӊ��=�rb5�Ή	�uc�21��P�����00�_��n�A�����j�$�u���෫�*��(�Ê.e��E�H�E)=K�b0�Ҍheo���a-/��Ø��,Ӽc�ۚ1�#����wt�I�G��4��,M#�%T���+�h5�G���;@dL����ē�Ƹ�%�r���&4�W7%r���M8��%��(8�u�Fc�`�k���_t�ɼPUpu������5��<�g�Xb�������-��ב���b83�c�������۟�c�,�q�Ѹ+�z�9��4�!�bIOn"�m;�
�=��Cvƌ�Cæ�e��j���{ܶW�G]�MTB�V�-��{W�'{T/�uq�8q����&�4k>xD �xK�XOb�1���hU�}4���L*�����86Sú��"�SY"V{d1#r�5��wl�,}�'�p��a�e�d���kUW����"Xd �E�nئR�Gr��U�W�����T^sQ���w��H~�7�.�V 9�c��m��<���IFгCJº��'��+�����5j�Ba\b�je���ܠ�,�Nq����gpU�5<�@�=xR]\�)�� ���m�\eM�w�OfA>L�γ����-E����/L���?�sE�ड�)�D�N�Y��j��	.�ᇵ�2CX� �[p7��p�mirR�*س�rWw�������(=k�'���nbm'&`�/���$����ԯi.+���X���� �!����{D���s���d��LЌ����4)/����tH
[l�R�����@�
Oa��d�P\�ح��ꆾ���r-p1 ~hSF�A6Q����vY�G+�9-������$o����hpabC��'���J����]C�*���=&���å5�"g��S���)���\���{B"F3�{���ɭ$�]�sh�s�b�F���݄���K�g�Ŗ�ť>���}G$��/ӝ#y$��,����I_i��C�.�{�QΥ)Z�p!̴�6��405j<�����V �R��(��T�8!^���Z���ȵ�i��Ӡ�+A�N]�
�d�<��q��0~�Ab�D�� �+�ӞC�U�H��/�B}B����VF�>Cd��v��CB(�.X��Y:s�����NUwe�㖄��%	�+2�k,i��
-q�,�>:Xb�k�r`.��c&��B49L���<E����wf�̹fUR������y_T\)f��T!:�e󞇑-vB؜�թ@8=�ו��Tgb�4`��t�ŗ_�&��aL_��b���c����MQ�m3tƒ�8(���v�_1A7�
����}����TOQ���˹h�C(���;�
���Ա:C���!+��c��L����h�N�ד��z�8Y��h���V�L��?Qe���#�jh���P��L[pc�+wf hg��>��<WѶ��v�G.\���#z�*��參��)�(���A�.�ɸ:�#^e��Ә2.*��:�%Н١H=p����m�V��r>��򓄞?��]eb=Ws��玙-�]�Y?߸2>͟K5;B`��ۦ�HU~ ��m���k R�v����W����FA�u��io�v