��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ;l�Fv1�Lژ�O���3��������F����Q?���b�V����Ţ� K��Q�G�D��i�o�Yʫ�|�F�V{:�� �{��LBB���Z��^sӽy/��[����I����k���'_hx\�Ƥ�?���ƫC8�r��j���?�[�b��Gk����s��$E�C���Iv{��Ϗ.��R+!9u@Gf6�e+~�7k>�_3�T�@�@����58fW�o$�T�h,|���z.yhb+�[��>���W��Oѹ/t7y����8�A?X�Xw��J~���k.W�$�'��(��ꉑ'[J��TF�S���o�z󷬓�I�UW���{�|�M�a���@�F�J�Q�tx�tEV��Z��i��lzt����#��I ������T0�=C��'1#"V,���)�r����4p1����Ɠ��LS�d�,BbD�י��)�@/
X����0�9�C�'�8�5��I��*���ŀ�К�;R�g2�9B}������Qj����F�5#,VF5~z�wY@�g�ږ���jbY'��&W���Q��p�>��@牣@N�#���Up��]���ߏ����\c0�4i���jK�tƩ�H-c�����d�@+�FRxY�,��~F��(��y���^�)P݈�k4<�w���Z���?4���E�}��_�á��š�0ޜz/B��Ѽ��#f�݌$��3��z#G �W�fĨ��H+hnؐ�&�,�Ɍ��9�ċ1�(ֱ�{��v�RF�T5r�����F6�}6��2l����Ɯ-pw@���
�O1���3��~1��І6	��v�A���@�e!����� S-����193��n���2aD��T�=����y7ߛ�&"3"�
)�Oj_�ؙ���J6��XFK�֟�� �m}i�/��������Y��+��##�����]D3��1M��>c"F��(��j��3HB�3:���Q^<W��K\�	���
ŉ{����`�0��MƸ��]z�����8n�H���ǟ,�+%[��pI��)Vdܚ�C����Y�&�Y>�'z�b8�T/�y�	�
��|�����H�ͻT� 7���}�"�
��/d�NY�(�'��r�Dr���J�)�re����q��j��h������I�xn��>s�h64�"�z ��d�-�윪;���Sh�qg;���Zi��0/Lj0ak)x��p�o#z�������� �[�YBwR�5�r���+a�8��찎�i��U�5h
���D�I&[���#���yY�O�Z��BM�H]���tS�'�G?���=�r
�u�k>�@SeI���c���oL�}Ɯ�u�+$�Z�+I0t����P[��M�`{jk�~�4tJ(��#
�,Ц��2�\��1b�n^XeBmAL��)&lxf��s�Z�����xy��zQYu
ؘ��f��~QY'��
�1=J ]�	<<�ByoE��:�~��1
'��+�p Q��^3��ػ&Fpw ����"A�.��H���8��.{�]�h�4;�7��U1������2��C_2�sӁp$c
A�l*J�T󥎴��靁������1ȋv����wOv�G6����p�)������jPn��\?�� wO��H��xN�mbj#�w� U�`�e����|�La�m�m�V%����l��@k�Y��鷳N/I���1����Q����-e����9��xd�I"߰:�~NɄ��U}�Ik_�Vm���"̏�+H�d��ڳ�iP�?Bޑ��j���Z	d�.d9.���@‑w�C�\kq8�X�t-�L�o4	邞��[�mC_�J�K�~�#��qv�;a��k��xpQ_���(�)�`�\�-�J\~�d�g�{�K��ib��K^%�EO��$c�ћ��x�)P�|<�|��<��ϯ��kIG�+(��O����>%���G��k�/Hi1�@s��g��������PC�����2�.�����ĔU���UR�ɝ��})��l�����R�'UI��̒��4�X\kG6=!\��7Q�E�ӵ
j5�'�/V��~9յ6���E�ffC���{����_��y�X�sRb����"j�W���xT���z�N��z.