��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$�ʡ��s`���
"�*![�S~ded,f�Z�?Dka�n+O��Ԟ�Om7�q�{"�%6jVlL����D�j� /���uM���*~�Яڏ����A�b�f�UQ*0u!���}ߕ�s)����
A*Pr!ӽtmY̔�).���Ϝy��i�T�������|ZQ8|�H�@�?*l�,t�<E���v��C�f�C�O#ON����M$��k� �M0������UÛWc��f)�A�e���R oov��0�WtbZZ��{.��Xt��s��'���}c^�4�[�D\hg�W��Y�n����0�+��Z����/��2M_�H�����N����?�;��+4��9g�S�.��W\
,]w���)�+�-	\���l-s���Ȉ�C��'D��:�β���>ϗ�V��5�����	c�l���������eY"�oW#��D�����:���y�=�-�V�B�?x$M���U���Ţ�<e=�Խ���y �uX�c4xj�R�a�U�ɵ���h� �����\S�}�#�Y
��Wn����J�� ���P"��x�\EF)�ӣ���Ѩ��	�\G�	���[I.^��ʛ�31kv}{GgVː�o�X��o���l��?Hӊ��`�n�V�uA���FI�PH�d��9���3l�C�;���̔�p�z��*v��a)�ed���l�jtdr�A����&�k�0�a�\K�_�l�W'뱺�.���QQ���kA��.ѳ��F�LuGm�p0O�H�^x{��.�c����A�Gf3o%+�[���R����X[�)��P�p�c��'��
=H�t0��+�X�z�l:sb������V$��/],��Z���c���h^��f�g�9��%M�|k�g����=�u�!'c�������s�#�u��E`ߚ��
��}�R�՜S�==�>/�@�ϒ��q̦
f^�|��F�<>�*�Z�����q#1٣h�Y"�?D����ң�Pnׁ�*����=<X�/4�L��ơSE�~�*��z�v���3��!�uFtȋ�19��a1�X�R1�'��8�5S4!����ҫ^�Z�0�%a>M�&%J�L:\ �:yVK.e��4F�m�-��)�5p
X/y�������v��r*\��_���R4�J��C|卣b���|]H¥��!��QԨ��á�{� J�h;@���D��i��U����R�����^�Kg��	�Ҥ5��JX6k,�������jv����9/��\�<6A�j#��JM��]�L��������ݿ�d��R��
�H'nD3�hR�8���h����s��#�7H�r��ox���7;�P���<��A��&��X�Y���P)�c��ٯ��5�`���pF�yj���f��${���Z��V�A��2[�UI$���
���ñN�0��{g%"x����{�_�N��Fb�Zd�����G��Ґ�HA���N_�؝��eJ|�AOC����3WÊ����{ҟk�U0#ta��`�\��,#�.e�l��������!��?Mѽ��:����k+u(%J�S{P��-���p���9�T߾����hi�{���%�7C]�������(�N����0S1�8���[��3��&���%�g� 2O������&��F����/ V޴t�=�T���i�jIʵc� b�g����]��5u!�`���a���曳���#Wª`��=�OcDn�����>D��XI�J�g�n��/:}:Dr?>5=X1S��ӎ��H���^�Xw�K�@w�#���N�\m���������٧�}$��.��G�F�p�"������v�pl�?I�`ӣs�����˙~m/3{(A�ĸ}��x�u�8����Z�h��"��.�dt;����up��}\�'�X�Y���읉ճ�ӫ,<^cAWa�.2E8P'
��i
ևe|��k�M�i����w)��`�K�!rR��C�m�Q�~FT��49��k;�����E���
h3L�mdt��^�2��%�!9�Q�����崛? �{��^c>��s��w|�m�d� S��<�.��$d�k����[����i+�n�z�u�B ��Ba����K�	J�:q�ףD
`�����<�z]+��;G�`�f�	��@#�!�ۦ�*���c���y�ok����잲ϑ-����)�	��p�F��f�^�����n������k��x
�N�c)��Ěn�&�d�a�Y�,zX_(�O�)�"�E���g0@�Ȁ��hI[¸~�@��S���)��/�b兛�~yB��kQeΒ`�`�����{Xet����HFݼqk�`��Q��
��Fg�G��)u���eYi�f�r��bR�?���ra��>Fm��f�,�hZ��å�o��Y� �].��F��Wdj�.s
�i6�ej_���ʨ��Q�?����<m�3r��"��EDۈ>bl~bM��W�����x����nF�B4����B�p�����O�з��3&�O��p���z���"T��hR���-��e���eT��o�To���>����:�x��U�5d�PPV��[�J���P�Tۗ�C�L ���
�G��/�-ʝ����a>�����HX��/���b	.ƧP�zñ+��`�zO �S��� `��I��4�	A�`��]�jg�1�Uszd{�6z��6@��AIb ��^�F���vt_^�j�,,=Lܬ�Yj�_բj�`��J��1uQ>�ם>���֊�a��.d���+� ���}�s.��7�J����A}�΅@�/�B�U��58@�~��k˂��r��Cӕ��-���ܬ��:���I�l-�D�r �P����F��o5ΣZ�a�F+ήښ�a�.0��@�o`5���2���w��v�mt��NS]����Ҫ:a�}�s���3>��c�Zl76�,w��q�G��]��!Z����81��G�w�^N�j$TƝ�7�	D=����ٙ��2\�+`7��es�v���W�g��V=��\
������z�C�e/��3v)�&[�j��x`dq���;�z T\�s�洀�h��@����w0�G�ƶʹ�1tJ'��b
vӢ|�þj
6�'�1�ϧ�Qk����C�l-zD]ޘ�;��#�����g�I��N��Љ��4� ����ȝ�3�{`H�9�yG��x�gM&nB�|����z�,��_�d.B�;8M;O�,�_(�0DC>I�ɜ��>��;�e#W2Gp�[7:�3�8���ϵ���M%��r88�$T�
�<4���6�U6��k��3�׫�>�iìWi���y9U�2�����P\�\���e���Prm�${�9ra��*�	]��7GMJC�X9�Y|�"�D�&�ɜ<��ɡ[�߲���Ƚ�� E樶��P��#n�<PX��]U˦u�<��vF�S�ڢr��8��[���y·e�gw��p@����n`<��L���lC�_6Ǫo��~DMf<s�z�=~�8LP����|XhyַDh��>W���"w��?/2�c#k�p��N�Ǽ��Je ���Zč<$r�J�z�nX7bcf�{��B��Y^ O#�;F�D�����;�{(��5�*�yҖ!)q+�A����U��J;+/���=in��:D앋Xy�+0�@$8[��#9�+�ԅ3W�v�L���D#w��	<��'٨+��K����4h�'`��/'�Qb ��B}	4)@H���jg[΢�[��vu�.�� �/1�5&].Ng�W��G�R#��^�s=/��j�� ǽ)c�G7M4@��Ox�$�H���ʓ�¹r�~ۄ��������|+��BE�y��;�ev�`v���H��'��z��{��8���ݥ�m���..k�_�O����/����[��,Z �m�{�-�^N�`��q޹N�w�n�����:���K�W��E�J`����`�����>i��{��pg��DJҽ�������)v^��X��E�4DlQ���°��Ǿ�!lGl��o�i��9v���7��{n�T��9,��{�pf�7�c��w���?��.~�\��;@�{W��f��n?|���o(���S�)\r��;B]"i�{�P�W����Q���ν�'�.>�G��Ks>��L�ާ�V�zMV�����8�^$���z��侟��6����n������7ri5�2��#�Yu�S��Z.������^�l�`���0�E{�Љ���E��2��7	˴>f�{[a�?�~�U�Qy��k.塿���>&�y�`?I\��	�=�O"�9��H_zu�,�]��
Ͱ��&�n�v���>�0k����q���Kw�����+k�.���[ʱ|(6����%։������(����'{��+�b�(��:����y�'y�x H�ߊc�-|�Q���Cs;ۥ�*
�\9�tX�ۮ���zb�xc�p����5�J��I���.�c
���(���m/-ꤎ	�D߯�ɮ���+�=	�2�_9 �Pi�]�Z�M�8��E���9���y�����+,��織���\��0zFYw-S���_�Eŗ�L,��%;��.�p�qb5o�X\1-��Q�4B�[j�V�90�Tuʜ�$J�����u����0�f��i�q|���J_#��0Lf�����[6�(j;�_�m�ozkl����]�c{m59��>���Vn冞�I�浔�&�5^�϶��[�m����ծ䤎J@ �r��$��hԊ�uߙ:��DR|�L
�6��K8� Ou�D0W6G�@�J��!�����O}�o ��-K�&(��'�Eg���t��B�q}L����{ע�	O��E�II�۩'tN\�$
�a��{�v��'�_g���E�q/~y,���:�D��=��ԁ����a ��SȜ:"+^�~�q�.{8���-ݖ6n\G%'�LV~�d�aWaG��p%�5�N�Z��C=�FmV�N�����rLm���b,&+u�B���U@'��Kh䩝:y�����g���.�D�̄m�J,Zy��w���D�m�Kl�)ec���I3��̢@�0
"�~�"O>��.O��kg@dl[6@Fqk��n�H���� �f�r��W�ŏUM8d1�E����6�y Z�G������.�t�ӂ����G�3�*M�����SXRrÇ����I���fn�c	w��)�#�'E���Ff~]w�0�=R�_��A�8!~�{�H�K�x������Q���oX�A#q����Mw�C̛{7L�*q�)ǒ���wW{��7�=?�h���OL��&���H=ǇJ"檫\#�Հ&�M щ{�1AeA�h.�~J����1��x�����m'��$f���1�2^.>��ˢ5��'~r�I�L��#Aٔcn�H#�F�!j��TB��=�8�24^"�"Ѥ5N��@��A��66[���Ⱦ���F�<�rx�m�F�����sq\��H�F��5䪎_BU{��C��D��,N�p�����}#˜T����)~�w���s=)O�|�_�`!�
D�ϴ�򟭑��tp��*U,���|Ȝ� h��:���yA����,
�j��Ί���U��mQ���&3�d��\ۓ(��,�x�����O�?�9�K�v��>�Gfc6/	���X�NT6z�方�e?w�qj��X�F��5X�y�n,�h[�Е�jG��1e�)z�t!���^� �6���Mt�?R����K�Sy��g�t�+wvʑ3���~�/P�ǈ�8Dk�p�l�B�����m>�/a0��=c<�cq$C-�MÐ:���
��zVt�A�ۄT),((7�n-=���tE:5jT �m�:�N���7�hv�Ĝ�B4Q����ӻE��[f<g���=��>���$M�m	}\LČ�δ)�&'"�]�Ǡl�&*��Q��ΔC$�.��1g�(%�e�HZ������$@��'�_ќ�.ϸ�`�l���\�D�'��?J�O�Ř���@�IL�
��!!�kG�q�{�Ս����ZlU����_O��1�H��T�K�Ǩ��3X�KQ�>j�5cdS�"��DH����?@ �S�Z����&�R3�Q���;�*��Fg$�S��v�cV.��h5����̓^ڛFɲ�6$!��,�m����6U���"�j݆��5,	�(D��u t��hK! G��Âxv��@+*��IⵙZ�Hu6=)�kkn&@_r���	��(�)'$1I��Է�yao��2�8������}�.Ͽ"�T���'��E酝U��=�9�<�[30��I����=�����*��U2%dI�پ��M�V	J��I�~X:�m�<4�sv��*��4�P��wt�CQ�['�d��B6q�������i7��2!��.6^�ƥLz�����xD�5C�D)��͙���0�.,8��;iE�.Э�{�^<3>���cu���0L�*��P����ZZ^� ^ة���%ӪJ�#��:�<���߬Y�dT��g�(@3%�xGe�%�̘��8c��qjE�l3aZV͓j=S7��Nk3y�F�x��m&X��v�N�e�$�Ҋ��w	�nxx��/+�~�� ���.�����Ho(R�]x�����1\�M�p_���|h��D��v�Z�U�,����b�U6h�:�\SK�ܥ��洬(N��0����gd�{jqp�
tr����=��Gձ\]�{�l��k��$�n����M2#)=6'��h3F'wi�O�6��k�Q"x�4�(lٲک�xgWЅ�P;�f|@��2J[��G� �8G��X���0�s��_�h���\$�����l;����]�� ��9�:��8q��F�9��E�J��׸�F�������*�fsC����ˎ�|*�O�l�X>��.m�����W|��D�E+���U����v/��2-}g��1��s��#,�mB�<��a���In[9�ϢCO|�v8z>}��捀�|����Q���.�/�����Mun�e8��(#c�k��O>�\Kҵ%{as�d_�^�oh�j���r���&�ź5�rB�6�קIR��o�Y[���Y���_���:��P��ì�?��(wſJ�ݧ۠�<�qCsc�ݜC k�%���e> �#p}^v��F���U�~ʭH��1�U��baX��>�26�O�(̋9�\7%5��հ�UZ��e�}&3��|HF����^��A�=;�,>'���js'xC�o��y�*�p�%��xn�6��j��pɫ�j�&N�w�0�������qV}�\���C�����w��g;6���`p�Q�ER7H��,�����s)��n?��\��S	�߅���K�m���f^�s0j�B#�6�wG��>u�`#�� wc�:˰������vl�}�m������*T�qu[^~v�hcv��u�X�$��`4�5��&G��m����>a
Lj�;g����+K���;�f|(�����0�ڑ�G}:��yzF���r����Ae���KLN��V�ɟU�R��qy�6J6Lv��Xdw�<e$N�鮕���-�n�^�z�#F���n�#��;�6265�N;.��7Xyn�R,i�n�gS�hD��Y�z@�ػ����_ h�����H/�� �i���3�b�7*��uuJ��{���X�(S�����ꃸ�F��B{|>x�z�����A��.g�!ɔ��F��)��i���σ+�O��@H���s��ͮ���`A<i�6d)YD�o�m���8|$�۞15������`��<�4�6�}Y�Q��Ԅ��)Ԇ���T�Xc�<�k3�F�r����
�?[���/�Ezك�O�bMy?R��R��4��� NN��|�-2غ�x��t��m��L�Ǝ}jR����=�j�	��+��ؐ��b�Wg��9�z}�o��6�?����o�g_�45�xy���¡���a*�u�|�U�������4H&��m�3Q�=��p��%_�7��!��sQ	��0�F��6����������iRO�w�����8����U	Gq���e�)+j�q!0�&�ٿ�P��Z٦]�Rݥ�Ζ�^�����$b��n�U���q����me�/
�G�q�s�� ���vyZ��{���q�!����̈́!��H�N(Գz�H��Jiյf�Y���i~�]f+\��Ǧ�{���-�>-L��"dm���c�R�Ʈ�������'���+K֖w��������;�&���"��]����k��n�S]8Lo:��y4�w<�j�\h:�پ1������P�E 6�"��ؽ?���f���.�c=[��J��R��Zu�����@��p���tFnK����66�$�K�k��T���?R9��o�f�?�ഴ�h�wlC�(���n�y['�,�8�"dp#��Qtc�ˤ��hm��&r�Tf��tm�2�|��}U��Y��9�r�&��'����o֜H��a��o�B\5+�j�+��oq��.�s	����"�ӓ|}f��}Y��������i>~Eҥp�Y������WqGT��"�dh1޼�U�Ν�!�f�g ĵp��|-�������ɱ�0n����&��wI��,-���� ��l@<�x �Rf�Ș�)s�)���w�F�]O��A�H�y����h`5������~�u^�[�7!#���Ŧ�ནv唐���������<�2հ�q����
�(�k�ܒ�����%�u4l��z�w�I��A6
��b=tu��w+

Z���T.5���OK&���&ӖKx��==�9ɪ��������h���*+�>]�~clʃ>_�Էbo��3��%4`�:�uF��U�P���2� #tZl������P��\"�Dsi�(
�`�NXU�ve4�"�3cwg���hUk+v�o��5�nʸfI�ܠ�kŭ��&['3|����i�������P�k3��f��3y~���!��N��J$)�a�i3Su19�mg��Ӿ�4N��J�	�����%{o�76gw�6����d20�����M,Ame��cl�� Y��?�q=�g�.�7�e�mV�4J
X�TN��T��H�S3\y�I��U���ǿ�;m��3<�]�c3�X8��d	N|���j��jw~eq����&�oe��n�}�u_�9�zЖ�qV��|E�XcauMI�-���^{�,�h8P�Z�[��|8�}<HV�g��.���`�{��2N���AY*[���aw�ʅ�.F,ǝ �M�Ё���1�U�:tS�:��w"����<E���KD���l�3v̒JqiA���@6���m����$���o�7���<�F+$R��U�}�9���I��3?��� 7c��"�'KS�ɢ�!ZR>(H���_�����s���\U�C�`��^��A��`O�6V���_(��������K,gjd�Mⳣ����,5s�t[e68�Ǵ�%yn`O�ѐ�����p��nX����_Y��q�rK�30�#��b��Ũe���ă�rC�L�-o�p�&sf�v�g'1�)k9@a6�}�����C���*��]����� u��T�tvӊ�_��8���>H=zV/�Ni����֜�nU�W�[x{��t��K?OF�(��e7拼Z V�j�O}QHy���	��8!ښ��՟d5�����Nmq)F�`��i�����I�)�@tQ�RPڟ������fC�~ā:��y����⡨ݤ=���KU��
����s[z,P��5�E���~��r��0̈��s�]3E694<c�F����r2Q ����޺C�6��v��<8�)ݷ��< �A��l�~�p��fH]�Z�!x��H����0��k�X:I%���zH�S�l@v��!G:�����dt/(I�|����"�֒F96ڕ)������S��.l�Ȩ�����}�]����\�Wif/�ܔ���'�T{n$;�R�KH4�g�nǣ�H��cVw����[���杜-�`�:ԁ,��jZ�7��y�k���K�k��\��@5I<���KYr��V����8�.c�ן��QK�\��(�ˋ�No��?���O�q2�����~$7*Z�9&`��`�3Y�d��74�p��
\pi�X�b��9�ȇ"���/6�-����	����MY8-�Le}/�=:�7?Ơ[RѺ�7q3��5�Pu-p�4W�H�t��K(���Tf�>.��)�n�,Xk1���ns.d"d������8�%7\��&�Ϭ�/���N�5w	�D�z���Yx�N]a�>xMG$Z�I]�ՉB���!ng�x�g��2F����Q�11k1z��y�ݘ)��C%��~��SoAJ�����X������%k��!�Y�m~����E��e;�k:v�<f	����`R���wSa/;���@��/h�G����<�1�>b��ɔӚ{ �G�d�{��d;�{͕��h�{�&q(�O�Q .=j��G��M�]�.\!�Z�.A(\�I&3qٚ�u�m���38��b|�Co!S��88�_��J��f��F���!"��D=�=Y+yX�����-�_�\(y����*Rۍ�A)���lܟ�ƒ�c	���dO�yz��ix���u���ͽKl�-,���
�,��غ�H!��KM���P�Hj�D�O�`d\������Ř �F�kȵƺ`T=�1<b/1,�ƍ�d�O7~r��P](L먊*+ɽe���icJ�m?�.���/����>H��)l6b�8��h�q|Rm�q�p�s��%!x-�4�����C@�s�5^ׂ�}L�Z���<���^�f+�)��u6��M��/��p�l2	�i�ί�b�_�4�P^�l���Tk*9 ׶��\���@�i�����}�A�|q&-uw�