��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�P�;�{��3�OT����n/\�@���V�F�	G�V��]� z�`t���y[q����a2��;��i�t��,-��1�� pz�jI;�"<i����#{���<�G�N�3�mŬ�#�:����(U-6��K��j�'��Y�}'	T�(L��ag�=���`m%5�|Nq�Y;�:�|���Q@Y遀 ץ1X�q��j�%|�H�����la�IKA�w��H�=0z �y���Ʀ#��au��#E*��p��c��>�$0i8Y=�P���(�]hϽ�8��1���y���*��V]�t����śvrs�C�������e��*э�L���?�������,W��?��z_��l��8q�'jt���N��A%(5�Uq��p��;;;24�2Ƨo�<��݃W�p��v�~��I���j��u7F�&daI�Ő�������xS��:uz$���[G��⪸M'-w��f��e(Y>��%�vO$�?cuH�g��G�����	d�F���^��� O2�_�M�#
 a�|[���.��Z��%�־��� �[��gTTg�u_���3����0l�B3���O��9]cK�G,�ϕ/�L�ոk|�w����j�O_�:Q�P��<3����?y~��VM�11�_���R�r��`Zn�BͲ>���c��ڏ`���N�V��J�`^ң⎊J�x%Aa���N����!�A��;ڿwD(��� �K��]�@�Ē���R @r9��UT	��W�3�酌N�j"�_�sg�1�H��2[�{�����=a�L��o�����Χ$>`n/��OE��D��G�P"q~ci(�i|0td�wT�g�����)!�d�>�ѥ�?~ �+3OZmX��A�j�R�d2U?��O@{g.�aĻ =�$����L�e��d�H���e�;R���� ��A{0�H����Y��{�}K��Ҥ��э�
� >�Ц&k�8R\�y��f}89H�\�^����k�mh�k5�y	HQa��ο��J?�Y�丏F�U���h֔�z{)W{�`��]���=��I`d�ɫ���j���uP���fH[��Ň�K1���"�U9�L"
~!.��%��I������|������t��vT(�,�g�ߩ����F��X� �u ��Z<C�H�W�Q��@ô\��1�2�c���r��51��P&������Yf�8��;<ޱ_��!Vm����J�hP %�&Q�m�!�{�ϤZe�/��N[�o	�C�.J���JU���Vn��w׽#��:`�,#*��T�ɤ�C�s�mS � ��$�Ś/�oe3��vw�U�]r��k���,-~����]A�AO��'^���L�RR%7�qi�ڎ�j��� 9�8%� �34���$�F�F��O�ת�ߎkO��#����U���iT~��i�h/��bx��,4�&Q	(q��ĹtV\ǖ[e��1̇���ܱ��X9��WL,��n�u�N8+���n���[����$,z�]i�A"�q�����M?b�`D��|\
ђT�$�s�H�I�p��9nݒ�\�D��//I�<�����.�[����Μ�����b���2�I6�:.�� IZmO"{H���Y��=�Hғ?��S���Z���1�&���3��!�.�Xv`u�Tq˙�	~5�vQ	VU����}~�K<�	&�M�t�8���&3�:�x�=D/�=HG�����|�yQ�>)�\n[ҏ�}�g�-�I;ͤ����-�{S�sc�|�u�q��I����QJ�f��^)˵n�j�}���=��K��i2[�� �3D�%Aj �R�խY5:�UFl���8@�����2)�NL��ș�PN+!���[cF��U�ₖ)V!��h��^���c���A5HH��� ��N���ޯx��G���O�uJ��(��	�}�N����K�.�y�p/�4L�ﰄ
��aE���Q�m������T����E�Y�XS��T���Y�i |�ԭ�]�X�Z��A�4�
˫|$eg�.L��'NҒ�������9	zBgeBp���"��9��X.���f0c p��)#�k^W�! V�C�@T
�e�(�N�G�P�������;��/Q���IR�5��F��ʡj�Ѝ�G�'}���W+S�Ӭ�GpJe>dx@��=�b�X�n/p�&�����"�����r��H�{��G�aE��Q윐�`	�Q���ԋ��8��(�s�JE��c@k������.��Ɉ�����r1�'�1P���Aǀb��n�7��?L���p�2�*�[�k�	ȶ�D�ꌣ�T��v����(�cl͂/8�"��Ok͈+�;����!�Ÿ����doآ�B�r
<�����[�W�i���j�0*UfؗFxV(��8�Fq���)��49�,+=V�����E��8�DgLG^�k�I�w�/�5/n�v�� L�!�p�o�GTo���<�%�[���gʊ�E�����.�i�v�'���`9�*VOX���eL2N@�s��	?���Ǥ:b����\�����+�������I]qn�|E��W�?RB���)�|�|�>
� �Ҩ5��(�1��S;�[}�w���_�mӱ��3�K�'ҧր�0WB@i��IS����"���cd��E, x�]-n�:ܧFV�t����B�Z!��w�����':,a� ����%�bW��I�4�����؂��=9Z2��xQ">�C�ө�Wi_;�Xd�� �y_K� x�3�1f��ȻQ O#E7
�O�ߩ�5�O� ���
�4�{�f��f��fm����dK�]��89��"�;�s��J�X���Dd B�xM�UgD8whd�W�?�X�����;��P@��m�+��䨃2!M�fO	�h��8�v@l8���SV��6v����EZp^�V���ts��@i�J���R讥>����Ze��[� �\Hg#��k��]��3�(T��f�˩�;�_N36}G[��l��7=�s���(�n<๷T����\���b�Rs��9���˧l���9�H�uk�x �\��î��:�T��]{����bZ�wX^��/	d~
��B��歀r}xW����1ײ<߹�L��)�1Y=Φ5ZF��h������D���2+���5OFP7J�ۄ���g�/� -
s�YNU{*�q���m9+���ku~���+`vߗ�
YVZ��,gǎ+�G���H�l�M�Q��^�������C>�<oM�̣��̯`6�Ar��N�\�O}w�REA�@��R�r��享]8�  DWT�.=G�h(��2�rF�_�M)�O1832�v��_��� �E�]$lp؋V=��m�\Λs���	n>�t����㮦�UD2r������"4���T=�QI��(��cL�$C=����(��y��	l4d����	B���8��6�G�L��ó1�Wl�|�����UAN�0ِ�;@��d�I�˚�DZNv��s�P�7tI��v�����Lv����F�W�n��� �C2����՝��B��2 ���$�"��������ӄ8%I4mǄ�b�Jh���*�X�^���(�q�"�$���{TG�-H,����>���l#G��,(56F�u���o��Γ����O���1	�׳N���/BG b���:��׷�Cx��G�-'��'���`B�R�Vr����@K#�l2�_R鉘ھ�Iv �a�H��裸n���K���˵���OU��븿7Gfa����9r�$#O��.�"?��3�g��׫�yv~}@Uem�&.��X�B?b����vC#�ښB��4��0y
}�o+�X���+8��a1z��n�V����Ȁ�jd�k|ktz�M�e¿얍vA���g9������L��+�M��a�EF��Z>�Y���G��o9g�\�;�C������ĺ�p$�d��^��V�N���C�K(_���N�x�V�>nMكE�9@l/�Q�؛X/5F9�z�0��2��|�ǐ&nl��SLӤ_�i��{~��p?w��Gt��]?/�SSAM�;��҅ \�s�J7Y��<k_���<)I������}�a55E#�I��s\�.�$�N&$"ݪ�G���H�d{��t�B�O���co[�,4Q��hTé��q+ʂ��w*n9.	1})4�t�m��6w�㗼>+ة� s#t;MI#p�t!�����;_���}��[9���M=�� �J�.��R�t80�	�C�a僡(Ll�H��GN�� ��6���A��+�-���UwB|Ĕ��{�ɛӻ��boD����X]0
��i��Uo{����VW{�[��c��5Ad+�]*C�0-�%�K䱑8V��T�ؒK�����>:����\$%�a�ڒ����fjӽ��6�R�@w�=��8Bvs1���J�>�@f�Kw�H� 9ˍ��;'��E�5��I<ݺr��z�uВ|k���D��3�m���yͯaV�}��z3��ւ���JX��^3`mՈ!�7�\��s?��� �_������A�+����S�y.H�_�I�BXt���a� +YtO\R��|We�ъ�'%v�: !�7+�W5�3-�`�F�����\����f�{��󀆟)��hi����q�k��F!���mX�-8��>�<\v"��r)��l��s/��!�a�d�����[ѭ�٩�;��S�^�����İ��g�'}���\���|p����tx��ZM�	����e>Ov����u�8�GÁ��j�56Q���+m���;o�2�%xFa�T��%х>,��[5z�Ң0�%|� ����6��d��}B[�Jp�l���q�*?U[�z��yN�d*�Z��IS���Q���y��Tܦu�M���TX�`I�qٙU��o��Wd��H���nGH��0u���	WD�4e��yG2�{�F�Կ�p��d����������Ϥi ������әe���/��5b�����A�[dbr��ug=�ELx"Fȯ�-o��UF�X�2%<'�W��U�ȣ�w�M����|��<2�}��|�?�#2���l6�Udhα��2��m����>L�z�D�6��}s�L���0da�v�����V:�'�Liv��RR��m��[;@��3Tں�`��;Z`��-w(�/*>=��(@n��۞*����Ě�F���E�q�sS��\���*A,�*fOxඬ�_�)�ӶkN�ǃ���ba�<.��!=�:�^.^V�J[�'��,����f����Q��&�.�J�}��ьHK�{��q	�N�Nh�ei<��S��`�^F3K�t|�1b��H�b�W�$RaB��Ί�9{�B��E����D�����7�D�����u�%��ϫ��%.�`�r�0���d/)�w�R&��O̲�b����	 9��{�9䆣�J9���rY�<����&�t�T0��G!�<~AW@o���y����(�W�2��o�3mdwS�H��j�6�Hq|upٛ����m��y<�Z%�%��ź��2IO����Yv�*��'���Ab1|m$bv�bk��%�:���T�t�YC�\*SEڍ'l}����fo��S�lH:F� ��v8V~�����*=�#�P�N��6a�H���|�DnM�°5��Ŏ�d���ܻ��"�A�d`�����X���ԑ��b3P�=8 *��;�m����z��ZO�g�#��ˇu��+Qμ�2?5�uhеĂ�?��Os����ph�~��R�{���)@3�P���P�-'�n=m�8��Z���TL����.���&A=�Y���>=P��@��s'����$��>�>��Ͱp����"xX;�/s&~B�Z^s��z���d���+(LC�'k-u��dO�;�n�s,G�c�Jk��Էw�V�����ۉJP<B��ݘ{� R*�)�)���p��~j������F?�y-'�n3
̿C $�[�Y?r܋ڐ�@no�r��:�����!ab�4���hw�%ZF���Ȩ�28�g5~��Y�8Gy�(��c ��۵���X�s2����z�"n�����N���$e��M�}��W�� |���B��3�GLt�� ��?������j*��r�n؈%÷��"n5>��\Z�6,�U�Cލ�,A�L�HH���(�5H��)���p$h��>��졞��������~�԰�G�����)�Q�/�vkأʸK��,��(�a��9֏-��E�9�h�H�]KAFJ�T�=�P�[@y��a7`:�y�qJ~�')�{g�O߆�B�^��5�*A��T�ԁ�{�F2�+�0�BF�S���]s�}��>�Cz�gr!���i�A��a�5��X�~HIcBK�$�Ǫ����x���W�k�@�ht���,�y��������*68����T�mW�Fp�1��Q�
�ҩ[�O�T �eH���3>C�/D��1��/9���A!G���ȡ�5���+��ݎ�Y�'��P�#�-�W����R�E�U��p(`[�E��i�b ����	d�2����#����e���Rv����6*&��,v�Ҹ�9�-K�#��c30�1ؙ4���<h'c�������s;�|����%�NR����ɡB�����-m�:��:��
0��`�XP����_���n�Ž'Ġ��Ѳ��b�������QԳ��-�8����U��V�Kj s1����P����;����3CA���+4Zus�s�T7Wwݍt�;�L�Ȣ^���M�O���nTA�����1���Vß`�*�MW|	����k����1�K���䈾��GA��r�u�~Z��śV��:��)��zsw��%�����.D1&:�F��hr�!�F{�x�2ۜRI��br��4����wt�4+��|­����;uګX �z�˳H���`)=����Ͻ��5T��e�Qo�N\?�*!&�q�cK	�
o����tҗ}�\	�M��5�4��0{Cc��@�&��c5�Z9{4�-�
-Y�>:�q�ߞ���Wjy6��L-}�7�4�L�A�L��̭]<�<��~�F�t�(�zϰk*�^l�g����T�-n!�O�V�+oI2�3O�~L�OB*�L�I6w�<s����g����y�E��	��hToi�#QʛD�i�t��X�ZH�>X.He���v�A_��$�ݑ����X���S�V��>��3���O�)���n�w:�a)�2�
�nL�8� ��Na���U�ZY ��I���r���z0)YЮ/W��P�ΘbX�&��Q�Fk!߆�|�)�g��+q��pG��l_P[�ABd��v:�����qX �3�B�|�PΓ�[�7ً��lM��]����;-1�4$Q{�۳"V�N-�>¿vό\�a��hR��������p��QN��.�ŋp������lꍵZN�{�Ms����3hB�7���pR�s�x��n��R6RF���Tol4�~���$�'���9W͎�&iMG^GQ�ҧp�$��R�~��]x�pο���"�7l�B��������L�FG0�V�����Rze}ZM$O	K�i"d1U�k��T�-~��W'3��o�x��\^�)�IB����#ߖ6ȿh`JY�,K����R�����E�LH>��:���e�b�6�{♿�.Oi��(kwʠ��Vj�W�B��r�5�֌Z�u^t�T[<��Cb�qg������&0,��j>F�{P�: ���y/��g};��x�R��-`-4����V܎EI�2�@���S��m�����������W�s1.ܢ~�����`Il��
99�(`�1���e�ܩ�=d�a�ٓ�?�Qm��g��Lɠw�/ǰ�[��?88�`C��V�Ɲ3+���D+\p5!��~����������q/T8f��P��&fWc�~(NH�qX��"C?�@�H�֛?�O��N�aC|��_�TfL�y��+�sDk�a�1�x��K��T1�X%�/�*u�&[$���L�L�-��U��"�~�]�&�o{e���!ey!���I�c�1zоM��.Yu��ר�)��C�m���5q0� �ir� �hu�����'���k��<r��D�my�Z�K����T_�;�b�%�F�a�.Tn�/Q�Q����	�}����J{jᴮ�+�����b�w�o\��({��_��˔�.��}\���-/^��z��H�[����f��>�������>�?��D�p*v�&�������[Fl�Z𘈥7�{.�A���VJwIàI=Z\�ԫ�z������V�o����FE�2Zm��S�&,�Q�p�+Κ�n�2�{���oFʣ����kk�i��PWV% t� i�-�x�^w��=�t��>G��|j�Q�p	��zѿ���&x�z,�� Qe.�a(�**3�l1�|z0��$�ȫA�f(f�b:�i�0D@I�:���C��>�.(qt�'���+rG�VYP.�~I�o����1_�U�q�PG�����7�Rm���f���l]��b�:����W���v���~�wݱz����<��~uq����Q���@�i��D��G�ĭ�9��͡���oI�I���_7�S�Jv�kL`I�{�d��ϥ�2u��0*��7�"<��@��䠻.�A|yv���$L�^�GS��������������p���o�k�O��+��i��@�B���|v9%i��B�o�����)G|����9N�+�6���RB�������m�Q���k3r���#q���HY�{�?�����d�
� M�h��(�#��:�;dS�]�4������{�(��Q&���-�+�Ο{1�Q?���:|Ȳ��l��Uf����)�[ƴ4�4A�/#�Q��}��t\�3�+1��պ���	"3�KF��;�CZ|����鰻.[��X5|u<��#J�V��f���R#�\��1�)sw]˻������a	���@ޒVw3k�u�}��ƅ��D�*̓�'��&ub0�� �+��K��N�zC��2�v�X:4�Dn1��/�pt�
��5��~��i`��7� \��X�$�$�%<B� 5���i�p�D����b/:Ğ�R)X���c��A��3l�Pn뻫�"�����[��~�8�'�"
Λ�,�@(�>O��m����=Ou-8�(���ղ>҃T�\��a��3�h)N�Ħ雞p	�ҩ_���a�^�}�a�*#VdI��{-�Ј��v�P��S*�å=��������s���ձ/�է�x8��)����vc�ǻ�|h���m
cn�N���;���y['�ױ�}���˓+��M�Uw=��k�ּr�h�>�ȓ�]�� 9 �b,C��L̵$uBw�@�`0ύ�>��}��ծ{�`�4x��q؛қ}���O�H?6�*'�s3�_��I�W��Z+�ϗ������I3"m�!��|oO�a�����@o�,#�\�eK*����}�ԅ� ���Ë����>�3��J>}v
�V�!��2X��2�S�Ny��*&45�S��2����_aG9���W����W��Żn%�-n<��KR�Ǘ�8&����jt �wF>@1ޡ462��T��I�����|l��Yp�N���sp�8��aۧ�k�'�lKY�9#V�<�@i�Ŝ��O͐&7��Fhf��`U޹U1����k�X���N�b�ۃS;���	�T=����,?E���iIU��G�n��k�@V�᳼�ƪ��r0[mL,�8�%x��-
�w-+%1؃�\��� ~��ߜ4A;���g�ɻ���w���q{e�%���,��b@,�;LS� �34���m�
i��7�E?���aȪ�U�Q=�%�U�Y�N���������#7���Y�������FS=>E���(v'���C����<��y/9��)�Iȧ��)�2Z=���]M�3��XB��I��uz|F���r����7�S�	�V֯NB�c/�n��ҤC�r����lo�f ���wN�Ө�*����+l���{SbA�\���H]yw�Jj�]sor�2����e��̉ι?��33l��
��e������.�|ɿ�YО�U�v��9-��i�U�Y�͡s�{p��O��a/g�<r��\,]�G��ʐLٵ���;�V,h:*�.�F(��[��J��vbg�cnb T��ӆxAxk��*������gٔ'(m�%S}����ԋ���"��F��I�h��l#��(�|�[�gӻbǫI*�5�@􂺥�_�n�$F�OTdk�*-a�pB��"P�ܫ��NѸ�ʽ2ʞ��,g�p]����Γ"�y/���W~�|e$��'��v4���v/#q����l�ׁFy�x
6���O���ݙ��>�^[���7��q-��vH�g�]�hHg� O.WC�OP��L�L3<fÀ2c(ME)��ª��Y6}$�U��)l~�^ǚ.�{/؝e��2�I%JT��L�l�IE��+:#(��.)�F*�y���j��z]�����wu)��g��4į�Z�1�jh��r
�^��`���Ȅd��S�O�ņ�R�!.���!�����w�Je=�����z]]�rpݙ�u�w��!R���%��N��UL&��S!�jh��_��¨(�ku9e�[����0K�.��=� ��L$�/O������Z��[��S0�u ����&�C�%
m½�-�8�@=�ZWV�2��$7��M8�Z��a�)눞xK
N����n��[��)��c>����'�K,A����	�d�4��YM��g�7KtmXq�5s*󞑱�0����;"a���Ī�P,�F�(��`,q�ȠW��A(�����4�x�4(*�1�9!� @S�eڴ�k�HU�����Y�yL>,$ $�lq�[Y{P\(Ф|y��Fի�#�n�j�&0��K��p��7ܹ��?�ۭ�r��S_�-|�d3��z�QU��[vnK�6JZ���2uRZ�����l���-�D��uA?P��N[.���ć�E��u�����<e���Ʉ����*�l��=Q˴�+m�ſ�2c*lY�f���H�$�HX:H��|Ӿ��R �I^�m��H��"C�� ━{sZ�b� �E|Y��?J2�a����A�*Ν�Y�
�.�b�ׁ+^��f�7բ���4ܢ@�B���ٍ�c���qTe��x��E>�P�<���noK��s@���O�����]���Sl3�|^K�#�(���ՐX����Z�T♝�^���f�A^;��L��n���c�pm�|�C�����}Iny,ޘF"߯����Vnb�[�ܖ��*�D�E������)Z��>�W���{����G�߰�}JȑD���>2�:0��f�x���.z�2W�:�޵q�t��A�lK��P�g�6;�hJpy�`��ǌ@o|pGp�/�L��������痮	x����#�RX�Pd�	��;u�����9s�A����Lٓ?5-ұ���=	��z@S����B|��Y��);�g���kQ,NL�r����2����QMzE�����F���a4��<FO��g/��Q�Y�ũ!�սYY���e��{3������.7�H�#� ��R-|��+<I`''2;��|��C��������/�.�"�����]x��� ���8��\N��E�5BGN���wҝ^V�(v.AZ�6�ޓN_����,�7�(�h!�4��&������I_���c	��#3��<{!c�G���cX��]�T�|����$'̩�٥������0ǼS�w��6��Ψ��9��P����[��Z��ht`o���6c�s��+߲g�����~$�tw�M���\C�t�d�U�W��IQ�K������5����&W�$�얇S�ob�� 3�7���d!���D�"���6���L�4��A��`q�-�g��!8�N`/̸��-y�厮�z.�l"=1��-x�-ƴՊ�*������%}�M<p����X�N��Z��FŤ���ӱ���h�K��Ѿ����B�w|Ic��~ʽ�:�����AF}n~���J�5�#�`݌jW}Yɧב��d��V~�[\1�I��I'���Y��LV�i2��w��;���3 �Y+F�]#�_,�
a �^|$��5Q�PP��lX�_A���r�v��x����a��|kѧ�9����Q� '�w�N{>}q����U� �d�۰�tN��r�RWm��kz-L����|�1~��z��&^?De=��P����!-��Ly��W*��`e�ܑ��Nk�z$)�,A�H���̀#�l�����ЕZ{�m�	�^)�+�o�q�J����h�LW3���Aȃ�J�R����K�Էt1��V�9��>U���YE��Q�V���g*�nZ�=� �K�<1�J��	;5j�^��/��c"�*��?�o��n?;���o����ׁ:�`M\������od��B-8��~���U��~X�P���X&c�a�1\�sp��%u�!:W8�4��;(��Xs:���` Q�o���K��	`a����e�ot�(-����W���P&5ۭ��W	��\�8ke�G!I\�]���^���De7��8Ƀ-g?�����c.�< ���8gYE@7
�����1;k��-��A�������8ۤL�"ϳ��n\W-�ʜ���s��*��S�!i���Y�^2ǎ�׫��Z��$�!�OW��(|q�ѫ'<s�:@)J������?W���w��5����;�wZ��F���m����tD�"��?��1����P"��ʦ 2���j�E�}�;Ϻ]=;�Z~����s)�M����UҸ��_�g�m�v�t���'��T���L�*��3H�	�~i�d%թ���q�y+|�:/�!����$�)�4T�W��O���2�w,h�ص`2d�jЊ	��Z)?�2�����6ߥ��[5�q[�\�$*��ʝ�|��^�P��ֹ�ݼ�����u��|�����eHV ��d�S����*ly�ߐ��@�����U�zV�t`�jY�8h� �F��6����K(�e�$�2MB�U�3���e؏�L���F��ER�l3�KQ�8)5J:�x�H;�l��
�O��S�u(��f�t�x[�w �gT�S���A�T�]�n���ڍC.�lxO�ɯ�NqV����]6��܇x#�f&�(��Ƌ|I��/2�oK���?ay�f��4�gC��Y��K�4W�u���U�C\����֎�/2U�ͅd�[���h%�����j��@�Ib?���R����R}ġe]<fg�DMCx.;��������+5�+ʜ���)�����.�j�r>���}��xT
u^�*a���!��]����t�	wM�*�����"+�|�<�Čzi[0ذy/ǔc+X^/NY�5��D` Ԋ�%%�*^���X��J�֥�ÁZx��h��Y�C
�{`���;��7�|;0�㎽V]o>\�;Y�.�扠<�-�F���\qg.�����S��N��G! =\H�.d��RZW��l*3�q�=b��0U�C(��Um�/�-��0Z8�����j��l3ե
�6\ʙ�#80�X�V�k�݄B��_uV,��2St��#�ՠ ��Y�g�K��!)&���ފ��(��� ;g�����j�Iʜ�פ	�F�7_���R�l$�S���k�4n��wa�lݽҵ�$�<�g�I�g�{�P&���rH0�����L��Ǫ����o�p�<ժv��$��+j��5��?]��e3s���1�L�����E�<T�(�����mF�"��N�'
8�d�Y��l <a,�1�/�jd�����'��lJ*uq��yb�Vb��_ S��E� !���*��r6m��=��n�E�!;R�z2d�P�uz*$}�m��jÇQ�;jN�`�v?�
�/B^j���=|�9�I^�k5��[W� "Z���9	�V���UUC[F���xj#Ꝟ[i�v�<^}�J�Z�k�S��t
��="� :*��G�5�CA]��y!�X�����i��~���j\��8�`�?,�M�3��e�h"H��x�g�����8�L7�C�n�ѻJ�>1S2E�T$���
�t�Hu�� ����=�M^����z���}T�@�������5�}(�4��hP� �@��ܚ}��B��#@��pM�UIH��S�D�e|O�y����&e���P�hIgM�]D�Γ���q�&�-�H�����n#��7u�bY�7~@�G��I�$��=nC���//z�<��@"d�^��]�[��暒��^�d�7��'>�d���L�Qz��ꮉ0�$��]�Do��奯I��?�V�̜�'0P~>4@�r��k'l+f��@v�4�@;�|�6���bJe֨��̋=(�;��!:	QxZ����gI�R{���^2����2@��s������Ւ=&�8ᮠ	4N����çH��!�9�M-�rd[���dݗ�OQ�W,;�k/�#�5�åP��L^���#]8�ˀ��?9�λ2VJv�{Sz�@��|i1xV6]����~�5s�*gÃ(@����n�mD[�wL��4��=��ܚ�{��S#8��x1��6��h��'�휼�r�K�@*�$5f+8a����~Ѡ�|���ǆ�p7��'K ��AB����BY���\� �V�uJ/Ҕ��!TV��iM��K��@A!�XA�9�%~e��{]u�K���J���En�s�ܳ@b��U�#/���������ђ��ŋN�����1"Ad�Cǒ�,��(t���vNl�P�Ȟ�W�G`��m��ǳ�s �+��I/h�L1���%4uƓ���!��k�Q�?[���ށ��G�_Q�%4�eD���?�.�@Ǽ@V-J�Bcu�X �k��u��*�e�%(�p�k)�-ߤ�/'�wG��{U��gԥ�N/��݀�V�hT�+<��3��y��߮P�
�8�X�՞lM"L�꣐~�����M�g�
�r�8�A%A��*��ٵNFn!���'��.&��F��#~0I?��A�����x�_��l�&�Q��*��O�� ��]�57���c���Qm���5U�4�Y/�NX<�4Iۙ�S�p9��+�D���T�j��4�wt�1�iW�^\���m���T�]�߆�e8��7A����p�A�Q@�� *x�*��0��_V��l�}�K5+�Wbm���٠Fp���{��;@~�S�E+vydݭl
�'�+)���pDIyp����ө1�����סc���HF�%�S���z�N�� �?=B�@��
o�B%q
�:��)Ϫ�@jv�a�K_d��5�m(�j9��/W��$8I���r�������(���$!7�BD�m:��U?�pŐ��F�b�މ���F(/L?�\���gҥ �WP�;&f�xM�=͓s�
�Ya�ᴻ��U�G�*�:�t�㘭����G%~w�ZE5>�u����<=9�k�Һ>#�j�_#�YV�trb��ɉ���o��;gt'SL��&sf� ↈ��EX��9�8:�-�7+n�Q������hz��Ɍ��q���_����o�0�0oȗ�Ni7~�Ъ�D�R�9IUQ���S	Ϫ}p��c��Ԕ�@!Y��.via��"�Μǲ��i)�R	���
˔�/ѵ�e�������w����ʳ̳&���0f�K����� |jH���������L��b?Dm0�H�����n��Y��k�P�V���YKI��1�$�t���M(��C�����^�bb������`�q�{e��G��o41�΋��rj%A��­�1�(9�/��Z��ځjz���ri"���'�d��:$��=xeτ�{�������C"�����*��H@�s�:6��Y�*
�5��`ʁ0=	Q���7��5�X�:�o�_��E��@l�(|D/�[�X�8�0�}�T�F�M�����8h��q�;��~�i����m�'����5m�zj���0:����v�����Z�!�5�����tW¥a��#O�z�(jB�G��I~�8ݴBe�1=���fM4�˪�=�[h/�_���U%n�W
�*��C�F�4�_o���e\C���j"�㓉��N���N�,�ZA1rA�E^2d�t�P��&@�i�� �x�1u�g
��;�� ��4��ە�h��Cs��ס U�|�)��R�Ȉ�CT���7��c@�����r?Z¦��!Jä�rd:�o�Mp�g�e��ʶ��^�Ӡ*�cVN�r� 2a�8����N�V7%;Y6nK8^���ĂҜO��IPx�Q`L63�\�GڎZ�� ��@4e[�I�!Ψ������TS��g��ޝ����A��!�d,u���T9�{�7t�yY^r"D��1���.�eم3{�Jf��PŢ��L�!x
 ��GR�t��F`WY1St���Bu��,Ll7�VK���w/ ηk��󕛹+�H�F�Q7�|�1�_1ОsPO��l�Y�B��Q3�u�{��!;Z�0���|տ��o|�J�!1�zM�Ψ
s1kv�H6����#.�i}�H��Q ���
�?HyZ�k�I���WU�!��,䡠��>uP�F��c�0ܾDcO���ȍs_P���ay)��$d[)��T�>��ݽ�b5��!�0%��t����r��JE���/6|*h	��w/�l��B|�+^�r\En0YQ}w�XH�p<�!�<�l��Й�_"'�#�bU��p�������+ҭd�Mx�vAcK�䈈Z��|�������F�e��Wk�ş�ɶ]�l��	V̗U���G�;ࡠ4�M����y��!iPw��=�/y�~e�턖>�����A �(�(h�J|fBx'�:TR�ȟ��d��K-����e���s:�#c��|U1C@� �T��- ��"U}.� �����HJ#�k&tљ[�F[��9��1�����=�NM摡8{��R���W*ӂ�g�=n�k߁/���XH��r�0�2��;L�<ӿ����D�CNx���B�ɖ�l���4rj�{Z�� g�x�^�=8H��)�T�A��?iJ�|����ܚ�I?o�1B/(�`����w�����Jj���-<��� �,E��^+���s2���S?��M�9���*T��[)1�%�OD�C��&X)����x����x|�_4˓����
1���'ZO�W�)����Y/�av>���d}Q���XČ[ bE�OuKAH�z���sU�;?����̷pT_�i�iGRLq��L�oІ��������b=��O�+ �^�2�3u�U��)Ɣ����/ ?��ts����D��_+��^����~��\�s�}�	w@,�-g�׻7�R��>(�NJIxzp�x�[Ӳls�Ƥ�E��~���b< ��b�u�6%;$MHԁ>�:�������ۆ�?������h ��nd�p�}��L�Fv�����T;;�ՙ�$Ҷ%JES�
�s�P�24�}g��MR��3�+����x���ZSa,�xa䯕��1I��k����A�&��c�`!�r(2�,�j�.�f%��c;ebV;.�D��.�q��<���K�7�
� &
%�ò�1e�KW��~�p��,F�[Zfr>���$�*�/I'm��ÉWP�Ƃ����PH�9\�d����CR�lk¦塆���u������O��n�1�����n��?x�<t��޳�y�$�ۚ�@��/����#�@O�����r"b��&IY���!�����n4&Ѹ����0���WYdÍ��S���sD������+��O飪⹨$O! "5�1��J5"�l�@�r�=�E2�*N��t䮯��(���\��2�~(���H�BELȊ
��k\sS^l���q�����8.�Ǌ��t!�|��s1w%�����>=��<@5r��^���F=��z�B*0�s|5����	��mt#��%�Z�Gk��Y^S�@C%7�
\�5�t0r�&Ĵ@Сmқ�J�:#; ����k�p��)�݉�^&�$��,���H��@i(`e��b9�qD�z]�F��ܞ�AM��L>�r�u����m�����$�1z��V�=:��x�Y�{��VIY�c�mG!S�y���.ip�T\�e�^	��2Cx�_�4�����u: {l�^=���� %�P����vfn�����5]�K�U
���8�:o��F��>b�bdH�I�a�U@M��L0􃉊ϫ�5�e}�e�p�E�+�" ���kM��$,n��h�t�np��>����*τW�Ӌ�C҅+ʶ�Z%"�1B>e���z��y�i@P�>�j%!l7y�*˗�|�Z��~�Hµi���^�L�`Tn�k��b?摜�ٶ�_�67-��C��#Y��g�K�懢H��o2����1,�Uf^]j�W��n�I��bP�
�_�R]�w;���FFQh�Hq�@L�6E��I�
�ù�=m�Nf.���z>$2_Gv�yARy��(�l���5���O�٦���N��
u^�I(�|�;�vY�Ҁ߯�~y Tǎ.KNgM5��09|�g�=D�ɕ){�T�f�O�g����X �*@�I\�x�Jn�¸/�2�<�*���	:cЮ���l��#'5�-4<$�
������<6���ܬ`���ysok&��b/���<%0�a.��2��;Kt�cF��K��Ԉ�p}rI�Ś<�\"����������h����V�e'/+���凳B��+�psn7��ܑ���D��Է�y��[�暹�`ENY���]���HT�O62��!���Wy����+w�|)�ŋ�g+�ൠ�wz�bJǩ\�)��'�imD�靭lmA�<��=Jʚ�6�xQy�U�0S.@� ��x��f�-'����KD3���{��)_��,��E!�� �TpA�	X�_�8Yڣ��Z�G*�U�*A���SZgs��k����w�a؞���F��� <
o!Ŕ	4Q�Kdr��o�3U�F r�8�k��0�-5MAe���͜0nۖ��m�lh^Z�#��z��A��������+�� �ʇ�w*�>��9����C^����)Uǃ�e�P�Ә�V��ǘ�bLъ���`�ܓiؗ�