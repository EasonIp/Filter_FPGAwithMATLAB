��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|n�\&���&��:�lQy��x9�5�A6�Nv;}PiM�V���;�4�ݖ��`PrڙD��� :�Z��O��^Cw�c5c����x1����T�d��5�u�n�3QҕF�s�s�9��=��N�<�{�t���^D��<���`F�\��C2`l[�v;�y�Wa;I�����7x���W|��L�� -�'�G����j��B���Zs�׃�2�3�B(Q:�����Pv��Āv"yw�X9T%:c����c~�M<R5[y�q|�d����K��E׌�ɘ�k��Ϝ�B��������D�.��b W��௸Lx�磤�2�HQ2_����RH���O`��yew�MBW�{� ٨$�dT�m�u*��*}�o�o׳��c�;�+T���O;	�綼����{+�}_\���}����O� �;hh�mV�q�ʈW�)Ji�����e�l))��2K,�����JX��~�)���N��.#nۄ\��M�>�䌸���W�Ź�f�ؿ��Ɗ����-y�Y�6i���]� ~�O�.�֑F���B�s!�5��{��kH�.(q�1"�Tw=ix~s�f�d���z�W+PML�T�ӳ��ەQmș403��u
'���؇��*�<8�3'B��3�Y���D0��ei��jAD�2҆���ʹj���g�3*�ٌ�S�zsz��ֈ]Ϩ���������� i�o�T������Y��R���cQQ{>x������D0�Z*��^�8�jB0�t��S�����)C�����l=��.�iU�MJ���ϲ������e�.?�3���X[�1>B'7Yy�4�4���K�Sdm,?Dz�W��m`�j�s���,j����+\C~ ���b+V�$A�Q:��Ԗ�$�ػo�vD���q ����؊[�k�^L[/6	ä������JKƧ� �SLOM9�[���D���
�3���a~�FZ^iϛ]HK%�K_*ty�	|�����&���\9%߁��O�s�c�K|�Sr��n6mN뮦7�=�=p��1TU� ��(#�:�{�[����'��.����^)�=�L\�~m�okN�#ڤ�|�'#]/b�]֡LR,^�׃QBkC��HZ�`p6�N�N}�N=��/��Y���4\��t����C:8l����`�$�6k���s���h4�r��:��x�§�u�&���D�`���O��`��]�8�`�M_4����W��m*?���	S9�ִ�t�;"�~�#Z\m���A+��]XKj$7O���j��HܪF�ܯ�d�7�"=�RȽ8�WR�#|"���]� e'���y��B��KX~�`��ŢѦ!T�%�J��ù�X�@F6[y��(.	������
�^F��ծ��&�D�t%ʿH�������J�����K�����2��0{�^�_�i������T�	��0W�xd�Zd�2���]������M�W3ً��m1�}쟏�_��Ώ�E��qCB���TF��u��b�u��iP�� :A	(�*\ˌgΘhD�����dd[<�İR�z�1��vq8a����q����i^m�&=�4����&� �'[=��b�#'���?~p��w��6�phK�P=�]b|c."7ۘ)�
?���6�p�!���FZl%���2�E���(nf���ŀ�)���F`�@�q�z�v�{���q+!��Z���*H���S�Ѷ`T�`��<�9wʣz�~�No�b��&hR5��ʥ~�x6F�h�~��-�>S�!����C��,׆���E��u�&W���u�ڋ��B��5-�/(�M�͑?z���b��Ϟ3�M	l,�8���\-D�<]^)�#$���U��=\%F�5VG�g��B7�6
�zd�#y��T�/B�xv��1��&Э�0��8wL��`�&����N��p�F^ZiR Biw��.n%uqN�����!վf\s��@E�I���J���:OMm�L@Nϡڽ��<�#�4�����x��?�$W������<�%���eR���<��ŋJ5YI�C%lԡ.��D�:��*�_K�iuA�`	��tb+qx�3+��m�ϕ6�g`�:S��P�����e�uC������P����G��/b�F];ʭ���^B��Y�n*Ѵ�~��R�'
�/���t
ʀ�B�Y��XG��7� �;JO��Ƨ�0�3W�P8�T�;��ڦ>|��� \���dwӧ�\JF�7d�G����	Rh�_w��J���.H�s؄|�N0H���k7�~TL� p�x5p����fG�AU1`T�	&��ݩ�{�f�!��9��_��6"�|O'�n�~r���b��+�n���8mT�yI:�����~��෻���)���Ǚ�#7S)���L�.������62.�/kϣH�����?=/JMF���$��(�^�� �`X2���ou-*�����7���=N���J�����d��G\�n]}�t`���FNY������4�}�� E/�g�ra���r�Dn4Y8�R����ףH�J擯as�l��84u��^{E���tؘ��	Ac�q�)<`9��݄�U�q
Tj��3ah��MIN���޷�Z��󟏨}1�Y�֏�XF>J^l�`�hG�RB�j*A�O�����N��L'��°�<<}��B�s/+6�>s��N�g4B�������X�W�H��$�Cb���(����=�,I�XX��SN�Ʋ��q������M�q�;]g�����K>���4���z1�Y��z�Q��5�^��d�SĨAb�?��c/�8Q%������R�WS�����FM��KS�7�@1���g����ܡN'�n7Թ���x�nCW���#�J�aq]���!%�L^���cTY#(RܮM��/����g�����С�2ä�:�#=�"�`��+���ı���~̴��ie>��җW�f��+�y���̶���Lnk�J�e��Q�eH��-�?*�(�N��ޘ� ���:b�6��3�₂-׈�����3�'kڧ��պz�O�r�J�4$J^��u\VՏ}���f�<fE�n|�k�,7��>&���i�ʗ�2em��I>cC�V?��ub ��FnF���:�ƛ�'Z��,�ע1~ T��~� �@x2_Vu�_�y�)(��]���Ok &�r繥��}��㨽^�>m�]g�8�Վ����Ÿ�Y-#�t�!�`�{wr:{�(���7'�q�@I�%?H���F�?��]��)	L�"u� ǇI�d��0h�8�R�����y/��8~�6M��鮞Z�i���-�Y���Z����1���ب5��22(i���ד������C�sWE8Xc
<��{qߡ"��Uշ}<N��h�e	�2Ш�c]���(?��l$%�	|B"�<��?U	KY�7��[�`tF`V3��ًآ��f���Ò���y���M�@a<�=�?�:˕�W��:�ot�F8���Y+f$��wk�}����B���?����6-��Arj/@� g��k�������#b��0�c2�	�gJd׆c��д6X�6��k�<�H��՘�wA_;W+nmJ�	5�v�.���F�Ek���<�q���r�^�:H�7��4j[���h�_��%&y#$�%��: I;|yX�iˋPHy�R#�_�2Qz��^��.d�����fց.��<�F�_9�(_�8�ǸDR`���4��n��K�Ί贶f�XL�٬-�)W2��� ��Ɓ�3� C;���m�7o�5K�)])����TpĨ=�\����{���
��Ng���Ȁ�AD+�6�W<\��V�T�i\(����3���48s	u�z��c+=���cm~�w�Nb����CV���2��������'�kX�0ă� ؝m�-��e��r�Hh=��2Jޕ��r[��m���+�
"�|2��F��u�m�8'�4�K>p&hwWB��n��%tR{"�BCA
��T�H�g�����>j�fr��~`L��q�����C�Ǘ�Rjs�q�vFBi�>�
�{�Ü͜�>�%��^c����.i{������=^\���<�F�����),��Y]Ս�n��$ �Hdɔ<"$�v|Dz'�3:�ݔ}5�\/�m���^t$%�lh��Ǜ}GX'����a%�Y���v�d+3��O��|���nD�sqg0h�2T}	'w��oj���I$݄QJ�n�����	�7�=6���ki#웂���=�
�$�B��#�pX���� Zƕ��J�	ip�F���Cꄌ6�Mj���㸨��&����@m-�X*YR��܉��e�z�O���b�'I�f�hF��H�T�����]�Y�}�0���[���Uoޘ�嚅E�H
X�ݎW��`7B��d�S�:�r��UIi�[�t�Z�\���|�;#)���I���va�%��� ������2A�|0:w��^{$z�:�z2w@��=l��$�L���O�4��zĂ� e0d�>%�N��G�Q?��M���h�1������F�gC!A�su@��y�@��A?�f��X.[,��p�(S05�`�{N8ZT.����N��ڲ>V|)|H�M<��e�B�ʮ�oh�ô��9Q�<N���7QA��h��!�|"�����y}�Y�Qow��*<96�]�($uh�� ru�L�7�-��0NRG�b���.�O6󀭢(����� �^8����w�*��T�ZJ��3"��3i�]�7[�� ��dg<�a����l�����$¿\���怊�f����w�H[ڪ'K�7ܦ�EFb�~Y0w(��1�c�����l�����;�|��$��h�g��A:@�i�i�.Z�'Ǫ�r�c�%�b�8�:�G���B=N+���կ�4���zt3��/7�����x��'��j�=��\ȏRa_1�y77���R�zI݃�2�w`�G�T�H�c�l��� +��{���o�tN1p)��A��e�y�$�$����C]���&��XU.�H���?!�kD�������)t�:����q2�`��z�T_h��������R�l�ơ�An�]ػ�&%ڙes%���j>)�/����l�v��,��up��H�٥�C9ƨË��ey��:��p(dv��C�6�A�sT�N,���w֗7a�!9=�-��j��°q�Ǖg�a�\ٔ}����a����d��"V	fF�5�����ޫ���.��n�/��>�N2J��]E��l���Yy =�+G��S�������ڠ��ah���5�SS?�9���T�Ը����q�����P����\l
grz�<T/�9`8����+��f�=�`Gr���i{�_6=�e����S,2®��o��%�q�M���Z\tTo��w�yd݉����.;^8�\yT��=h���`�uϸ
h��������vB�K��~�!k�K��L-!�h��56wq�.Dr^�(3qHv*���i�m�2�3���,2�u2�3(��Ç!�!y_^���0[�3%��e��O��?mH�.	���g�C����i(��@��+;V�O���k��:@X��e�`�U�uԅj��l��d{��Ь�X�]���ˡt&@Yjh��eg]�
�k�u�v2;��[�YPiUg��q^�r�Xr��Ɲ���~��Jz>}�����-,VL��éZ��݌s����	�l��f�$�p��( �i����ϖ�#�H��`�Ix�x�T%��x�-n$�Y�����&�?��Ɏ&�3-W �13�we��w~�B�8��3��X�24��;>�כXnS�Ab�mV��iJ�Z�N}���������2c�oZa���d��*
���u����e>^9�����̓~� qT�d+�1Xe�"i�(7E���z��L
9��I(b3Νڡ����?˒G��'�o4��k��Hm
�5)���.]��6&�`/��C�����P�J��0���⸟��m�bj:Գp\���V���)ҙ΅5��/J������[FsP)b���!^�`� �p�jĞ��kG���qr�OSK���H���;b+�+�[����0���H{bܽ�Ro�i�mqN�m��}�V�/)s���#!&~^hp���˺X��t�]�=�����05ȵ���=iv�"�#�����<֛�}�T @k'r����_�4Ff�"n8Ɔ�mu�"e�lx�%(f��f��QliZ������bɟ�W"�t�OY�[�7��/(~�������A�B��%6L��� ���u~}Z>(�;û����}a�G�����\�6�GI@G�m|(;���/v*�EzFqcY������Y��tG`�?�u��{ǽn���+��f���WQ-	s�tU�ߜ�޵��Q�QN���D�x�Ӿ_�h��P/�������6�:�14>,��vڥW��b�N�i0�[�e�:�@k�H�|��r�@���	��$/�O��2%4Fe��&T��:=�+�z�C���8���*���d�)&����>�Z���n��ǥ�]����5Q�=�e��E��
�s��Z���A�����9KO	+��K���5�`+���%2���r!Y9��8��Z�w��r�\s��M�1�I���ȡ�Γk�5�y%��m���SsΏ�`�)�l�j�M�����~��1\��\Y#=q �2(���	_��c<a���r��xs@��Q�>�t�K����=�ɔ��MV��E�w.�%5̴ʖ���T,��>���U���L����<2����;��ＪS0=N�,��m��%Bi���s9�=)_���uTEh��ıBb�P���8S<ze�e��QD�kA��.��[���A\U�o���P���E "���H�����d�m��Z�Zf�Π�����L`)�+m�V��s�]�v��Ja�
���):���_���J��N�Ph���D,���k �]���~cf|T3�$!{yV��`_&��z�ɇ����xS,16��Q+- ��دb�E�<�%�SgA-��W�qcV�r��Y��6H�n�}�ezDWX'&����x��w�����Jʘ���V�-�?UmOp����F�9������6�?E�!/�	��5�1�:t�wp��6k��PH���tv7�n�4�A�"�Z��Ou�'�=��+6�,<�l�7��M��U����(Y8�쪾���e�eR���v�iү��ɟ�SG"[��N�����h�Z�*�!W�\{=-�Q��0?9䭝7��}�����K���I� +z��G��솎W�����q�,"-iu�)��C� �S����@�	^4�~�`n#��57��-��f�4��\�$�:�J�G�y���Vri,�2�W%0�f�$M��ٝ(x�r���"ݒ�S�lu��>޿^��*29���B�p�z�ī5V$;�u6xԺ�t��H[�)��`�~g�f*�^��A��^�0& Č����;-�M�>$%~��ݎk�L�	��"u�FZ�"�q{)c�`%�ZC���Q�x�%��8�6����X�HM��2Ȫ�!;09��5r�q��ŉ��g饚�ږ�7��L�J	���Mo2�Q���&]c"����k����Y;S�"6h��'IC��B�=k����Hs"��y^c�by��g��Ee�1�)�ٜ�r��+�(c�Y�ˈ��oo��n1��4Z�bP��cX��j̆���x�͌��OQ������,���Ep�����`զ���>K�ok�pT�� ��f��YOe`���f�h����6�JK� �d�0��}�&��?	�\Ѽ
����~&��q3;�N+*�HGI�^Y����^�֡3��A2�6]�#��^��@I$k%˛�R�_1��� ����pZZ���DP~$��_��?��s�%+��VcOm�Ҷ�q�C�?@��]F����6�y��F�y�W�������i���Л��jye�V����}��^H8$���2/n\N�5���Tldɸ���Z��t����摓	��[����Lr�1���r�C7��Td�a}1�*?^o�Њ4Ӷq��O��6 4R���^����V)�4����A��k���Qrk�HJf>�!52enZ�ľ�!�9�2�K�*�2i�b.J�u����X`0�[͉Թ�&�����]�L��
C-�����"�k�M;>���O瑄�&�)F���ʀCO��2M)�[��%��.�%���y����<c��V�W�_n?Q��������	;���Umu�
Ή�(U�o�s���IͿ*|����
ۜ��d�vu���}��Taɼ0���g�����_����?}�܃?y�?���q��C�L��I��Q
�����I��([ܟ4L		�ܤ�IӜ���Ev�>ə�F
�l*l�bd*��[�S/e�,B�φt����#��Z�¯V%}�y�!��Ҩ�cdg:��~���=t��G3�;:�D�dSga��>:[�c�#�-����*8����$��ApNC}G�H�&ȥq#�qW��>��f��'%؟������F_v>-z��r��Qk�)��?�-� Ld^�=~6i��T�9�݃��I�5��0b/�s�_of��AY+Fo��sR
�8�0�!��dV5���C�KS\(hW�F�W�\|mS~��&x�Bt��6���8�ry.�L��
�KX� ՙp-�{�vU�$��3�[���=�fM*�ǡ�_���N�}��W��̭@Ƽ�,YF�nɬ�������^h���[!�C�ǭ�P:�Oi��e��f�K@�=����qq��^g��;��UZ���V�Q.M����?��i���Z���1F�r�/�
:5E�^^�����C�ҿ+�^��)��+_k����g�:�B<92�(Z�Nȇ������_�5�a������rҪx�bj�h:��0$�`�f��(^�Y��M��)_����e�WB���:+�5d*1���+f�} ]R��e������Ű(H����ǤW����3a.�Aݤ)ro���,I���Y��>h���_$���t3��M�0�O�k�|�4�52�!(���qc}i�� -��eO���^�R�J2e-X����>�)M����������I!ntXbP^s	��:���B
�3f_!�aU���/X�F�g>g��@���`��3?M�`ZJ3K�	��r��~o�w,���ʵ���¯2w"�!WDбN��yӇ9-Y��f�d���ɲ���*�g��C�������pv$�X�B��䎁��gFj)zD\�qQ�	�w��m�x;N��Y�t���^Aq�r͕pY4�%AT��u9�0=y�7U̜ UB��>a-̒��(�r�
s��¢�c�m�BJO��O��}����fs*;Z�Dw%�J�u���%x~h5"��k��f�v�,DB{������C�>�%��L���s����mң���hC�6!�.Xw�������!fqgMZ߇w ��UMt9�j����t5�Vmm��{\�+��Dኙ��c��[��]~n�3%&���of�᧣6�Z����omLƆ4uՇ�����d��9��$���a������Z��4�8D�סy�)��������ȭ���%�Q'���Ÿ�h��P�\2�,��� *ל��-5��0GD�X��ә��Sq�y�֑{�V���`�g�]W�'�Ľ(�6+s��Ps��qK�y�ڈba8�DU8,HB �ͫ�Br��F2V�=�r��Z��g�lI�HƧ��a�e[p��S��H!��VZP�aۭ./�����~g�7���p���$+��5�cY�PJt�F�7'K5eYZ�n$�%�� dWb��y������v�j�`}�h0ʅ�O�$�D�؁���`\M�Hɭ��wV���!B<v��8�Aj����HU+�TQ�($�!�D�Y�9�����#W�����c�}�c�kɦ��<�u�8�f�O�($C6�r�i���{�a �����~��&��E(^NR��!�ۇLtq�D,Ơ��� ��g�b�wo�eN����;�>�yD�:c����
 �t6"k)fah�>���h���̀d���%s�"�i&��ش0�qX��P�3O���P}�v;x9W�1�${c�S�~�=�ЇX�+�4���e��_|R;��{�kC��ԫ/T�����&�������UHs�`����o��k�,�νd#�����H/�"ph֮�88��.:��F�G+��6�&_�W��b-�bV���>`����Y�~h�iu��h��|��_X��۵�Z�X?�����[������7���D���ɻ�R�>��ؕ�&�)�%��<�{��~�(�%([8��^�P�g U����=�����PH*�&d���� ~�9��T�r�^p���ﺾ�O~R5d�_8#��tn���,8��T��g;{光��}Cه�x��?,�X��L:���I�=��R�u����aצ�k:I�IN}L��/�N�#bs�m9;��6���
����<�@�I��j/�6��x́��8`����v���rg���~o�W��޽>�~[�L泊xVJ� ���E����e��LqAi�Mo�����eA`�g��K�6,e�3��b#���@���/{*����k&�Ϥ2�Ԩ��0j��۬�!q���"��Y��KO��*�@n
g1�!c�������4�u/�=�Y~8�Q��޳��@_����Rm������ë����`�}�Ő�m��W��V-�L�%�_���@ڌ$��� 8)'�l�R��+�g���:K����땉�^�p��},�V�hc�_�Tf��S�!9z7�&n#�ɫ7j/����N��Sv@)Eq~m��v��8~�����"�T�9ʪ,�K����K�C2Uy7����,Ϩ�:��.0a����#�Y�v���L�l��(up3�� 692�QDd�{�=�(�fG��A)�Ay�I�����R��_�\����s�{GS=Z�K�Лo��9@��yG@�2��K(��|B��z���8�c�F��3�(>���%������V~E��=EQg�^�F��*<$�^���f�W��m�$�5&8mRȅYM��Qa���8Bsn+��q�NĮf�[�%f�ُ'�����!�4;��9A�]�F��ln��cޏ�z�r��6J���R�B?���Oy"�p_�9b�͖q%j��V��h�i5��ے.YQ�ҵ�_<A�����ݟϦ���t"���mv&�g Q�jR>^��|K�9T�6)r���\S�2ş��1�����yq�8?g$M��io�q������g�����g(y�C�]X��=k/Pr�Ga��lM�02%>b,O�$���\�e�m���4�����4���E�~Ɖ� !����fѾwG2U���A��d�:\��H�<������Q�s]�2��ܱ��P&yh�~��}�)*��ij�!NIc\W���Ǌ��i��fr��x�er(�G���~�(G�L�]~U����˗%ޜ9�J+���gɪ�V���~�1�t=��sĀ�Y|�g~�suDkA*7��|M��h�g�G� ���Z�Z3����Rs�����FJ?�������q����PC�+Ǥ�2U�*Op�<�. �?.CFs��1|w�����B��@�*b����!�pdh$�޽5����FQ��Ca���:a��	`c����i0勂�oT�z�'��*#^.���'�<���������Z}Q�Q�vyT�~�غ���.�7-��S��Y�u�d/����9Vx��Z0m�[G�4kY:�n�@2�Fd����@ƘA�x�P&�]�̨���_]Ov��du�����2��I�2UΧS|U�K���.���!�X���!�g��"��xp��oǛB	�E6���3���y�w����v�9����L�����3�2�G��՜��!k:���5ϵ�E��ݻ��g�,!�7q���l}��'�'wЙ����z��ʫp0K��+g��k$Xݮ�z؎� ��+�R���Xn	r�e�M�4�E4P�I���U������b|�V	�F�����~{���C�J?&g�y���e���a���l�5?�z�'�]uFdd�ȁ��.KŮ}� ���96*�=��àk�d�����'����l`�?�Tb�c-�M��B��	�O�f�0�:�/<e�����(Q�Rޘ'e�Z�{`-=��ڛUI<�f�c��0N�(�թ�:)�T��&R�A�H#�_+�{����gkP�v���,�
��	%H�����I�Ę%�V�V�Ә�����8�P}�����VW8�,3?��L�����K
#Nh�ָ�o�����B�K��]uqF��(�sft��)�RT��!v�c�o�?ֈgq֎���z����c �rvE��׈��J�c������b�ғ�멞}}3�J� �� r����3ՋV�{xh!��|��n(��p�h���a����A��E�oM��ւZ�x�g.��^�#1�ϸ2��}[iqZ�(��pc�>������_�<����?t^�D6nF�qC�����]�ƫ6cMb5 ����x��l����p���R�>�D�H�P�pi�ˈm9-�ΔE�b�te�u����GEI0�2lk:]����ȸ����CЕK��3"���o�GŵRk��յ���$3��U񥲧N�1(P��ޘ��FCKZ��_��������@�� B�q�q�F�������@G���d�;-�-��:2ħ��;{U�Wv��6�$C���M旦�t��r�	����!D������q�y�!;/@W�LA28�W�&�(3&$�EE��J��HQ�gV{���-K�N���z5Mn������o1����k�K<��fc����@�@�tSZ(�?�6�3h�#�&�p��[��j6�Z��7R������
�c%��> e4`�b�{ԝi��E�7Eo�:-+;]#���.�NX�C�0j�d"��HIm]� ov
���Ŋ� �=6ChO� ��i��p*`\b��"�ߟ3RM�M�����>s9x��Gh? ��b�</�J���r(I�TƧ�������*=b�)	*��ư_P�����Q+�����038Wq�Ⱦ>�_Mۃk�3�`Glh<Req
�(�����4͔-�b���=TM�A��2P�B�	S�����"�X	N�������m�V��"�e>[d��K�.�u0���ŕ���5^�Ff����1z,����xFMF��x���j��'���tg9ذ��H�Q���ʲU�Ԯ��@_���n8��즾��e?:�<���}9�wW�u�Y����`�R0H%�)ㆾ�.L�� ���GoE���ǌ<2W/�)�ҩ�a��j��I�$¯�M*�
��i�e�+�N�T0���z���B��a���M�.o9�|}��B4�,�3���n�P��GhKl�&s��Iϩ�C����rN�+����ķ�I���7�3�R��~С�������d�S&u�v�m�T�-��:��s�o�[�;��9kg�'���-���%���g�K�u��M��`��������
��;v���ӽo�M|N9��pi1TW��*�+�OI�� ���T|4��,��R�/���5ֺ��o��^�Zn���}ԂB6��Qy�1��
�&�6���cq�6�`��u�P"���yj�Ce �ulZ��e��}��ے�߭�dXҼ�k�D�8 ���I���CF���q�s��W���lհ(�36�b����C�Xx���]J�	5.��Z"���EaKc�nւ��3.�?����Y�v|y3O>�L��Ē1#F'K7W�_�?*��w�.h�²��qD�������I��RA���o������4��������[�¬�])��ruQצq�^� ,],"��/�1��e,���>%gX�3�V,O�ٲ�`�7wy�`��.� �|�,�GP|����$���Qr��+��<��A��M$���o��בL���+���#+�t|��9Rτ{�q5��^������Gzu���ׄqel����&����MG�E�@�����C�rTu��w��v�	A�D�{A@��Ry�g�Ͻ7_Lۆ��+���ߓq*���J\�!�n�v��f{uТ�}�2�o�خx��Aٻ�v��W(�j
nx�	��LG�JvI0=W����=�dQJ�T]�2q��e���k62~���|�D����w6n1 ���[[D���6��E��<ax�T�)�	3���3s�/�*r�-OQ��(3�(�ᕉb]�~�Xoy#m_L��R��Hlg��`�wM��M���D�<�7���Z�]:�E'�aW�����X4��$,ȃ[AO-� $��c�bp��������f���(gf���')\�S"|�I�;D�\�d^��=�hA�Q�XseoS�~Y*��©i�7�]������Y0$KHx0��^ٚ�	��)B��Ϝ�K6��#jK:�(.����s�B�=ι�w�ه�Z-d���w��.����o��NݮU�d���̂��3�G��k�\sh�a
W�u����	M[0�49�,�0uz��!̤I��ӎ�)����];f���k&ă �ou��X`��(տ���
R4[�!���ԏ����A*�7d��;*��q<����Ҳ�,�L7���sDKO�0� YZd��hB��ln�}H�?�HQC�}L��Wm�@�?�C���g�M�P��Q�7���7��'X���9�t�#�����('PS�$Z-$P��}�uT�O42���s�w�|uX���y�,�A6��w��|����j��LK0�P��%Zn�-���LC�Fr��H�Y��_�?M��c�M:�M
E�?5�B-���z�eN��'HJQ�g�V  ��Sr�H��1R	ɏ	̜ϵК��Ί3�Tdw������G��p�������E�a��sP��Yx<َ�s�#�<#c�h���͏;��
��	a�;!W����"}