��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
����Tӂ���^�2����+t2v�g�VU�r�H$�\%8/�!8�1���1,c���'���c l	�� ʁ����h���z%����\�?�;�=�6����w͸>/Q'\p�~����|��k﯃�`d�C\br��a��D�z)*�&fV��X�v��H�F���i$�MJDK6�#r�n��'�>ro��K��[x�?���IÚw!	�K�D=2<�x,�kx��s,ŷ�v�QplC����R_)�|�m$�L	�cߡPX���:�zI���H 
"k�6C���O�^8r��	�RؠN-��~��-���5>�*�hbD�c�D�Ma"���BRҪX�F���P�wy�"��=�댣�����
��KY��Nn��o�o��\�������-��'�'�?9v�i|b-��g��R��i��x>����	���Z��,��G�э�i�ʫw�mDT1E#(/#<S���c#E�E$}A;F%�K<��`�Ɖ�o��<����9 Q�ӗ�vg���$��zk����顛�Jt���>���.����U�!B��'o�{�18�>���ƽ�:Ӛ��������!��(�!��`X�2�3?�s��;!��f�	�ɉ�jԷ������o>2�c�z��v��
·�{��S�_XSw�h��e��o�o��߂�K�Hi���mb���ܣ��M8$ő�V��B����[_v��@u�ԔV���.J!���H5fG(F4��d��ثeS
.���T�����V3��[{�7a
�[[�wy��e��^^`�2��� ���j�9�Ǥ��O�,W�x`���f]�o��2��dPk��ESq�O����Y�mM�Z�r�<oȯO�$`q�z<��VN�, ��C�|�����jt�ė&�0H��6n��������_S��������8,h�%3��l/�f��P=�q�_����X����`�4�(��D�4�}/��POXR�����Ɣ�p!�Ù�́RD�J5W	�D��'YW�L�˪��z�C�(.�X�5Wa�f�+�T^��A�P�.����� �O��M_�=����C��C����Y'�p�� :�;b�k���bo���x1ƽ�7/ /��֢���HӜDÉpw�	K�e�& J��ӷ�Of���.�� hk$|��W
+�L��$Ff,�MxH7�ԇ�3ٺtrӺ|����\r*+�\@�g��������W[�ʳ$Y.Q�[����h�)�ҥ��(?9�?縒�M��l�\ҺO� C|�|�oC%��3__c�e��X6�2��)�DW1��U�<�q
����U��
O|��p��f�c\�����������w����c��6����'�5G�޵�������/k\_�FzȜ�N/:FTc������a���Ӊa+b���3�Qs,C��Þg�O,)$���h Dpin�XEpT�%�ָ�$Ϭ�QaFZ i���,&�<b�e�v���C�t�^>{��%ar-o� A��T	��Hx�Yv��s�0�ʺ2մ{*(T��z��#Z5�E� ��c�6T}�N��h������)�桂�t`��/kl���>X"� ��e�k3�6D���$/�����idR�#�OIZŁX�JmN-��q�ۄ�a�SL[طh�r�� �2��*��@vͰ�I����`����ɫRN��#'_����4N@jŏ����v%J�=Ed6Hə��z�����K�lP.����r�y�ߺ7f�7��D�H��yB7=�Fx5X�
��E��P����F�;�\���S1��w$�v+4����T���s
M�9�ƌr��������/�aCd�N�r'��e�1��E��vy�lN�粃Ķl���Ƅ5)������FU:s��Nњl�g2m��8M�uյ�8�Z3x�oɳ�(�?���`��T]���`D����U>���$�'ě~���ɞ�ݳd�_�kJ_mM	�oV]1G�5�����F�sK�Ҟ^����	}�cͲ$F�����NG=�TJϣO�����g�&H?�c)rdODO)��C'e)>r����	cQ��$���B�����8 DXYOI弜^A�����܈��Wմ{j2s}�sv�Sh��j��]�L}�q ��갇�m{��t�=C�XFNӛF8/���B����CTXjg���a{��~t�]F�<G��3���d7���T�i���Gc��`�;;�
;������UP�.u���[=�ϸo��57)I.�r�z���	��>$��S�~q�QtY�U�'��i]^��Č ^Z�����%H��V��<�����D�A4��utTK���U.gg7�vh+{Hf4���f	�=Ä�$��~':�D�.���7�bg��e�_���;iD����N�	Y	;1K��G�B��)D�]�}v~��Ė'A�l�M��A�c8����7�h����E�tfn!X�_>�"CK���6�nJO�_|�=���,�M~���c��ύ�t:1�Q���oRN߲=�� ����j��!"�=s�-�B�.�������'
�~jw��0�Ⱥ�26:e��S���& ��l��(໙Zz��|R��Vw�����e���\"�)G�Ζ�	qp��
3�ĒkD�2�Ȥ������\o���t�M�04��S&�)P�P)�n��U��Z�o��~�׌J��I��'�� orc���P�#�OI�_Q�Iw�v�O҄�,5ψ-��ԼR~sY�������t��a\��o7� �q�냌�D�B��y]�^�0܉#+���L%��A�Ce��~?�ĕ��Hn�N�I��h�����|(m�^�O�v4�"[�e��.�,��>�!t	��!f���9��X�O�����u����,K��[�����x�y�������}���.������{����j�JUմqmx��ɵLB!�۷v�8M�����Z	��MF��m�~y����)8�obE�������/��ty�O�On��[��U_�Bp�S��f�����h!��n*;�����t4�s���˼bo��d4�*g7��pG̛�a��܊�A��#Ѱb8$��YBR4��3�S~C5,0]�OK	��v��j��%k�������yy�� |���?Mv����M.��}�Νh���9��V�.-X����X{	��߈����d��_��I�H�ن(��
2�L�s<��`��l��0r�&��ש��t`��}�P�P��M�h�e��D��1B�g�Q�
�����&�m�r�a%d���E�*p��*��՚��B����=RÓT�K8{L#k~Q�̫�t%1��,�(��_�2�|o6�/����ڟ�#��� gιr��C�o�g���#!(�K����?��$Ud�ZGՇ��:�݄���
x88����C+�����4\�|� T�����@����M�Ȱ7`}|֗��� H�����ϫͩ��#W �ZO�J2$=�~1�7��,�_���
��l\�~w,�U�;?��Z�9�����mu�z���~gڲt�Kȧr�������^5|�a��c��>7ZṦEp�\w�=&� �ڽ�e�1��T��Yi�S�&N~17AB�՛��/�8��o�����v��ˀ֛dC!��#����%�i��W�Ⱦ��n����4��q�MU3�G��s@�W٭-�4���S�fc��[ع���d#��|�4v�.�٧#M��_~NZJ�vS?��,�4n���.�!�*�I��}�S~hOho��xEA�|B�F������X~[��4�|�]d���s����d��<\��(���4K\E�9q�5� o�\dݧI��f��`���0�WfadG���jmr�&!Y�k��Ό�cGe�ke��w�7����!rL��6K����v�(�0��^x��D���l�.&��B]!��c���8���\����z@��G���̢���4T��0��-�?���
�Q���|��
1�٥�$�K��h
�k��l��/gd��y[�@�g���BK�g��\e�!ac8T�ıP���`��9;����'�5�����xIA�O$v"����,���ܐN���6��Km12YbQ
:=t��1��X!�G���j�>��=Sd`^�B<
E, �sP�%P�ƒL>Z->0m�k23�u��(�݁:��ʇ�n��j�ƂDE�b��S#:h�d(�z��
L;�Ζ��L�����B|��|Ȣ�?�"z?��)TZ��aFڝI��h�����H2�����m#���!#k3F_UV�,�+��Һd�pZ��U��0A��
9n�L�v�7�jy����ƭ��������a�<Vz�KS�tWd���}ADc�����͊��u5�\;����i/�"��S�t�0P�k��p۟*�'�r�d�
�w�)�m��F�ݽ��.*��$��QuH�\����P��m~&�oԵM}�c�o���8?l�^~��VIKp>j����K���Q`��'3���/���j(��b����O[B>�|�f��~i��4`��X��-ˡ�"�<㉩�`�����t�tr�(���:�<�5�wRF}Y�l��A��;S�@FO�eЂ76ɓ�����(T;���'��Kɷ�^����¼,�]H�ev�,M!F���{"6�"����D�g�0�}զq"�4�ق�~|���jw�
Z�Lx*[�Ԗ���+ů�af��p�����<k$A��z}m�:�p��ؐ{(5�[��;pG����wZ��M2�]~��Gw�8Y}Dw�}��h�ʊ&�WI�wj�3�G�l�o�8+�y�9�&H�=��te⣗}3�KZ�zE�VU�l�3���X}b�ை�Ȏw�����`\�BB�]$�@/�����H��ZI����&��7�2�E�]����V��Jc��0,�'���1����<��"7b6��K3杕_�+������+����pS���3�,��B�ȇN�;q��悙 �Mrj�ش�!�9��υ�a����6�p
�|�8�qc�V�"�S�( ��Z�@�G�M7�'q��èp��}EX���J��c���QԈ�@ߌ�
\�N�B�R���h3{��E"b��z��z\��6�Qb�/L��[|�����H��!�xw_�m��g�����Q��,1z	��T�gQp�T%WM�~ՠ�7Gi!����0�~EW=�+OrQ/��]
@����O͎�(��cl^�m�Ґ yp֖��=�ڣ�'�ǕR�̓ڊ��e��g;oةw0n��jN�����g
�#����R�6ޟ71R�������b��˾����C@�Y�6��j��b��k���z��o ?Z�$�=��n��C+
�Qc=�ݯx�����EP��� ����h��sn������ ލn�����I�5u,�F�!7f����uC�+��d�g�MY�k�5����X�_�	���ؠ�B�*�����|���pyJ?��ӏ@ܜoAh4��Rq���+����Wv���X�y��wO�<��	5�v�ޜ�ʶ~t�s�=�`%�ξ	����8�`ƽٸe�ʻ1�J�X�[l��:��B&���ˠ��ԠO��gγ�#��W\�W�o]7߻a)Vyw�UUr�XK�{~P4�1��e���:L�h�G�b��`�&	R�ܬ�9v��Ϋf=u������l���:�h�ˊ�B�UD�'��l�0�z[�~5lv�9B���M�\�t�Ʌ%�v|T�;a6�n/��L ���!������G ʐW��V�:�5MU.�c��SB�� ��s��rՙ��ͺ61?J���Ą7o
Z���PT��E{"OXR�;�ԍ[����r]{���1��Ų�J���o�c7#����8�-T~�2� �������8�W�&���<\.kH��������
QƱ��:�C�8�"v�Q	6rTD�y�M	$b�q���gtD_�`+�޶*���A�-���tǉC%}	
��n����`���@6�?��v��W��f�kKu���g�����ĘmM��T�)�ߍKp#���gsy&J3��|���AX�H,�RB�q�4ɵ��=���,&Ɵ6��՛&#�����?�}�g^h��LSظnʅ|�߻]W�ɚuI���ڈ#�e}^Z�)�U2`$���t�Y�k�`�+8g*�K35R�_~���:���+��������+��T�e/�̧tb�h��	��|�N�T\jk����2OCN[{i�(l�P��d��2���L�[Y�Va�S�~f-n�L�}�`�������iSD�㩂�{���	}��U�0R��T�W�  ��`��vE	Cr�MR�ݲ.Ҋ��?�bVat�Ե���ڥ��
�������)�s�6xDM�h�vV��,���di����H����;ǖBL�ߪ�p������A��pu$��&}��g<��\��,��B�,��:4Bc���U�x�f=4|��@�Ĩ�мg��mC�j�ϋ��[��}>Ǹ��ڶ5���%U31�*��Q2�;��-�wd�N�g��$�D	"�#^��(8��w��*����� ��M�gC_-ɗ{�scQ�GV@�r��NQI�)F���Jg���vr�kA��T+اbΰ��I}>�I>����̩����p�D��P���,9���>�=W�m0Z\��#-����qS�J;L8����n��x�l������oҋ��ף�S3�����%w4�Ē1K��H!n��Sb@_��$��BZ�/��6b�6-i���4�3���]�s�SM��=��y	�R{����D�91[�F ���n-���
�&=A9��4��c�s��+*�@��@]&��XUF������Y
k#?�LA��3Q�.dp�PuCbXy1��.�J�`��
�2�������G��G��DT��᭣R��=<��߯��Rpp���HdO˱w��^��	��],5�]b�i�(b��#6o�M���>�I��gՖ���Y�)3�OL���6lrEy�`ZA��2���K�f��-��o��ڎ�MV-�٫�'a�-��lWT�o{��K)���gE���'G��(6@%c�����͌5��鳦ڔ�dp��t���}I��ɦ�9b�@�!���˖U	��h���՞�Oa�t����i����?e���4?��"*T� +�)��[��6����ͪ�5���:��p��x�G�ic+��k�ͩF�YG��b}y.}e+q�X�~�d� }�>򟕭�wk�O��(�;Ku�>��Y��������&�$o�%�;�B�ӅN���ܲ�o��V<��ͱ����u_�n���l}yO!�o��*X�I3\ʵ�5��]E�fy3�����<���|���G���z��)O�'��j�\��o���O��UA����ľK�;ҥK>��}�ZIF5�I�5 �]��(��>wnup(9n}{�&�]߉����F�� ��� �/3�T�'8�5�4� )�L8qz�~����d�ts��m�Z0�7w �wnǈ6z��L�)x'/]�7}�k{�*�l�L��h��mN����/&c�=�Ż �/ T�&�^���a��m/Ϣ����6/�ΰ�=d0n����R5t���=foH���y�8�3�c�����8�X�d���ݒK)>S�!Shd	ˉ/L\&ۦ��b������m7��-�O��>G�I�M_[x
�������W��kد�/}[��=��r]��)=�t{T�����6����݋_B�(_o3��\d�c�WJ8l�q��w�睵�k�e\n��x�=8�DP5_S��B�j�G�KZ�]� ���8����+u�AW�u^���!{��1�̓@W��r�(�s�ƭ6�X"��)���:r����Ig��"n��​F�ι�d�1�ؘ���ɫC䬱=���\�Yu������Nm���m	ܼ�P�J�����il�(e�*)O�@�ܹ��wd]���X�p�3:����>B*\DT�5��6�������7�����D5�Xbf��_d��>�Cx��<�&��Uě�:�,�W㊙���N%�6�H#�����Q8���T:ɵ����E������CER������'��5-�(���:FoTꑁ雖Au�Sϸh��*ț_�@��_0ʸ��eܳ���&�p1���
�]��=�y����WI�0i�a|&IB{�vvb���S�
���i��E����0rz�Q16�@8�spŰ��_=�/�s��_Q���g�>=o҃^&� �:)��R�4�x�?�J��2�����iD���)b�Җ����v��e��wKVh����b�e�(!+e���n&Y\HW_�z|U�o������Zb`�c����cǈQ�t_�½�d��ê"�T}e����ʗ ��켛��������(�.�InC�� �P������i@^�pږ��vΣ~p-8$��Y�k�5���ŹT��Q������,���)���jؽ��C�e��o[�Z]���yd�g;�>�IQ�+*Gz]��(b������zH}�Q
D�k#4Y	�8|��0�ھp��A�d�$d4���=.ƅ��O>���+�Q�/k̉/�7�E�"x��:��HѶ30*#�<,�B%;��Ywr�M���몓V���?e^�#�7v�=��K���J&^hf���w�\!��A������|:r�L��G�o0�Z6j�^�*O�o���t�]s:	՜2E��w1~9>?�_lY�+�K�
�'����
&��%e��QB�a����A�J��~gҿĘ>�5*^�h�k��U�0��5w馡���d�Hܛ;�L����V[���E�CX��
'���^ܳ����}_)�6;��`�7*��4��ݩT> �O:�B�� `��*�F�����+H4�!��݂u#;�U����!��)�*޼�Ѥ���^[�V�0&jtF�Q���H��M�)e�/,ބƏ��@=�莣t/x_؎�'��g�&k|Hyi��"x9��S[pSE�*��ۃy@��;k��e�� �(eW���B��2�+ͤ�ņxF��dA��]Ѝ-g~2����ZH���x��/�t�Qb��K0(^Z6����OC�T����k�uu̓���S'�Nt`ˀ,.-��<���ƜF\���#Fn���{]��c��K��p�d�4���|t���i�9#�������;^��܈7}�3R-�t�T������Q0�H�@�v����z���*)��=�rO�e|'o�j$�f%g^S�tW@v?���x��zdZ�RKF� ��r.u\��r�Q����6���+rQ&�s���!=9r -K��UӇ@k�������� iE��Y�^��3Ũ�'�n#����o-O��v+�_�b�x�\��g����Lb�˥���0�������$%|a�@ʛ��i$`U�[��S��U*�&<�Em�!⊡l8AE^,;���N�MAh{A��ϝ4<�͢E��|�h��CRX_��)��rL���P�:ۯ?� ��"�|f��y�w�^���a<Z�Q��'e3�n�I�a3q2��� _Jw7v<q�p"̖$ EӅ9�rsǿ����?h��V5�<�R,ۗ�`1�D�����q�9�	{s�3c����+�y>�k��w���9�r>xߨ����� (��{AP�4�?d<�x���L���O6ʐ�J��sT����h��WΫ����J��k֐9���H�β�䁷�`�;̰Z�W5R�H�ҍ{A!�q1�Q�y����h&N���}�,�k?�V���U�J,%}ZD��������4���f�|�Zv�7��,+:ٽA�Pڌ	���o��>��)�� 5`/����V�X�y��HZY�-��U�H1�����7������H���qT�x�z� �M��$?|P&���$ǢG��,����a��s����h}���;�ākn���:U��ҐZ������C�>�ay$���z���
�^�b�]����A�C����_��|r��f<�%�e�FIqi�'s]�f�A#�8K���Epb�<^����w}��\V^�^��Q9�P�s�eWKU��.������w]�AY�qL��f����_gޝU|�70�i���d�]��P�:o�툂�w�\�!8d�J�_x���L7A�R�;u�_���U��[3��TK�̒ۆ2r�$��_�[ ���3�N���	�fAh1�_B�D���K�o�Ԍ"�of�;�� 1���/}G��A�9�x�yuN�(�"b��G�Nԁ�Kiد1J�POLTk�\ �0;�_u8��'�7��>W�e��Z#2��݂<��JP2�\�%C	%���8�����kCӳγ\_�(f�gf�Q��}:�f�����%k1;h�C^|vC�حS˷OԴa����]K�KGc�U�S��@r�f
S"<�P2�����3����=���r`�RY��hلi��������$c���U�9�ߺ������^��bN�_��.���&�6g�P����[{1%��
��h@�E~����PD4�u��Z��������W;t�xT'��@�� �s�/UjL㤊����o�{q��-$6OȿWt�������j6T�zhrR