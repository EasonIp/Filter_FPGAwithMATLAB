��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�J��"4�=�7(�T�JѺ�ő��,\��s���ӣ�F�؏C�_e��Q���#����OE��y<�HT�X6,�V�vq�P9\4HƁ�գO���@°��3�۴�C�G^D)�����j��g�w��{��&j51P����2%�t��u�/0�Y��ݾq�`V8��@Yy�<1��1w\\*D}�U���iB�ݲ����,t�jE�Ǿ�d�Li����RwE��`��:��Z|�6n�<^�:�0U����n����C/��B�pe#��`-`W6�`�a��G����u��s<C��(DAy�;弉��Ij�|kl�Me
�w>\�����0`|4�v��w�	4,s�_S�:ƶ��VR4����<'�����I�4��T�b�l]���i$���e��W��F������|��Թ:>F�A���j˧�gS!�S��̓�� 3g+΂uW�U����r� ~���e�W�d������*p��X��+`t8k�P!�ϙ�9$�[ʠ��?r�itx��a$i1���(�]�pq�(�+6��o�W-��4�M��Rⱹ���Ϛ��4�9��2��N�@�2_��ңz p�;=��ʌ���͒����iޚ��Q�+�+]�3D�7XQyvƟ~�]M<-��IN�>&��
tEV#l~E��tUzctv�0�"E����j�������Y�f�#��A��%�
`'������J켜v�/eQ�#Y\�/�^��L�-�n�k_��d�������������߀q�����:����h�6���i;s�XP��az4��* -.i�&}-m�b�ߚ��p��GI1��H8��R�j3�|	*L+�Z&�)�� �_���޸9����T��I��� &mC��G�&�;�F
��������܎`�h͝�����=p6�Q_i�g2\�oOI��|u�+Kz���.,9A�7&���Sz��Q����=�"*�e��%���iF��:j	ˠm6	?�Z%|ì��+�����cmX҂�IW��c��-���>�:�X�x�T�N����K_`t
4��8�Sl��y��S��a��?�0'���:��d+�~����Vd�M(z��U���pش����+�;�Ϊ�ϏE�$iƶ�^���h(5{�ݸ��M�f��!��J""��=7ζ6ȵ�w�9/�WG{��CA��L�N0����fqEb��ƽ��.��"}�j������wNTX�����?,�b�����gF.@1W]��O�x�m[J�e��e�����3���io<�j��G�~2*�ߚL`$�����w��Ğ�NENn�ڻ.T����5őh�G�+J5��F+	�z�e`>Q9LN�N#E�{P�!8; �D�6R ��X�7�D��Ic"-3��3Zȋ �*#;GҴ-�8K���s�:�{�8=�n��w0��*M�&���������V42l~���V�K�S${Df�tb��#N�s��#�����~��ϑ�+a���f)1�.��j�zw�`��w Q!��c�g�
<�>M�t��{�{��<M�O���K����ް4�L�n���\9 ��j˲����=5�A��t�����@k���9�h���Q_��=*Y�=��Q%�^�������~WW1J����v�Rs��A��[���b+�H�=]�+�Ǟ��`J��åyD��=�ԖA�o��8� 5�A������}��a���>��4�޻e�����'���Yd��'�Qz��B��%�p�oXk�tJ|�۱�(�|"h@�ntm���,���o�J4��q�l	{��H(W���������L�v��S/h�66/��[��l�-κ/{�`B�H���A~�������'����_:��!s�h"_���gx�`���0�G���}~�\�� ��&������+�cY[3�DϜ�}lq|yȎ*Ϙ#Gz��l�V�8����S���9= Ƭ}�����p����-PD_��F�f<cr"����u#Q�7��q�w�g�m���a�S>oU��Oo���
 �E�� `蚇������E�F(6��
��n�[�-S>�,���E���
+?������u��&��X~"��R���V����z��Tӻ�/I"vs(�bgzn`pW����d���m~]��;�)�u�I��V���g�ԘA2��ȸh^z�@%>1m�ԂCF��3�����Ŷ5�#������.i_ku��`�5B.�h� �}�y�L<��9�9�s�Ԕ	�9�a(I�s
�Dj��~�����_�&��P]i�|��/��� ���KB1A�,�6��YWs4V�V��T��P�ŝ��,)�	��)�Q�pz��� ��N)/ݭ4c���cؖ?�����
	��}h@9͞.G6��Z
n�&�'�ů�b?����h��*�`��-�QЙ�����B����mM_�7��|�F�,u+����Z�%gA�ϊn�3p&��P���I2�H��K����v���98��^̨���p�;:�j��%��?S��FU�Rba7,�桝H��h���+k1�*g�݅eu�S,N��R�^�h��Nj��6��MD̻��C�_j��w�7�h7�2���Q���dU��JD;�R�
:!�
�np ��{���.��TX�*L���7Qf�_�%���:���잸6�@�w�v�_%U
�j㛀�M�i|�A����By
-��-�K�ݫW�*��v����Zo�%��Aյ��ĥ��2��[V�����Ru(Z;���o���vU���7����
�`������9ۖ嫹fݘ~"<D/������Ð����)��_��5,�k�[�<D	6h�<g8o�Ϻ�qdpw!ieB�I�����l��ȡO���-?LBx_(���qe�I6JL��y�6�2�8TV������m="��_ĄʸV2M	��\�#4�|\���t�����Ȅ�?�zO��\oХT~ρ5L���s�9Q沿A���m��gٿa�:�{��Q��f���3�ȉm=h!c�I��`�*��k��>����⏢���Cy�W�I8o��M������pQ�%0��wJ���6�%-$ k;#�fe�j�8 &gUi��>�V1v--I�{o���c�*��[9�0q��z.8��j #��v�+q<�	9z/�Kt���@\�1DA���|�&U�W��.��p3���SH`�p:ė���gҨ5lw�.��_��gS����xki�-�E���\���v���z���>��n�i�ͥ;��P.�~�ǡ��>���c�G�����}|�	������Ȣn��\��0ϣ�ѻ��KOD�Iވ�jG�}��p6�T�J��
$[%}ě��L6����r��$Z��rM�HГe��KG�'.�m8�輠��<�tu�2m�p:<u*R���I�z��)zj�� �"�	0���J�t�q�`�/�I�s㉈��r)'�
��x��?_>�k	��\��r{�6J�z���t��%_�����}֤?���9�,���c�T��˘�{*�5�#.C"O��r��v����ښe	��H�Ic	��=�5�O��E�9VЛ@�!�GY��P�8U܋���T�h�Wf���'�.�
K��������W��]�4�f��<���Z:�&n>���|d���J����ݘ갢=����!Iui-�T��x-��2�!�{ML!f2��DN�bSOL�7c�A������=�_9pG	�v��"�i.� ʁ��
��7�7}t'���h��,���s���GꝦ'_��ɬ4�x��r�sA�y�t��x����G
���?���@�|�ѳ���g�B�MِʩK_ˮ��3ʐ\�TKC�N�A��2����tVxp&)y�z�T�s�.ˑ����;W��Vڲ��y�Kp�%=uzg� �l��Rw��dr��{��9�9��4L!uu�}Z�^��t��i�qSf���� �E3�`�e���;C�zf�����2s��A��i�bJm�E� �so��Cû����R���:8$�Ɨ8�k�/ٖ���k��9g18R�Ѐ��ԡ12U�b��rq��úU���盲��V��zρ*����?V�x8��	��x8�S�ʘ-�(A$���:�º)7#�VEk����t��{��^�!zn}��zY���c�{�x�}(�*���ZWr�T����O��9	��h��qR����EM��LbF{�_�K\��u�cµ�]�E�=��^q�{�]I)��D����Q4����Ī�T��'}����c�����2�������W��v
��W̻�3>��m���@=�	����Yv��l���"� ��UP���~�*�G���Z<Scj���Q����d(����Y��ԹJ�>��?�ZXc�WQ�������i/8M&'���7�r@34X�kY�B�l�Tr��Μ�b�hn?@(:��7�m.v�˟��s;2�r����$Bh�F�!��x�rt���GӼ��d��t%�[4�X�]�|�V�!�.����NpY�r�%h��5��BA�.'�&&+m�3�p����ów�v�ic�]��;��S�<��B�x����P�"|����bEUƿk��R����mwO�R�{AQ�Q��E�Ps���2���7H7Τ	LEO2B/%�Q�yZ�5|B1�� _��G��Y,HXڎId~�[hJA	���'$�R,e��1�{-N:e��q�34~��VSU��"���&c:���nnP��v�Iu���a��G�D�6�}� R:��]
BJބ4�j ���Ր:I.���=h���vu����)�˜sĸc����9�S�y��2$w��7�]��o�-���I�<��K�
����Ѥ�)9�JT� �Aӆ�O�C�v
�Zv�<��R+N��2a��+R`qC�p��H<L��g��u� cl�n�m<�DA��I�R�Sڊ=�6F}̒��t!j*��`�M�Bx��4q�����m����	P���������}��T�+G2�@ZK��q%��Z�_"��)� 'Sڡ������}K�֬f�y���Ԥ[�u9�7��A2�qi��CR�پ 5�e����9���.�38�A��\��n�����Fҋ4�|���+aӨ�D^温�b5�_B����%M�̋l���)��u��%1���4U�
b;�:�B���F�@�?�/����&m�S!���?��tG��ɮ�jX����t�b�v8ր֦��L-�)6���aS�t�qmz�^)��"������%w$s�`��IqD��*~!F"ξ%����#�,t�щ<e�sX�l�r���R�zx��-s�c<T �1��̎h�Ѵ�.�	A:�����2�M6r?9c�f����{7��4�����Y�˙����־+RG� �����v��R�^a�c�D�BTj�Gդ�7�z�\q;�����Y��ӢE;+6m1�1���9�9wJP&V���:k%E^|kT��; �B��n�`�.�/���"��S){+M�r'��^�:6�pF��z�M�*k�k�<�=� �wX��ؠ��Pӓ ��nbNM�>^��W���$W�s#��b��O���Ugj����,�:�nKy�Ib�H*�͚����j�Ur�Xs:�=e��%O�"�Q7��	%���LW�)
������I�ZH�ar��_o�S d0ʹt�kҞ��o�f�Y��f��t�۵F\:+"�hLC-���/q��#�"��`/�vI��s��dS�S��Խ��P��Ӛ:��#�1�/O�U��О9��?ft8-q�B9�����B�f��m� pdE�Et��
$gמ���r��Ǜ�:�C2�-!���I����q����~Iu���0�dq���)zQLc���ubQ	��'��KvToqVƊ�9O0�7@�~ ;T���,�,�4��O�������g�_��=F+Žm3@����R��/�,N]hm��Pnmj";P����{Fs�ڍ�|hW���er�����?�NJu0}�Aڱ�yin��j$�"�	]�_VRN����F�����L�7���S�{���&�R���(��D]� P���\d��A\.ՔV�q�[�o����@S�S���oH��=���u���r��q�3�3��F"��L�n���Z���w���e�\��h��2���$ۜ}�oTء�n�- Y���iLևcG������r�n	w�� �0�������t��7<�p��Usk�h�_=��jH8�9US��q���^Yt�o}�̄n�U�Dd�R�%��T"�̃���ڦޢnK-��㾫�j���>kM��L(,��-w�~�@H!��x ��mb��a��w����S ��(��O��|�����[�%�-Χ���J��2����������ze�dÂ��?�������V��w�����I�k��B�!U72gj���xiC����h4��ۣ\�Kj��A9��^o�g�X3p^�z��FgWf�T���'���B�3���Ol����bĻtK�.4hK�ݺ�@��>�ߋQKl�'*b��<�LV�Q,5�41��v�	���������y�d,Ȩ����:�u=���k���=kB�j�Jn5�"�F�n��0z�A_Pc�P�:�_{�孱�Ur��A��"�)������*�`.펚΃��v%H�>6���j�}�~��w]�ٯV촖%��G.P�Z���v��R6��p�lw}oE�8-��i����C3�ELSY��S+� )7w�DJ���t��{��<�;�i��OM{/\(�s�}N/Oȏ�L'dB�����ⅽ	.0�P�'�d^�7���� -�fGx�r�6#e[!(�N�Hs�	c?�R]>���r�|���k ����u�V�S��5�|�2��!��pR��t�����TZfWH@.�Wk����<t��h/��s+�a�M)�W0����VB�W�H����Z�I\�9ëd�H��v��R�e�������Ȃ���m�0W�u�,����?��G��0���B!�G?��QN���r �J}�>��ƚ�{h�N&{��U����fS���vuW}hЛ�h��ǂ��	nŇ"6ZP��^�V��l`�7O9:�l���Ӱ�c\����P��V���52�}\?ʘ]©*�8E�0̊��A-d����X��L1�B��-��fX�'�Ȟ����R�E7(e��ރ{��F�)���g�:ic�����~��H�)As9WE;�d��\�^zۑ/`r!�O�%c(��N_���K�^�`?ի�۾�H唔GQ� v��GC�D~�����Y"��a���&ޒ<�G�f�Y��j�k���T�u��5"�'JۓBn�&um�~�!�;J��eύ��	����Q]ʐ�GjԄ��Ok�i@AL�86�4�3pR!���D���6���Dre0Z��&!E�ɭ�ee�^��
fN�/�)ɑ\��&/J�����'D�Dg1�i'ߘ̾o����FG
GU8(�p'�[Q���q�����r�dH��-x��G��sX���YN`�n��)�;N[�z���Ji��&�Ü `�����H�I~�ֺ�r�1�3�[��O����D�Y:�8���MU��U9ﮦ'v�!�i��P(oK�#�W|E4-e�O}�m�Ea<f��+[J忎:��T6��Q��?�3�dq���|�'R5{���iNY��l��mUG�K�}����.�D��yL*YV! ��KXG���R�t0?���4�]~��N3w=m��|��G{�������n���{�p�u<��WRS\��x�8�"0��,JD�'lC�D���H]���'Ј5m�u�?�@�����=����E��C�ڊa��`�𫞫�W��DV�*o�n�~N�T�W��F��F�v�oSl�A�o�����@�\]M$]6Z&|�	��$]i�AR�H�7�����F��ŷ�!a�������{Ҳ*�!~Ol�%Ij�O�	|XO9��Ŭ��|��G�?dj0Dv��$z���������� j��O�d*^�f�b�p�����ĨO})/���Uڗ���)��MlM!�.��WeŖn�&����!N��sݐ��F|.�D�O����EDM��	2�ypFi�XK.����&�aOl�]�����3'�?���u����[~0b��1;�+�?ũ��N˅\t2�M�v-Aa�����X4NN�IC���b�����~W&k�`}�Y��1��>�*3�J"LnN���S��C1��J�/Y�5^A�g燚^;��@���z�Y��q40��
�0����?E��T̖v��=�&�9Tj��:�>�_	��O!��F�#�k�u�<�j���'�%������\M"m���$4(3�A+5�޶��>�$~��6]wW�}�&�+ Q�ŒF��Q);ӷ�*�	Mm��+O��ۉ�Qq���ԾF����珑��?r���QF.�-�3mCJ��^)yo>�1>�a��Ƿ�]��Ҕj���B!J׽)��(56��Mi{j !�M#�tH�V�$��S��$�@�1t�	��Fc�_Ë�}Ӂa�	 �ґ��\%�%�x��e�rF���k#tČ���[}f��U��)i��I����D��5_#�\��<�!��g���4���η�)�ֽ�,���gfLZ��ݏ��s'͵Z��}uW���������� ��М��#`���������?���8TM�K��L����R�i��Jܺ�f�A��Ӯu���ik�O���_��D�9�״��W���� p�����1G�$'M�7�֔�߃V���*��#��2,�Ӫ>��7��$��p���x�`��
���rKH(f�K��1��0�{�����_���O��" �l����!��3p�w,�9���<���|�2]m��#���8�2eo!mQ+�dK������¨��z�MI�A��b	z���ۮ�Jt�E1@ՙ
�M�0�.��^
��m�_���}&��q�T��sB����<E0�XY5l]~���6d�\!�a��w2X�q�X��t��j�]-�)�[�l�	R4�K�M�<��:nF$ �lo9��q�<�ꂧ��o�<|S�����:[K��I�v��v��|N��������#<.y�W p^_�j��8] �HP������5�8��L%���-�	5��C��f�@p��;�\�`�MMn�G�d�3mo^���R+u��tI3n.�#@gO���ג0_�>bTe�'P� I�=-2]����*щ�i�W�(����xG)Vɧ3#�R��##�a��8�WE��sC�\5��c��7A�NF��3l��Y=�M�����c)�� �}Pw�"�k��)�Q{��T�i�\CH�d#-�bXp$�B�"����Ms2s�.�s_�y��^t�y&Rj�ԉ2a�)��������l���фc���ʂi��`�fY�f�$���S/>�}E�l�܄M'8Lh`J}�<�̴�H�s�]ì���&d�/�H$İ�MK�X����Q�K��^+ ޜM�1M�\���#X��?(٘�g֡��3���R�*��@o5�@��g������ώB��z)��pŀǃ$�<'��(�M�jf��@��r�K�Zd2�`�?w?	�_4�����J3��k(ۨȪ%'������emF�1�t[3]_�=����^�1��>'��H��� l�G����sR����̩~�i�QRk�c�� �~�Œ�꟧�u4�3O{�ZW��i]������N�6i
���i>%��\�3����C�c��+�294�����QW*OX��[�B�`CϞ󭊄_4?#&B�Y��v3\��HO� (�G�ݸ����o�#舻'��i�,V��:��R<	w�8
�E����hta}���G==Ɵ ��u̚��;,�����1�b:���]��T�@��Q��T�WR&�J�/��r+y<-Û<�6�ʨ��C�Қ�_P�����eZ��"��B|:�Cmכ���p���th������^0t��Y�� 8�u�������'?]����;���*��=�nQ�K/��S�W5�ʨ�`m�j�Ŭ9-���8��4e�wP�ÿ� �f��e����P��t>��	�s��
r���eI�Ü��-WJn�S���U��Fx6����������?�C��S��zࣁ$E�nf��W|�!3��w������ٯ��|�� �w�	>w����\���-���Bbц�4o�/lK2���S��ޤ�P`�t���K��i�Yu���<R�"A[���;�N,毥4���P��w�J�]��l� �&�`E���"ٳ����:c�b\���e�+�ʢm!�}��� d��˞�מtK���D=-a��Шoʻ�"<f�]3��>�.1x�_v�j�މ�����}������R:I�� $<�Ώ!ڈ��y��K6�CɈ�ѓq�V�.�\f�O�"$��h�n��$�O�m�Ҫ��E��!�%�������o����;��F�6�|�Jwt>ڳ�S��
��a�@��5��*U3B�ƋD�;WSPcf|)r��j���2�%�-�௘��8JDڅb�2���8�(�����H*	���O�-OS=)�o�]���v��2��Mjhtn#�������\M��n�� m?����ʔ�8���-����3ߜ;�PK��\^�+�/�σR����:m~�I��+�
����S��h��m��)'vYn��P�6��Tm2/�)N9��	l�U��\s	�.���q-���h�'V$�o�GA1�F<���5)�b�6�6hST�19p�f?�l6���� ��V3���E����ŝ�n�:��.iE�o��� �R��x��>�����g��Ūf_��"D����'�g�/9k��^A �&�1�qy
E���R(X|Uv���(���D��v��p��4J_[+x�����w|��=n$-��9�g�g�0^��u�&�"����o�=ƚ-�Mh7ˈ�>5!����{�v[aZYB��/4%SIM�s�'p�������\�����D%�kkF�>�pD�V�/���`�n�B�Cb���|A-sF��\ � �<��h^�r�<���M�Z��U�?���1;$"@s���K�������T��ei�bӇ8�6��`!�-�R�$����ԍ�!�p���5� ���C���oC�d�j�X���#(�PO�4yx'��/?  $P�5GaπZB�Q�.���dI�qk�.�Oܼ� ������\���O6j�_��r�kb��!� �!��?h�o�^��5�ո�n�2~�Lu	0�T�i�$�|��p�����+���QU��xaWe^��4`�x��_k�ӡϒ�9/�و�|������Ff�oͩ7�$�/�����wr�$�"F�{\Slw�M�:y��ߏ3K���I�@�f�6G$�y��r$��ֻd2�� ���]q&l�#��tKQ��E�1-.D}\R,��������=�d�G��\ ����se YKz8��ߛ�Q�������|�L���������s���ٻ�S'�.�x��
���roρ����nzl@>m<�+�H*o-�LU/G
����;C_�0�<����z �����>��s%t�1�>�d�2^��4�ᳶ8�	|���G�~
i��g=4�4IvH�۟�d�����r�s�O��Ե§4�}��.�H��a�:��)�loGP�S�j���1G�c���ɕ<p`�E����2����-NKF��?���+�ͳ��1.�nQ�s�k,�lQd�/�3���/Y�Sе1��2k���!��3�&`N�k�������t�ϠUZ;�y̩�v
T��|S�^R��&-���^�p�(C�D��_��� ��K�^"2��+�/[�"W7�=!��y����W�N���P�2hd�@�I��zK^=�:�v��Ļ����M	�戕+�͸1m�(YK��u�F��d�/�y�Q�L89 �zT��11ޗ��_Ӌf���A��UB�䕁H|�S�*���x%��]� qj"�֧�A\�4���R�_���&>ub)4'����p}紃���`Y_CnR�������{�K$��T�H�-� � - 7�<b4c�:t�#bPUƂˬ`��uܖ������t���ʿ�M� �y��^EؔQ�B/2�zT��<M˿B�k�9L-
a�=�˼�#�
9{ș�+k[+���w1�B �H�2��=mЙ�34A���.�M7���!x`���twvB��Eh*`�F�I��u%<bd`ۛ?�A�l�݅!c(��0�P"6>^�/�W`톅1���E5�W���_@D��p�/�![���ThR�$�P�ont�&��B%V�F���Ru�J�2�#VE ���$j�#II�>`��|�]J��Vޑ��N�,�ht,����s��[��@ѝ��n� @�T�޻�I�^GL��/f1���JT
�![W�;ٜ+]���Q��T�z\��I���iެz�|�R�y��?�� �q���J`���U�vW�4��0�\Vw��}�D���p�ݾ"���B�H`�xw�S"I�g�����B'A�.��	AC)�݂�-W}�2~8��EMW����>�O_����$?s+�hƔw�U=�ҏdYٔ���!k��!ҩ�c�@��`����zÆ�A�����"���z���.�"t.��`� �SRx��x]]�)���J��9l�q���D��U���9'��\7�;���