��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�J��"4�=�7(�T�JѺ�ő��,\��s���ӣ�F�؏7ޑ���LR���SӞ��&7��+1����n�L����[9�.1���P�y�I��v�|6�3fuN��s���S�y}WѬ�=�ֵ��S���&�_����G��+ǃ����0k��g�1����2���t3*�7�S9���0�Ҵ[�j�f�������S~�}��'���y���D��1����.]��� 8�u��$���y#��.�"�8��1��4~��Q-R�Cv����4�| ����`�*�0~ws�JF3c��4D��������Ϟ*T�h��$�sQ8F���=��H�]2��>
E�U����b�f��:�s��o�A�ZUX!>�H��{o*�"O%p~�
<X��)&�aI������W�K���A2�Z g(!��\ǘ`������i�HF)��{���7��
��w�� �i���'���i�f"Y���W��Q�t���9"�3�2�L! �F��%r>��rGsG��&�F��(ҿ�w~�?͟s%+�%p@�[�;V��H[�ŗO�Z�����!�\�bP<�o{���������%1����-͘WS�k��Y�2��spז�1	{y�N��M)��Χ��X�l:�������Oyɑ�Tx�Y�/$_��`g�]�gw6����e��r�z�\�������N��������vg.,c�� _Se;;Τ�Ne���r$�-Mߌ�1];�����L�����i�m��@� �+7�ũ�K1����U&�7���n[�^���2i��	<��s��c�����U�\'䡡��1��2�L�Ί��KP�`���FQ`]��!<J��g|?,��G3�i}i�Z)ԏw�.�r��S_<�`"�n�fd���CH�]�.�%h�6�w>hH�J.��H�d��n����b���q0�ȾU���Y{�1A��Jy��	<�����t��8.^ �������h�i�`�n�(��]8��]G{GiC�/h��-�Q>�i�5�9%5� �V�1(��xP�������sm�������rsȲ����y��/X���_����ٍ���2�� ��$�460���ɖR������b���2�HH��y�!�uS�2R�S�����b"��9�k�ߒu��De�H�r��}���q�:M�"k�Xl
0T�Bzu7+c+���>Ձ:�q��w��?w�^g���݇3d����LN�jXJ_
;M����.��O��Ç�*/[`��G�ƺC��P���孏Yf(�����Ǐt�����~���F��Dl��*ӷ��~��T��PK]=p�N}�+)xYBc��_�[�Q꥓��Ȟ�+�O���>��ѿ"���,HUl
�	=L�{�Kwy���f�4$�EP��f&'a�ȩ9�4�f�9 w�O��5�w�q��Gۻ)�<D;Liǉ��x�of��8��W�K�Դ�uq=��i�i�=0]����gަk��������A^YPxs�ߕQ+�;�l��>����w�oꬮưr�;Sx#mxH�BI�ϐ����c��d?��Ԭ�=e�&����+�US�=�2�cD`�05��"��r+Ɋ�>]�1��'���+�����G�f���9Zw�÷�qP��vsW�땻z�BtX�<���${�w�NAq�9"�1P�e��S��G`����7�oݰ�"q�QՀ��ս&���q�	C5n�H..�Jb:�l�d�����R���4кg's����4I?����#��-�Z0���=�{]�~W��ۂ���̱_���ax�s�Qn����G{����RB;�Q����� ���F��CT%H�0C6�T�/��*f�_|��ba��C���	L��U)���C�Y���S�o@���b��c��z� ��5��h_�7Qг��09U"�ѩH��^A����8h	B٪�pQ���j���a�M�1btjΦK<����P�Y�̽�E�����@y�_E��T] ����ZS6�ߍM�����"z���)�TC���rwz��ׂ7I;J<e_ Y��g�ó�v�ɻ(ke�'��QP	��R�s��.,z�3���m3��I�{ye��"�m�M�Px]|#�g#��?rtH���Z�)7�-�?VPx}j�� P�~uOY$��E+���ַ5�p2�������g�DNV��Y��)3��Yr^Uݯ�t'��j�4'K@�L�Ǭ5�nK�o����/��i��&�ůA�'�D�<��on~)x�6��n+���nK�)g����aڦ-�O ��$�ă�̏�+~��be��Ld���"���V��Z� ���l8��)c��(єRIeR�ҀD��3�m�����SM�Z��%�Y��P�bfg:TŽNH��Wm^e��8>UZ��8.ϳnY�GU��� �5�,���,��*st��W��s�ߕ�Wl̤+2AC<�"I�� ���ϵ�j����	"�M�C	�FR����.׿�V8�au}����}_B3�!��Ff�r6�	�&v�ha@ �D��V�}��F>��}���C�Jy�'�_�]\����I��w��^F��0P����C�U,���.�!O)R&(Z@&�l�O��+ś�ɚ��*�T��	��hγu�g��+̤��1��1��߭���B���V��܉�-�!�0i~��Y���`��"��&�;mğ���H��y���Mނx(���� Bצ��M�A���*�&��h�a��r���]ԛ#���t6�
�\:�~��^��r��"���N:>���Ű&1�M?+l�TD�q|��3<I���xx�!���(dIg�"]f~�C���*��Ƌ:V�s(�i�٨Cnp9Ӡ��b�6��}Qc�OZ	%�sG5�ɫ�\`0n--�3VZ�YQ�ޓ��8�J�{�� 5�3�U7"�b)Z��_B��GW�r�"�ц�Z�GR�(��,"��S��ŴdP~��r���k���x�ck�Jm�����wDhΰ;8����ā�ޝ�4�m����%"��n�z��e�I)),���o16����R[@։����ll��/�j�)��l7�����ˉ�(E�^��&ńn���b�Q#�f��҅R���r6�#!��t8��>�IyFĤ�}����܂T֔�^ri�&�+aCƥ#Uu��Wx��d������u,r���0+�����~fa�7 �p��1�T5o���;�?��Ӵ7��PW#���xWtMM%[&��l9��_q�"�D�4�Jc��b��mm���2�[���Ǜ{����^��3w 	�J0xV��9A�D�.(<�IS���Q�( B�NLrX�&�e�dV:�W΂�G�����%)���v�\"��~�7�Ƹ�v�Q��_s��s>tA���A��wY�Rc|��H[�������_�g�N�:L��-��Daš��jǓL��X-|��&���2͇ִ�s0n4�,����Q~�c@�w�$�b�0A�wir	��HF�6j�1B9 \���a�|���TrR��,�]���u�67��9]Y�B�Bd@8���b�����[Mu��y1Z�TR��F�
3H���c��i�*Ci����mdOE�=��×���*w��/�"��0�p)j�o��&#��u�;�A~K�
�h�9�F�m���S��@}�5��*fT�}�=u|ԩS�}����!Ws��^���~^�E�h.+_���u����̐�7n��ǋ�o0�2|\Íd�w]�C[�*!�d����d@Ad��h���{��>R��K	ޘ98b�B�!O%{���1R�Pm��3�Y<�u~G����|l5$��C��Ħ���sI���K�j��� yw%�TK�g����[�8=��pU����e����ђ�Ǣ`H�����f�<�L�M'����2�|��u��B�����j9`7�C��m��������iR?�TW�����I�t"�O͘��桐��#��r�;*#���T|b�1��U\7�u=�B���d�.&�T+4�v�8��+�H���;��!��-�A*#� I�&dG�"��>��A�J*:�$�d��z���$\���d£(T}�.��5�FÔ��9ហ�U5`���;H�<�i�72�v��6E�Pdi��oSB�H��v���a�)A��Z$9Ox<3"}�?���Yk�Ÿ�-�2?�<B _V��`�L�����\������ܖ�*�ɹ�o|_}A���߁q�hN-��ݭ��;�8�����ם��\+T7l@�)%L!ӆ�C]�
r{v�4�8n0���Y��VA}��E;b�E�Z���֬�t�B6܎yϑ;��\�J�U;Ld�Esb;t>)Ă[�R��P����S���EƉ��Q�f�N
�^�ä$�*������.8�4zi�ҹ�gxjG�P��=�$��Ob�\钖"�z�9�_!=W����
iC>Ya�p1�h��� �E�L�_L":1r&�-�i�Φ~���+���1^o)N�4����6��b^�;-�\����`��)b���r[L��>�ϑ1針/1E�Y�(�`�F�H�7∍f�ސ�$ �1C�z� �%^N�،����]��ֺ[��<�6�a���vn��� �$�?���U�괊�c���.�Ƕ�-x�olb�.J��Z8'�s�A�ή /��G��s�1j����4>���*y��O�����_���ڷ���/4����PF.��6���(9.�1�u7v/��u-ұF�P��m��x��	߃i��;Vfgԍ�:-}A�k�*��=f�`}�)Ce�)r'Ԏ�,��I�%L��GE��/���}Uf�E���ݏ1��A��>�
�qw�F�;��������o��Q@!
n���6<	�t�.e��vՉ���v�_��
�I�/Μ���̫G��� ��׷�f�D��*��iRI���nf�;�f��;Ì�*v�T��*V��6���(���U?L��/�MЭagp^n����0t�a��׳`§�'�O���̓��\�<��8����o��J�b����2.�b~Y�<L)_�.���؃��7�=�b��ˣ!�9�鳠��k0�E-���(��,BY��>��`,�;Ʌb���Y�b�T��w7�i�ԫr���r��6�k�ΘkB-p����������(,���ĺ!P��ۚ�BrN�fts8�HL���imu讱�8�'��>�|�Z7����o�D����CY���B(zS�.�-���1�������򨞢���P��W�ת*q����$�:�,	���n��`.�;_ If��<�ƺ��{ 0hòJ��������Ò��L���*ߜ����	�7"�8��]��?`o LU��p	�m;�f�oN,.��}�1��w���,^��X��2{�z
��Ϥp\�������̎5N�P��J��r�z|+ܢ���U]�[�f�4���Gx���!{x����}�R q��ej��L��_Ǭ��{�vܱU*q&�t���=znw�����2j�=����{�)2s ](���\�;&�\��nqw2�� vb��gj?����a`ȩ���g�P�+^���Ǌ[�����.$�D�
���D*�</&�����%k��K��KV���節��]��s���&�0�|�P� "�+�1��_v������A���F>�H8̬?]�&��e:Q�����uΨ��F"�G����/:	�;@,���V���!e�4I)@�틟ꟁ�%�$m⁮�+h��q�%�F@��B'�@�^@E	
�B	
����X��4a�4��ƹI	Y/ՑD�i>d~���n��A@u�Q�;`���^�A���� ȕ���X�h�4�օ���<�R^˲���]l�yT���ڷa^XWM[��{������O�ʯ�ȵKTagQ�E�pǐM>�H�5��Hij��)i�{� @�]�ǽ��Yl�"~�c���jA��hB���E��5)b�Xa86�v٣���ߎ� {�;FD�փc�������0��.�f~�K
���et�銾��x�_!�c�:�wb `��&��N;&���+<�څ��Y2Kӓ��
'���`�@8u�g�K)O�K;�غc�#��"�b�Xޑ~��
�l��#���d	�Ć�
0;�C{{ill�c1AK��ļ�pr)f/U���Lk�.�lH�D��.#�&oN�=������o! N�C���Hw9r�C0&^�@0|�/�pnfh�>qq��s����	}�ѯ�2��1�E�ޅ��I΋�E���Z`���á��&�<�a���(���o0&^\J�b�ဓ'-;��t��#�2��������ײQ��y�I�e�;?�d�����,_�'���prZ選鹈� :��Z�њDy�ˇlů#@��{'����i����VR[ZirR�Ԯ_���bɹ�w�ZBpF_���x���L��Ǿ)n�T��<��
(9�\�E4�S�a$(��L:�a�*Gb=!�U렙����2�U�����d�0�K�Xی6���Xq�c������(�i+ -��NL۴'��bM�[�ev��p0��)�08� 2����qS�7t`LG��� �|��SNu@��m����4��LVd���[G���NW����b�nY5����ټء��R��}�.|�>�.�"z��"�}k8����� �@}p/b��������؝κV_k����J�q+�G�&�v�7�(���,�i�,b��dOD�,�n!�qx�䚧��~��.SL���A����l0a��u�/�P<��u'E[�S0���`^}�G������DF��9Q�,�S����ƞd�ِ���7�
;c
�2�cMS�zo\;|7�{�$D8�fvs�	8D���'�$��>^�<xE�����\�e�!�%�n��BŜ�y�CĚzI�W�D�O�ݬ@���W6P0��c`ǔ��x�m�\!ԕ����g�|�("�]ԩ�,Đ�n��0���d�7�6f�*yC~����#��&d���rF�=�������v�B��Tsؾ6:��-�~����<uy��X�hE����[�'���v�z��$6�%7��%��yJ�����֎��(f��Mp�6SC}y%/�f,֌���̇$=��[z�n��X��~�[�=�l��F������
�ޑ��o��D�H/���H;I�O(�uη����_�|$�f�#����h��!��v�~o��7�Q%t'�ȇ�:ߒš��cKm2���4}~;����|8=C��Ƞ`>��=�;i!��E5��&,��.4h�PF�JjQ���k���[B�ͮ�3�t���N�Z��Dx�lg%��W�(2��P�kԆ��y*/� �S�'!#��|�>��8'k�uP0�٧���a���L��N��K__����\�4T�R�:�P1�ak~�^1�����q1��
���F�s=̶�L��>i*�Ag�o�ʹn?���(�F�Jr#ˡ�7����r|[�Zj3L��m��gaN�A��Z#J���9`����j���$s��R�dr2�Haî[Y��^�f�>���됏��骟����~&��u
�:�����p�ů8�o����&3���YSHZa����YP�t;���iz���y�U����pW��@��h�0������B�!�c��oB�@.����gS�EтKZf��K=�4�w�ЂS��vtA�^��K��ZVVmC��_�ş�ٕH!_��m+�k�[��/��B��"����f����B#Ewh�����ڳQz;�ˍ�l�0��2�n�A�념���p����б��?�7��^��j����X���J��4���W�����6�0\B+1+�.��:Q�;^u1	���d&髯M�B�{m%G�{��{.�W�ZW��_&;0FYa�Ȳ�3�j��^.���)��EJ�B��^��S5��R�H�$�(��`'�MN�>��ɱ�%�����9jm<@@۳ᰨ���o�6yC�yr���%��ݱ�l:'wt�l��o���g[t��e�#K�Hfχ�nh!d����8�FiS�qW���{Ƽ��%(�d�Bn���=.�/��Y��T�f�']��¹�͘��dM�1{�Q�K��@�
�s�A�{[:GF��3�ȿ�'>���p�I��
w��d��W���w1��<}��`�P|�qcCOS�O:���ZIRc���=���͵�K��?�!�Js/���,�j�;8�~�z�Q�Vu���V3��3�M�E.�\
����u�2��+�@�徜5s��3"�&˩�
:Y�х:7	(q^��V�֐b�%e�pK칵¬+-b)M�R]�\���%���8,W�#��hg�Hl���J
F����8�ÑV���`�.Q��]�ZT�T��0od�;#��讽2���\��t
�/����=�l�7��K��tn���]���ӂ5y��1ty��[�'M�t=^�B�����w�?�ߵ[N��.g�!�q�H��G	/h�(�z@'EŴ�J3�����Gm�⣬Z���Yl���ڜu騰�7|�5+I_qaK4�q5��8��?�P-�4��vU�-�m