��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$���뼣mh�5��\���N�-�[A�~}Ǝ:�yLcLM�`ۙ �!,��kVY_�Clh��Z��)�$|�c15�A���b�nJ�U���[-n1~����d�/��TL�bh��"�����4V�ΰI/\ʹy�7��X�8?�V4�z���f��Iw�]0�Ů��Ek�9���8�H�Z}��R�yp�X"�*X�jx���m~�~K�F~���f� �
�6��p���іs��T�lvsA4��ۑ��u��N��G���'����Y Yj�!��$��{�wg�݁ �Ʉx��Z[�L#p�ft�Ϥ��X���'q�Z+��*ĝ�+�5��?ưrzurWR}5����o����DO-�6+�}(UD_�E�-�Z�<�;4��V1<�Q.\�-�ԉ<��T�^Q1���؀��9�>�~-��zpm�'Z ̪�"�E�Ix��J�����9�Q�UF��j��l�>W�'tM,*�^'J��N�}D ���U�慷�MF���TY �D�,5BC�^��ؚ̮.��ۡ�� 0���4�����!�s��S�B[zI�,���[_wՌT\&DmW�������=U��2��J-�%�E���*����I`,�e����n��cH��7/>�����ǉ�b�\���o����'���E�!���T`~llJs0N���������R�	2P~�E��ΘmD��}�0��
0�v-|���(��\%*)�B�����6[��f�W"����sڀ��[~W+����7W�VnG������� �W]$�[և�^C��Z��}׼��TȒU����=��/ �l$d,[N��i��_�����*gfn{^��g�B�X�ւ�~fޠ*E��_b���xF ��e���vOWG�L��<d�9`u;a{b���~�I�9�
�'�d��Ϯ�o��
��ʰ/�eX���(�uz���~�g���?�8�`�9�p�7Y�����K^�I�=�����K��#�]oU�ա���8>��L4 a?" k�/=��Y�k����d٪O���ڶ�� ��l�k�H�9�q7s�3Ĭ��+3�����-�}Sǁ�T���QZ��]�X�S1*����$��m� ��Bܠ�4�C
@��N�);j)�cGJ��r�V�=��"�%��SWa�0���P�j5��0[m'ܝ����FB���]�R[��ެ�$���L��*5��>cI��Ŀ��^�#��)sU��T
�쾢�Ǹ��G5�+�^�����yV�����L�ţ@�j��A֝�~"]A�n�Ǟ �`\��-�}MJs�����-^Ҿ�&i���S("B�<M����H	�I���`f	�_�ֹض��'c�̵hgBx�x-�|�Rn�g���E)��^	��_����Vѐ�5Nf�,�)v��`��I-J⹪��c��V�L��|��]��E=��FTjnAs
#	�U���+柁�HUy{et��x�:' ��{?7�h�!C*��r��ǫ�e`(���+[f3�D�Tґ5V�O��C���&QD8��y�b�w�;q�8��u��?
l�4����,��n齑�b<Q�WM�3P������w��[H�@ԻY�
v7�� �ϖO��Ї�w���[���d1u`��F��ZO�3	 ���]qc�˭z��	D`�P�'��_�H'��
�r�|=����F�Ý�JZ�(
���"Z���<�3��VҢ�>��d�ٔ�݆IfA}�f�(���D��L�gTO��� ƥ�^j}�U����%�����V\G�֦��[��s=��B~�?�5kf�C��;g*�W(agU��Ϟ��a.�x��q�xFn�-9b��Q�dsk�p���:�Ѡ���'@Bd�@��<8�n��a�<`�e�`z8����m��^�iD텅��àW�����xq��d-�;�*`�f?q�����֐d�*��a��Y}>x16�+U����������c�0�֊���T�1�a�AO� ����F-�m����!Pgz7�B�V�Jdd������E���~����I�5b����p������Ƚ�i�e����:b�?}cx�E��������	��Ь+��]�jՇ�Gر&ȗ�����8��ަ�����]�St"E��4k��l�PN�H-�?���Fxa��`�+��u?DP�����U�]�iӊ��1���\s�93_D��K
e��q��~<�*�gu�\��O2�g�A4n�{	.�R/4���'�q�o�s�A�%�љQe�O��$����So
����v%%��^H�E�����:ݲ�I8(��3�1��t�f:ϵ���@W�^�--B��S@�E���.�v p��՘�"��#�P<�#���l}�IX�4y1��5�|�Y�n��ZPd%�����Q$~DG@	tS�"	<�Ev`>lVK`Zg��� �� c�"�'��<�����)Y+TþX��5իtԁ�lPF{�Q����C���T7F���[��z,��T/+��,���{���9���V��J����c#�qר*J�w�[���45[ņ�̱���J6{���M��P��;&���Y���<S��_C;��I���Hs����n�F+�:�/W��4��O^����B��nG0 /!i�"��f���i�}��`�8��{���Fh��S�vtQn�3�P���Zs��XQ�#1Q\{+1uR)�	�s����yⰫ}#x�87��:�вf�r~V� �
[��gM�i� ������k�t�mj������S�"�FG���Kɓ�e�g��T�J��g���0��*E�����ra�^f0!�h�qۗ�\1e�K?����;��E�e�g��m7	-�ޛ�/��u���!c����ų4�:1��&�>o�u��7O;Dtr��@�������0~��צ5�,�q;.o}��2��lt��(���X[:̃Z���<M!�n�~͝Ҙ4̀P[�{���������s�Iw��չ�Y?#dA����L��ɻ������%a���ZQAv)j�Ԇݖ���@�
��l�ǀ�2�KگOT�����'��sk��*���~�&,Z�I[���)����f�-;�y�bo7�mN�Q'�[�^7n��FΦ�}o(�}�A,Yr���CД�՚}��"��K��4��O�?��йٲ��KTx�]78�δ�Vc������U0�<�H�H��0��S�I$���gK�����	iν1���`�
����߮.ͯZ�!v;^PE"ȏm�n�x:�שX��:�u�[/�2�敯��D0�{�s�����o�u3�:��0����
�JH��U!�sH�MZ����O��[�{FV(���:K)~�sF�Q�|	5m�{(̗#��4d��|lrr��K~�D��6��&P���[$�W��n��q�4���4w�*3���q�\�za(�͖e�w$��e����Vf'�?f"I��w��t�|�T��2�fKOi���0kz��S-%�#nRD��Zc��yﮍ![kk[�<����u���c���}���Fi����mZ�h2/����y+b� ���R��`TL��M쩻 ��-ً�E_h��|�Q=�~��ij����F����tp��R�k��dtz�-/���DA��2[���nl�;`��e�<��`��3��4����y���@�\56s�Qf|��d"2հ�[r��Iշ舳��Xv��F��B�K_j�þ��vc�Rp�k�5��Vmf�'�l}]�˳�u��cP��&jbxE��GO���&����z�↑���vDu��T"uw }N;k+[��
�]�mT���G��=�_�b�󬩸�Wp�#�1��4Z 2Tv S�ߪs�^�Y�%I�=�Ŀ��DV�K���gm��:�����n뫚�l�H�G�4�0^���-�z�%_Tn�i�X7X�3��g!v �j��k_���ӵw�d�J����>��d�'�\�s��M44d��R��m��I8l�'����`���/��M%.6Lf���0�p'*8�`�k���sO�	��d�?e�-~���V�M�~��d+Y��U+��C���υ�m y�m����q!qIHb�U�rO��3�W�r����a�/��2c�Ajq*��}�Ͽ������@�I��;*�+rL�&���FNUV3�j�lb/g�z���d4Z��:6�MԎ���Z����`[�^m.8B\P=��&��������e��q=�k>�A�Չ�Ψt�x�qXg dj2�mz�z�/�_mw+��.X\�kN䌀d�"�� F9�M^�(k���1<��/�@_�֎���	�t�U�
�@ԉ�ym����À�4��\�&=�b4����SG��t���в���!@`@;tE��:�Zώ)��kX`��f˯���9�E�^M�Ѡ��d���uT��#ޚ{y(��\\c���v�i��=9����`��G�s��k�qN*߁Eٖo�{�.1�6�U�����zAZ���JT�.vx6٘�v�k���Zal�$�C��r��;1X�*���_�;9�w
b**����̓��t��eHx~!n��>�~���,�Lˌc_|�luZ��љ��)\c/�5�RJ��r�?adֿ .`���]�)��M=��2�>�'����֭�dнk�U�BT
�58&uq]w�I�,[Fi��>�<0�kƑEkᖳ���)Y�K���ς���R��<I�ӭZj��1�'J"��a8|��e�Sܨ�ݡ�5���X�v�l�綮�/T$\��(�9�+^�/���=N����WQ����!d�0 �+M*�x{&�}��x��ț�F�;jcb�G�j6&~����d��Yk�C�&f�{x�I�\"�/	�~��^��b��K��E�E�9�� ��!��d�3Z�?��6~\�6?�ig���qe�J���ܹ-[�����={� �����P׺����604E�N���:'�.\c�����e4_VK�B
�-��������M"�J�k�K��
��[U��~��|�;|o��N6`��� ��'c[ ���vk�����L˕��hDS9fǃ��5�'�y�|2��c�=m������@��^�M+�V0�ROfWe���£H��3d�=.!Z/�!�_C��vo�괰"x�էKHI�sВ�� �����M�Q�lD󰭀�`�]��ƅ�h�ݿa�G
�2E�X���w
d��/��,j/ �=Ȣ�^l�w��J�$��1TT5������zg�����SQS��eכ��FUB�R�F<e"!�nW�2�"і|f�N���e�"Oy}dO�����`9�
�)�v*�qR1&��<-���Fyr�7O/K C����q̇�D/Z��<i\�y��=�������(�[���r�(�`�Jن�u0@J��'�!�%Z���ش�@8�{���.�O��7r\:(%c�6��"l����Uw�X��z�`��r�,i�'��٣�w Zi9Vpq9\�d����ݨ���?[z�<��Y�_��P�3B�8�.rR) cv+�+�5(б=����l�_��`�ut�Ye�\Q��p%���2�֠/FB$��$8��P'������Ynr�`��t��9;��^f�!��k�KS��(�J
=�Y_�twh��������7,��G�����n�9����J�dS�����0*W��V���O���)�5��*&v�o�h�1�#z���֙ali��xX�2�̸`�H���-�Tb�� ��l ��Xr�^
ƀ���;�̦RUer]�I�~8�y$�Ju������ye�8���ǵ�}���#��e�x����#=rm�g��4�(z�1v>L�v/��i�¥L�t�y��M,�������1�)�t��+j�8�p�K �%��"�S~�<�L�^c堜�b#w�Mt��1g�O#���ݜS��
��)��.�a�e��`ū�20��A&�/b���5G�D��9(�=ɭ�dՎ�j϶�ݐ�#�-��{g��S���r�l8�^��5��t��:B�v})tMk
�r.j�ǆ]|���݉�C�>�U�����YJ�^��~;������-������0'J��s'5�5��s�����tiDؗCT��w��ĭ]�D����!
 Q�5��U0�cW���.���P�����Wyh������Eҕ����)��~Ҷ{y�<Q%��,o4�"�_��3�<���"-��_��x�W���`ˤe`,d�Њ��4A�L�@���g3R�%���M������?����uY��o�$7�1��Z���K	�h._�`�hYR}q\�	��K����v���@�CZ�0�IX�{�vJ��_��K^���}��n�����p{�Ќo�{�͚ި?:�؄�l��ExpىA/���Y�i��H�������϶�8�'h�ʚ��Z�M�#M%�:T��:
���M�2�u<�
�x'�	�P���W�l����%��a�o�?��U|�ݒY�����A�x	����,�+�;���j!ќf�ϓ�U��yO����7�(d�����4F
a���~����Q+�y� ��f�C�������>����<V|���{�}��Y���)C�w	���F.�����/���(_n4-#y��*5��J"�d��Ue4<�bY��+T�7��橕%n�sO0�i�|���ٔ�P9UX�� �S����ީ- ��j!"���q��	�}Tښ��Ya�<����a�(�e_E�q� �)�RU���^ih���W��;��!"�#T��b|@�n[�O�u��+e�(F.b�����|���2i�e5�n-��~��1���:��U��[���.^|�GW��E����#�K&�7x6���:=#m1Z�����K�ud�� �% HBn�p����e�L(����.K���hW��샗=�Is%Y�8}���]Eֱ!͗]�1;1��� F����@td�����6�Fg�*|qq~���j�D��Lk�2�y ���/vUG�{����=��u
�R�K�}�[}�ĐH�u�Yius �h�i�SuPDE��OG��R]z����P48���>�_;ߣka��B�?���a�fJy-�{�F+�JZ��.Gd�o��Ck�]aվ��d�W1����b�m���,I̺ʤ�ؒ����Ga8�c�_��]w�4p�h�Jzu'�4�x\cN��c�U�V)�מ�P�RI,ƣ�a�&$N��;dpYzY��@-��Lv�$��+�VX[s��S[,RxP��Tg�Xu��W���(�:���k:>�O��Th�.p@�Z}k��`�4	���`��o����q^�=�ʡD�@]����LǱ�H�s�}k��	��|sA�0�xvD�w��B�]tm�t�1��T���7! ��C��L#�3%�hW��[��1�����6�KY��r�{�o6�?ř�5�'�iB��4弦R!�&����c�#K���� ��x��q/��JP�
tP�����<l"�NhȌ6ϓt�a��@��<�3�RA�K�Z}03��;��� �a�f������X�
��g	9�	���l��C�F�V��-7]����Ӻ�~`i&|�ʿ��2)�*>�=!� )x}D�G�x.�T�Z �"�)~��6����T��|�@vҼ�lI�;�Ȩ�}�L�^����)��<� �4�$��+�#�:9��7w�v���1�����NƘO���J��]��AT��Z��ҖHe|��֭���kƒ�=��S{4�U!ʦ�b+t\����_#F��:1T�wx`��[�F	��s��_b���M��?�����qSC��(�St�pBa*�����`��=h��P&����(w޸K���:�?N�P(���
L��Wf�=V��Z�z��Z�r����ޥ5S��я��O�݀����t8/gC���&���t2�)T)sr~"T�RQ~����x�4�ʗ���<�����"�xE���>��0>�Ffc�Cޢ��U�d��A��f�0�EL����D�W׽h�����R�0�M4h�0Z_;�JB?��a��V
}�μ��e���*K���'�"S:��/5�B{��6�~�֔t��3o�6�D�?��`��{;v}	y21_��\~�-<�D� �W.?"55��2dP��s��D�p����!f�l���n��[��ncma=�8�nM�pR�d�W�\��$�=��->�'�!*VoL�KCVo����d�%:7��	�8�h��%؎E+���7H>���/ۢ�b�@c��x�i�j޾�ݠ��$�8�KJD7�X�ݒ�[�����������#��*YHSz��&��<�Dp�<��q��4��m�;E^�/��M¼K�L9k!�t��'�d�b\~��.���?��B�gJ~����^.D�u���G� �� �A��P\�K�[L~y	!�UF�5[�o|.#��$��{|y\���s�C̨r?�Sڄ��Z��nVE>����(οoJE�-g��9��O�(���*��BX��]���0h��Ƕ�8%�z��k�&��=�R��y~
9���*{�QL�s/VLx��.�i��dQ����A*�%�^]����:��KM������y���4c^��wۻ�r��:hZ5C�8��=�"{.�$^�F��C�7,���"-ӉH�urx�3sg�&<=�o�����z��2r۲~:KwY6mPU�J�3F45�2�'+��@ӝHz�2=�38��3�EɃ�YX�'U��W�Hg����qJW:�9�����7�S���c;�93+*��9��ڮ�R��Ց��V�_T��������LH��:�6�y��Eyd��俭�?av�-ǲ�^�:\����:��
aE�V=p�4�H�7��#��o���3�T �����r>ѵs��Y��Cwkujs�� Y�,��a�o4I&]�*�h�nB��^P�����\y�]z���C�ߦT�:�