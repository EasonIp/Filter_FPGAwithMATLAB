��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��S}�_��f�`�߃d�7VH��Fu�M>x�{z�0$��c�\x.-�M��h�T���Exp!��p(�}dR� �����m:�"��)u�,��||1.�dn��=��qN��)�tI�ؐ�!�,9�v�2�Ǌ�$w��E���c�D�0�:'�8����Ȃ9�=�Ǣ�0,!�(`�h�h�����
��ݬ�i�U��'�u�JR-Zt��E�wW�{�|ݱE����s?ԳmV���Y	�6���ŷ�T'���=���c��3��g�ɥ�c#w�1?�k��X�x��ƺ)#�s��3s�%�0�R�
����O0�k�GN�L潝m��M��`=ǥz�3�4���d]J*+�BO^�A8�CK�Z��n���J�=�V��w/�ͮSUҔ����64�N�%U5�G���$���� 3,�A�w�wr\��%��>8�F���{LvO(�����l���rK������8����|n��C�����jڠ�Y ]=O�
z�T�m{�=���ׄ/�H���ب:�js�Ű�U�[D�a��'&��4W�ʂ�ף��&���Ԇ�v֏UI�[�g!��A� I���8Xuc�`*g�,�ԶԈ���@(,D�U��L	��D.�K���:y�y7C�n���]� �D�&�?Ƹ��#�L-!4�M����w��u��8���[���+���d4��>�گLX7�[J�ƨ# F��s�0�Vt�������\0ݙ\U��浂G[��|U&C9/����$k�H�'�7���	�2*�e�+����m4�����%U*'�T�n����A�bϋ����j���S� 0�2Bkc3�.*�����-bw7�����b�s ��r���^�or��lO&��݀�;"3ؾӺ�I��2���j]���o���z�"Y��#�#'3���N0�ʥ���
o%��~��. -�J
e9��i�`�7�p�:�Cd4��b�sTpyg�\�w��D,,L��!�J�2{y+���W��8�*���ޗ��_W��DHZO�.g�@��j���;"���Y�e������6s����x���T�cمѮ���б]�Y�}p�_�Ӆ�F��UKs�l��̙�N�s��U���9tw%��3��ץ!E���0�����hJ�y�g��>q�ɲ�lBCrg�1�7��G�� �P��:��J.�����d��V�v1XG�tG-���eV 2��!��/ZMnXa^�+]6��]E��잊��9-��w`-�9���k&��U�r�����y\�+��2�QVH�dFO%VcP���P������)�'s���3�<�#{�����e�AȘ\=#�Ց۳�W�hG�KbV�>��V_���H�2�*�T�����r�S���PK�e[�v�	�I�L�����e!� �����Z�٥e����H+ƛ�����T��0����핒Pk/�lϋ�I�r�~L�bzv<��Iŕqޡ�-���A=�WG�*"<2�\+�B�r]������W�J��|��xހ#y���+Rs��Ä#$y|�ɢ�׽�����2nJ�e[|6Y�t���s����,��N�����y��~f��z��s\bO��
����ܔ����d��e�]�v(�Y���{mt��$�$ Ny��$
��44����o0�q�C�JM�L�䂍����'lȓ�\C��R}�/�w�f���f5�����Ij�k����V�i`.;���s��막˥~@AڠE�!]���@%�=m(���45��%��{I��\�p��O�B8#>P��sN�T.-�Q��j�]"�E�7T�#�Y�tIly�T@��R��宦2r��p�{� �_���l#�9�˂l��a�Լ�9$)f�O���Y˝�G=޳ @벤YAD��v������O�ž)�r=�RS#�x|��\ t�|[Wq�j������0p�A�X�l��u�Qk�'	V�~����.J*��/7A
w��!g���ãe�0�h�k��7)�	s��X�����S<�/s�-L'�*��5����B�)�n���eF3j.���wN$�����.�R� ���3n	�X�A���r����4��욗�u����[V��F�r�Ri)Q��H��srU��d�ߢ�Ϣ�"���P���h��dA�Ie�Cx��	�k�r���^ ��t��t���S�&z`\���w+E9w5Jj����"f�կ}��^ż
=-ZYS��q�i������*���
�Ğ�,ۼ���č�_h� Q����ݵ:���k~�P�{�|���葻���DXm�f��B���5���X�9:���qD׹ۿ��%.a��h�_|U7۪��4h1��W'n$���Iwq���|2��������j˅��қ	�m#�.X�τkg�|��7��d�″S��"��F�ߘ����<�֙���� _wj1��*�u�%(��X�~ػ
�pkBsY�4A�u��j����=kQC�[ȕ�"V�ͳ l�;l��]�!���-�4B_D��J�nO��$��Yp�u�U
�2�A���՝��ʰ�c@2�S(�XzR�J�&4�B�B�z$!� �I�G��BT%9x!ur-��ۃ��:{l��w%Ƿ��H�0�B/2��F�6���bh���kW±�z�S�g�}�)Dh깋|H���Ww,�?KU�^��1%!��j�3��@�ES ���w/�`2�y)j����-��N���;��QU>���M��C!"��;n*n�ٌ��s�|��P9by��%��\�T���a%�!J�^��ၕ��fR};Έ�Q�Io��nC@X#n�
P�ʟ�-�D"�]Rf[�Z᦭1*,a�����K]0R�Tw�UF�nM��z�$i��W�L�䜹O�0kQh����'u���*�-	4�.mC�B+�"��X45�%�Iu�1�̉\y�Bv���$_08k���_��o)��qk�h�崹��4�C�M��p�Xb�����C�G��5��ў�Q_�ǁ����)j?v8:�ɳR�2g�����%X;��U�I�Is�>2[��v�>"�׷V������i"�Pf�1��'gIuo$X�*��C�NS��=A�{lG�۷z}�(D�e^��q��q�|��60CO\�ژ>��B<��8��?	��D�.�����h�J5�0�D�]m�%��؀\1���#ra"�dN�a����C�P�Y�a���N�U��[�C�K�'j��_PZ�(S�)v0���l�s+��x��h+�nR� 4���L�N}aA��:_�Ф=x��d�T�A�\xP�����o ��*�5�$Y�TO�?�B���=�9����n;��p��4�r�5��� Q�w_�I|��'w�'�{3�"��U?�o�У�L��?�%J�?��2�l�T����%�	S�޲uS�䕑4r�m�۸�F1ۨe��@e*PCɅ�����,{#Պ�%�02��>�\���LQW��Ob�:9�3�u��v�p}L��$���8"�^��~�G�^���G���SK�Vx��Wf�wiܗ���)�ԫiQA���Ѿ%�$��J��H.�p_9q�����o�M0�µ������$�8��Ҹ��#�Q�f����	gYX2:D.�#�.��A�}VO�j�<lA�2�v�tQ��u���Պ` {��ϖ�u�jHwP������_y{�+���޹I!ITl �:3My��Q{�X�c((��u09Ql����@�^>�?z�(�<�mse���ޅ!��)�\*4�(7P���3>)���A�nT*�+|nn<���!'��$V��n�U��)ˌ��?j�S�垨W!�#�-uM�*M�3��N���J>	=!�¶�\�J-J��PU,��DMKq�C����ej$D>�x��^k�枺Upmm�<��݀�Q49���U�:¥���� �m����ʦ�W�Ko,λ��x�F����8"+��|�+z�)��3⑅j��sO��ҽ�O�$�i�TЈe�ⲷA~Pqu(�H����c�⿔C�As��Fy�Ҏ3�l�T�n˃)$�	��_�1;i��	I��M~ �b�̉��juu���Z9�hc�_����.�K8A\��x���K�\k��vM��Оr�x|� u����' j��s �����ߟD��>I[T�����2b�ptW1��`���0XhT�(|�X���о������ݭh�q�\i�H�I69)�t6� p�}��X8�_a_$<�b"4�l�Bp8��ͽ�KL���T�����Q��tm�
��Eq͢~	:�̥�������y_�J�h)��<R��s��Х"�G]̼�B�ܣ}�&vw����ɆƢ�hS��kc)��CE�RX�xf\?�Tz9z�pS�'T��j�
Rw��陏�A8�$�U�GN8r5���z�>��Y	���9�W�zNxh��h�1� jҶ�:�![�0�[YGI����3�<��,n���Gi��l�uR����Zi�1:F�u3��kgi{,Ɔ�ɞi�^^�V�u7��v������oA��YV���?G si����L���gq(;������,*Ӛz��Dr��z�.;���F3���2g�sat��Jhb}�� L�L&���C�F�#���&��h3T��	�2gc�(�7HG�>m��~̴�%z����w����!*j����n���\�T��T�at��1�R�6[�3��YB����1'��u�nnj�.�]s�I������!	0Gx V%sr9we�pTq/�N\)z��*�P��$�O�5��Ԃ.��o�#f�39/��gXf�@����n�x��y�A�P]�ol��^��W�+�� d�*{{�N���x�x�&xcF=T��Ż��/O��LI7J�).�����LMɧ.J:n��M�����)!��6W�!4�0M0w�0���څ��/F=��ٚ��W,{��f�c͝�*�  +�8C�P_�4�-���ﺉ�-B��=n ��^��o6��L�+H����e6.N���^v˪�N>�E>�OR�E��q�F¢@��)�̟�K*.��UÊ�j���������� F��X,*�X�]i�^�RV��{�3����㢿�[�ө�wԗZ�W�� �X���KF��MZ#���F_u�R)i.(:?x�+� ����r�i��E�ׯh�?�+�+͇;��&��͉C� @��8�ʮe���}��uM��pH��v U��L�*Tَwʒ�����8�I���Ca�����Xh�
I��_�[w����-A7%��-�$��Z�9��sY�5R���r*nP͛��ɴa�#Ul0s���F���sm��3�ܑ��D�T��S�Tjծ�O� ��8%ĀW��� ��Y����1�r���c���L���}E,��Hi����;=����q�ʈ�8)=�<^�yk(
X�� O0>+��Na�7I]c�o�t��1=���x�$���.H��G��gwd̳��!��f��]�����*�d�~��:�*
܏׸�xa�I{󛾍���;�n�0�7"a��2��-Є`��P�����;)���D��j��u����u(�ޘ��}�	k����?]B�����L�_�݀Xfb�@+�к�"ѱH����rH���wЪ�I��5��H��r�\�jY��'^�n郢"��p�N<���#�\�́QjA�<�k�QUjx3	�J����
q�0��ƧQ�J$��*Jėx�x )Ea�a��[+� R��ft�՗�mA^�k�'r�:@�`~�Fp��3�sT G�MHuM�"���:Y��=��QBأo�� 3��V����Y�ۖm��cV;]{h]�hi� ��l/Z �#�i�R��=+�c�(B����Z��T�t��!���Xm��9j�)�(��%#��u۬jr��"�,�;C�xX����pRnl�B�Q�p,G�3�(�%��OH��3����V��˽������s�u ��� ���v�ʥ��#@T����6U0]0!nB����i�VH(p;[��r�s+@��]uh���h�ħ��F��Ua�D���ʝw���~@Z��}
@}p^'+^i�y)�y�iq�j� _@�y�Uŀ)�)��a>�F}烔�m"���_I���{A��Ε���3�2/5���6�:�}ă����}��ݟ6>'�LvM� �k�YR1@,Vs,�腵���b�+R����3�]�0dN������
�'*�� o�E�=I�F����BC�0%����:�r��u�р����E�ԍ� l�v��� |.����9�,-�v�?����EC�Eo=R���z���9�0���!�gRiL G��YkG1×c��!N�"� }����)����(��|~��Zŵ��{�O��Vy��ޔ=7��=���C��}ʐ,�[p�ADu��"m(���!���"��O.�5�� �|��=V�n��#t%��{zm� �|��5]�g�E�)&^��!,�V��p�����4:.��C���{Xa��7q˰�:��,m��e%�.��A���v`����U�c�ˣ�&z����NDU��PG���?��v��g"6cp1	R픜�]����0�}z-�brq� �6��?���~���� �O(�����V)	&�E�6J$�O/Q��h 	ymE����}(/:Q?Ci�����՜M�B�����}m��\�G�#7��5O�[��^B&����a9���L�47���?,��-�7�~U�xt�I�͵����_�B��	������u� ��u����aH���?JI'kV��Ug��Vl%{�2�������\�F��,�2��Y��(�ցǢ{qNi�8y�z�8 7lV/B���$cF�c�߮��X���YU���q��d�d����gO G��;a -����p �r9;�h�a�O=�O�׆c��"#w���/��5�V�N�?A���#��g�7���2gFMp�V�.�>N���3$;߹�6��X������?jv]-�\j�%Ia��h��$��ېu�%4bS�O�]w�`3M����.H�{��EXH��%�-���Q�/�d"B  H�Y%�ArE"�qOu9�&=��]e_�f��e��{����z�8t+��Pstx��"��9�9��Y#~�'��NB2�/	��P�˸D��$�-T��u�g�ԣ�N�}��W��-d���F��KY��8�Z�SĽ�s��Fsf����:Y�$N~gd�6Ł��f�/��tَ���l��-oe]�br�_��*.�1}�<g���㝽��`�(H3�$jqp^B�J>Yt�e��oc�Bc���y㓷�	��^���	o�æ�fq	X�fy�t�likq��������nF���i�)�k
V��$�aE���&:_qB"�V/�������J�cC���ϧoi=$��`��xƏ�M�uK�e�����@�T��`�o����k$��em�0Ml�(��1����be���~"0��A����spέ����g%�.�5���S�+�n�Z�ԓ?`�$����-�y��4C.��T�E?Z.��\(��ŕ�G&K�4����M�g���e#%Ϳ�#�ܧ��&l�r�{�Z����ʦ��l>����H�BP�T��O����}$0F�~����@#^��L�;�'Vb%�PH��|~5�SK"�O�+�Q#N����(Y�h)�?btޝg�;���8�d>o��にs�J���ٟsB,��<�#Nm�L�ܮz^b=��5ٞ����Z�s�q��"�EKШA r�Ɲa؂T��1��M�W��,^�B��ǘ�:��<G�e� |�9��}a����|XY{���>Z�.��0��C�2 P�Vp�V���WX)�"��%��6u�f���7:]�K��}���{s��8_3��4֔7m䙟�k�>v�
Ud��:#:A�� m��Ywc�B~�3`�މ��$���iڳM�W���>n)Q�L��%!Йq3��*DK��֘�s���.��2V ٪(�̢�4S���|?��Z�N(�Ҵ��簇� �L}��T�$��/}|��Z6P14�@��ɓqe9h���_	�:��� J8HP���0 w��>��M�.�#� ��Pe(ξ�tn��_-�т1D~}^9dݫ�����ʎ"��j�[1H~�� PF�XK؇Q��i��Q��!���_8�oz0�����J��b�������Py^�O+�lK��IT9�h�c����%�5r����za(�ʳ��ڍ`�J�-����$O'j�ZV3�׳EG-�0s+��Y&�1�o��^*�[i�K&��ff��-���&l�����+zө0 $����`�RfWY�����#�/���D1�@̺�:�����x'x��[�����wgM沎�X�1pZ�g������v>�i=��|{>^�=�=/Y�;�������.�,�i�.����'�%���WS3��ɵ`������4���Є3�$�R�o3\�ɥ��<�k��O�e��D'�x�o���m�v�?Š���*&��[��%aV�:�*2#�{_�N���Y��6��1�?0�7
5ՙ��?��4 ��w�PJ��d�w��z�l�hf�������F�z?��C�ҧ�d9YG�lu،�x�n7���،(�|jO=[j 6��#�����^B�Wf*�gzh��x<9͆2r��r-Z����<Db����8��,�a���`�Aƥ�<e����	*�Ջ�o�$�C��@�I��ǧ˿�oEc�XNs=�~��͌l��7�_R�� ��hǋtiÎ0(���҂��~H��cCg8����0[��?�=�f�V9r@��fE}�����*D�{e��w�C7�a�:\�1�Sr�@�
M&���^(t���n�(�6�����[���rߞ���v�W��o+�1��@����'O���������q�]k��N(h�� ����a��O[!+/E!ї�c��&􈅲,�!
(=�p"Y�z��(�5>�fY�~�e�
��qP����?"��GtĲ[���։���8�;B�r��]�@�T����KHF|�Hi�`z��;ND��/kaG�Y��q e�S��BH@o�N�1��J�܁�N"��"�d��z�Yq*Y�c�Vm�X���k���mw�]J�>1��%��ʯ�k�
|%tO�th�(�_b<7`�q�>�� �QK�㳰c�d��ŭ����k�Fw	�ҳ,z8'��Û�L�A��e�x�N�y�M��"���
!�K������QL�l.�,��}7�{�y�Ʊ������Y3`	�33�i��&����k���� ���N�9B,+��e�4��A0 �G�ڢ)�t�d
���v�fr Gl��#$�\ݏ�d�pO,$�����]�)��c:=�)�����\⯙�5�������f�o��â�䋃�Ql��G:
�{�h0�Hi� �#�b�D��Z�!ֻ�s*�}t�4+R�BL��C�H}��Y�t��F�_sA�4���^L̼�ۣ��fw@��^������*�NV��مkSGjۉ>jo�伌������L��Da�X�u��w��(�a�o�S�&����ݎ�~�?g4��x`Q]�og�����K�R�3'^��杨ψ��H�{i��|� ��~�k�*O8���z�[T�7��n
�+���H�`Æ��"��!�<��¡mܑJ&��&�iZ��KroDqe�Z�c3;>��+�T�d����g�*���rZ,}*���5�m�����2����'\���qs[�(���L�k)�d���\b����f���&����n�O���~��r�$8I� hg�}����/��V���ǫ~���
���,c,������Z����;_�a-�.iA6���<x��1��O9ߤ�%w����H$���y$֡�s`��AL�m]�
__4��"�{v��������:`!�̢�X����.��F�MRA�7T_��Ӏ0����̵0b�{��H��Ul�I�%R�X)�V	�#�%�&D��a��^x���޲��Z��.���MwC��u�bO:��I��
��SY��{�*zncJ���c�9��:�F>���XE�Iom��,x2�h�^�#����b�c^���EA<zY0`_�X�� @A�`�����X����r� _G!L�O>}}ц�	�3��Q�d��� G�5[C���V~��B�w14��jHC��u%U
}@c���"����b��=hSf�cN.�
t���h)���q@;����x�+�[c��|n��B�E��kw���߸��t?���n��|alf�3X���MM�N�j��W�̲b>  �;������l5��W�"T�%��ЃSE/9:t{���"/�$�<_�H��1�Kdv�S���HT^���%k���@�B�'�wFb��R?-P���?D.��N.Z������+[+e�J��J���.+nÃ�-�YuZ�r#�"5�74B��)-�ݹ�@�lz�X��Щ/)
���z)2�df�ƥ6��B�p����-�*�uכ�r����Kcx��Z	�ې��p~����Q��\Y����b
xT�"����i��~q޸0���Ұ��� ��1.��́��-3�$-����6�Ij�<��ɤ ���	,Mm��\Rн7�迓�)�%�\X���=��m��Ҳ�!�Ke��o���w�z�4nJ��<AT�O&����dK�)�㌧��G^��Ʋ����$�n�Bg���=��#�su:���v��fU7*�*I�-3�`�����ʌ��5�
H�#�y�I�±�f�!'�m�N3)�`�����vr~�%�Z�ث�e����4�Q���B�U��JH���h �9�/���~)���ho-�g��ԟ�	�g8���Il��?�e��d������x;�X`&��3f�a�h��^�� ���9���6�!>]�z~ahڝ�����,�$Q���՚�`�5��1
��+�q��� �n�:O]�1�_��r{?6�Ո���d�-H�<����+�U� �:'��ڻFj,���Z��wF���2>�*��q� L��ع7��k~ʪ*�%$�>ځ��Dϵg��WJ����-�Pu��]��M���4A���a�G+T��<�R�2?vŐw
7�|���4�<k<p[Nn67����ïr&�$�7��G���B���P��*��J�u���X�Y�6]�M�GJ0��.*�濲W!�6��!j׉������	�car�s�vf�~�hr���	Zlχ �	��b�W�5��+~�oQPǋOZ�E1Bֻ��l��?v�@&�Z��<[}���"Hg�-�1li�m/���>�M>r4��3E��̡^�q�,e�r�,'l Lx��=d�@�q��P-�oj���-:cu�_O�ظ+{q����-X!@�xj�{(�����n�~�\$��W��a��@��_b�Z���SU�v��VB
�6=Z[%גlO��{�K���I�4��u7�Axbq�9jc��S�u_9�H8�/�B/.�,tR����9�-}q˷Mu~�^�S�:���W^������DΟ�؅>OSvo��^rAꃗ{�[���vU8 q˖�؎	w�O�P�S��u��Y��%����J�w�� �S�R?%�u�P���dn��k8�2�;���9O�G������p^��u�1��b��3@�4�WVq�O��}M�溃��񌓹�xbr�©�Σ}�L�t?2غnj�z,Χ�r�����@�(��')�u?
^:��|&�w�p�b	���o�nB�M3��bI�	�]�'XЭOq6�YA�����V��
x�gk?���h:��˷e1;Teegb�u�W����>�3�:Ap��
�Ě�l�RI��,����>;Fzi=%ܛ)�|���-X��4�D�׎����@�2I������\�"7u!������I�'��fAO���Q�(�ۭ����A�%���[b++�g���Y���Ἃ =�a(�V���ʧ��yZ����\�V�~@xI��B�+��V �Vs��`\VB��W�WϮVķ�ģ=��dͺ�����ݎ�%v9aFn5�l�K�A5�T� )���e������X4�@/����0��D��nJF�8�VN�ڞH����Z���3f�}7��Z����òp���
�x��o �ٴR��֪+8G ���0d��F:�[P�w������\=Gi�F�,��$Lw������!OM<4�lJ�L��I���X����.z����O3��8�l��]����(�ҥ�l0'Z�u�<ꯞRd���!�D��&�)�gu	�bۦI3m6�O�r(],r�P�w \��_�e��zTt~6�S\���#(�]�Q�H�r�̩d�U2��1��8�������Gd��}p��� �?0�����SR�Vs6��},k%�uT�.P]ꚂT��P$W�}�*4<�)��I�+����0�	y�O}�|P�j��y7AKR�q�t��d3����*$�$a�d_�JW���o��Z��N�������x@�ھ��4�Ⱦ2�� y��#�D87�� �?��ު��P dr�=Nu� �4�6��'�ȉ��,j��0�IS�'K˔	������Qs����v>'�» &^�2�6�h{��ȃ�zZ{;�)-u2jĞA.�v��'p�a���ʎ���ӾdEW+���&�:6Q��^x�_�͎E1��	~�L���8��o�Œ�