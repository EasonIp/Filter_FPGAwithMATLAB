��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�w�tܔ��@��zATe\��5Â02�}���iL�t�F��������T�NY��y��ti9) j'�A�&e�U( p���9��C�z)N�`�+Q|�w��i��Q̍%�i$NzUC�ﾕ�z��v�K,g�%�zI�_�N��X�:�.g�VZ��hL�_�k�O�P2��!x+�(E��Y��&��3�T]C��`�/�]X/݇��-�q9�%�q�!�g/1���!4@���鲼5��s�^���u{¼Yi�����*�Ev�����Fv��R�?��Ԧ�oY��	_�u�>:��%������h��v'��N���	��eg���3�#[P������dnLG2C_DU!K����A������zGc��,�v����������0y�9ByD
c���v�����/�{�X �Kfͯ��`��'`�S���f�t��河�)^��$m�T*�����"��1j1:��O�U��딾�#L3ɀ�Pz)�Cb�C�<׸�uf_�Oe������X�mZThe� ��3|�����Z^NOV��4W�e�������bJ`M.�KNh�#��u�m�#���S�l��,M�Z-4�n��EM�q�V�/~K�ɶ{�)�q%��Y"(h�ߥUv�S%c{��t8)tφ���ji�E���,!3�5����S#ag�>�̫�yGJ;�Ϧ����֛�G�z��%�7#���L��$��3O�%q6Z�[������pL}'��Yb�U�s�����3t5Ga����M-ʹE�������HnV�sSV��S�4���Ǆ��mm�O�i[z�	Jͺ݁%<B-�lVڮ��-��]�XE$������EA	�H�Ob�]o,�\�V���m�^w�]l�o�?	�D��)ʢ�8���¼J9�ھ��MѢ%��x���N˨�x��VĊ��.��D���11L���om�i;窼�'��(U���C�}d!�<��ջ��*���
K��-�/���NΛ�3�{�&�;��qV�X���/�B%�ؐF��N�x�|��,��:�߾����<�[�z_��C�m ��4�!��W�/��w���M7OI,�eI��yØ�_ݟ���I����JX�:�hW6P���w��Tk&�F /�hc`�j B���.�"�!U{ݤ�n8�I���z��ųK^��A�B��������S}~����<[��2����8���l$F�}�T���Z:?E�y�)�Q����]�,�C噌�όB k�P�x2@
��3�7�m4��fv$4�Sx�n'���dm_�>n���H��M%@�1�ӗRz\�3���g��\��)��� ��7���a��T�K/-[�+��&�DEr�_ן�ȯ�����? ��䣾����(* �(i���]W�:�B3�$�Є4b3���<�O�	�-��Kstϟ0�<BkgXJ2ݱO��6�t�O!L���* wbX>m�BP�W#�.)EE`
�eL�!1jT�̖�8�r._C2�ay��R���9R
�>�̺���Y��kJ�(KKw���(����zlw�n3���4�lP��өca
�4�'R!ÙM�(� 3r��m��s�J)����|�Cv^f���v�