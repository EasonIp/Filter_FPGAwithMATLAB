��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L���"WYj����i� �N�7A!�@<e�]ң�;��5D�監p�.� ^+��Rk0;Õ\z�7PF���p�e��	��j�kdD/���1M���(���T�e+qr)zD���FWkV��������\���mk�*
`�R���	j�' �� m�cD���9:�DhT]�����۶�����i����ޙ%��d7ܷ��	�:���U��(�����#���wv�pFc�o�m?���<�δ�7P����( ��(�����1���o.O����BE�l�pSX�m����
'j�ߑ?�a\����3!����� �@��{`�'�ĉ�FQD-+�d9UUr/�0�A��kzJ����3��º ���i�\1�nn� ��z��S�9 ��j�l�l�jw�Z��o�Y�ʎ��be��Kƿ��4���9:���M	�ְΜI%-���P��N>�r&]~=|�4����Q�{sU����ӦP!1WaO�����5����|��E�m�[��Ns���'��Q�ԧ%�t�����T�+k��^��a�O���lY��E�-��w�"��;���S}��F��l��8�M�� ��K�|{��(Q^�����ݰ�GW2%��M8��!����A��s�B#+W��{���_�1��t��Z� ������'�/����Ԏ�9|�Bzbo�;�a���ɼn�~�G�½ԛ�Z5����V�ܔ���Z㉤¦' �Ob]�߼ƾ���*ӡ,".JK�ңϛK���k�K�c�O����X�=�p�p�:�^7�M���o�8*8�9`���i�YS�-��F�\:�:�꽏�����^�~ì VQ2�Wjx]Ѫ��o)��YЏ����ט�Tg +�����F�-�-�u��|�����Ա��n�
��G���"e�Ϛ�󬯌�!A���]�m��ǱkA�S�MB�&9 �q+�M��B��v&�[1�X3Lׂ���q�T�FcV���XՍ�#ͤ���\d�Jj|��F)���݋tzm3�h�rF7@C�kpT�S�)gH�v�0�Ԍ�������QH�� پ� )$`��5A�Z��y�l���L��$�2���踧�����/{g,�<�M�MA������.^o����M��U~���`u�؍j7J�㓢��wa;�Vqc���ԽD��8��!!�h���w\2D �S=}��5��B���% Td��Q�UU��2��>N�?��!�x�|7I;a�{.;����J�`�ἪT�'t("���c�W�n S*�����l%�d[)�N凉`_�h�pNï��2c��] gֈʯ��h�^��M�C��9������Wp��|�q"�|�����Sh]��RHl�T��l�k�t[�iZ�T�����j��#F��� �
�5�5P�h�oҚZ��
��C��>2�	�kl��-Z�x:���$�3?tm�b��H��}9�\5D�ףj)	��/�۴��5A��M]w�.���AI0E4]_Q�~AR���@�ٕ��z�f_�����eW1��y+��X�],!��Cݒ4����L @̞M��gS�M3[�/����M
�3�U��2�t��H�"*k��<7�
���fY�舶؜��b���t!��_"KHqp��4s��c,�.�@��a��mhj@�.f?�~��k���}!���!"�F��J�;�>窅� �P�vc؅��WhV�LB��!�� �/	��C<�?�����T� j��q  �g�cσ�$����\øf��m}�����ړ�РyM�-��M������˴���ju�&�|�ɐ%'�ξ=�\�����g/RWP��'£���q��E�O�y��ڠ�ԁ�P똝k ��W�zM"k�Oe�,s6��[��l��Cv�6[<2�u�(���e�"�h��7���s��$����|�:��OAꆉ#��Z�S��J�����¶ͅ	�G(M;%�j��<ז�k��{�^�5
�$���/%x]�����+9̛��j2.R.:����R`��<A�_g$�*��9�
�.΄�7NRTu����֗D��z�zyD�)�ً>A֯Ix�v�C����v#���c��"��MѶi	RXv��Qt����F��O �"���s��:�E�T�7�YC�L_��į���p6�?��}
�?EO�KzC�C�_kyxG\��C_ݫ4���1�hT����s�L�Fۢ4�]���ܲp����\� ��V%\��n1�\(�?|f��N����V�o�L��e��k�_D��y�  O������Х~�ˣ-��2N>>�##��h�p�j\��c��1@˸��6����[+�M�Р��V��a:�(JƧR_���#=^R��z���}����E�%���]��T�E#�P��1H9B��b���F�
ɇ���]��/S�_Y�,��h�C��m���+��Λh���Ք�1[��AA@`�K���r۶�f�%��Kf :O)7��>5�Q�ʿ/�Hi�*uP�4�ǲH��^��)J��p�� �nA����>y(��l�{wA�0m �o2��Hj:C�Q�<0�r1���F�5��)~7��}¡����w/@H-3k�Ŀ�ۜث ��Ol��dʯ�	=�h���o'���pP#8=�Pg�-X]�-d��RArvXl��xh��fn�]�[�ޞ��	J=���m7�׶�(������`�χ8����O�/�|
ou���.��㨆�Xz<9�?�@e��:� �G"����vSԼ���ޢ�+k=�,7��<�G�3��/q,6q����*]�=��0�0�2V�u��=��b�J����*X��C6	e����|��4-�K ҿ�ϭ�:t���� 0j<�����o)���)���H4���?p��ă�a���<��F?�4҈4�'�:�Y�8�Z�b�������v�Le>�Ǡd&���y�����r�.S?h�?��eX����%���zsᙋ�WS.��eép�J�9���w?����k�����:�T��vߑ�W<c�������c{(r�{����T���Tr�@�u��qXP�7���̶Э�&�μPI�����5E���������U|���U��3{��TLe��>�!".��!���a��*��SE�祲.d�K�1���-����*]y�1t�+���&��οw+ȡPmIn���G2����yڂ��*A{������J�|Ҿ�bY�P"vx0����p��hk{���F�
Y�7��,����uOM���"�C���G�)W�S[���V���waC ��ƿh��xK�&��pCȥ��n�.
$_��c5���qYZZ��_��)3��F��&��\nŅ�6����d�zoEQ
'��9����^eE4x���FV>*+-{�0VX^j} �ƺ�� 3ިO�^˞a�n3W�l@�E���*���� ��̀�b+`۳�+E��!�ёb8o���|�W�G^7Ý�Ћ��F�|�	y6jb��]�ҫծ���5������|��L�K��؅3����5����'�)sk�Il��c*��YQA�Up��c;H�}Vt�z�0�w�\����)�l����M�Ԃg>A�1l7j�`_�*%.%�?��g';
�%
��������G��y?�t}��*�8R�w��]n�nj^�kQ��w���J����mX�N@8e��7��8f,<��fx��vH�$�E��?Ą	5$s�\]ik��#
;������`s#�������I��
����}��c+7����uD`@�EOa`?���Ř��}��ड़��F�9��S Y��u{�x�;s��V� F
S�@�Xȇ��ل�Y�~���Fԋ�%��t��s�O.��o�8���*������0G�V��U2e��y�Z��4����B�}Q,�lc�=��u�Q��-_�|� ��Y�D��}b.�aZ]�����.16�Q�g�IPoJ-��y�������@��$f�6@�͜M�����~�#���P/l�7���JS��qH�l�H�^�n�4���˲;���u<��e��9h�M{�$(���}�NS��b~�(�|���GZڀ�`�*:��E) +M����|��������qH��'E��O�"V�
���Z��j�&A�5{�D��<���fN+šP��7�Խ-��S.�w�DK3�(a��qV;I�y�L��pc8��8�B�1<��q�b�)�����Թܐ����q�*�F���袡���F{�,��xs���2��K�I���K�JB�;T~��/7� ��N��8e�ƀV�;�"���gƯ���_��޾�C��b��فun^BN-�3	��pFXp�ǅI�5�2掴[�M(�X�d���|��IO���kb���~>k m�ވ��M/1V��X��hol9�@�k4�yj������x����Ԟ�Ѩ�0�-C�M�<�-��M=�|+�Dr:V9s���˔��-8Q�_"!�Hk�}��#T�2%�����Kk%��B�ѓ#g˭��VӸ�ctK4��lX�����(�E���ܰq���D�P�����{R2�U��+YE}!
ܑE�w��Fs���Ie;�{��m;6.�zg�V0v���Pw*��,ͭ!l3�f�Y����|ȇ���O7��1�Y�5!v�\<��
�2��[.x�8�C��`��_ ?l^U�L��h@�BV�~��LD\j2ýG�_|a8��HE��u�nLC�SBU�3����+z��͗����V�Ӎ�c_�k}�8����D�w�3�#H�U�IhMg�YO\�E �vߝyb��$/{���1�^��K�������$y4݋d�Y�M�LYDSڷt��6�z��_�7���θ��eV�CZbt�4 ����f-_F�i'�k��'Ȼ��qmVㆽeS_S2ɯ��H�%�� ��7}����}��0{��U���X��T�o&Pگ�u�tơP�4(�%=	�S���r����`��D����������C�Lqg)#�-E�wm���A�'�AS�}��]w
x��L}<�0����2L�'�
 Gú:MUTs�x�#�Y3+�:_�ď�7�AU$�%a2�j1JZ��*N`�
>$q|M�a������~/|�eU,��h@�ӣ��qCLv7.QF̓�q5?�ߗz�g
$�ǟ�i��ǿN�n��tt�e���~���	�0"¦���f!8lSӹ>d#��sS%*�-ִ���8��cǟ��w�'��ӅG�H�5�yx���f�撀���	�+WM�Q����_�"%�}�խP�zi���ʐ����wl@�#�ʗ44�}�����$ӍE�⧎-����)ƪ�`���Mt�q���i�.B���a���wV1���>���(5��a��C�:�h��g�ыAJ#R)�޾�-�t%�U�<m�3�ٵ�<�9��������3"���]���`��jphU��n�̱f�KSIY�ۿ��jВ�z��cG����@vj�������l6�����T?���1w�S)�,� �er�7T�eLaK��M��X�f��ۘ�}�D�nČ� ���بN1��k�D[wC��:}��$<�^�F9dq<�EK�5��>�9d�`ʚ�E��  �l������E�'������C�G�i�b@���@&ggR�>�Fr!h#��-���1���ܮ��J�'���^ڼiY	��*^�\�����m.���C���<�*-z�\�����C������b��*t�_�REp��V8�`��<O��m�3z�p���Q<eȎ��AW������*O�O��+-���)������h��<�n�zH�UL�_U�JF��$�%[�<Q��-,eB�U� P���Oﯔ+*����о��X���Ĵ�g��q��$���(�!B;���lк�x���i0�� 9^���am��W,<��� ��̳@.'ڡ��r� �߆�x)��X�KVvD���b�=��2�5S|��ǂ����c�p��n�G��*���5O~���XKV~����.�8?]�+d^{-���h	�t�<��ڞ���%swRK�$�� �RZ0E��G���U;2�RQ$��֋K/{����r��g���6D2E���=�A�I��C�	Ja8���,�kQ���=;�$֯5%,¡����:)�j9~�D}�k��Z�Jt����L�.G���q�/dB$�\3^=��'iK?�o:lYIQ��;{ȱ�{�'� ��(ܙ��:�i`��Ŕ��@�jM1�]j� d�(z�+ʢ���`�W�NZ�K�P��u'1A$��lok�J�͐�ͤ4���0�I�0�8��/��:#XZ�Y�Q�&�^T�0tz)��Mnjj��〙
9�^�Aw�95���!�������|b�S.�i�1�6�H�^�`
Cu��6�(|b�f���y��db�Z)��S����Ķ�zEB�#Gxd�f ������xO�|kY�?QȽ����Bm�T<��\�=~e!�D��N3�;��9S�>�N����˚Ł,#�{��JG�.���wfpG�!���l�x��U�\�k�d-8b�����qˢ$?H��x��'�����ܿ��^��I�
�����CPL��>�	%"k�����zc��6��6�{�'�t�Pş����u�E�	(�;Ye<'i�8ş�7�RHI����:r`�1������;�2W�Y݋����좣}�;wQa0س��i&Yr�9�1k�WL�����$o�����b��׬�tBx�B�&{�n�����Md�[���?&�:�gU.m
Y��q��AYm_ۺOK�����#FU�ԵUy�1o����l� ��.\�c�n��s'����b�'��H�j�BA�.@v)X�`};�k�oV[]�tNlK.tF�YPʡ@�ٵ��ͳ�(��#~)#�u�C��߈�Es��{���Aq��3��l��C��ygB�8�6j�$��勜Qb^#�9�(�}2�B��1��#��3v��1B�K�g��E�;�]��G��]�\|�2yP�fH-U�6�ex(�u� �}�6��4���̆���ˮ-d��烁�c���i����A�LS!/o��mf�؃9_oS���-�5Nd����ΎȺ裰�{�@b��������r�;	���j������)��7���2��dP��*�k�W �I��=�Ң��TĬ�kz�>�ٽĀ$0��CϞ�V��HY�X]f��s}H�o9[���3��y��A�K8���V ����{3p�q�c�5�J���h��,g��+�@ �˝����g��q�������ד���PZ�*h�ţ3�@�D���a��}�B����Q���IS� �R���+7�A�����,��3T]@�'c�@������j�_�l�f�1��~I�n��l���v�E���lK�_T�8�!H=n�om6��'"���۠C����$[�?W��v�W���Ą��&'�;q� ʗ����N��T�~a�S&�9<�}/8�/�<��v�cрL��@�k��LF%�E-�����N�z (��>s��4��BD���TS� �؊��&�Cq�I�t W:Ķk�w����>�lm�m�;�G�7=����`�S�f9����^�f��4��I(N�<�z�����l�,U:F>`�q���;�Ք��٪%�s��H����.�����k���.����)�axK:�{[a/m�_}�%��fG��O͚ݨ�G�J��$�:���"0d/'��Z��
���8�KC`�tN踿_��띮��>Q"��*���hm�
�w��-�Ɠv�R�����{B��W�G
\�i\cF"疥e��+F;C�.6�\����pNK�A�o*����O<�]��z(\<]6��k�ƾ2G@��_Ũ��ūmn����6��.���rT�Ш�K���� ����Q��9�cd`��y@�@���þ|(p)���̯{V�)i�yԑ��C���_�$�#������G�;��kҞmgQt� U9b:p}�\'���L2Q�-'&ʕ{�?Q2�5��:"�J�uhz�X��(�N�a	L �V� ���N#dw}~k�>������A�
�]{�x��?��"� I�G���$4,I[#^�;���io�_�N��L"v�.�%yA�������d�NAl���'�U�ݣy>��z:�����u������?�k��S"��!G[x�j\Q���҈�
R{��*�ֳ�3O3�S�񔻪��:ڠ4~C-�0���xE3���:�j���+���.З)�X�.��w���D��+��򭉻�������.+�K���0|�í�v{�uh�;;_n#P�Kc��(�D|�(|A[|�[C	�������{�}>��RQJ�,SN"􈼀R�ND�$����S'���� ��)N s�K��Ё��� ���Hj�~�O���0A�R�k�:oΡPPC��k�����*fXF�Z��T��6�A��1�*��בs��S��y_���{�o5^��*�e���Aq9�)��+e$���.��>�sߎ�(�\����TO�����{�t�}��,�-�f�΀+j���3�������0	r#��WbV������^��)��t��Tx������o<ʙMl�&��-��}��/��)rPE�qpK�67�&LWx�w�\�uغ�����oV���?��VY'Q��ʑ�(�ҷ��Ҏ��"���l�@fz}�0��Ö_������$Q���[�E��J�mZ:q�	�[n1<7���h�9�x�PuymKkn��/]dM�b�d���	L�GMh�����K��Jn	�|���ʹ�9;�c�z�JJ���f���k;+�I��p	�D�C�q��MK�5]�k����W!�`h�N$�� 8��E����u�}?�"�WO=�x�xM*��6h��L�k4���9͖L��UWh�"S!�"��v���ڟ �����ߛR9�>e8~���e*!���#'k@��5|ۂu�.
-p�"��3��+4�+��0vl)�\@z�#]A�,c-�خk~ФE��	 �X��AÏ�[2��� �����?2Ihx����5L���b��2@^X"Z�ל�����d;c<�
�߾�.�
�r�O`:�C�5e7Z�`���N���}��1'��|�4|ۅD:��i�AbD��	X��7I�KƲQ�(�C�i��\���ݹt��P%�h�~j��6�r�V�;�@�_B�<����״H@����P� �y~���B{�H��K�ZB����7�^y:���Vwv*�n+�F�O�̏�`5
�����4�5���#�@*���U�������+��k �۔��ae��v%������K�=�Y�W��뢳��e�7 dȣ�qdg}ʚ��槗P���V�n ^h��XH U
�\�_�	mn��9��Zne@6	2�{}ִ��ӭ��hY�]}������bV*�蒩
�9����Ba�׎�����&Y�!�p�Q����}N���B��U8ljy��82�z�����h)�S����g�*vE���.�p��W�D)�ן|����\�����T@)D�k�Vy��&�L7(�(Փ��I�ҙFs��4O�-����w"xn�J��4�����,�I�� ��	J(*�"�W�m��� �88.iъ�b�&�,27�0�?���h(ݝ��'1$˒�P�SV.RZ�ۭ"^o� 
�	�S:�����mM�3�]�j���UF�>�"��F{��^3��	"���uM��TF��.,C�ds���@]i޹������ƛ�ť#�p�l�<�~F��i�rX�͡BLf �8\:�1���>�Y�tEL�R���w{9�O6-��e�7<x�ܤ@+]]͚�?hz�V�_�y��f	�џɲ7��Ԯ�o�g���?��"R�����I�\�{�pq�K��PU�AVV���U�lƤh0��j_aO�%s�\R��ʲِ��r�IF��uLѶ��(�԰�"E/q	�ݗ.A�e a��݁���ץ�\��q��S�4N��Ҿ�yʩ����?0���y�HR-����)�Ua�U��!������8�|'����l���!�I����	iO�k�hrjgA�gi��qVg������F�0�9��^���Q�k>?�����:��7��dW�#l�^XM�*E�W�;�s2�v��(��.�P��n�XgJ|�14�SY�C��KBy�+��@X`o����)��M����Tt�:��m֠|�s�Ԩ���t�-�8J_���(��8�!�x��m�e��F���rȱ۶9랃����cj��J�h:�=�~q����\�'; ��
ʹ����O����3:+�-�\ԉ��
fk��?X��сEn�N���_ oD�����v
��Z��ZgN�zP�ӓDu??q{�HkN���	�B"�(��S�U��k�F�6IK�0��s:���D��te���U8�nJ&���>8��t$��)qdCmf��s��M�D�CI�Mxu�sis��΂����! RRl B]|2*�e��������� Mc'i)X
 P5�~.�7ZP{�n�FrC�t?
4¾!K���_�2��Þ�³ �M�-���j��ϖ���ʧn3*��ב�n`�� X8���6t���o]�'�����:au���#��~�?r9�n6a�V�['������<����c�70�<�4��D�t��:1LZ	㺓=��,�m�~�]�;k�r-5���q�lQ�����+�b?:���Ə�7��])
���	�^�ʌE0�	�TE'�~['jqe��x{�P(���o��T�[Q���;4Y�f�y@d(rh�u�2!����;P�c����dY�ꃽ��>���@Ӕ�X�'!
���w(a�aݪ�I7Q{��i��{�X�K���D��nm/IWZo�%_J^�  ����M̛�-r�[��D��Ŕ����8}j�g�,�;(̅�Ʀ�N/'kd�l���;1r��Q|UL&$s��u�Rg�>�!H� �;�)�ӣq��J�s������+n7e�>�U�@�`�X";��Y��1y���Cn�G����`�����-�l�	)�=!3�J�wT��fK���񒼜�E
������C��0�T�5�
)!͡�@���:܉aE<����������ؒ�]e��26�y7�L���m���c�@fu �$EZ�/xBK7�AwP�� }�<`������ Kуd��GB��;��ҕ��$��J�q����G�q�jϤ&/���	�5���w	�k8���n��v`h���u�y�z��&��7�PJ6��]��-���E�^)#����,���8��ר��h�3��᷌0�B{�
�1^��#Y��w��5I���6T�-��S�9�NiP�ɮ@�A�4�]�����{�𭴢��ڜIk�,:K�'"��I�S���J5<���5H�j,5����*�z\��J�Z��xқ�7hr�J1�Pl�k0z�T^��La,y;�|�귽�c��(���Dč�y���E.C	'�9U��6&�k�Y� �/��t��m�K��[y�Ġ��kNP�`�����	��-�^*���:�����6����*O���x>���r�E��|n�!���%رh�;+�&򜍁!�ǅ��2SYȹ �+)����q�k�@P�ޏ�W9���P7�V`���J�vv�k30��_�Y���a�X�V{#�)����h��-������-��U��'G���Cr@�t7n�54�#a�i�����B�f}���B�%W�����ۘ�v�)c� ��eY��;����8�^����'I��F��o�e�8R��J��V����d��pԵltK�M���:,Z�z�D�E쏡�����?i��?�CEl��HC���c���1I%ks������]?�����+3#�Mm��֔�rt����e��
���	���E�ot��~Cl��*���N4�!�l�<���m�8��&~���_��`G	%cI<g�FM����ƾ0�����{i��D��X~ӆ���W!�k�PY�b=���;���c��U~L+h�o�b����d�:鑐t�NpDP�u�s@vQ�l�O�d|Vۋ6�?~z���9w�1KV)�fQrGz7���	�Vy ��X��S�M!m��]���A��zB��*�h�L�0�!F`K=��q��_a���r��EKٍt*_�8�d�N�����M\:�ނ���i{5v�	]�K�0����И=�"��?qw�)��a!�c�g��W�qV��& L������(�f"�<��B��m����xȻ�s�}�
��H�(z)���I	=?:G��O����P��]C�J��@@�@� ��˴�6RS��A��m�DxNl;�6�&b=࿍�^m�)�KES���:��� |F�2L�� �̀���t��ˮ^{IΟ�Y��$ȈBKh�U�����r1�T�m���4
��W;�W��Su�c��ڀ��n͈�4ʻ��$�ԇID�4����=y�Cf{��0�x���"X�:ى���|v1���e���|�v��m�t� �i ��֦��s��cn���@9QAr�LZe*Ci�����`:�H���
�����.�����ؽ�$V�J��3��1 �!Xn��� ����Pvqǔ'L2���TM'��k�C��F0�/���q<s�MY�7��F�V|8'K�:��d�����U�W�`�&���*�8��$#C8Og�ς��"$!��U���)E��N�J��t��Ī�$pU�zL.�?��;dv1�l�BK5�8�j$�:0��~~z9��8	��;:�]¸�{�	�1�N����,�-�]X8�>��On9�4���2�� �K���= ���ћ��u6�XC�C���p$��֯��b8���E����1�8�[R����"��c�.��ޣ�jS�AN�;��2�R�7SJqP�hB��[/�~!ЧmJ,�/H��1�.�x�CC�Q���B��r�o�`��]cpdj���h+1gNB���r70b�v���tKjW�u�M�씈fx
{�2�pj�b��Fp�a�ӳ��ѧ�T�N��{�1�e�ʔ�EX�~�����ar�O��JM�ct�����G��JS�9�7٫�Re0V}=.�Uh�3�O�������(-�	#{V8|��i��庇��z'R��wu�ܜ��|mN4b�����K8��9��ȡ���4�'g:�{ἰ;':���T;���p�,�&��/��N{s�Gmc�Y,@+�GLM�ǯ�w2�aν�H<Y�}4��Ġ�;��� �~�'�}� 7]^�譝� ���
V �U��>��%�|�o���N���)'��T���8�.:�O,U���x9^g �Ar�g����%��Y�Dx�s��R�Fu:L��u��~�{�HI�qZ��ʧUjGm�Aag��.�C� �$�G�Vtn�Q0�<�8��jZh��(u�e:2��i �B6�u���M�G]�x�>	9�g���n�Z��RLD�W��T�[X��T��0S��<.���#�[E*�]�:��^-���Go!�،ЊN�3N�$�]/){6�|/r�1H6 �+HWL}��jO�&��?p���p{Ӽ�(�qo�3=t�-���A�=�5�q֗�}1Y; �l�yA�56�Jf ��$���Y9-���H ���;�]'�,$􇟏�N��:����	'ܐ�Qnz�̸F�˕��ҿ\��M�;MO���(�%�GN&zxߓ���������	��1��=�Ր;S��'q,�4-Y|�ѯ��T�AwO��(�c�a��*�����7~����#��4�����8�x#0��8�C��F &LŽ̻|�qhz#�_����hI�!T_�Sl+����W��mʗ��)�޹}�W������:�R8C�!��+d���>�S�U��4p�8�t"SPL���4M��2?��g���db���vi�S�T��ֻ��w⒌���|�TQ�%�z̺�{>��g
-Mb�����d髝4k���E�!���F��ʻ��B;8M�bE�p:j���h�U�c��VN�!ب�1y�%�0��(Ʒ$'�����&a���P������� ���Z��r'�n�e= ���n��!t��y���f-ӈ}�f�|ed���
��JD��q%DƷp��v� I'�w9
N��E�V���]o��X	I;h�)& ���=�\�T�5��v	�LVM��Ȼ4^�)α��$�L5�>;u*�yܬ���*�IR�-_�;n�@�c`�(e1D=Ԭ��{�F�*f��k]}���O\&4n|���z�fR4�;#I��ջh��~ a0��o���O�,���y���=��\����cn�Ap���+��8==�Ń�)�&��>@vg���vr��	1�Ж��_�?��O��n����b���Ȑ��D���y#3~��H�r�c�iTM�e�� %iG���`D�3<(�Ke����u�$)Ȣ����E���c�i�z�L�e�:O�L��˦�R �亯�[��f8�e���$�pe���f����9��]����ߛw���-R���[_�j#��nP6�%��]:o�s�
��3h�����=� �;�f�A!��SiA�3�t����h;���3�I���;f�owt���R��م}*��BS�>C�
-�U������Uad��-�Gc�Ș���v"ƈW��k��g�ٰz���Cb�C��6e�>�>�ւ��D�i�D��D��c���pl���r��b��p��Km �8 ���Tl�Mj�� o��:�c��A�i���̎�Sp�Fx:�g
K�w�}��`sfӀ�%�������N>��y�;��#S�q����������n�V���p�3i��|�UX�>l�WVX��
VT)7�p6?��g��}oEdh��0��_
<�
�_�U�Kp$H贐��a����x2[$0���<1�D�{�O��@C_�wV`q��5<j�v�� ��i7fn���� ʁĀ�8W�;o�
$�#��\&�c�(t�\������Oo:�����1�F�7r����s�c�2m�!<�'�o)K���{M���g�f�n�[AcA��@B��J���W�7�>U�GY���������G��ȣ�Ln�g97��1w>?!=�v�Z˴�gB;L#�ۉ�h_-���7��s]��P��R����د��O�GfQ*M��$y?�'v�X�c�22�[!zyY;M��- �?���56l��1�W��P� �]C.^2���:<" ��ڣNq>P���w,�m��p;�(SP�|��[�o�IU���e�~���6c-���B=��&^_
�`}��¦����?RE�+�]wKf��S^�o ��uq#�%9�RY���Yf(ZO�;��w����9o]�g�E ���iT�u�W���1��\���K�a;�|"�Nj�&f���,�B�çj�Ȏ��VYN읃/~�Et��q��6ޮ�=�@�*+�����Ȧ�k�w���V	6H�X���,�� ���j�] �E
�ξ�$���Ǧ��P�N�~}|5Y.>�	�h��D�u�.�s�$���-EȑƗ;����XR����,DΒFq�@e�%��/��<�V�3�R#�Ӻ�r�s���0��9�$9��vK����\���#���+��ELu�d���"�U_�u��ٖ> B�T}#ݔ.�uz��0��~�v����2l�;h�J�w:H��E�|�w��7�����b�	�ͰNS2�����i�+��#Һ�S�ז�[4� {��#�h�gN���V\��$|P�����ާYL��8�^�b�N7�@��|{��4�a<�(2��9y1�;�Xq4ϳf�����GH�b�O�'sim�|��Jŉ���ź�ޭ��^Œ حU�u�~v	��A[�S���*-��w�O�g/�Xh�{ef����ۇ���i`�5a���n�	ι��,�2���2��^ϔM�� ������=c�Z�x��;#���nbޠǓ��c@��aO�OI�������c�����=�o߫ ��a�h�����9˳���D��JD��v9���m���{�)>0�G�yz����f��k����X�Sz�6Jc��VE�U�EY6�/�T4������U���Z�3��׃��d��+�
��+���y�W6#��~3�}GX ZKy��K9��.�;R���I�L���v�H��0P�2�
����dk�i^Gb��(��Cr���������^^f��gv�F}($��P>j⟄ƕ�?=�����X��U�W$��o�gD�K9a���t40;�2�����L���#�H�B�j��B�m�DD���X�p�w���5_
�Ś�9�ݵR��R�m�B^An�L��کvw�N��[/3��%�����P� Y�T��CNQ!ˌ۞/����2ץE��\RP�+�4��#����?>�Y�ֺ`4>��S@��a`�A!]cn��$�^��t�N�JR����ިZqT����a���ʭ�T<���E�ęZMm�t�Ź��|�3�������6vr���#8�R�6�O|����l!�Co,�/���g	�ة���,rOͧ'%L��P�\�?>8�Ξź�ЁUx�!���xa�$�>%i,I��nҋL:��!�!Sܬ2g�Sw��}A�rf)C��v��盽��=�`���~��QQ�+��E���ݻKӯ+Y�1(�1��� �-��^q�1�oL��J�a�w}�'lF�[��%vm�l%�Kj�ŝ�	Ep�(���ɍ5�Z�2alWՠ���e6,�����C}���I����r���N��/ƹ�z&_OkFz���$�� zH,X�S�p6�_Bͪ����Dw@!	�"<��,ܲ����y=߱ \�Z�`���b����7�L[�[u�J�I�0uV���QbX�>�5b�uK��}wg���+%![����x!�G���b!z� ���e1x��'�^��P��gFP�ɁW���j��yth���Va=IV&t�x�����]XH��f��X�]��l迩j �c��@���d6�J+m�����'��!���.��K�h<JN��*��!����dш���4���
��P�>?�(�U?�FKz���.���#�����d�x�]����尒��+h��R�d������© 8� �(�x����`�UR��6�E�Oè��
�֐Uf/'�L���!��}VRsN;وN!��h.q�e�y�Z�@C�I'0��%^��xb�A:��پ�u�Bگ��o��H��E��%�����R�_�"���P��ܮ�=n�����Y}�b��A���c�#i�NH�P��p�L�V�� �Xc�H������t!�����C��~��������%�Ӊ��?��G�`�o�:�W*��Y\���h�;(��^1�( ��K�k�`���V��Ș����ԖW�W�w/�i+�U&gn�nt�%c��ha&��C�@<|Q2���el�3�=�h\祿�9* @�h��P3�͎�� H'q��y(�`9JpQ6Wi���z����K�qA��~{u��XVo���G��Ͼ� �Fj�.d�M�Թ����7u{���3����3���+kFp
�p�H�݁�1��j:�.Y
38>q@���yT�ރ��=G	���	�W�&&�6�D�MB*C�����a|d���I��D���;�1L6z/{cp�_c�����kt'�)�(%��]5�AIpȭ�#�8Q59������~�d8���^�΅�Q��G��w ��%��X���S��Ơ�v�B�P:g7�NL�_���xA�8�a�t�o96�k�v�~�Ҧn���w�^N���=Ub�z�|�ײt��]:[��`|7z�	�2<)�M�b2g�E�W�0���-7AȴX	H�-Jg��w(x4ki;�%�c ��z�m #NM��G��}u�X�s��R���[�A���X�H�X"N�i�����r:N�v�fM�˥aL�#>E0s e����Q���7T�|��k��|{[ּ�mA��I��n���;+nm@��c��N��.G|�����6(&a��V�� �d�}�
�|� ��(��V5ҳ�
�E���@&|s���J��5��$+ҺS$z���~����ʑmы�;��G<@��ϵ��^����|a�BpݮHumg��3�0K�0�����ic���i��ȏ�$nGe5��Y�*������Z���O	����I������5�o��Y�@=�[kq'��)U��7He����r��&�DA�dn�u���=�-��:�j�p�A�	9"pS�&1A�>وw��P�P/a1�ԯ������FwD�����M!��[��M��=��MU����#�
��*�yx�S������Yw��+Z#��#���o-�I�K���S��vCg�m�X���̔��I���c� 5g�.�Fu ?+�M�͸lJ.��fV�ȅh���]]��
���;WG���_SX �l��u33������9�\&�������{	9U���	���ݷۆ�q8��s��1�	&��U��?s�ׄЫJMb�uLV�	l��Fw��[ORT�Sa������;�.���3Nb��*�s|�|WM�	q��/�� :�t��"G��|�qU2�}"o�@i������V6�3���0�� ��̴Bp��/A<�g��x6��ݥr�_����lw��]5��x��������W�Si�����4�o.1m��-=���&�r?����a�THؑ2l����������g�B�Щ��yo���]��HV�y�!p&Ǻ�P��o9��s��h�W�-���꥓�{>��՜y���e<Q���S;W��-�ac�Ck��)h��Ij	d��J�"�hF;�B s����i�l������㮢�/�Vy���.�^��o~b���He�oՍJ���G�����qw�\��1��C@�� ���}Ċ�V7�nKL2���t�F�y����m��4�y��U�~�G�Y_v*YmB5�|b�R���%��
�FQK�n��T����<��Gz�����UT%a�V�7�������0�O(�I�`4<c�6�S����Gc���˧��fz#�O���/��]i{l��\�]t���Z�RB��g#uԑ�w̝$�\a�/|{�CNZ����e'#��+�u����+p�g�.��<� $��.�A�<�)�;�rE��+��L<�>r7����L�1o
ڹ�z<$q���5OP\n�;U���J@j]�W�E�¬t����mdR��p@�#�G� �.H)Ç�`s�NH)%~F��ˠA�J�P�Uv9�lxz�Sq�`s�iȚ(�ۺ%O�]�~��'tC�TO9�1�0���E;���uM>O�kc���� v-�ȶ��	����S��h6 8�i���N:
q˄�^�*��Y1�f�>�'0�	O�)�C��@e$y��&엠�2�(�AiW�!���P�1�O�,8����n����w8)|s��Ҷ79=�h�%�1o���@�4�,CF�V�� h���E�g�9��i0%	�5�*>�!�R��@��+f��P�@�3t(����B����,��� �b�,��f�e葕0�S1�7��{�U���	w��-�� ���ndל��p�ۿH\mP흋�R6���G{P��˔�L��:�پ��t�6�9�4+�"�?e8�G��v��h�^$���,a�}��A1�?��OO,>H85�Kl� ���
ts$����)	�4TϚ�dy�MP����v��yL�:O�گ8J\݄��	v�uQP���b��zَ�yws�v���l�j��7����q�v�l�=$���i�IΔ��w��� ��\a)d�* 銥F�$���H����߱�Z��8��=��@&��65ç�9.
�6��i�X؎�d�e�������O��lV�7��&�9�B\��G�X������0@�]���G>�V$�P6reJ�^�.}_�8��"S���zq�77y��+�uhb��v�N�~�*�;ݹ��.VN���?�� t>Y���>�+cw��Kо�6Un�Q㎕k�q��@�y<%����.���؎]�>2���p��%V����7�uR�9&��cV���3��٬�a��[q\p�ᖨ.�*|��v����yl��޲��Om��,|��2����P.|ӿj�D��,�e�6� ׸�n��,8}���q�ŝR���DX@LK'?��Z�=E�3`�ޯ��b� �yDr�Qh���am�U�O�h3r	$?�	H:@�&���~S�R]�u�{�()���* �?6��5��/s.��?���mn�x?���Sy7#�dF�fl�r��O���_�����U��"ڐ9�$�LB23��^�]�=���*�AA.D��g����{ۢkf߹�!}�G	iK�)��@��L���}��7�����y\�+�1#o��Vǒ"��I���"�N�u)��������/�1�b�&����̬��c���Yyi*f�X�'�BB�-`����[(	�����Q��{*f�ڜsp���;��k��ꖮ�y���-9YB�)7�7[p����	�r�k���Y�' Ϭ���`���q���r�I{�:9<g�X�Lp�
��r}�$J?ySݫ�5��~Y�ǹ7�'.3 �yg�8E�I��0S$�h�c���Rfv,�3��'ti��MKН�hO�}�L�Td축ޥ�+h��e�tq��_m  sƬ�o�>U����@��-E)��(O��9��ғ��]n�a���Y���Xo���JCT_10�$��������Z6�e���9�1�R�C���r�f3���#�[K���_�%���J��`��C�62,YkAN�/��Շo�,�tn�s�tꙝφ���cJ��g.Wbe��"���aB�f\�6/��yQ�8�4��^c'w����J�N�mVp
X�ǔ�jk�hs��.���rB!�`a.z�Ѡl����@��uJ�� U�`JF���
���`dQ�ve��^e#>���ׯ��8�ɬݙQ��zW:wX�+����kGEz��;"�Β���T���E���v��''�l�/Y��Bh�Ǩ40V�x��_v�O��q�ƪ��a�F�H�B1]�U��f���S�-whO��&=��y��8�j��t��d�{`���,Us��l�"�1-g [����.0���-$���"5�!�&bpҾ8�?؅�Wμd]-��0� .�M{�����R��#B� �;Fu}P�ƽ��}��1T���ID��[1�4��1%����r��^Db���Y��g1i<�N/T����hj)�^dL+��(�#K�W��l��2b���v@���R^ɐDkb/C[�%F�w��S�Mh�p��^L���8wV�8;t�%t%�H
$w�2�G^%H-~0���zI_��S�T[��_&���MOOP���'��T'	��t�'~���A�����F7Y��{"+�h̿�_���z<�;�QIW�;��:�lY�&c�N-vm��r��C3�°���eY��o�DW@ߡ��}uv©���Yl��)��Cy�h`_`J�|`T��gS��6H2_������5҈�&cz�̛Aë�=S�b!���q0�����(� ؟Z{�[bz�����=@3�Fo�@ٷ�m*�e�z�V��l>�-8�*k���1�z,JA=�i;oL�!��~�����x�BQ�	�sPʷ��G;���e��'�$�ss��_�S٫f�~���x��M+�}���P^_�| �ZX���`�Ϝ-������ ��2����h:�B�=*^��H���g��@+�"�c�lq��;���*p�����;H��;ł��ۥ��S�ݤ<�%ڜ��A���o	:��A��u�vrD_�vO��M�l��;e����2�ˬh�ͫ��e�g`ƦL�tk}��Ŀ���T"�ܩʰ��:�Ik$��y7L/�L�ny�iSʏ�zT=�/�M}�c��C�N1t�����dS� ���E-Aҡ}6�L��Ff��e�N#�!��٥��$S���m����.������e.��~��XO�y�@wP�FN�BC��uV�@i>��'4�g4?�'��ez�܊�W��;&�!D.1O1��0:�9�>����z�gj2f���+|�롧=5�]R�X������Q�|�<@��E8��a��E�@��~�