��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��ʻ�X�՝PW������P ��
�f,w���U�/�|p��Tȇ����/O�����7�$�.�>Vn��n�m�x����g�v�����cj�5+j���ރ�L�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�z�b�&��R�'�F92īQ�-��r���n�]�9}:���=YJ��N|� e��3�
F2��w�*�3���� 2���1h?�vˀ�m,0��ZR׻Q��Ѧ�l<뉈���[g�Ђ�JR�M�I������?O	v�	�� Ψ��{OZɀs3p(���u��>^*��:wK��V�4w��	���h��&Υ1��b[:%y&"f�Ou�ɫ@�Ʃ�NƆ��Y�t�@bw��nd#�g�u��ys=�]�$Z��ev��H���s��ީ�{+������蜂�C8'j��B�;2��w��@Z���$ԽTT�K]��q�rx|�e��`�9��
7hm�GjH�Zx����uߋq��
c��z�B���G�*�Y9A!�A����[�|9��]8$�aژO�d�hl_D����Q1FG��A0c=+��ʧ:�[��d�j�k�K���G�������H2LV� c�'��_ �u�������0���$�⃉wX�v��gA0�eq��ʨ؛��jJ��`g|�[ Ԑ;��"�ߦ�F;�,�c�H�H�Sb�W.��5g	Гt%1$�R�k.qS��ܢ
�h���=9-��7��B�_	�D��A�H�����j���������޼�_�*�)�� �U��ߖ���wA?JLh�;����p'2a�T�4	�ǽ�+�����FިU�+*x��ɿm�e�����N�@ͦT-B�]�g�=�\1Q���2��\�c��k�gѿ��X�>M7,e��w� ����&�Ν��?ˢ�i�+f�8v=��%޻��y$��)D� �̄>+���3��4-�$|F�T]��Fn��&�x��5,�}�51�
q�Z�G����/3͞�O˼�m�%؝����#��_֯�&9��9��j�,�2���j�(Q��M��ck3.2�U�L�棸`��������eǠLsu�>U$�Ր4��IX�l�;n����U�o�o'X��ơ�0��@	G�\���=j�������R��@Z;��ܷc����=
`��'O%��G�إ������M�c�f�*=�Mzwd`�i�7�X��%�Z�`56���D��R�	l����y�خ����1e1�>�c��3T#���G��he�
��'6�):G���_��6%0��z�-�N�Dp��2�x�Ҋ��ydx*en���ɒtx/�b]�sA�t��r|�ˊ?�ٗL�sY��?�w�)� "�4���D�4aOC��c�S�@���v��p= ���n�Ol��(�;#�5�%��^6_LCp�{�ZϠ�ȅ�7_�l�Ǉ�3O@z���G;����*�6�co�P?�x�n!��O
���(�)��	�i=���mǝ;G����4��I�4�׿�v�9�ʂ�I� �����I��b5�n���r̈́��j�5+�m��A��*��IB��])��럈����}+�IW�JzJ"#��[��-#N�K��16�ϬM�BV�O�O���<�1T`�G����7�P!�Ź�0ݲR]޼qE�{��X0�81�m�+������X�5�%jK7ߓ{���i�IH[-Ƚ��o���%�\>e'�3�i^ؕ�-��� ]7<������4o�I�Z�w�[	���V?�t�uG[�x��B���L�7�@f�}V;�r��u�2�?���N�RY,�V�7� ȕ�pL��4��q�s�k}F1�Yϟ��+����	���&<+�ۤ\�mv�FĀAU�܆1�!�\�}��Y�FM����{�)��|�?D���`=R��q������{�W�#���#�'U&�c��;E�`E��M�㝠:V��#�ys����Zy����N��Z
z��]b�.ho7�1�H#=�:����'��4�ޔK8E�{F��G�C#xI��E.��g��J�P�FFBSc�h�"��0��;M6�y�gy�nMq��WA��J�-+U bo��F���fq�S�L5&���)l}7|��w���D̚�r)ԃc9���(O�[b�Is��Xj �����asl�b+7��Ƈ�seJ��� �~�����K/T��0�3y�6c(h���껥��4h 7��!h�ط�9�\��c���Kc?�'7���=0���uF����^q|����.������t�xEj�%��]�t+�a��&j�_��;qK$N�DD�m���L�FD�z��V虹n�-u BPI����tө�/&���V��sΣ�}��#�P$ڗ�
]�{ྊ��T��F.%9ykq��:?k��.���y���U{����"�Q�(�t\0nSV8gqN�ڨ��Z�|Q{��������.��$��t�� ָ�%Z,��ݟ ��9�O��M<�T��4瓚�t�]�� �����Y�u�r�\;h��RW�i�>��IS���sV?wo�����;5��ז����B�Z�~Dۊ��V�.��a��	�Đ�li5A)�q�1�
bkl���ڔ�`��#��Xm��<Y���f>h�e�Mx�=�V��E��u����;��ԍ'�ج\��9�{�N�7w�C�ޱ�nS���N�[���!C�@�n���g�o�]�`8Y,�qpL��s�R���Q��0��F��".ՌS�Z"��%ۿ����Q����W`�ˤ��F����_�ԓ��#����5�u�Uw~�i�n&���K��O�s6�O��9�a�����vkd���S�L�]?1��ژ��	k�9Ǟ�-Nd��D�V�ng.畁�V���O>�����0��QR��3��d����L�ߓ��ղ���/�	��A_�ro��jX��@�?��a](y�I:�Ș�;�{��*�@��zX��eϓ�W<$�p�R��'�`"��J��f�ۘ�W��A��-��s�u�Z��g(������]�hB��-��{����������-����IqM�
.�J���R�������H��
�aW���v�*�K��ee5��Z8��Q_j�u�U^����kw���5���}�0���Kq-��.��Zz
�:�42�Υ�<�"��Ko�
;��a��LN�h΍�����]��?b�!�&n^z���Ø���G%��S�^��$)�/�w�S�+�&q�@�d����S<P���	؃g "��7��ͣ�/N8ⶱ-T���n'(:�<���
)M,SeB}i��<H���K�R��u��t�E��\����>�ȩM�G�E��>��Lur���aU.ㆂjB�?��{�-����^`N!�% �����=~�5\�A���T�Q�\[�6�_�/n$�W'�D�<��i��S�&��P.=�_