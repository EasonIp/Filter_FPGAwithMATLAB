��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,G��U�	�oJZ�@�z�����>*Q�p��~!}8~��m��sDmN��3\��\�A,��y��,�y'Zs9|�v�G��Z��J;����`��"��t�������UnRt��8WP�Z#+ϙ���\���~��/M���jы�IFA�ާ�z���"����ĎKY� Ҝ��Z$��v�̥_���b �V����2��O	>@2�Ĭ��E!���m�'���)�\��P9L}K��͋M��a�ا� �F�Ed4��S1ϗ����i�)���T��|��rf����}?�6a�"��*�'�6 -�|8����>�6y�m\rNY9�k�᭽�; {�D��m�B��CW'��t�(4���ga�뿢��WcSRof�O �|���S��� �<����|y^`w%�_��Md�f/BA�o����h�VH�4YQ��M6Ó	��U���$k��Ln��XoA�G���o�YE�ÅP�rM����ϰ
&an_~��){S�Ϙ����Q.�|)��7(�~���m�rVhn�����k���{0B�b{�R�z�J�L{�.��,nN�OG�}�Kcm�DT�Jс	�0����\*���eG �����H-$c�}3��^?�����I#�F�����E�84)Ю�@�&$�r�?u�����Z�����tY�E\i����M�w[�|�x�r<=�(�#�s�ͅZ u35�%������^��x�M�%n������E&�N�FW� ֠�Qt��=�O$\81�	*�=�k�jcR�ş�U[.�s��s���g�C:TM��b�	bCqE
x��u3ҒօQF�R�7^�ͻJ�9��_`�e��Z�1�F�qq���	ff�U5'�K�AD��4*X��zΗ9�o"����kٝ����>���h��g1���S1[���Z8�P;�]n�Qz�f;0��b�̞��}�5N�`6}}�u�n��㫉���y��!����'���n����&<d1��K�gU�Fz6Mt�}d�߅G�SOe�Zd�=#�=��cPX�l�8���g���
,����zG�&kTģC�ꪨ��Ϭ����OjD�<hk?���O���9��/�!��06��҄�I�9�%�YS��b{�}�5|,��R��R6܊�o��1lI��
���?{�h��(]F3��)2������Q��1��������#��j�̧ؿ&̎FSu4+ F����GG��4��T�,|7�Eՙd�jn����5Ϲ�q��P�'Y�6��Ii�f6�}�r���/�:�����Go�lK�Oe�.5<	�ً�Q/
�w���C���"���<������7e9����8�����00� �����X�d/2w����t�J�6���s��O5Fdp.�&�"�&��nj5u�q�|�x%-�>��ݞC����WP�L=��&R��z��S��91��?}�[S����22�*�X�i�ʖ�����,�fh̻�R��
���8!�b��G^k��#�0��ϟ�������XaxR@ K!8�f���aLEh�X4�Bz�Ʃ'��v$WL�g�Һz���1�#�$0�0��/v:M	�����i7��ng��%��J�D�%UmWW���ӽ1�	�_{��`��|~8�=U��q-��۪��in|6���p՜��z%AB��I�D�Y���9 �8���e��.� �&>�!U��I|z0����IE(ε\����t�`�����O%�Ŋ^dN�vr(9��2� fO9ྀ�w�~3`,�(���R��!CXE4����!�^��7!�"�L�E��[�`Y�ү�6��e�D�i0a��X�Zn�Q�H�������LR�����+���x����w�i~����%?!%�`���d?�ʄ�xL�|&����~3�կJ�WߘH(o:τ@�Ɛ�����`My�\q�0�z6u�^�]�X�L�{��ybs�'�{3�G(��e^���/�k�񎄅z�`����nҳʧP��f���x��0�jO�?*a&?'U���r4g��P�<$� ��8uR_<�ֵ#��`JGm5��o��38�,W� �͉=V�	�x0�)�x/ڝ�����n��5G�}�^y�L�b
��w�<�#�t �Y�^���q$gQ�RH�{;>���㡷�>�C��<}���P5j۰l�Z,�9���`&�z}�Δ�0������AyueqE�2�H{t�Q�4'j2����Ծ�������8����z�_**<M��wߣ�vL׃�{?�p�;@�G�ꢜ���������;��t��w����Z�ǔ��b�g�^ϖ��wpk��j����[#��d��v�i��$��j?j�9�~O�5����h����K�������h���-��Y]2+x���E�5�X�$�KmB��Y��M��>���Nsp��R�;F/n�s���!dK�q�
��-*ݓ6�Yw�P�GP�6	Z�/RUD�M5�j�V����@ѽ�̩]E���ְ�7��j��n��[k���� /�B4C��P��f4>��yW F��˴Is_s>�A������͠C�\j�v<>�מIӥI�@��M.�2�wV�)�.���F��t�v&�����ҟ�o�G=��̕Z�9��X"J++#�H��c�|75���n��n᭸���e���2�MM��2�~�( �x���++��=�Zk�ϧrW>uD����I)i6��:�H�
���D�mX�w�����٦�`5TD1��\��7��h�Ö6ӣK(H\H�l�F'��/ՙ��`�;ħXĝ�l�%�I��4��q��X�D^r(^w����㪞�33bVD���y���V��|���gHe�!��u�[��hҟYT3x�n����1�:SV|"����$�I:�����T�&#������:���č@(�;��qKۇ��X�+�g���? �g3`u��q?;��չW���nf��ON�'����S� ��Ӡ�\F�������2"ŵj8�Q
w�"q���Fk�uh���4��B1�[��!����Q��$<и���ZH���E��1!���~�Qq\R�o�W��TX���Ҽ����|��Zxڙѝ�w%���/��}�����Wu"��c�'Ӂd�d���9�	����HZ7����w��π)����@C���^:�J�QO<��;�[������������KJگ��ol�U��rb?x��^;_����Dos,ا��x`��Z��UH�$ы��a2��Z#����3��H)�2��L�E2�a�H{7Q�duG�*.�͂�������^�.�1�d�bT3g�lQ�~+\ue�4ͫnI՚�������ALl�J�{���F�U����7dԲ�l��{&���Dn�ˢ���sq�C����!�:�8�RL�\f�p���kG�������r<R/2DCAh��k3���6����n�����u�N 8sټȝR.�Jۆn.�&h*�#t:;�A���٥�y��oK���x�[>gZ��|��� �����K"��M[t�ǎ?��1�$�L,7,_��p�'C�C�aA�d��Pl������ҍ�>�	7�\����C�����Ck>��~�煫-R��f���i[�
Ϻ��>�Z�����6x���I�XH����F�h��$�BYa��ѪE�]�*��ۦ3�`+{2xDՑP��s�;C�»���XH�_�.�K��2�cO	AR� ͗��*��D�R^$G3���4�W� ��m���`�� ��}X� �"�g��-X:�*BP��+�$��=Q�n�X������&��}cs|]0��1�հr���yK�Ew}�c��/H�6�D�	89��5!^.�~}���}un	)�^pl�1(r��:�K��b��m���I�����oS��i�E�.5�sP�|�[{�ݙ�gG'bኀ2z�D��ewuX��.�dK֞Ћ$�����DzJ�+;GP�(|���Y��9���šz�m�_Sº��nƻ���|�vz��k� �̢3_.V�G��=Xk4`E�f��!�0eZ��#�`$��9�y4e=Z���7��hjL1߀B��y�/�E혝�h�,�Q�(�U��D��r�)��p���}ñ�yD@-�Xd�����9r(RaC�:s������̻�"+�t�O�h�]���
��/�kZ����\�L�\4ә*G�W��|�n7���q�I�p����/�y�i����L^���ޢ�v�e����n"��ۺ����r�&>�6��F5��� j'0{����D���(2q���f������>U�2/��4�������t%�d���/�g��
��e��u�-l���8��.��z���Vׅ���}�,�"�8'%&����i��]���i
�{b�Xl^a�[���ѵK1��<8e�%ΒY�=Ʀ^權���f��b�B��I,y&��|�=��П}�_-���]��uAۄ-��==�O1���Y��m����?>�tQ�J� �s�iW�b����'�Ė���iT>8��Om�'m��&��c�9w:��?XPm�V;��du�H�2h�o'�/� �&��`��Y�d�f����TL�i���kN3�:U|�����NZ5�b��Ζ�z�Z��EQ��� ǵ���=�z�5�4�WѺ�PbϏ�£l�}��"��9X���&�<DV����lT���VA<����t��I�e-6�5�9n|Vk)6Ԍo$R��S)K��8B���������g��F��"�"���Y�%��!�r�l��,7�NU�u�"5��/��CTn<�v��X��R�F9�����>K���5́�gT�Y��"0қ�PA|JH2F�?��IГ�r�ҳ��X��eOf�&*|���#�<�3��L�Y�/��p�瞲A����d���Ep�hr� ~J��3�3M��)���b$��n����� &��U/�{� e.V��b��@<]<G��`6H��a�l�H�Ӑ�h�jX:x�t57whÃ{/�	�0%x��p���_��=?�m��%q4ڻ�ܫ�ϻ�p����] nfC��H�3�v�A�J���_�L�(��֫P�&����R��J��?�1z�C�1}�Ba�׎`�
��$��PPr\o![ı�BLHɵyo!���+6���q<cP#4�m`�n�	L�xΟ&���f,�AɎ�`l�oA�����yr�rGD���A�b�;ʛ�B�A'9ˆ��_hiػ[	�{��5��"�V.m���jae76��%�(��EM=��tS�p�^���2�^�߉�84��?�5���lcC!_ҳ_���FG|�@���Ac֮��w(��w�p0�u�P�B�W��K�?7��]�d�z�׭Clx@Ns��H
�#��ɢ�Q
� j@w	��±B�9��"�GSW.�����v���Y������
��ay-�̱n�E��D���B��z�{MB��⮦������g�A�R���&�d�o�cwl� р6��z\K��!y"c�z�=� �����J�:W3t|�|�E������.�|��nd!��PQ�D��_���>H�om���oh	���Gᱫ�9 �N�S����<�Y	�s�]*��-<93*�6wMJ��~Oh=��n�!����>*WdF�,9��1}�Eg�~��ۯ�)��79�������� ���_�����K���	�����*�Ҥ�Ө�&]����E�;�j�ƣ�?���<CB�@d_0�yˆ2߂�nN����G���{��-n��"]��>c�y1��L���SS ��d��㡲
:�a`�djz��Z��?�^b7h��H���tqf�z�׺�n����d;��7�PU�i5e>����n{����*� ps��ۢ�3�G� Z n�*t��*3��Beƚ�Q�hc8Y��i�ҎR�Spq�p��޺@�F~�jVj����-��ƛ����T�IR�VT>��8��iS�1����\W��:9E�y	OP��Nβ�d]�$��CÄ���Ef���;U�4eMq���H���X�r�(\���lŖ.���^��� ��jJ^y� ����^�ɬ)޶��y�߬nˬ���_֔1:�{��W��E\�bh�� ּ"�6l���� <��4��H-�5�g�p�� ]��M�N:������:�ȕ<qꐼ���\����0�xJ�];�����L�t�7waC�+���s�4#l��'J�G���b��r+�HoS����^�Og�F��1�2�i[�>[�vA���͗R�\�>L?��r�/�@Of����E�m�k��(�ӫ�4�OJv���|��pd�1�4oP]M���������Ks�Y��R%?���]5
�P�7�;{�M�+1{T�
D�����ܵ���fS~.j�b���\;�_m�M8U����b����ಓ�'΍9�