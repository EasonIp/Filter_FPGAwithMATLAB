��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�J��"4�=�7(�T�JѺ�ő��,\��s���ӣ�F�؏�
�N���8F�CP�Ҙ!z��Q	�{��V8����G?�5� 9�����c����X�H>P�E�}�.L�-o��ŧght*3ٜ<�Q�;{�0ȗ�`K.�pͯ��A�%q�{i{�nwYF^�)&���w���ӊC3E@�p}��$��:�+0[��ԭH��<��VD-ь�N��((��(|MdS�`N��X7�F�7{��8�c���O�7����h���S)����Sԑ3�q\ߊ���|�*���in�2���w��7ok,�M����,-kٵ�By ��j+Ɂ�nY�V�n�gV'�]vÌX���^������I�k#����{�m凼0ʻ�#"p�Q��Y.ߊ��~�x��yM%~��#�Xƻ��%{ǽ�mg�9��a�N��l�r��`�ӱW� �`z)ɜ^�~���{}�A|4�y�_kT���N�Q�,��X]��C���2���\�<8���!�Uf��[�*V۞Jo�,��n�%�fnX��5ql_���Q_{Q:'{.>�V4�� o�ηXw)R�/��Gٷ�<̕E{���V�N�M�?/|�D�5Ad�{��	N�}��DF����ʚ��B* ː�����] Ƞ��O��~�k���<�@�uJ���:�N��v�a��"���t��4��(�X6����Pu�iWL\����Q5�G��#?�?-W�lc�@c�D�rmA�AiO3�]"&��ގOċ��e�M�����R_�{xo�,�� WJ�3�C�P<�)�yq�mR�8��Gޏ[ߙ�G��G(m�ج�3i��� ����V?���6�}����J�IE�P�Ú��t�*2��> ���F� ��	��v�V��RO�C�=����-��,zŞm<��1��M>(d���>��_�iy���*0��H{�G����#ˠ1t���0E�+)<~W���N�u��4P�7y@vW
��Ur�</���K�=&
�q�iƈ��$��2Vk�Tʋ��Km�e��P��~����L�^�0�A�S0`7Y�$�����#�q腭���~�T"���JS㧧�U�矢P�n����b�5�b�J�q�-�h�y��G^��$�_��-�8��H�Y�t����CT�ԥ�e:�.�$�Y2*c�(�q��O�,��"�d7N*-����Sq�߸�<�sǐT�6��l�V�ޒG���t�>Q��"U���9�tz��[� ����W"�#���2�<j ���yTt���!��9��l�W-y&��j	�1S��ZN�4�N�Y.�t䄯�)M���L����;:��4^FԳ<5�Q%x_�_&jX�@��u8p���o@	Gp��:}�!�P6w�9vF�4$�f�����ksH�l���9�*KN��֞�)�O<���!����VF���l�����\ީ�@ϓ��Y��˫�;���ؤ]�
"����QLV���DC;����e��|K<)���c�[s>&���{/Z���c��ƣ<SZ������֠��rqp����n�@���zs?+�n�� ��lL��P��~��wN��(Q�q���z}QI�������2�#���L��|Q<���b8�Kp����BԌ�S#����@FX�4/�K��g��NcS�&�y��K�"?f���G����_��_� �g��#�<ce��A��� ��DPv�^��r���M1$ B�A�UK4a'̯�U*UY�����)�_�ߞ��)Z�)�z	�����Ĭ���a�̎w9��<�QԦl�<�p�v��O�
	�A�)��C�W��⬝�͗��@����(�:�ƵM�A͏PO�Ō�}�Cc�!uh�^�h���uIc0��CW`��� _��Lt���%��=�D+�����yI���C�T�$�����>����]�l;ԛ�laP#����A�AQ�b���}W1��7��'�[{ZBb��I3�f�v�}�-g���w2)��QΈ����������ͳ���9�^�A���]��(E�Yy����%s}��߶��,����č��҂���{�H���'~{{���,�-�)���V|��o8�ED����Ј�<�A'ğ���_u��M��z��'},��ƌ-� �pU����ÖħP��ۃW�<��3�{�Y<��k�c�P�@kهN�:��+��
�A�Ka�kg&��1�m�����1�Y�2�CE�褠L�J	��TX�<`WT�K6�?s�,����ѫ[��دQ���tRгP4�*ӛ�{�J\���A������}�Tgu��UlY�,/���M�dq�cT�cé�u�#|^U�U��xn�F|¾e�����.l?#��5A�Y9_�iC O���/)I�&�<�u�z?c�e`(*�)�=�h���
�Ul )P�ka9z�L��7�{�d�e{1�f��O����5s�g�r���G!��=�����߸�d\!����+�M��g�Ӊ��U^�]̙ky3,:@�+�2���))���鳒"s���l^Q��r����廒�������0����Ga���{���f�Z՟b��s|�U�7lp?1TCD���b���gx���,�Yȕ5��
Z�E��g���9b���@�_��^�$C)��M2�����A��0/h7��>��;�ɜT3�A��[�h�1�X>�����O��:}ĸb<s��]A@.���b@ ��rwح�s7((�Cs9�L��� �<R�������?T� c��M��+Quꋤ�L���Q���m �8GF�|�TW�*�V�:���M'D���6�A�qT	�ꝗР�_>%F���~]�\FԸ�#^�J;��S+(S8K��6���{�$Ggt�[:̄5��vY�|��l��O��������2�3r#�*��p��<9r���ߛ��9����c{2�̻����m�jB	8��SX;QL'�'m�$���7�v���c��@vۓJ���I5^��*6��"Z0�U/���ci�glǌ����m�j?Ș�zr��ykpi��ƙ�p}������@`���]3���QJ�>���.�G��	�����H#�o����x�%�vs�f{�=����	y�x%��=��O<U��=�vC������	��ψvT1��u�3�7���������%��)���d��3� ��~ ��C�-@Ҍ���^�}z@���J$ٖN�t� 1ї�JG��{\�)B����tC�d���7���7f����I<A3=-���ą����c(^��m^,������1�u��(ꎔ�8�t��'�d�H��k��k��8���#|R�rb�)M�U\k�OC-�:�(� �W,x��i���j�R����6,�A��I>��F�a�[���w��H��jr�9�T�A Z~�b����l�{��SǼI�e��B��+���1�1Q�Ca���dA�$�(�iU��`嵔�Cne"�]�ʜ�+ݺ��pظ��������L�u}nYuCI��۰2G�Y�N��.�U���L(�V�<HƷE� 	�x���+����&��|���`P|�������D;;L�N����+`���E�{5�fS�8m�-�8�N���o�^LW���ڒ<�K�GS� ,CRCoI/u-�Dt��%�S�YS���A�񄀇���2O�1�(��f�~��o�mys�;�5f� I;���s4�x�	��B��(\祊 (f,Ke�����)#�pe����:¢r�U��3X�K�iѹ�vD##j�c�Fٌ�Rw��J�����ǹ����I{(�u�S�.�w��kn����u\g^�B�.��Yq�.:�>���^z��pHs6�3�t�7YHҮ�3Dg7%��܌���D-�BY-ːo�
�"����)��d��V�5�s;@��i'o[K�}&�F<yM���.T4�Izx�H�H��y@���m
d�l,�
�Ϲ��!����|���K�+x��&rj��Z�<dl���/!��t�-U&�İq�Ϟ��xM33WX]�F�I�"���U9}휳�����R��ak��U鄡_�0������ 4V|mPp�����l��~M}����C��V<JV:�lH~b��;xn8q�� �IuZ�8x����(y���Ra
I%e�_��P�[��kG"�>�[$$�h���bX@T�8&��,���	������(D�u���!/� �ν��6�`9�t"�eW1o/Q-wAЂ����f�
�l~ӻ����[5�zLId�9�&�ç��j��mu�Q�U!V-L/$j �anT�:�D�I��]���11(N-v�c�|�;�̏a�=[6>�%�}�_� ���&ui����kMlW�Bճ�S��&P�fLT�A�fV�nP�^H����zqG..Q�Rr0�7nu9'lph����2�g�D��x	��(�����'hTױ�U3�(:Z5$�jhbJ1��D���2<��@n�8&��:��`G8v�g�1� �Ca �KO*�8Z�:h�T�u�Yxm���»���>'.�a"'>|1w�t�x:��n��j�Wt��f��J��ܧT��y��#O�y"PdHe-IXң���.H��[�C�j���h3$�؎C��Fa���rL��e�PGfl��'��E��V�!K��lN��ąI{kz݋��O�ZkPv�hx1�����>�EI#�fO�}�퇢Zj|2���7�ѥ�t����v�Ds?:j��̡Q̪�=Y��V���WuFh��2I�bۀ��{VVS���$o�
����n�tυ|1���Ƨ��iq+��ۏu��ͩk�d��R�|��Y8��wK��l�8�S�	砳������d,r\;SQ�Jh��r�#��#��I��s����o6�|�6���H�oJ��lh��b������r����>��t���&�	)�V�ɡ\VP)��M"�5��ysӎ�[�O�3u�j���ŌD��e����5�CH��FB��k:m�_�Y�O�N��sap��{kL���Q�Csi���u��ތ?A\�6[lM[���k6�v-���!Szq!u��luCT
�
����Cl��+2��4iۥ<�,�P:�����[$5��x2�G��9e������>���� #̲�G���t�"���6�qL`WB?K0�w�j�������ж}����}h[���Tz�T�j�������	���[�u�f$	���h�u�p�+/�҆-���w�.������3�)X��cHj;�)m`h\���*����)8K	���^����1������cw�_�A���P��+��Q��u�ح���X�q��>cF6�,��ʺ�F1���\��Uφ"��;r�!�;5�Ҍ� �-�^,e*tC��Ce��w;��{y�\�3��D�(��.#��oTV�U}]�Q�+շe� Rl�d������,�Lb� �˒|��U$-t
h���~MJ���W��&��O�2^�h���É�]��|Q�{��ro�Ш"Yg2�`���@%�{{O�&Y��B�NmvX�X���k����l~�x�d\�Q�������Joe�lR��v����93�FO��`d�\S�~�ģ��eղm���E.�%L�ɨ�"Q��5�y~`�<	ݞ?�@�f�i���8���Y��mo��Y����S�6��*1���R1��{�t5�xӸ���\�2Hq����K��iM9�W	Idq|�dg]}�'���B���A2��諳G/Uv�{X�;QR#�m@~���2U����{<��_<���>*�q�@O�F��hylI�K&��C���M���yx��ްE�ca m�ITw�'��d*��]J�;m:����b�\���ܵL7 ���`��'�q�8pG}�,2K�v�N�q�@�t���D�cs��	+�%b/;�A���>�e�u�5�]����;�6^S���j��Ce���
�����O�:�\�b/�� ;�C���χә��aEk�d2ٓ?}���|l���k]��T�{��U��:�����Wm�'�e�ܬg�7��8���(�f6�e��*����ݽ91���`��/x1EO��3�����mp'�iVD��2y��
JEZ\n�?9��EwCd��	�P�_�:nɘۤ/�8e�� l���Rb}�Ձ��Z��q�����E����[��}�%�I}EM��crexD��%q�x��9ԧNO��D={\��	L��=����X^��s]g�<�H������r�mFCx�KR�,��8;S�篢^P�p��kgy�9]�£lzCĳ�mq�wC�#��V{p��Gג��(�7릊3�u���P����B_�J!�/R)~�X�)B�8�7�4����L���f9�����(|�N{��fܹ��� �S�ɊZ'��1)�[-s���n��$�ip�2ͺg�Q�^$B���]������R�}�M�2��[0�_�n%�M�Rt�#t R<)P��K�;)ʢ�Ż^
Q3=eC쎈<�� ��^3��q���1�ScJ`�%?��5�>w +べ�̐[*��y;=v^�n.Ԝ�w���uK����RR�nP�;����@V�1���~��M"���w�y�b�a�|�谭BA��q �-�xj�V��M��0�jֱ�P�u5x%fɷ�x}>������H�������}��:m����'U��
� ��<�`���҃�Z�?PX�BW%uR��*�D�V�C�H}w���<���	qCTy�v�;֘7���{<	�o���u���NL���49�Q��V#�����]|wi��e�;�O��Nf���xUGB�hV�y�P��`ܬ�yL+߁g�S�Y�9��0G��π��������-i�?5�����N��N��a�zG"ι_2��&�T��&�/m���ׂۃ,˵�B��y�@0�^$�����GE��P���wwP�oL:�-�Zڸ����Hq_ǫՕ+<�\�PPC抧U+:�ڏ����E��'��\N��ٺђ�@��-�#?�a�_`�R��O�W�hH�`�;�94ȴQ��+�#V�]�I{��r�]��oF����-O��A���a�_��KK����jP���}�mxz`�y5eMػ���e���%��٪Z����I!�L �
�/X��ڍ���X9:E�!���T>'v � 3��؛���a�ͪ��N���� 'n��%���!�/��O���I��̺ν���ʯ�MXx͉��\w�ɎT��N���@I��8&Ө�V����`ى��5"�v����4�c=���2�,�j�:x�<��ǉճYYԤooW��������)F4�/k����
t7���Ј���;*9�����E
�"#��w��GQ�l�5Ȯ$��|�Ξ4δV��헝�����"g��^�	�t�F�
�Y}l���~�-���(Kkc��7�t��x����I�K"��<1�(>d�5T�Ouu���_���SP� F(�u����އ{adgg�a ��$d�ۚ_uE���S��^fv+׸��@�·Պ����Ң�BD����R=�Ub���j�O0{j�{�J��M}v#7�w����Q�D��%I�������d���P�W$�Gٕc�i�lo�{$��6�����,�P'�|�9�hSST����S8�;�Q�k�_�
��
����+�,1��6g��{�P����׻��ʄ�tv"��)���fsc�2����{�:�όt��l�ݧM�n�a!5:YW|���'����S�,pߡ�J�|���N��M�`��Q��E"���P�:��YY0����|�EI�4�:�X��S+ }^[-��I�e	>��f�]��ׅe���G�֬�0T?a���i��=�Y$6�}Z�^�u%�xtX]��e�n~1�y�6�W�:3�٘$�"Ĳ;�b���(4�Yؘ��J����n��s�;���Ŕ�:<���WC9�.�)����A���.m�ogUa��,��Μ44F�Ki��@v���ź�A�c�Sp�c��~���q�9u��?60��:&k���Åq���!Ǡ��øY��Hڝ�|Z�:?VE�[��^~ÄP��8;�{ 
��W��H6&^��_u6p��}�T�D���m���V�i0�MsME_�]Mg��w+r
�_/��e��c�0�G�������6���K+�c�(��R.G�Ǭ7X2�/��L�)���P�
vCK� <P���LZ���}
Ķ�6O!��P
�
F��9e�D���!�����*�r�[�̕4�|f� ��{b�<��w���T�<B#����ё¶���c	�� �4�X[b�,"JM!�R{&���1�cn'fn���&���N�g�e���K�<�Rv}�*�B�бq}�I���R�#E�ܳ�:�O(ʺݺ���^(t�����G)���Ͻ��A��)(_k�d�|��uEl� �M�����=ф�w87���=��R�o�BV���"�S��mP0���6dmDE��-96ۄ�
�^q尗
y��&5Ƒ�}e�z�����&v�ˢ'{��̈́�؂4���o��'cq�~�.�y�� 9�'�3�����x ��m�B�{�d��	)�)-�qn���o:��_:�Bz?�3w�� �uP ����B2��82C�ǆ���#��>�s-Y��x��O�i�Ccɂ㨞�,��&�J��c��iT�&�O��ņC�m,�N���zܺ(&Ͳks\���9�S�#M��V���۹f9v7��
8O�Evt�c�);�#�� ���R�@�3�~#D����y���)�NZ��r��^��sF�}�=��0-�2���{.�D~�+�I{�p�62�!�3�|��Wj\(�)�;�E�d�<P�'7�������Nk"�S٥�O��beĈ`�k����.XXP���p��s�nL/����T��R$�6X�~nO� �� �Q5���:���У�"C:�����&���ς=>�����X��bM �&�NYf�5��N�|��"m�X���"+�I&��/.�۳̭�E��{pJV�֌TN3{�Ȥ��o�h�C����g���n�R�P��ms��W9a3w>��l�ӄ�^D
c*^���D�oT��O�M�z�'TV��v(c�y%O"�~���c���a��Bд�{����E;{���eՏ���I
�`�����51f�rl(��ӻn���E�͹~���qNO<�������Cѱ^݃��l������t~ �-�Y�t�!���ʜ���k��7F�ܵ�doLA���钋VR�0I˺j5\~x��Y�
����얇%
�*�F_�YF�R�h��\fFJ��0_r�½�ӡ���
�Ƞ� ��1��܃z������ ��K$�^P�T�� ��Z!?j7A�4�)aV�xf�J� ��.����	�oz�{���]d�����S����/�����hM2h����Xg:�&��3Q�X�pn����O7n��0�?·�nѺ�D���_�6u�_�C�iYjy����=U�C�$1��yJ�P�}�m�׆�N,���.����CuϗN媯\�=Q�2��At'��&^g���b	ɔ��v-�J�
����Hk����jmY�#6�풾�?6@�{�z��K�2��K��D���>�d�5��XZS����^)(�#_X��%���B���U��AU���Y��[f����d��sC��h���X2��Z,\�U~�d�����CxG�HM+�V���F[�1�����/�&e�҄`KXTLbg ���Q�5@�r���~�C'�}�.�b�ғ����mF���i;S��8��~VY�O�~l��n�K��B�d�X%ZD�*��/�C�39�5q��$�D�da�SYq�jXdy���*����[/��Ґ���M���Ӎ��U[pjlg<�����%��s9{Vhi�{X.7VN�	�:N!L�]�.�tK�R�p�V��f� @�����˂����T�d�P<�i��0'e��jd��RA�5�6��*��g���YA�=f�k�}�)IYq��vɤU���6�d��,�f6��_���:��I�/U�xx|���0��X��.���ѕ>�Y��~��D�=:Z	F���"d��
��/E��0��+-���zD���̴E"�������P����$���9ġ��oV�l�ȿ#���c�����܀���� �]��R4{)U/EiwyN��%ذ3ua���9�.�s������t̐`�d�m'-[�f��%��a=
�)���!8�NE��^�J�Z$Ʋh%����o?ҊbY�� N��{�*�e��g�`Cmó�{�-�(��<3��]Ҭ	��9h㤞�rIԵ}�	��gP�cO�v����]�
�R$�(��! 4�.ӄ2��Y���k�_=3��萠�'�O�J�/����X%���� �B�ҍ֝��rr�×��m��b�e���la�L>��v��q>i��tHzj��d��wol_�r����z��KR�KV�W!�_�/v0�ɵ1�J�����p�LԢM�e�öy�yN��\QIUM�-�OЧ�uc���*���ǜ=!���7��IW�U!Lȱn\'���Jк��|c�G�tɹ��p;9��8���ˍ�H���l�a�u6#�:/Czm氕��J�?�0���DW��:��D6��j������e�3P�t4F�ێ��K_���M ���U���(�׈T�A�h+���7=��E��5y�Lɧ�96�)�F���n�U��X� s�"%�Vd<���%+[X$Z\����HL�D����3{���.9��8�ޕ;���k#��ΡB&�ڊ15��w?����+�|q�b�\wF����'���Dl�6{�8�ݏ�}��K��	߼��2��9^qZ�����τݭ�Q:٭yRo��&� L�
�	�k�Tzhs����X�h��812	A��S@;A��1e r��x͠!+U|��C�:�vZ\�a�!����fhK-��'���jm8�.}?\�c�,kff���sś�EWqW������Aur��B���;������}�����@�4�G�Ix:@
[�Z(��V	0cB�[����+��m� 7]P=;�`Ap�5�mk���~	f��0
������f��� 4�b�"��6�98A�U|�"�rK~>�����J�W��)K=�"�t��f����~~�J��-��N�U�:V*����&�nԌ+��\�$)b�]��͒p�����K��eǮ�	����0YjBK>4�lk?�Y���C"�c��j��g�_���V"qz#��a�ò"�%Q}M�,�=	g�D�pY>�`P�TE�M���)�C�����L�*�D��1��w�rW7���Ke�|��6M��|$�s��F`�M�X�f� QՀ�^2oĠ,n�3.>���Y��vv�p"�����z_�}���������=��/Q���L��=HLR��]�Q�lMփ,`"�/C���1�����8�dT?�W�6��u�#��|�p�-��ij�!g������h~_������N�ߴxo|�� T�Ő]'�q��#�Q����2�OQ[';<�x � g�",-���ߦ�f�M������6�e!4��
ȯҙk8w�R�s�q��[����]��l�}��sG/����xPz�n�|�j�'�m��M���q�a�����d��a�a�턦��w�e��i�[��,��%v�֮W��4/- ��gj�\��3޷kֺ�p��#��B��F�E~��A�=�<��>�=Bz��Z����'B\�A�1(c���W�1x~5���5��9=f�}S��^�[�'0��-/��kW0���p��m�
��zǛ�<��e0�,燥�4	���/�E�'�fi[�>9݈.�����ǦĔT��E`��!MHr;������@�Ĥ���q}��*A�M�l��I�@�/�
q��O�CEt�N^K�A��z��li��]����f]KA\������@�ú���!���o��A)vj��ͬ��r��.���Y��P�J_ x~gk�	��/u#�9M4kp@?���z�����܏�#��˳�����gk�y>HG}�ʾţK8�g%���S~=�9/��ͲU��8H�߯"T��(Ѽ�i��'-P,�ln����ım<���E��!z�]�j�h81-I�H�9�J�� �P(&�)��G5��F�y�;�5�@^�ѳ����������-d%hc�zۊMl[Ɖԭ��' �������U-[���Ǻ�l3�`^p»��ݭE;���p�G���}�Fc�o����F��a*���_���~�k�����
r_�w֞�-V�j��=ʍM(D��pz�k�Kb<���)��=�\�Qf�|A&�;��q���Be����hT��P�kn���a����³y��|��5T��iIx�"��L֏����*�e+HW�&Éd!����a)�\���òһB�P���O�4��F�o���t��47{'�#�����Ϡ ��_���t�ʳ���m<k�������f���nPjѼ��и>(x�7&�JX��-�N�Y���Ϻ���C��g�xV�໨���c�&U�J�]f>����%�O��ĸr:��2I�J���%�k��{��q��xU-0��ZB��#���՛ ����HYS�0ub,�Z��^��cI~S�-�8�;�5zo#8���OX�}�?S�9G1���g����JTr�
�\��6 %`Y��̾J<��u�h�ι�����.��n׈��l5\(�\����{�2��S�WX��6�o(��@�� Š���O��L0	i�0'�?N(G�?4��w�Y�9���JDL�_	c��6���,]4�<�� �w�=OY���������*"�6��=	#�T.����9n=4�K����GX�[N�G?g��E�����~����Y��k�d����C�:
��_�b�K�'i�(7-n�z�P�,�Y�_^A��O�Y���!��'�M鍑|��g+FT����R�dEܱ�����q�O^��\"��2�)�pm(M*��0�uF�M�K�zH02ǲyLᏤ �sq�ZFz\��ZP���*9������b�'���r�W�c܂D㮼+� K<@��� ������O�5q:P�*�OT��#�6/�E�T9�6�3����p�n��[4�ߜzW/r^���!
� _�j�4*d������6����җ2~ZIHC���n�A�\�f�K"X�)���F��~l�L���Gd%�d3�Ȼ|T!�`������R�Q��.�a^hP(��r ���Jv7U�唝iM��5��2[CL��qʩ��
�vW�f��\�49_��0��8Ē�y�S����p��15Y}j��?= �Q��i�� <,ڮ��fz��x�'��s蓂�O����|^�ӈ�=_Ļᅿ�"�	m�Z���Vg��y8(C���Ƭjy��޿�t^8#�����Ds���yIȈY<'J`��4f���ӱªg5?�|~�sE�Sy�$k�ȋ_PYb�ي��,~�?�������H7�!�7+�'�����L�F�}�2��Gw�(�f0�d]�%,ܸ��v���YaS��A&Y�5��h=(��c�|z��	���s,��i�m��;1���u�W�/�M�̄ϧwx5���Z��):Ay�Ŗ�s��+�q0��aM��i}#sH�>$hE%m�FQ@�'��	���3�Ұ�H�����"���[����Eg��{Y+^ZO��<T+����Ș�c���c�Ո�)rU���X٨�6�rh�;����7�k��ᗖs�Mm�����!n��3}l�# ]ia�Y�����CR�طR)A���$^�U��D<?C����t���ۑ��PW����5����,ք������)*�`4�^�@��͌y>m���V8Iv)��:��9>�ė'Xi@g/�8���o�i��:Z#���#$��n\���tC�I���E^s�Y��2��ĳ� �t���^C�_�8��?	�ME����:Sk � �?�M��+W�;�<���dQ~t��S�x��kK~�<�a[̠�@%����\s���ii���w��^F틳�_�R�[�L�L�<y�7�s�V��0n>����#�4�G�+p�'0uǟ=,'e:%��z�i6\�.�?� %�s$��@:��oS� �)o�^�~~U�茹\�wU�[�O�=�}ur�c|�*�03�o)�eQCT��|��e��Q"- ��˴tH��UNF �4�a���yє�R�R������=:�['U�-�	����x_Z:p�M݄�J�;�.�ߗ�r�f�c�7����t}�2s�<��PK�@;b�u"�X�;ɛ�ؾ۝$�t�{�����F>��
Tv�"�+�"(����ß���m��YӲ�(�m$�̱��޹Q�����d���d�4����{���z�������"Nr��F0b�s��z����ۡ�,�8����~���������i�ȥ��H%��[iZ[�Zˎ�ԍk�9�1�6���zq~	֣��_3�G'�!��i����w)ht��W���ci�>�`�P&[��[-��u3o���̬5���M[Ĭ����Cm$�����2|�}8��ܱ���&����K��W!)w\���{iW}�@��rdו��}��������.�Ni�m@;���%�K��t����r���4eTdO�:0t�����~aL
�W���x$Ǳ�Hemw�r�������� �k�P烆k�ަ>d�n0��B,�>��w}��jy�Oz��Hv֛3�:ϸszW�Ln��{�œ�?�`�
�O�l|iaNÖ��*�X�<��IZ�(T]�h�{آ��\z����'���R��qߖ��ڶ|0�����%2�;�6�qxkL������7Rٳ���������@W	�G�B����_d���ZΓ�w��
��9Kkv�\� bL�C���)�T����.�xJ�� r�A�e_VS�c[�rh��?+�)�ȴK~�ˊТ�x*(�u�#�T/:V�qt�p��B�`���mUq�/�P�{��x /ʯ�ެ��`@����^J�~"�����������7�Aj�5d~9����,�]�����  ��f�΁�b��B
�\�tT�������������r���Pm��v����a�g�c�@���ʪU��m����
�&��2.��L�VS�U7������ISEóK��-�ŀU,�+T �I�����Fc��Y�{X��Te����f1�g��ܼ=/'�n���ɲ� &�M����{�9)oJ_`�.�ey�qT��^�U� �����.�緑v�{|�m����X~����XD>FRx�����uu�A9`�'B�h)M���!�``f�����ϭ�u���ʭ��� �nr�(;I�ė!����� �Q|��o^��)��F�o#�Qx� �˨�x	-o�n�x;��mJf�{Q�\���^V�g�I��r,�q�
��Y(���
�.��7������/Զ� ����Hd�KҢ�I��\:����G�V���px���܏�6ՠv��������]���+ų�u���f׀�e��O��KZ5�;� �CƜ��z@s<�Z#��� n6(�~@�T���8(��gԞ"�Hm�@�]�UGD�,�@p��j�Xuo NV��`^Ѝ�!��K����E��{R�M�f�ڡ\H��}�zt�E��ո�5�J��G���tsj�5�a�j�+��A+{c���>�"�{V���ջ�E�l�r��_V�1�]	�L/PGL�`VUh�B��!N�-g#=�6*��0�� 1�+�B�"&+s#&魧�&�R��o��.:�>�7Me��=�%[��J��;������*���A �����D�Μ�o0m��t�^��j����֙B�	Z����C%�-<&*'h"?��������$��e��#�(4�(��W�'D�̐}�` ;��9�G��OH�����^7D�i>u#�s��s�����-~XL"mw�)�d4�|t�:J]-+�j� ����E;�*l�СȄ�e6�)�j=�� ��Dy�tV�mi!�,��)1����
T G�─���d�8oAιR:���4����!��I���E}Z.�AE� �M�)h�1�e�'��/_/S���|�>��8��ɭ���i���Y�Tq�`Ì,k��=�Q�=	������$�fH��+k��M�)�]�v�1p���[LP���Z�C��ɲ��@j�\P4H ����y�	��yL�>�ؐ���)VH�I��>�ԭ)R��NC��4?y���m$!6[zl{E�I�N������}/��rᙙk�Q� k~L��,j=�^6�B�,��qh#m����t���Q����֦@��IrNd�"X��$t���T�+�ǚ��C��X�^��}����3E�2����3�YQ� �M8�j]l��ڋEZ�����'~E���ǈ�_[�ޫ��j!���1���Ɔ۬�|��X��a����>������ƣr�d�+��S�Ζ4���aI�b��:��* u�T(��T:�>'���UEiHJ`[�5��IE:^�轉<Z�����[�@�6�%XA��_��aQKg��2'�D��i!! �Վ� |��o,#"���#^Yk�)��L��Sh7�l&فO�<�=x��u�r=P�Wh4��n�R��ᘠF݈���Ź��)�{���Gm��4T"o��/��\��0^���&pY�Gp����l6�B���Do@[eh(��T�s�薵��iDQ@��ޮ���mt��[���YH�����t�t"vE�<�Ҫ�/��"�@��"��s�d��ږ�6�� �N�	��4�?����B��W��� ���eSU���ͺ'����+����ۏ�q�' �g�!�e�g��������^hҏa��\��L��5�Xɻ��t�/,�A�p����2#v<s2�߈�j:�K��$��h���j>[�wF����"��?�Ԓ*������Xg �j`����J�x��a��C��M>�v�$����oTG�|Wmg�2F��[����V�z�SO�h�P�R��'o⵮bŸF�3����4�&J�kD�[7����m��JNb!�F��O5�Lv���� S�7\����ߛ���v\p��n6~:C����Y�] %�)-wW�U�% �0�I�KY-�B�Y"��o �u��Ѡ��:%K�,YN��zJ�J�,��m�_�J�R�{��2�e���}�k�-�W�=V���r��q��Sߋ���P���@�s3�,���	�R��-{EW=���+����%)-�΋̓�Y[�O�b����Ғ�Dgj����=	�0��0��4����傲�5-+ ӂ(	�
,1�_��O�p���O�h����3,;�=��=��J�c�M�A��
����.\�w��B�3�#^��Ů)BP�.�����Q<R�+.����tGD��f��͹~>�K9�i�q�D5����|pW�;6$�B�<3ɓ���-~��g��X��$�Z��	�����,�V�S�1~d��S\r�b^�1�Q�?��g�L���A�$szu�VF <2�~��8�m�Ec#���8�R�wF�5����8���Y�5t�BA2U@G�⮊ԲZ�n-�ˀ��l�`�|P�� ����(�؈+U�J�*�p�T[��2�4C�fW���^�L�^$�A�e����v(����C������ܦ�X^�R�HwF	%��o\'9��	_x��n����#s
��O7��OkM'��E�^f���5ȼ�|N�ȑ;��"��un�QТ����v�}�H�����FQC:������Ӂ�n=9E�����%���r�y��+J��N�g��/2�2b�mnZ?�m��*�ց��7>�8�B)_x��c����o��s�p�[d�k��B.�z�^YmOɈJ=��k�WE�`��~�w�����$P���Cx ���yE�|��u�a0B�V!R��{��w*Z�'���X2���]F@��⃲S��@�A�<��$��K�F��S�e���"Q�=Ze�D8D��X����b�mr'�P�	h�9�
/�u��4c�n��MQi���H��س"��3��P�p'��֋�P���+�\�m�Y�#B��u�Wul���n �=�ie�}Ǭ��wC�=:(�;8MUCq�v0]DR� ���S�D�Vgk�K�<$��͵��\`��.��%�%Pҽ��Ƭ}M<4=�0ݿ�v�ʹ7�4�y���qr�$�=$u��~=�LʎZ��8�0�0r!��U�f�p�I)j��c�mM�(�c鳶"zE�fZ9��k�#m��rHJ��(b|�E/{��lZ������o$�L�)"e;��d��D�L5ْ��=�j]9�)�A���+�eMs_�md�n��w�l�s1�7�����/R�)�ܷ��EZ:�W�V�-������}�sܥ�ex^��c`����)~�Zy���;�|8.i�("g�'"/(�۽%T��K��.n�n4��D���ݕe���y�i}�q��G�0k�mk���کa��!�K�.��+���D��~����1����<�����g���o�!��9��G¡�2�CP75�q�)"I���Q2��U�qk*���d_&�f�x���=1g�E�7m�eU��O���6q�@t3v�iYm9H���o//l������_Ӏ�TO�=P��]z�(�ׅ��5��̗���r�k|@�ܡ4�J��.��͸7i�N��!3+�d��I�%Sq�]�M|�9�HG���O#�swhը���Z�=���v
ߘzngJ
AMs]r��T�!z��������)�%�k�F+Qm)�԰��΍iNc؁?s��o����}�d.daH��Mm��-��Ŝ㭱�eN�Q�۽�d,� �WR��r2mL�=�J��%\W��co����_f�w��DzU9�3��i@�F�����IE@~N��-7R�O&@����;	̳�0�H !���M����ƚ�:���P�Q��cG9P �V�;�U�_����땊��{CK^]������yx]:���M����3����"F�B���)� ��C�2w=r���� ��!xQx���hO��Ж�Ev��
>�ju��)��I��њv��&�J%4o@�=P-�o�^����ӌ/^B���=��Ι�6'��%�(������d��'y��F⊰o�Y�� �^�T�\��,���#��L��� �;V���DJ<�W�|/�Ղ���&6��Gp�Zc��J ]%��AJ�q%L
��7J�(Z�S j���	1�BS����C#;��A�F�17����j��Z��y�0}� 1�*�j�O�Ϗ�������+��`K��Z�է^��l�Ww�a���
��xWN���{��Ǆ��S�NL��so�r��K#��ߔe+�As�]7��<4s��|yb�J���v=.7��)n�����x�%{46t+x;0�Zw���ێ�%��õyp%��y?}��S�G�Ĉ��<nR.vͩ!�H�|�u�[Wm����R����%]�{cn��߅Ll���<2���0V6k\�~�o�2|B��)M3�_�����3}�Y�7���}�Λ��CM�v�{�80�9���v����'t�?"�t8,�U�eq�/{U�1v4W���5�;>������R��~xjq��jX0w�tD�$�Z���KRN�J�x �>��	���v�tA9؊�jU�\\��!))h'�fҶX��do�x���ԣ�q��=�9��%M��5���a ����t����d�C�H��s�����]����\�[�+~�b�b\�����n?A�����=A܈�tK��u�_s>����#H���	�$�`Ļ7+�exlp*�_���_��{P�`K��A��j6{�P{w�dy��%�/�7��a{����9 ��>��Y<��F��wϿ�����E��u���H�ߨ�q$���{�[�M��հ����o��'���޽$(Ƌx� %��	�	�=T��#�Y*�a:��E�z�p��wZr9k���p�4V&�#	�޶Xņ-��$�݈W�ʓ|}W�M�Y,"��0��\��>�gpct��7Db�6��]|@$�Gxl�+��3
|Z�j���b]��K���+k�ϯ�Qrnf��Z�<����+^�Yӄ�$���m��u;[b���4�d6(�K�X�JC�\�S�),��tk�:'�|�U�@���p�%�KiЍ�iA`�gF��~!��wL,N�H���#�_�$�{�AK���L��Jc����f{$i2U����˲���H=�dhj� nBF�qqmӍ0�T��.��왒O���BZ�Q�a �x�kM�ŵ�Qyc����gJn�+4��~��g�%O�{�oT#�D'� aM���W+��T��t��" M}�p�'+S�=��!s�����&�`J�f[�W��E���C�梈}����^�b�`���*r�'�"� ���D��o���3���ߨ#̤<#b�AZ,�.�1����+����d��WE��7���w����j��^�E�Sj�>��A�ꄠ�<�%�� ��e>el�V�/��T9z�\�S���x�g`/�	����w�������Җi��$��� IU��z��s�)F `p�Q�L7ɱ��L���Lf�G���ōj���b����1�q�����p$�3�:�0O��#FQ6����j�Ye%0ۈgD�;sS�k�.ģ���j^���+����p|�@�K�nZ�r]F�غ+�L�l{D���>g�D�����P��6ea�"ǲ@L��V�(�����t��.�p�7BkL��ܑ3{�8�g3U4�J�/�n�R�CA�;���9-s�Xc�$�6OL�ܤ+$/�A!�eZ�7�Ao������OE:���3l�'|[������DhA[�K��]W˿���{~��&`@W�/ �M��`Ϫ�#(����T�2�U����y��r��NN_�r��;d�*��Ĥ�B�|,����I�D����r�0��S�����ѩR�����'���/f�eb*��"�S�}��0��9�i�s��1���ԗeǺ	U�A�Nv+�;����plX�T��B�	�%�P��P�q�YSA��y�?�)��]4�n��"O8������^�Z��:�@��<�Q�B
;;�E++�~���@O��4���\�oW��?@M�cE�F��<�p8�Cց�z���?A�Tp�MBNAj�Q�!��K�Z4��·J�͏<	�%�,G�h�#ҏ�x>�c)�fu����`�����&:��������u�`(��w���@����7���k��a��d��ѣ\�@���Q���4�n8�.�ߞ-\� �T�1�-h��z��^Vo��8Rb����Z�+R%Q�C[Z�ru�[�&
�F7�ҞM�z�,���<��ֆ̕r^s�\�6�W&JG�xU((B�|y8�f����>�׃TnExX��X�}�a��ep�4��{6��^-���
�ρ(L�<�&�s�`U�Z��d�%��
+�$+}�Z��o�F�|� T�.�QI��^f@���⯈|���$uT�e	�.@:;�d��>���Ug��YV���VD���F"�O���[!$���ܵ�?N;�C��B�mQ%��L/Y*6�X�&TrvOn�-�
����
:��*��d��q4�Xw�R'��~J�8����[���k��~.�׏ѱ6fM�Җ�J�H�\1IOz�]�_�O�z�jALLŇ#���1|��г�I�ſӘ������)p��|�V��{��=�(EY��`ui,�N��c ���"+�bd�xf@�l�����Ⱥ��Y�ؾvr���$�-M1f?�Ϫ��5gQ�ʩ��?�b��A��!�\��Í��/oR}Z��/��n��c�<V��'��M���56�� C�/���!$H��>v�F�sXtujN�۶���_/��"m2켘���3��
l���P8���j�#ջ� "N�r�~�����}�wq���mhm�����s&�y[dB�q�k&m'E���Y9�87�-0y�ː$/R�����aÉ9q󨣒r�-*k����"���
�g\��偈MQ��˺谱��F�ܾ����!���7�?s����Y�~�G�9�(<�]e$g%,`�N��?X£�<� �/;]����`\+֓�׾-[ȈVځPz2��V�Wa������~_D�>�����.��rR�Ìicϛ��N MHӝ�0�Mm/ې~5M']��i(��9��!$o>��'x��N��6���z�z�.����B �}����6��HU�
tpI"�O�x��7��Θq\b�XY+�y'�{���.����~V��B�/8e\ ���`�&rT����"�Y����Pb������k��BHIo����6�w�����z_���c�����%nM �۰b���J %"�˔y��{�ـ�ƶ�՝k>R��7]�\��3:�ً�i��l��	��� ���{ gAԯpe��񲧎�����%Xme�(#�~m�P/�w$�ߨ�J�䰈� �O�����5P'$z��s��!���i'��u��qrwiXC��vؚ5��h�$�l�'���}V+5��x�qZ��a� �H�f�-�LM���x�bZ�̈́C��
����b܏R����*�JK
������I���;^��@	�'\1���_<���b���>[�:g�v*�j�!Ww"��i���&�����6��OJ|�~a;|�[���+(�q��TP�C�[~!��^nzS�
B����s6ʉ�f�u������`x� ��p���e.C�����bc�9vɋ�T�q��>A���1�[ K�z�a�N��U�:/��J��<�� d+v�����ֻl���f=���S8���{׳�d|�ץ�
�[���ݿ���L�Jf�1���2u�M���SϞ��6�3[.4�O�z�n
��K�
����d(���Q5�='�'4��MOFFJb9�X��U���u5� �i�ǯ�ie��q��\�'LDʷI�Α��GhC���Qbc��Ox!�z8b#ϛ�*�K�E��+�07�=q�BwI�-��兞IQ+Q�x�Qp����/�N��$쇺�,0�b`H'X��|�W�0H�'��A�{e-6g��5��4�}��Jɖ�(��;���	x�d�����_����Q�Ȼ��o�PD��V~�q�u���&b��s ��oГ/
H��-|��=����kğ'K��!:F��kB�L�r���F �ťɺ3��`<�S
ӹ0xU����o�=s^�6�٩G:�]�[� ��3o��k9y-yAb�B6��T�+������N��v�[}�;7���(���̮o?��������F]Wy�B�60�{֖� �*���]|�{]w�s���z6��Q�0�*ԑcR��W3if+�*�Q�O��
�8-s-[M�Z�+Xd8R�I��JR;�Ӡ6Z�;�g3���AA1�xK����'X||����)'�i��f�GMi�4�D[�'O���ӮN(\>�����_��XQ �_�5����˳��d����݃�Oa�b(
��?뭭���dN�m!R�:)J���������8��F�m��4��l��'����1H���
L}r?���{u�bd��ĀJ���N�Y��7��_n��knn��6nE�Ҩ&�-�v�%���^�ʗ����>���e�7%����~&q�N���~mq��i�uY,	�_)_�է����'i��sG����J�B�iO���Sf>"GM�v�`�b�`.���Q��>�zD+�`-���uc��f�A�>w??3G�1%�`�0:ж�������qp�$���/r�t�H V�r� �@�i�ߢc+;Dp�8�>��$���JQ�gƘ\�]lUP�t���)ZQ����K)rR���b��f��P�\Z�'��QC_a��x��z�k^��1,�C;A�r�.l����0�A��oe��!�%��WֻƎ����@J��/�85M�9�(;��3�jA���h$&4��R< �uX����%#�`���O<�9�*\�װ��:f��'f6ڎ��*0�|V"�������8�tTj�y�*]J�J/5g�V���֣Ͻ��p�Ђ����FĩL�>Q�(�����w�b�7ﳉ#_�>�O���-�:�p�����q�M ��K��E��G������/�v�TA��uh�h^���%a�&����l�zw?+��D��ܽΒ���4�����dw�%~BQ�Y���T�_�+'��ۄb�˕���k������ݹR�2�ዛ����E�'���9����� n�*X�L���%"K&�@3��`	m^��q��6����J|F�J�� �c�D�+̜����ޓ�k�4O�H�;8P������B�c�]��mE�uh6>U	��<�k�MuI�x���ZO��B����욋�{D0.���WP�C���}S
��(\�����\�P	L�,)k9�D3��.���]|��w���ȿ�(\�,�A�R���i�� ����S��`���#!B} I�b���8�z�b���� ��G
	.�ԅm��u�b��2�f��e6���ß��R�5�;��BCSg��A9G=��6��]��C�x�n�� `)W@�`$'�G*f\1˳��6M~��x��n���1f����z��F�]eg�YS!6�<���$�&�k����;��W����ETf�ڞ��b3ᔑd���,�K�y@0ں��<����w�B��x������Z,�d�Y�]~R���xK.-ujq�eȅ> ���W	�Tx���]� ־�#$ƒ���=u����r��|����p�(�67�vT��o�j�#��Rq�?��=&���G�<��rj��%�,�Y�`ثT�Ƣ �ZA&��G)Ws�ݰ��0�ߘ�1�^�<$J�>?��,�l1'���+ڶ-������Z�7��\��*�C�J� ��P�>k0��0��b)kJ�����2/�Li���&=�%��,7-�yp6������K�]����8�`]�] [���{X��vsV��Gn�a���0)}<�%3|E�
��
�M8E���` �F1W������q��-k�X����bj��:ڝds���.�MS�j&oȍ'ϙ_��򂇣*U�㬒���z �5�Vaքy�:qr	֖>���q92N�^mЊ3?���&�ŗ�\�Skf�S� ͭ2uQ�'����������xm#�H�	��˶崷�ҩ<�����Й��?g$x�ddA1�I�b��+;��P��zV�{�t"b\��<N�Բ�AV�~D�:y~;VǨ�z��.o�GQI�	n�a�]� �6�*<U<��,���6uod�:���0%^����B�f�?�|�m�E�,��D.k@�A�n�~�	ƶ�L:��ȫ�&M�!�u{�<�'�\3G�mQ�����ǢOc�M��[�.� X#�j0T�"��)�yU�PN�c�O8���.��M7��`��+�m
�){���u�ד�{�B<a���,2�-8��%t��
���8�nR:�+���>7&i&�:�no0�v�y؍ޠ�.��0 + ��������04��Jd�ëԦ�$���W��*�m_�<ϧu#�� 4����Y�KIB�����H�m����|�Saawxҹ���䣣�8�<�̙�3c.x��>���7�:5�S��<bT�ҟ4��YP��U��N]sz� x?�G�V���վ.a�0�yD^���+U����1���\��<���]�E��$|:�6ڈ@02�X�9gW��A*�2�{�j�%�q�Ҍ��j�����L�QbB�����Vɸ�����Bߪ�x�O5��ɘ�f�}Zw6 `}0W-��������ݤK�2&����Z���%T��P��]H> ���)�fLPaD��:��0|�%&�6�	C�IGD� nz�6�#^��C��Xn0��)�|����#�������Vſ��\.z�S���PȈ��<����-�*9����S��i�^�*gҐq�t�| �5�w�8b��L�_?��fb�"h�Yf��:`_�����Ogl��9��S����џ`_V8R|j��/��97L:����AO����&�މ���m�e�:�O@s��"Lrp �����(�9�)\��g�XSU�1��:��su�Hy��B�vK�l����#@ 7
-I%�2�xs�J��V�$Æ)5b8�|}>Ձ��E싕�3?3r �M���:\���IAQl�#s���i�}�� jZ�s��o~��D����,���rX ��9:��I���ɔ�O*�n@�.��`i���:�����������k_�7k�{�ܤCg�K܅��e!�[��������r4�H�C٬�eǙV�	K��HG^U#�K�̳�lt⒲��cI�!�8�Fp-�&����q��yn�?:�Lɀ��3+�1߱`��.9�������Hmٸ���0�ɑ=�y��=
��\�)��K�Z���h�����q>omoz5�VT '����(����@C*`LBȏV�8*D,X���Zb� Y�?'�M�����|��r�:l�-I�	�2�������m-��U))7
�+55�����B��;��� �7�:���q�D�6'�Ub�w_b�N2kJ�H�uғb&��|�1��G6  �K�R,y�\2ʢ����otx��F��M��l��Y�[e_`�Ai�f�^���{������P΃3���(?h{���ҹ�V`��ʵPEc�b�WK�.Vt���Ȧ���@�+��H��!A*C�'X�M�
	kç�5�l骕��(݆LyU��c�k2�X_�fy��<���No���^��R���U�������e|<�3�����T;��9B��+|���o��C��p������,��S�<� �،��y��Ϝo�xк�,���N�,��7[l���]_���� �5�ưsv��r�Q�>XoF��c��|Q�+EE���1IO}m\����ٺ�b���Ij�^t�Pd�&ɪ�o�.������宾�������6��c?˙���!-� z�%��6/�C��vH�-l�Z��5≯���Ec�V�\�xy��.���|r���Q�a�'�`�R+�ǁ&;1z��A�m��<�i�*�Ǐ7۩6��(
��푸R'M�Oh���f�K��g�2�����L�X�a�QX�Ccx��*�6��'*��rڝ��d��ʑJ�+N-�N�PI.T�0f�ZH�ߘ����44/e9u-�%K�'����ogzV��s�j�S���.v�	���˾Z	��P����zcz%M����Έ^�K?'P��=KU�,�FB�&=�L?�3.�2E��+(Z{]�z2hu��9Vخ)�����p7B`��&��t�!te*_Y�d�h ����@ݼq-S�v�QC��jx��v�M!����
�=t�ԯ�;�:��Eq��Uҧ��~(��j�׌k��r/j��厛�0$@}:��t�)_���^c���nE]pW�g�t��$�'������#��4s�v���ѣ+��ΰ���g�Ϛ�է��� �º���HLA��]�E�l��u3ga�ky���E�R# �ʑ�xt��#��XvOUF)P��VF��1��p�����j&��=��(�i<u-�B"o����nl������|'�VB��6��,
"(E���_ݥ�Q�O�E^e���*-�
� G��������>�5!�d_|,�v��ѵb�j���|Ņ��KL��3�,�Լ�+�����y���PP���I�J׳�n��8�VƎ`c���؇`����Xj����:�X)�褴P]ߤ]Ǚk�p������\/���s&i��
��k��};��&g_[Vw�Ib|��&��[-)�������X^\zz>a�P  |#p�'�U8Ϣxg0YQ���S/]�� �5,bJ�c���3/�̵Tr��遍2�G�����5N;���،�-��:�#�G�C��k�����RC��a�vB�k���`�[�Wע<O��K���G^�)��5���	�Z�����n��m5/C���e̉aI�F��ì"5�n�vɡ��M�#��M��\�=�yq�W�����1����6Q��0�"�[��{h���C�u�i���C귞��|�feg�~|}����P�3���j!M�
`)�͏1��{�����,T�f�gA�?�^>&�ۅq\����;Ռ��H>����ǤT�[��A��C�5��/߇,[�4�;��!y�ƸεT��z�
�����Sߜ��A(�0����5�,��$i���mM����X�<�F���]u��̉���ܵ�[ny����#s��B�8��w {�T�Z�$'��d�.�*z�U��6}���)��& �t��G�:�gCG&��Dӻ�����X�?��77ϕ�p���V�Dp�,�
t�`jՒ�g�vT���zVN�z�������$��\���N��i�ᲦQ�X?Z��E�)=��ś��ΎT_�PTg���e�I�-� �jY�Hޡ�@��:4��ba?����V<@HM����i�Q�L�B�s��Gk�X�/D%� Y{��8����\m�c��M��Q􂭹l��=�>X�'�[q�V^C�V�eʄ���}�s,uϤ��k��J �z��=��%��>m��q��l�d�R����^]þ��H�����UI�ˉ�������E�4_�Z�gF�p&?a�U�^�9}��ܪTڅ�H�ϻA�s�rۙcK.����J�P(�S>ʨ����y�������|��t���@9pi��{ R�'�Ł{��۳�����p�V�1�ft�Ul�����z��3��+Tl����r�Bեr"���ެ;%H9������|1����k����$f���f$�m���!�zn��2H�,^�g{�aD�+�@��ٛ�V�������5�`5�H9:�'�?\�����q?AC(_@XE�X�K!B��f����{���X���v�efc�xp#�t%�U�����	
a��9�"�Bƃ�	'Cg�JoRz�B� s�n�߮%q%3PD�yh���k��/G�[=/w8A*|��D} �r��b�l!W�s'������0�+`8�=�~���#�wJW�=�.��'�^I���^)v���(x�.�&f���_��{�.!j�����/�R�D�����|��
�+y�����`��v�@�iz�u�j��Cx���r� ��L%��0]x�����1uS1x��&����@�%5�
�� 4��}�ޣhﳯ�}1[��$�湝7���Q+��1[~�*����¸ć�S�'�P�
U�V��t�Go��o�@�=���sk[�/؊E�u��hb�Րz'Q�2~ޏ�1iO��1^�!R��.�4t$B�q��0�cڄ����q�1�!�ƥEhi�h�.�|7)]9nJ"J�|�|����I}z@��Or��4�]�����%�S4���
gC�Qp���i����c���sOI���m��
Y��4����"w�SdFN�>	�d�ͯmK{Mn[�T���������x� ң��m�ۘ�����"΋b�qX-:� ���~����驚�hA���!L��=,�&�Xa�Mk���a
�ơ�ۓ��L��>6+�Z��F�i8���pБLFd!�>@�6k�}��G$���Q4��~lʊ7hHI��1�c�$�*4�<\�E3,��������J��܅_��ߕ�q\h DX{�|�|�n����۳�Ax�^��C���>�P*yDA ��4��s�!76H<�����H�̔��.A���Y��,<���on�0w}�B�ś�k^)�"��T�Գh�x��.7?��bz����ؾ{�X��t�{�)(��=�}@��FyX��B &�R:
��8W���fcGz�jSޘf��G?��ki���{ޗ�/���1A�#욼OgAՆYSQ��	�^	�IMϖ_W�3ޅ-�@�6#����0��e)�/�I���F�ߑ���C?L��R��D��ܐ���4I����м�{�B���3B\xb<���$�B�ۚ�yo�K뀼���|�|�U0�_��V�Cgm��Ų��Tj0wKX�������6��Oݷ'8�}�~GB%�	R�o���\s�I�:��2���[x^uF��d{1����޹���o��*t�4�oM���v�w�����Ն�w���b,g�)��n���i3��?�����D��{OC�`�fÇ�ɻ���Z�c��5=�q�������|���kj�52���^/)�m$z6��/� ��B)����ϙ�X�w^�_� �i#���z�*Wy�3�W����&hC��AH��?� esl�y�׏cC��	+���������5k���F����w=�Ä�Hί�?��i&.��h�'�1Qa���@v1���ڱu<m��&�z��sgD�q��9��v���B�d�nXT�sȵAV��3v�ft�J~Őh�[�iW+;�X� =p���dB����C~����ə�T���l�s�RU�	��e)��+^f%��DY����5U5L�§��Ybs(*�+/,N���R�ި�'5�m�������8m^陯M�'���!t��Y�7Փ�L&��\�&�>���ڮ(I�,�SO�D�{�H�1��9l�be��>��N�Hׁ�,�h��C��s&h�U&��%�!��NT��@d�Y�iL{��o�u%�P5>�4�Ҿ��vOZ@�й�c�*:�K��@*#1JT�4�k$p�SI�B�0���?��L4��z���m�e_�4J����ǐ�1f�,�.��4g�ђ%��1��,Z������2u�JL�KN�N[~���a0 ��B	������f~�>Σ��WJ��Ui̵���*)W91bc��$��-�8�������-�ղB�n����Z�{��`�_���e����<��U<$��K;��ƫ�>��w�|aǿ��Qؒ�Q���A�Sg_�Q.� �Rv1���S�^�Xk�^�RD�^�:��������K_S'���>��$�وG�R�6�K*"1ZW�~��ʓE�rk�K<z�jK��ȡAO?ˤ�S�h����0�M��,�:L�O�5M����KT�<��%����1R\�9&x^b`S!��0�������Of����͂�>ΐ��B�B��j7���'o�2s�sl���}��������G�3,�E���Vɩ���GC1��!*+��6�O�EG���1�K�ˆ���������z�|���_�ٕ�X]��P B3���h��i�B:�U����ݸ$ m��H�7��~F��K�`9�x6�T�|��]�1ʃ�`�P�����Ot�
��71=�eR���0�J/�DO�s�2�Z
U���[6k����/q��Q�E����;a�4����L�:����1��C�@��Ĉ��/1ycBW)�NRV�qݝ�e���*�~��#�k�y�f��fξ�5��z��S�g�9n|K���]G���>g��#J"6�E���Aؿ�2R|�˰�C:�D�?�Yc�Pޅ
)J3�*��1�=�0��޶֟��/�$���d���-�K����W�M��{W��
��y:[=	0��I�(�.Y�Hx܆��QIu�P�T�!}�@�Hu�NXYAwJ͒o��c���,]�"?pS}Y�N ����\���o3��}��9�߽i%j�Nz��f=�f�~nT�����7م��-�X&>\3��*S�a�7Ԝ_ ��XL�܏���<�|5�qz�T��uB���;�����5jB��0�P�={��e���l�,��X:b/����5G��_Ue$J�[�!;?'�XM����Bb5���r�6�b.�y2��7��d�"	�E:V�fs"�h�+u��a��D�ҁ�
Չ0zq"�[5�3�o�19�dÌlo�4�g�~�{��*z��X=��]s@�@�T�e�}J�W�"E�����D9��)�T2�!k��것j��9wm>jcp4�����%����U��yyFw��qgd�%�Z�2	��u�ÛߵeG��d*Q�A��]lGIy������2^��W��Z{+�z�6����α��x�Ə\��mE�4�n��
���m�Ef�Foza\iX'��g��I4t���{Hn��@�.�h)�wl�<�]˸~�w�Q�zh7�#Hi4Y\�O�=��%y01-��X��f]φyT�񲊈��˵]�wF&�$^6*�ț�rMx?Oz�L�LL��HE(	pr4�f0ހ������E4+��Y�:`�Sn��Ӌx��!�|�7�Ul |�b�#=H4�ధ�D�*�7�#/�B�����$���ۥʉ���0��vB*M9)���֎��Z���ؿ�HCE�nq0����z��b ��Y)�M�b���3�j�|W�CQoOW��:�W�����o��֓��"�Q]̔\z����ӡ�А�Z4R�نE��uS �ﶤF?���n��s���k��>�~9����.����@�r-��t!>v�t�!����M�������"���@`��%���iX���*W���x�1kk_���ܔN'>���u�Sv�1zT#k�ys��-���b�#���d��q���U����ԙ��[�r\Gq,��^��<�g�O����%G��'�
B�Z�:߇^`u� ���m%8��������-;�k# _6��82��R� {�6dJv���D6��MJ���\��Qf�Nj�4?Y�Cb;�"*�[��#C������T�N��VW?3th�eK�Y��,�1�$a��t�8�:м�3
�sD`Ø��ñ�?�K\#�A�J7"VH���o9��� �k+G���4�`���6p�\��v.$lF��om����Q�^�i��"��ï.y��������f�����m��H�]Lh��F�ۜ�6�i�N���mA�ݾh�h��0���h1ͩΒ��yW�&���-��m���{XB
�qlz�B��&��`�Å��nBX�7�	���U�aS�2�}�K��jz�"%��������@4me���n��2~X�e(;������C/q�������/��j��Do�"�}F�%&{ ۖ�H�哸3Vim�?�{�2r�V�kno���}՜�l.;-�͉�PF	����?@��j����O%�O��Q�N����C��:5�J�1�������[ΰ¾~�4�ET=�A��-��ǳ��AX�A��MI���q]6WEF���H�(�W`Vv�eΚ�]ţ�p`wP� P��wT��MC|U@b�{�gs����R�\!��X����*em�0ro�~�, �=d+y��-&NVKQ����:�?,�%�ga#�Q6l�3�y86�75%���N�����Sw5����WW2ڶ	o��ϼ���J�K昻Ի����;��2v��*����7`R�z�L_��v�k]��;ĕ��C벙&O���a[��~����(��@��˰`�g�*:���p���}�� O˫A��'B���p�	�����&V�����:�l���8=��(qh�,y�k0l8�c�d@���/{��g����W���"*8���K�_��YW�/=�bu�Ɯp#�3A�g��<�Վ����qi{�Ąg�g�s�x̗l���)�M��m�y&Y����3ѤXX%��f<D�!Đ��:&���~� `���T��`�HӐ�F��)���dTu�o�9��rSHa�Q*�B&Cv�z�9��
��d�}3�$���FX*��D�&!����'�����[�(r���CY��p�2UuU�Φ�@!1]�d5��!Ħ��mog�P(�:ɕ)��n�1O=h�b����zZ�<����$$�d���m�Qm��q�~ɶ��cJ��A���&1Y�j���ΆK<�����[g>��v>d�O��(�����>]�ÅF�x�p�_#��k�g���A��_� r=Z���g��l��9������̪:�(��(�� �OC��E ����R.G\_����t�rW0Չ9Ĉ̳�b�L��.��]�=��xN(\�3�zDl���[�tT/��1|�8����?�����sd�'���4A }ԛ
V�P223�C���_�q��Ƶ�ه����8A|q2��0@�'ug�`�=��dV��R��%�j�=|�K!g.�I�\��G�i@�-�:��T��K���r� ��o,<��s�L�4F�x������?�*ay�!n5E���� ��XX�C�
����������a�as�����U-p�f+y���o0�g��;W�G�E�J�P[�
��!t�����g;* p`m���/�P6�2
]���/QH1F�{�t,�n��Ѣ|��My���$/�8k4®��ǀ`��U3ԛHtwZZ�
���I2	��{U~�Q#�Z����ƽ�y���� T�ʩ]��)n�=y0�RES"ݬ��Wt�H��@��<O���zΓ�<`���P
pr��SF�(C��dݞRs�LjZ
ˌ串<�M�@�f��"��o�v�b
���0���R��u��{�l���X�,C�fiP�c���_�G�B�% � ��jeLT�Q����"���'vy
�Y̏]������P��a���鐻�6�ʩP��c�C��g��"TS+�TH!�ܾ�y�hEdc� �^�N(�N��N)��i�.��[�;Kc��VvV�kB����u�*�mf,��꣡�/B��bԴ�!�}Y�gy�S�Gӊ��c�f��U��(
IXF��m����y�~�b��9�x+ǵ��B&�	�?P}�\�fЂ�eq��Bo#)�vAg7�Zk��z�Q����#y֩��%��7�q��׾�T\�)9�2򿢽E���.�>�|l�/M3otRTP��x��p�8�T}!�w7u`t�����[=ϓ}�����>�^�"ʫ��<��+O���{��qQcC���Z�;v��j�4�K��8�좌�'J@�j��\��5�;�	�������c6-��2��|�^���h���Kvr���Z��ġ���MOc`>4*�z�<�Ds�ͺ�@-MJ��:d�\ր/;��#_���� �t�Kh@���W[�m���d�&��gYO@�U��������3�|�s��0��u�F���I���$�Á�p�X_� {�K;�ΟZ�L�70j�(H���t���ƴ�ɘQ}W�:����5���+b.@L���(MWQ�]�m��L����,��a�@�Y&R�mrA�wC�Ah�����X���!ݝ�Fcc�1BJ���R� I�rj+�������������6g(Q���A��d�mJoٳ��{O�:.(�:(�b\��X�[3�ۚ^�n�V0��x7��v�K�b�I�E��S=;]t�����0������vB:T��U1Iߧu�%��g@h]���c؁S���N��c��/p�ֱV��ns'M�l�T׭,>LA�h�h_�zi�>>��uگ�B˶��`��V� \�~^���9��4��O~q'���9xd(��+�d����[k��ML��.
�\�$�Gt˦Y�Lg���Xy��dbٚ��޸��$թ���&T��<���z� �"����}&���#�-(�AG���s`��{�K=��O`Y"qa�	W��ݜKZ���E��0�Y���UB���4��1���B���2��(U踡?��W�t��N��-#�f� )a�]8��c�m8a�ϣ�����M�3#/��%LЧ+f��?�NR�_�wl>4c.��u���'ѝ�X�CC_3��I�"p�%�ޥ��}��]i^�:��~k=6-���E[F�e�����uXuVFe�^˘h�a�_�
Wڙ�R��������7�t��Ap����x#�N�߿�/� ��6����6��	���)�b6�\>n��t��f��Z��fIs[���#&��6����l�9�`���I����B�Y�4ϵ��[�� b��9�fm4����3�S����~|z�x{��\H��:�w�JP����Pj�]<<�"�0Ꮲ�]�ؼ,�K����+�;=iZ��| #%�٢�����c���O���M��A�1�X�ֆ�`h�H�N�ř�����!'���6���yZ�
nQ�	�j�tCMl�p繜L�X�ij3�/��^,��Z�J��2����Qx �r���1첈�*�Ӡ{��ލ`���d�˜͠��U.�E�ۋ!y|%N����QA��3 )[�lR7����>:�A��D���p4ƉzT�C�T��Mxdڅ�r��.�8F�$Vµx�	�:İ\Y��|�n�%o���ޖ���w�@m���-��}���,M�9����0�J}���D��,�8�����e�d����#�������_�ǰ�83#2��AN^=q�u!��$a�^rC��鑦]#�dy�N�!�~� J9 O��E}��n��@��j8�_�'�����v��H��Hl���K�� ?q�ɴ�t ob/��"�gu)S�>ֺ�>�hq��"��`��{q������o[]����̨��vYb���3�M��x� ��[q^�4r[�T��C��GG��}�ְ����� ���-S*�m��4Zs���/z��7�
�υȜ�-ӄ@\�&���O�F���C򨞻�*�����-�*gk*�
�mO"�s�Jt�l����v8X�0.Fg�@Ր�x�f�9�C��۹����<�I�f{ߒ_��8l/8 |��� ��?vп�F���v�ظ,gÂǾ�=�L�̯k�b�]0����-m�=.~i6�H^�
fa�ϻ�a�#b���Q���A������ߪDu�,5^�t{ġ��M�t�?� 
|��
~��n >�ۃ�W�,L�Rq�Q��nT�8dX)-c���T����{��k�^��z͘td���Ѕ��G5?-�%���m6`қi���'��!��E�v�爐�	9�X���ϴ�	K�U� ���ؙP�"��W��gA��)3��A@�#B�WX�3�H0(�'�(%R��}G�����ɾ�'�Hkn[f�8��5�'��0MT�P��l5��K��3������'ۚ�,��5B;@�S���""�MR�%�yt�]��\�՗��2߬Ė�*++Q%�:�8��4��fq^ē�M@������*P�ۨ���M��/G�=�J�f��tz��Q�C�6.�<.t(�G�Zb��J�X;�%*����O�9�ר���U�%�G�gn���d�� �n�_�O��N��A�`�I����qX~q-.�W�V������ڒB];!,�]�lH�1;hcp��t����W.�ٯ��� �������R��/��ڇlJ-@��Y)�̊��:Me]��G}�	#�C#Xﻒ  *��d�g��6u��T�+'n�,�5kJ4 P1�����q�9Ǉ<z��p{�!LCeZJ�O�D�K�˟3��1\"���lϞajv���?K�=H�����R��GĈ;=گ�i�f/�J�?.,��Mb<�F��c	����ӣ�KJ�p��)*�9l/��ΫUҎ�ЈId�#�}s��~.84�~iڰ:Kf������^ЄR���������P�!���7�O8@�f
C6REE�+�)��;=.��{�)n̜���Fck$l����Oq�9aTL�%���+l$�����O꧘�52�G���#���D^��+"�tJ��~�w�{U-|8r!^><��O��[d���9 о(7��I@��2�ߎ�\�!E�<21�3affQ{�7v��웾jC6���8����
�������N.�Y��{=����{�O6�7��~���}ߑ����_����;(�e\�ɯ,.<�x�=j/���c�i��y\��n����/�zKd*� ���BWC�Վ�Vp��|��^�_0�v$�n�t��||W ��z��zN��e��:Vox:D�jA�y̝�!y���Q�iI��'q��=C֌�K!{�\�/������,斠���{Z�V`Ւʖ�i��n��Ax	t��J�Z[�}��^Peo�!�N�w�n�T_TrԽA�tm�nSgpp�|����9~��|���\s����6`���k��o�쒙Ҫ��S?�g�`�!�-��;1h���@��X�1	s�VS�]� w��d��?���@�ʱ�H@p��s���F�|Z�9A�q��-_��E}���p���).��[�� ����+}�k*��:4v��y�0�՛K�]Fs����J��6
q���A#ٵ�1��G�Q��v�4R�g{__ل�Iv^&5�z�l>�B�X��'�O�*u��L��C���:��o��c�#��
��u���s��|�xp'�7b�0keJ��~�����&l��Q���T`h���'�(g�!J��^r��d�܋�X�k�Y��A�H�V�AI�Sw�	&�{�DGd��W �Xn��_�T�oIf�H�\M_5N��$� �=)War�Ec'�
��'�p(SY`p7qNeA��`��Gu�G�[����ƺ�^�r����������k�n�q,��3��z\�7\�^K�����aR�����?1��B���^gi�����G��x����O`.���4X��Y+y��|����`��5ت��K;D������20�ފ���M]`�P���q��U��~��J�����R��7��9�������A�(��ag@�0�r�Fȃ�
ؠ����}��zNQ�P��<����h�-� Ï��G��PA3�8�n�䈻���4Aj�FB�9��N��_2������z%(3�x��>o�2�'��	]�	������^?F�cX�z�o��-E [0���EX��a+�� ��G4��X�O�J��ǰ,�Y�Fx�N9�a���4��w�G �0�Iu3�pz�E�������A�UBq����tmg�!��~��;b�I����5�}��)�|!�G�UH>�w���Q�l ������N!u\����ۧa���Ϗ�3�M��&��lH���)rs�#}��Z�	�Q�}8U��޽V�P�/�����H	jBp��B�1s�ɰ�e���S�\H��Ǆ�C����(",�!YX��}��J=x���䟆��@k��:$�)�1�Œ;E���a��$9*�e�x��p�E��G������v�v��ЬU�Î�n��V����n��W^) �tĠHM�NP�w7��� �&z��l�f�҃��U��,��xp���q���JЇO	�_�jk�x/ҏ���U �!�t^�hY�"����×�;x\���JKw���g�� �ͻ7 ��H�l}/�E�\��R�C�;�\�/���7�_u�ZN�}O����v���o��c���pW/�z9�<�e���#FR���<,� �}!F�5E�F� 'gدR"���A�!�\v��z��A�/5�:�����q.���h�*�Y6��s���1�o��h���}�U� W����0�������=([3�Z'�k�U+�����`��.�{a�L<m�~P��ʀ9�؄���I!z�X`�����*Qu���f�MM� �f,���
�^o��u�;�~��'F.{\\�P�@�'�o�M�c��Yc��v��~eXE�=��'5<�t���SY��˕�����,��l��b�ʦ8��
��+xGb��Q����*G������:u΂���t����^������%������I�Ŵ�٣��Ƃ}Iy	c���-�갶j�������]ȧ-V��[���g~kh��|��t��8���]�')�h��c�v�n%�+M��@�<|�(�����#�WR]�)F1A{eDpD�b�������I�jy�7��D~�y��['�KB�[��2�$R;m�A� _����h�z��B��z��;����%w�I�P�8�$���6̈́۔BW$�b���{~��O.Ԏ0�ھ�t6j'�n
���2*�����i ,�<�x!
5Y��c%�ay��J��VE��Ė��ha��TQ��)�M-�4'G��fu<#@�Ni4H/��l���l^�Q(�t�Vr̵
S팺���2��i��R�`��#����� 
q㯯�o�TsmhJ����n�Q|��R�dQ��[X������ǆ 
�B���!*h�/'j`�0˼'��G��cL����m�ȱX.c�S���CR�zu3�V��6즷E�d�tY8c1 N:z���+��_�@p>h#�����h5S����O���#�F06�#����Iu���6�|���Q�g��/5��_P���!/�{T���V����+�{�Ͼ�FNr��\@:����*�����:p��^��V�W+	I�ĆDi����5Pm0	��z����!���,�󱤊+������i�ƹ�WC��CZ�)�s�t�|L�D�v�5��].?*�f	���ő0�ƶ��WB)��<�
��xk)L��0�'	��o��%u��O�p��cP0��MY�Y^E���{�9$�0@-��1oٳ��7�r�'���� s��8�%��w =uVe����>�'��Զ����w�0y:!�&B����ԮZD�K�8��˹��;⹇�n.HT*xX�^��<N��i�ɵ�򺅂�{nL��S"߇�w,�EIׄ�\�Ø0m<�n�ͩ���8U�HV���R�v.:'u��m�lY5Wz����]moK{XT��\�$?k��L�I�#�K�{��3Fl���G�.g��|�u�by$�:is�4����6�͜I�0ZB�8xFgh2�1B���J����ډO,{��{�C��\��I�o%W��Z������fA�L܌K���Qb09Oc|���{�YV];�����]�;��q�Nؗ��R��2p=F@wKu�K��6����*�~e��3cX�Ϗ4B�;u��۩��d@W����;�dJ���oe[�4XgT$_�^N"��e��a�ɫR6���h�"�}X�f�Ze�Ůʲ6߄}5�XX@�p�
��e0Z��^à���d��2�t{,Yb�0�A��a�Q7�@p����M1�4U������1�"�J_`�y����1����a;�|*��Gl�c�&�G���ώc; ,xFrW�����μp���^��$8��k3+eCE4[� %�Cˣ�Kt�O�5/|����чY֠�Dhd3ʰ��yɕ=p5���14D\u}���!��]\���=�Ĳ":jCv�4�<v��%ۤ�&���S'[fs @	 6�(�o�&s�S2}��N+������\�Mm�z3
�q��o��?P�#���Z.��F(�Lqc[�,h
�̒@ǫh>�p��<i�=~V?�C�`�[I��:kc�-L�CN�#k��v�sG��g��N��M��d�'����jy�D}��l�o�\�8CL X^��"n;?X��K�! �Zc{�t�uL&o�~`�vӯ%V1~�B��u y�|�^ucQ'~��_r��V��m)-�����%{za4y~З�v��t}�!�e�cID!Ԫ:BG���d虍��]�����
���D�i�鬀��yۘƝ�2�CZ���3��9�?PŜ�3�Q�x��\��Ľ��!��:�QIE�Ue����{#��?��gP���� >��؄6����)�����~L�y��j-`W���TR3���2��)J~���0U�k�0e�_��u�ۣ�M*͕������y��SH�Y$b��- 
��,��S@dV$
��L0f����e������MJ��{��ʐ���� _Cz1����p��L:Wɝ%�æ��c������>�^���]?a�]='T�%��ke�T�f(Χ�24�d��¿�K��� ��-����r�}
��l����`x�ΐ��c�`� w�M-���1ĭڍ��zn��!ұ�۠���Ͱ+L
n��f��LE�T�D�9���<4��և)l#���� 6:�z�۶Ԏ[���NSLK������GB�t��V�x6�u�ȇ�J�ȌK�W�W*O�Q[�+�]�I,O�d/���k�&1$�{����	���ȓG���qB�h�Y4�	���̨3��MSO����>�8�v9H���פ�q�i��]<��kg�
ˎd�nz����f����:���R��}��؆#:`����D����i�o`z��"�������ι
�]4mMt	Uc��}�Y0^�ڧ�zp瀮Ws3Rտ5�ƭm�s�Ԝ�4��3A�jo� ���֚}
+���� �tk%�O�yd���X�b8f��@R�zf �+�ۊ;=�7�b0��Yct����ce��?9��e��Q��VVV��i&i�WZ�-n�ȽX`��%�[��!���rl�+�q��9�����cٳ�E_�s�ؚ�sKk�����ߵ�b��/C"JC\yV(���D�y�%�m 8�Z�E:/��]�|E��,
��}�����lG�c���t|кcGQ:z�0~�PLM~Ip,8Z(m#�iZ����A�;� n�AvZ�t� ȭ�-�4�x���*�V��g�����K��s���U8`�K*'��g��fSrR]?.���ͥ}2�0��Ɍv��� ��9n�#ڦ�r$��-��N�Gk�Ɯ���2C��O^�@���&8�-	���\ ML]�AW�������nΣ>���m�&�����0����(~���JWW����z����>�(�s"Ł��`$fՓ���9<[Z���k�8k�K�E�62FNV��J׹��ZN�J�l޼����,>�, rɹ{N�@�ċ^Hy��Lòj�Տ�ճ�����J}�E����ԃ.�ʐ���JN8^�[�'NC��M�&X�*Q�}B
�v0��c��]&���g�?�[�V�W���av/G��6�MmyR`~��8FƺA�lƤ�I*߈�l��4��X���S���?�y�C3���:mb%���9`\��Cn~M����C�2����4,�r�(��X����$�?����:[�"勛�D��+��e�У������z��z�6 "kY�F���⡇��;��3Iu��S��^
������D@-����iF6�g��B��r���O]��cT�XF��n���@�(S��H�_�M}��ǨH��?����n�� jO����j2@i<�sno�k<��K[׃x5��6fz���V�-��2���+윮��
n|�g[�
�ϡ�-A�sv�MU78�pv�q+��(�.+N������Z�)E_�
��a2�f]����*���˚()�^P%`ζ�����O��Q���W�奰�\�O��(�#�0{�@�c�8}���Q���f��Iu,uǖPO3ŵW����R�g�kl�X�Zb��p�P'9���iO,��&Ɇ�H�Ԉm��rtd��	_��E��`��q�>p2dz���x���a��/+��KuS7��q�ahE�i�c����,�u�:|�&5��4Q~{ >��k�O�w�nQ�2,_*��G���A�Ո��I�ju��b]�o;��L�L[��A�e��t���k�7�a!صىv	'w�cA�[��D�� �z������Y�ݽ0����{�������hD~	#L���*f��քF��=�.?�� )QR+g��G1r�(5�t�J��=�r/�P��f.��c�X��gD̦Z����	�G��˙?Z\i��h6<A�R�]�Hc|�
��p��s�s�/�W�Y�I\m7hv)�#�<68�*��K���Y)&��>�J���-jc���e����/Q �8:_6�w�Iʸ��E�r]6���SܭUu�j#�`���0�-��>[A3�b�^%6����^x�n�\���Irn/����^��:hVt㉴�k�z�.��H�X�p��u��a�U c����0y�:����*����>P�~�	%	>�b�[��#Ji�^�}�K��ЈT�a�[?�s�ȱ���	;t���f�!�P������+G�4��c
K�%�A�Wds�1	��ָ�X9pud�VZ����7*s�{)�O8/x����P��ċ��A�.֋GA��H#��n*������
���6�Ƨ�	�i�n��mVGע�3��)�����ʚy��F�E��py>z�}�PS��{�T��uOM �+w^f�1��m���l��<7^���_ԭe���J���k�j��/�qb�
��
�O���u=j�|5vVoY@��y@Y^��ж���d��9rl��=e~��M��[c�������^蛷G���ܛH��/ ��L>ivܧ���n��\�>���C@l:���I_�`Ы���l��Z�S2��lR�3:(��LP��;]ϡg�6`�p>߰�yܯu���_NP �nr#�sF|=��l�@	������u��F���F��ȃjSlp���'#ߎ���$j���s<[��8@�<n��;�)��
���i��1�Id,?i+Qa(�GQ���>s��qX]@%�%�������t,��x܁�U{u��t�"t~uNocJb����Y67�R�:ܦk�O�2���>r�)l�Hd��AB֥���/ݿ7�Y��f�ðy�up'@&a,��9�q�&GA�ab��0��n���xpF0����R�Tl�H]x�7�?�܁#�G��>8� ���g�qM�/�o��19�w?��t�Ќ>3G��� v�����u����LM3���pɛ�9�g[%�;Z��S�U�N�J�S~}y� ǒbƲ���܈�������tV��rM�'��PX�K!��Ɵ�*��]�?;ڡ� ~��m��!ZK�G�`��0�3���.�19lPf#*���z�>8�1'N��٤�_��F&r�_v�Wj�Ն���A�3B|�� �*�mp�.)��5�����9Ct���$�m���ֻ��R��#<"П��Y(}]��7��Dd�s_��)vOm^�"``T0���<�<�좚��a���z�ouꤓ���.��U����M�?)�p-B�lI�#�,�U@p�5C�ttE�v�$G�*%����k&+ى��Buv�;�j�.=��|B{�=w����H*!�Z}W]nr3݅VI)��Y-�|:�ގ,yҶF�7�s��F&C�v�ʁ�pk-`Q�����O�~?a�I+
�LDא��nl��k$����F3:UȲ��A��y��0��*� �$�jteW�W݉`Ǎe޺��;�mQW�'��,1d)��<�H)*��KqA���)5�|�/N�E��*ȭ��f��~������y�����*�L8ms�����t�di���RM\�i�cJ���Vb��\@o�����+�x6 `�x �I��)�,� LU_Y�a=�#�Pj��R2f�ѐE��O-�Y)�N������)�R	
�Ǩu�+%X���o�R��8� ���������p@���~����Q�bxؿ�֘�MPc�ʏ�8�qZ��m��b�~܃؈�]=��kQ�k��gYp�����$��u��9�_ۭ�����}�B�!�����a�!2°#� ��_�)�S�5ˍ�+>H�*���ف��}��3)�f[�K��.C���/{#1���T\�A�#����5�ug�t:��_�)M��j���;^�����To�L�,Ρ��@Ր�1�����j��e�W�ۀ�E>XWP{k=�B&��ƨ�Dz.P���㮏I��
S~h�����q�u{�!`1vpRU����"\im�$L��>@�\D��d���B�PҢs���M�~_���i�ܿ��4���l��=^%S�0�Qng�b����$kk̜Cɳ$�s�K����P�Ŋ	%+ {7�+I����?���{���������e*��3��M*9�N%�߅���+��U2'����Sw\S��o)EC��7�u}�'�%��?`�>Wy:�I�3��8�_����S�\�LQ����i�P_�V���~9'.Q����t��L�3W��x����2��֫��f�J��%bߢ�jh��Tv8���v���R�x����z����D�pf[56P����ϥ�rA������ P����L��%? Y�c!c�SjY����l�Y��=J�d��ߨP�=�q�������51�"y_q��t�	��M��kޓ?8�*��	���T���U]"�p����z�G�����=tg^pZQSӉ�D���D�E�W� 2q���r�L��%C[�]��@�?R��ϡw{&��-�a�ܲn�T2*!�Y��W�m�8Y�
2#�a��P"ē��C�����Z�NGQJK^�Q�<LO���6����ڇ���o��>�VR� ��LY=q'Zy������n+��d@z�[�ݻIM����n���Xtw�Ă)qEW �-��<Ot������1�v�[�PQ3��S������x���9;e���H�lU�!�0�հ������;T�w�D<�<q�H$h����y.4�#ueō�#�\� ��9�1�ey�@�7����1(�Qn��L�h}�0��������v1�4�����5���jU�*6�Y0��/�?V,��>�!J���!��V��:��V��c���+ilw"Ӧ����	6ؐ��?I{,Cy\T�� � ��DO̮�����p�8R@;�f}Z��T����C�ŏc��U�
��tp�ȅX����Ko�i��O\�
o�����M�]��[VY��i`Ӵ[��c�����7��ɝ���.m�Nܸm/���Ze�F�H3�pɮ�2G�N�>fE�P(�I<�q���U�wYWeu�.�!;���l�5#s2��L_�u���z^o�L���㎟�lz�����e��4�:���K^4b;o��İ��~3��{]�P`��%�Q5�V1���G��CM1�✠F�/d:���+XC|�.�Y�r`�;=�g e�ܵ���n~,�Y���]�s�U]PM�u4��%��ki
�y��ޞ]�eU�`j�����W/�<�+�_��]�ϪPq���}倞�Q�y8��%��B&��b<#�.�<��M�Q�KW��+-�ng|��"4�H����m�{���f�s㯏Ex4Doˢ�E�b+�#!PO����A4r	���ֲ��� ���}�i���!���+��nf.�S��Hj��g�
�Ifڿ��)���_dsM&��뼤��
�?%�Mಜ5-��uF��!��X���lBx��,�9��z۩���f��|,�e�P�a�������lBt�X̦e�A���n���m��ѷ�?S����1[��㲄�����\��a�����|�&=]�F�����Nck�u�g1�	�HA`p@m��f<cR��t&�Ǥ�m�bL��g�<щ��}_��p���J�Lt�
6�R��Vg�goW�ڱ�%���6?Z��_h
��3N��ÁI�a-��fF:i���F:1���)c&�@m�%�x<�#��=L@Y��7�(w��d\_���F�%��Oq�@TE+��r���YЮ���G�N�F�Ȅ�bx�x�>�����X�h�b���(�HŚ�'���wE�k48\5� Ƽ�6�TA�1 ������n� Zf���?�$�L&cnx?����w��7�r2{���P�ĽgDW;�x���*bH�//���#�]H3 ��ⓈCĺ=؍�@�Gk*�%CaGv��'=c�^�_d-~��c��p"��Т|����5��)�<���|fƿ_��w��3=
�C�-��u�y�]/�ɍ���fE�F�"+��-W��E$ݯ/��f~GЩ�DM#�)����e�XEl\k��
ط��K���,%>�&��2����Og�^^��զ�ށT�榀Ð�E9I3E��1Ā΁=rx�ȃ��tW+�*|~>z��?K\,@�����������=�&eyqT�U�bLo�Ae�q����v�C�_!y��
��eq�~��v���3L����Q|��^?�e?�UL�1��n=1C���7GV�b?Ũ�7m'rvh�*��ي������� ��"���q�1#/5D#�H�}�{������AagL�\�D�����@����+ύD��X��,��x[�:��O������� h��#��� )t����֚q0tș綹�I�������>��J\�!�Ƙ_M6����ϫ����$	 �+�ӗwiWgNe�lI_������_��[�	K��EY�hV��a5c�6�M������m�
آ�Nj�N彪��gҷ�Ǳ벜�%�EF"j$�t���u���c��"��U�^�%�6PN��P�j��{h�	h�cK�.m聶; VeE�z�t���US�C���Gj�dg��k��K�2�j����=jZ����Ŗ<|��ht�.bIܵ*:�pH���'6���l�ݹ�_��G"U�&ݗ���̔�$��8���ej5 c6���4�X��{,Kd�[s%p�z4	2a�'��#%�Wk1��>ӓ��l����aa����L�/"�̶�&o���:���G�W��b5
�i� =�!�n�ԣ07���¡��} ���Qހ��(�i�T*��� V�>�6����Ap�E�>%��y|ԝ��vT�W��â�@��Hf����g�l�W��\/@F�4w2(QE/�������~y7hP��	ہW�U
��g�c�Ja��{$o+o
�;��SF.g�m=]�i���m�n�@򋨅��)U�����J�gh��˵���DW����)9R�)Rε��=P_PE����Oښ�'�vt=Z�<��y��)�[���K�r��=�Ȅ��d�b����`������ԯ���BZ����Ø@�Ӄ4�%˽m�K�^�����6�~!aa~st�tYk\�"�>�A��NMzh�4fW����|����e歗 ��~�� ;�X���v+g�iB�o��N�C���x�޳�1;����I�⤪�7b��$[������w�s��T���ݦh��d	j�@�_y��T9Խ���uE{F�9`�v2��ʃ������>EM��:t? ;�Z���bX�V��t��X��'v\�EJ���66���t�ONܾ�B[�"�׸��de��d�\�u�h��c�P�~�� �����.�JE��3<Z{�&X�q����dG�ڰG���F�ɩ����_�y:�� RX��p��wk1��-�3�?������U꥔�P-�IUܷ�R� �z7�o�|p����:����x��|�62I,�c�ak�Ɏ���\B�WN�pH�#�Ww�ݾ+���mVR���{���)rr�X���w��!��ۜ���Z��E�B�
)��n%�yWXl���∈ak)�+��˷<$==S�@ТEj7��7(���I��a��ُ�2���!HV�ͬï�ѽT�)��-H�ܡ.��0�U !"	�c ��EY@������;�1`tO���"z���^O���i��!:� ���;���#�<M{R��r�9m���-Tl�)$�����e6�����Fe���,�S��=�
��_�N������[���yAuf���e�8�K�C��)5�~���?D���[�K�I�����Yk7�)e�]���	b��`���~7�Z2�4��L#�P������?�<�ȷ'gـ����~*�HD=��I��3��SAl�[ּS{B4�����j�pL��1������r�Ka��޷p�ly�s@*��=���C V����5��U�@v��/W̅��nU��,�lס�>g�0z$��ҘNs��ܱq�V�Z]u�U�G�sZ�%.�a��{/�v?^NYD�ǢΉ}���S� >T�+���F:��!��~�����<�� Y�uńu�K��'�3��f����q`�MT����U}*
 �g�ߣQ��|�+�z�R_5s����5S��Ț�o.N�jx����+�/_�l�!n03�Z|����[����"�v�&$��f�~-�%	�ō����R�5�¥&ա_%p͐�˶�h�ߐ̊��_�ܖ1���]�e]���y�����`��!*[��<�}����<Ć����� �+̐� �@ڡ#_����6w��Ifv����u>iH�t�u����.&���բb�VV$X"�]t����������ޙ�=�i�ˎ�5骅�=��r朎ϩVW���=�LD&�2?�A@m���U8��+	�W"�#w2�2���Q�/*~����bk�B���m��>%7�5���𯕛*%vG��hz
� fR�	xօ�T�%M���K����������V%��IrK���Cu��{�0M];��L�j?��2ib鶭����C��e����	GDB^���������l�ҙen<�.䏂�!��*���]�b�J��E�0I�wO(�&Ԯ�]C�]�΁fa=������J�7\�ǧj��$���!0~ bQ��G�BK
�ΘK���(���ӛ}�� ؈�����aV���6e�:���Y�&��8�B-�/:�W����(�f�۷ط%f'[�m���cF��#��yת�Sy��y����_r���hZp�nJE�=��BA1�n�
'�/�*��+Z�껲E&/��{pǝI��|�L�a]�A%/>h��+�:;���,Y\Y�,B<̒�O rj���K�T�29����-}��h��)?����,M�s-}�*���Z� Vo��v|�|R��Z��a"Q�r����h�?��46�\.@\;���C�?�*���6g7['��2h7�$l��m�_�@�r�6�!V ���fy��?S��a9��*�J�L���6ZqU��U�X|g���O�	�I�uD��zkȺ�5Ld0y���UF�XVjGfB2��5w�~��J*.Թq�	��W�6����_)�0���X������B ��1�c �-�y�"&��g��k���_��tǹ�`tmF|�1Vc����=��K�v!�#h�Ψ�k��P�|�Kk,J�\_2�&�O�)�%����N(A/�y���Ľ:��
���J��r�4�0�5����&�܌f,5�<.�uV�[�\u�}Sw����x�������39�k��P5Aeݕ���V�2�і���ɯ��v8�9��sI��8㬨"�#]" �#TY���Nh��bQð+4������u%�rݗ3��G��jsN8��O<٪����A�2�ˠ�;A<�G�#�ʝ���j�*�B�g��\�*�xT�ˎ?�r��-�L<�˂t�ȓ),��<S���DY�)9F��d)���Z�+G��*��D��'O�8�Jnꁿc����DXN��*�1�1�\zX����j}*D�i�Q�Aqc	�B��LE#�eS/�ƁSn%��;�k��h�8���F�0���1��t?^�mV\MR{�Ņ�ѧ����ﵤ�" ���[��Z\y�Pf�WzS)+�.�A!��:�'=ﭲ�Mv�IFp%ٰ���zF9-'���,���������\)�0�N(=T�5��U��A�M�`h������w��7�: 7��rcO�^����6=XTf�+a�c`)���a�R�~L�����(W��FGe/�t�	��HM�U[)���e}W���cń�i�1�,	\2<+.`���!�~��Du�ڛH�I�K�a*��_V"Q������B)�F���g%i5&�7���SP��wl=������镁����YS���>���zx�D�1YB�E��r���ޣŠ�
���1YJvYx`�I��|]��_9�p���~ �3��NG1���I5'i՛��ya�)���yК�X�7��k�S�M4l>W��H0y��r����ᛖ���p7�D �-HJ�#J��7��P]TR;��`�L��
����Z����oc9���Ĝs�=�u�DCA"lj���Y���@�/Bn�
yJ�p`�&]����p�0'�]��}���t��ʡ9��1�!�Oێ�:�.�������?I,0	���:��(q�r���,�P^�v���<�^��U:�`�ӫ����x��0�2��조��4C{v����LJ�[X��@��2o��=�l
�~"o�bF����QzS`���gfa���߱������{'�Nd4��M}?��9��m\j���-�Q� &�^j�%h������r/���YIⓒ�~(�hƱͶ�9~9��_�o ��Fg`OO�*H�2X��=F�+D��bn����IL(�V* %<�}�ט��<x^Mx$�S��>r�;��g�(2P��$�=	d9UTA1���۹C.�Ԏ��.���a�־�Q5mTS�x�����hЙX�{�PP��Q*+[�z���:c��AK�m[�i~����ԭZ|���z��J�������Rit"��G�|1�`Y+ǍT4��[�a �:Lv��P�$�*��C7�}8΢�.�;��za�~#�Yt�~��C��*q�1�jS��7�ć��Q��7C5��Z�#bG��~��,W�{:�$�ڽ�d]2tGHB�K�Fq�΀�"�6f��F]h�xV�BP�/.L��7rh}ŋ`��Nd��J�Ey�:`���;����,�)G�Y�}�Y�f�ɡ����t��ek	�q̧: ӊ�H���/]�*�A��QV́�\,�Vmm�������e#q�s���6y�mJ��E�`B�XX0� �	4��e|,2�aVD�E�B�g�"�׬��ѿ]Iikj�I<!����,��b3'��ï�55A���{� �Lc@7L��9�o*��n�8�NрrZ)��O_������&X�P%�91�_�1Pxe�I��mk��X�&�p$68�_�T�` ��X����vה��2����W�'��asie����BT3H�x�GS�˼:V���xx�+^8S]����|l�w���,�Ƃ�*�?����GM!B��4"`C�	:%rПӝ���A��D4i{>c_	ѻ���|�q�Z[�q�F]�L��7���ؘ�3�.�GPx�6Qؓ�f`B��wH�"EG�a#T[�,~�L�����m�2��C�	}�l�V%>"j�b�u
���s^��es�O�:ʣaѣ�*l�
#op�$Jo��!;�9�>*[x=:��`-��k��(��GR��ZF��L�Шd�RRP��l�BS<+a;b�'rm����W J�!|l�p��U�b9!�is�v�6�����_R��[4##J�Y�Y7���}�XJ�K���j&Ǝ�^3c���ގ��BL���9/�UV�|໘���[�'(5�B������у/��[�^r ��6��b��Ax\���}.�ƔƇ��=a��#���XZ�l�c��L��L��\7щ����M	kIZ�)�{�n��P�hO���mH������.�.���dc7u�XNm����2��ye��3��pi|�<O��1
�׷�:������+?�����U���3�c^�2d��
��א�׷�:D�<�=!�Q;Fr�?�����N�y��"4���^@�� �`��ɹ]�\�(.ǇQ٨��)�m��cc��
 ��'!`�q�鶖|X�c^��2҆����Œ��}��ڕZQ���)�����z;d�J�g�VtG���3�kD�M���O\�sU_���N�r�,�qr�Ί�7G~@�@�&�Rm�e&�ٓ���+��E]�Ԗqf�{�''*VH"=�L �>yeE�T>�zH����]o ���
�D���#�=�L9����4ħ��o����؆���L�"E|S���=څ����q-�~"<��'6ū���<.�e�����9���!�D�u�j}1��\#ȘTl/�T����@m��c�H:�PnOS)d�Sd�e��&��>
�4x������[H��,z������f޹�xD��_�v��U|��!J�?z 	4~ծγ�]�tߴS�ʿ�{7e%C>��)p���X*ޑ� ��q�}/�(�S�B<R,̓��X��`0�L�9ǵ4��i���Z��t��o�y�v�� �'=*n�&��m��E�}��ҵ�\"�s�u����e�U����q`4�&�'�����`�O�I΋,j�m��!�lZIu�U�Y=���m9��ْ�A���O�i�{��Qܓ��H{S��e9�ϸ�����8�%H�`����cMWڄ�-���"����F�����j��y��.O�d��S���y�x�sj^�i#k����Z7&Y�P8#B��ȶ��̧�î'�%y'���!հR9�C�VVB#�l���AT|�AAW�!������	�zxn��t�˓�rq�C�v/R(�L�����j��� �r�@�?�G��R�u1$�t��g�6qջG:��Gl�5 ����>��f�K�:}�u�H�ѺO����G�aAw1�6��l��'����8�_��-�D��	u��ށ�d�*Tj�#�8f��k���q%��ӪR��O��;���i2��i%Z�	���*�]�r
���0���-Qt6���t��BF]Ywk�y�KvȪl���x��=�K�����;����'����>a;+���#�7�K�&e�5�p}���ݓ������N�'�o�n��B���]��@s�\�nvb/��/�m(�J��)��1�S�W��ʹ��:��K l`U7�I�M��
��xcl����S�ES�E����a
�q�.c���8b8n���-�P"3�%�	Ꮦh�0�H�Ī.�?'�<4��<ʴ1�6��ư5�^3�>�E�g���^���N��C�;T��ڷO 9�f�ጏ�sn�!�uq�)��P�pԃ�J*t���+X��j�Y����pɫC��w���"q�e�g�x3���Z.z{�D��>k
�����灥�)"�Re�-D�gv��@u�X�q2��I�ΰi،5�9��C�D���{gIQo����.��V VO'�+x��)�n�|����t�rjI�T��	�7x����\1�	��r�0곱(��-�E��[�%"��?��.�>==���Y�]�Bʰ�o>^��9v�N��lԢ�3�_4��˹�)��e7֦�oZK)D�^�gC�F�Et�٬�"`N�yS$ݥ.[�Y�!�j��当��x��-U�\�o ��\�j4F�*)wk�4���_J^�Ax�����>k��w�[�l��·�|�ު��/��m)(���nS�tC"���)��Ii�_ �}�>*��5ı<���t�˟��m�`�/SX{Q%�z�w	q��+�]��}�%c/��{�:�sҦ3��(;`Ob�&����X��(�T�B����yo.�EĞ�pt^22��!iP�Q��q.�́���l����j�F��.y�~�6�,���?���/RH�w��W�'�_(K�S�����'�[�k�]���
�حz&=b.��X�������_���Φa�&X#�m��8�Uޏ��
c����]���HrX��A��ɕZ==�4ܗ�����ɚM0�%}�A��ͺ�����S-�ҿ8��Wa�m`z�s���Ma+T����>���ѡh�z�ƻ�x:�mF����������.$� �*�;���Vl�`�5��
Օ�� E+?#��t�{��z��႞=гs!I��;
jo���3'�C�O�U�C��Ò	ں�/�8�V�+e_�,�Fi�9�^ǖ'�Sʸ�FO8�)�~-�$ZŊр�xuR��0�h��,��+�M�F=`K�y�X%)Z�3�"-p��s:7�1aG�:6�XR��&`��$���<�tߦlaQ)�Z�T��B!u��jݺ���_2�y���).��U	���^�2����3�W�o�{U5�.�N��ʊ�OrJ2%~L� �6�~�,��}vɘ&=K�Qa:sD�دb�<�h�q��ᗟm�}�rzz��o"����j��x.��^m��E�H�=�U�?���Q���Pc���p��h�>@����ſ���7�/�.B=�lv�⠪Vg��O/�:�a���N.�L�G�W��r2}�(������ǽ�F�� ���-��P�^��e'U�{SU�i?�~��K��N+�yT� �����9|���Y�ٴ�H|b�V<�]��{#'��%���<���K �m���?���f(�{���bĘɪN�n��xA"�ox�l�v�1��y��Ϗʛ$�ħT����n�]<|&�+�>(�X�GS��>���%%�+��0`u����--�o9���= �p���s�_�:Z���u2Zz)ɱEʭ=����c}��L?�Lނ��P\,MM�>�ǚ�c�$ d8���hk����sU�ɀ��y�s�@���W�Έ%�?z����!�z�n�F�|�4v���Y�~%ץ��]�OՐ��wJ	�[�/Ps���}mt���M����N�C���_���j��á�=Ȟ�eElV�' B��ъ��|d���y�F�=#������ �'�˘.���7q[�B�y�v��~&�xݰ����'�����^� R�{<c�j��N�L19T�[�ƭ?f�Xk6 %Z�h��H��j4Eǥ�$0�� �����-�.��_�!���u�"ͼ���YQ_���-�߀xe[D��pӍ_](�a����?,Pխ�[E�)pH�D����Q��ªR���s�0��2��o_i�ڟ�����7��5���>��8?yC�}�t
�& �����Z�^�m}-n��1 ���x�"���(ʗ�K�қ����~xe��ݝ�Z���*0i/M���|�����V�2�>�ҏ_D���#�Æ#�B�������|oR��ĆXU���a��,�U�Vx�;�Z-����q��=b_;��|&9����;$�7$�8��~�'���[9��۵��%DOb����u#iMI��[�{���G+مDi��X��v�ר�o��H��p��ۙ�rܙ��Z �r��@x`&d��s��r�'�-D�΋�'�rM&��U��W,��n����d-��(����5�a����l��ٺ�k��__�����]&�P^�FO9?]��ƃ�����0��W��Æ	W�+	)'b�#�����Z�cU���4bV�'��G�^��KO\7 �8u� B7JT@������D�&��8M�!��{T�X�Q\f���`�~�L�����t���wZ5�5�sI�B��W�|f���<�i.�Y�f����{���-v0��)�iL�Ū���&�'�CYxђ~�DaL���W*d�W��Cʙ[S�_vP�h��\���X�sB!K�I�����m�)g��f��nt�2h5�!{����ɺ!���>� ��=I*�G9�1�pNG	��e�Ax�~�O5� �H��kU���*͋��	�\M�y�v�:���0��)�j��pU�����'͇�e�����苄��V�K@^��5��L��1ݿ6:����K����O����{��;��g��I�k_9��UA����C� ����i<TX����j����G�?5e�l��	��2��5(+� �t���^
�WF��c졙9l:�P�o����nc�Ԟ�#�iB£!��6��Ȳ���[������R<�ә�>@�{����͂�3�q{7�{An�c 	�\�}��$KZ堳�h� ��o�aE"|c�B�����@� au���CH�/<�3'�Xo�H�¤B)6�\�'���?��ŏ�X4�Wi��l; ��?���q!��u�=��t�K_�����:���Bq	�<��̷�TdcXOK����_��aU+�4��zG�@�b ��6�Mد�k,�l�P�b�`,���v9��Tb7`0����9ભ"�a �K�Gޅwʴꛮ�}���#m��]��9���11���h�l� �'��`B��3{V ��V�{�R�����Ia ��u6��~���J�V̏��*03BC�:�i�>�'�*�n�Ã;�g�	����n6B�!���p��n�	ߜ����5Ɗ�[�R�X�jH2ݝ�����EiS�:<3q��G����a��5�1����V��?�b��N��P��(*o�)~)��M�Z����Ӻ��bG}u�']�Xe�#�WH��<S�G��f���'��9u��>r�_LR*7����5M�0�f�9F�u����0������,I+;Q$�xMz:rI47����R �'�5ʿ�� �z�~P%4�a�V~3 L}����ss��w�):�j�#8s����҄�788m�5n��=@egո�PM�.�U��q��������5��(c������ڕ���]4AkA?�o�8��ô������e�p4���r[;C�nt��`�e��|�))mtY���7�Y�\�'�UT�:�S{5JL�'���x�`�w��QF�;%wM��H�f,�u�!�n�=�8�ԼƅDO��-�'�T�[���k�b����X��g=�m� ^�Z�jUs.���+���m��>��I�~�wV��H�)����O�3��6~^�mj5p�ʍvR����=L�~��^w{�Bd4m
 (�es��CuCᥑ�^�Iy@-p��~( ȑ���	G��ǨJc,A���������z��	�7�?��P��7��Ш6{�o96i�l�a����Jq6a�C�1��)�'��T�Wl{����گ
R�CiӄK��˭��:�Y����J�nn��tZ��#6�%����.�`��8��;���y	tC�!�	.�g�5�v��Xi�$���sm,3xO3�ꮌ�~v"�\m��{q=��\g[	��KƏ����:��0�r\�Z;A�n99hdC2bF&P؏��I�Gʴ����	Yh1ISc��`ߠz��4�I�m3�n���L���E�?��	�;:�u�opeic�q�w����S���]�9���f=ɤ�O�7��#烧T4PRe�&ݯ	XT�ȷ'�^���YL�Ϙ�X:4�<�ksO"'sPJ�]� ze7��<W׸�*��$���~����"��
,"�H[KP�62IM�4�*�ڴ��c4��p\#�ԯp$�?�GyJ���_�^^6�)��-����z�J��آ�5Y�w �y}'�F�SkO�NUo���N":EJ��HXx�/].h��0Y*�CN3���~�^���qQ������&�\ey��-�9�NZV+���lwI5��h:J_��6����9�$����������d�0:�w䡨Uj�ےޑP�56V7�LA��Z/�iN���-m���@k�<��ԱČ�eB.|�;;����~HA�?vq<M�%�-=����F�S���2_IWڦ�]�yp=_[s-��a��f&��G�� Qa�b[R�sr������
��H�)��M
p�d.;j/<"8pC���8�ns����"D�'L����ΊY��̉�MI5/�|�
�tJ9β����U"��	��wś�(nY�Q}���ku�Q��L����B暵1��irIR��L4�)I��PFL�"�L�1݂�:��
I��U�[4ׂ���R#�*�7�S�G�a� 6�����~�Ɵ���oؗ���s䘬�0�vr�;�>/��(Ҥ�U��i���ƻd�~O�D��PPu�?��6�� ���=���@f�c��:}�TrJ>��A�?T��o�49s�6ԯ��;�z��O����g6������c�<0��o��+�S�{ Ӈ/|�r^��N�u5�@1�p���,��E�k��1���v*Ϧ6C���J%�RVD-QX-@�"��D g�s�/����Y�G` ��R�⡋9�c�_4����)U:֟�D���;�`�.P;{1�ކ������h������C�'r�I0�*?��3���~���	j���Q��Ӥԋ�r7�Ir@Ā�6��S@8`'��1)��jE���@Ğ.yB່8�!D:$Ԧ�6�����i�ZBz��Js������
��h��6Wyzq�b֝HΓ~{��8Y���X�.t^y~�<�kb�!���"���I��)vy�a��@�[�RC�	`x< �R�'I��f�WE�A=j����m�#�ȝf�U8@_��D.H7T#���gѧ�WW}@�o��ُ�Q�~24͠� )�t �\u��\��Kf·fV��㔅��b�XDIu��I��9]q�;!�UJҡ�����I#M����_&�;TƗ�a�3��e�ӻ�/DsJ~�����r����w�T6�Ch!#�������EG0m5/E�o:��b �D�� �)q\D��:���ݰ�?�)�ڗ���v�V�T�nY��%�hԽQ��wSI�t^��Z>�Oq�1�ٓs�-��B%��bE(auS�8MmW�`��O�~�*�Jݵ�¾����b,��Hd;�T��%��$���t����>���̚����	4��P��rўɧ�a�CѸ��g����0��e�Ԇ����H1��;����tM��=8�_���2���� >���|f��4��٢�B�i�{�W�.�t{	�T����kI���N�VF���m�c,�R�>��(~B`�:�`_Ղ�9p���V�k��mQ�Cn]X �PfJ$����W���|Ϥ�%�M�X�4��|����ē�9'�������$ �Ѩ����)"��?�c}�v-�u<1Bp��C�T���_Z�H)�uF<�%}�Zlە�����D�@T�����x"m�`5.H�ިg~\Tĵ:;�]aqf�>��C\��F'�a��^ؿ��\s�D��o�a��Ko%�;�I���A��Ć������YYm'+�Wi��f�d�ǣ�5-�G:�O:���JYΞ1`q���r�i?�c����^�B�q&�p���^�Csnwп�7Wd>v�dc�f��/���2�l�IBR����`�!�⯁�=�xWK��W��B���ʃVi�Fz���:S�XIuS��>sC����rG�K�zv�G���y�9��e/�T^6!\�L��i��]j����_����X�M�)H�Q�R	�_5u�,�CU�A*�o���w����EG!fj�4�#��h,�7t�8��	k������]��V޾ ������|DQ�ZgLA`6�d�×�F'T�l(��x,! ?��P�3��J�F�U�Z�_ ���<�mB�3���#dt%7�t�P��h���Ҿ���Z�Δ���N�����
��=g�09��]7�u
=`S@X.�i�@_�/_+��86-b�]���_#:e)��Fd>�v�֪�2���b�ӴՖ����j��E%j�A����^����;%A� ��X�Ԁzg
�։�jI'�X�`�y3�s���ȷOD�~�+�h�mRCij�����M�eo(_.�O�*��m*/u������NE���<x �C��
Lŧ1a]`�n�i$�9���4˨x��f�Y�xk_?�������ȠW%8����p�AGb3�==\�4��i=B�6�!yf�ߐ>�33k��e%���ց&�#v	+��1��$����!�Yc�1��)L'�d���M�ZL7"���:���?��(��9!z�.!M�[$��s��N�)�kw1��m�2F��Sՠ�����l�Z���P�MqI�~�7���TM=��y��\��j&��Z�Y�a{|�-�N�ށ�m�d�A�����s��Λ�ȵ�q�b��5)���l~6!ba����`eYv@wڥ�q�Ωc8����O.�] �C�f����r�k��2�@*�G�'һ0y&�H+9�x����j
s�����*;��\1�s��OBf���8[�L2dD= �J�R��I'Xt���(/��W/3Lܠ%��B5J�_�: gp���~���a�"��ʏ}�bY�g�RD����VB8y�U�8!Ź��ot�FC��UHp����sDӏ&�d���zq�Ԛ�kZ-�N���� tuT�V� &~�|4����{;��:��
��iɀ(*�J$ӤkTbG���/l2D�LV}�M��_��7\%ٰ!O�1a�M��JE�!�*��"��m�@Ŭe>��5P;?��Bz�4�YL=�'���SX��&sV�C�ٕ�uC��L���KV��}2�:Pu����ǿ*��/֩����ׂS���m��Q0��o��V�l�s�:ȋ<
z8qݙ�i/f�Z�c��[\^2�����Fe,��\�����4�eؔ��^fT�a���	�a���b0�D�����%,��C �k��mX��KK|�o���Ԇ6;�.�BǶ����*����餒Y �@����M��S%v����1��/���%���tJ�n.y&_�.��~xeF��?),3^�����6YDg�*A�O���^�?�3Ӡݔ`'y��%Zz��1�2�_7K�+����@�v���zO�5tjn�żW(�%^��8B%	�Y�@Rɲo����� �]o�<,��ܰ�����?H�Ö��^�c����c�<�����k����v�M��D�̭�?t\8�U,���,<��?,�;��d[ �o`ɭ���g���H\Q$̌��6�K��{B^~F ap�b�����UΌ�V�����Q-��5(0w�U󩹾n: W4ӱ7�m��8G,��I� �pyX�쩘D��-{ާ��t�G�2�K޳���?30�e)w�Xe� �1u���gi�O�d%�1�l�s�����h~&��{�}r$ͻ �Ʃ�~g��X�m˰<�:1��[�9%N�h,*w�8Be:͔�TfyY�7g�x�2� rQ�R��Ղ�1#}��]����2/���\{�ug��M�`�JE��q!��U�9Y�5��vD~\��W��f䆂E/
��\@V4�9[(!p^?����֯D<��:F-�&,,�B�0���9$�/1�9��<e\�1a]s��V��lQYC⟛>����XI�|�@ �tu�Q,_�v|�E5��Tf�L����!�L��L�q�μ�)A �(U�(G�G%.��C�B5�\iu�����B&)���������-#&{�'���Vk:�Ĕ�W�ghUi� nOB�y��%7YM�'D8�fk��'RQ�,���+��<&��Ul^�4��ie�c�	��)ph��2,���'q�5.�Z���/;�o��nH}ݪ�
$��	=TnɡL�CZ�!!&���^*�7$:�$����nJ��T���m�XNX�13�Qں+1�utA��f9wtM�"c����Ѷs�����~�{`8�o��e��k�����~q� k�y�>�ڬ��h��?Kaul��s1��w�RV�P#�_|ZW��@u�c�'SG��|W��K�\���O����C��%�iv\�2��XU7�6ӟ�0�G���GU	:A��#;�;ۻj��̒�19�Hb����?b�U����������OX9)O�FIY*����N�B���9���̛,��9���:�8�'���Hkp���yn����D��W�w��U̂���.9q�c����t�Ե�t ���o3Ȗ���ZN������ő8;*��*+��$q�{YYr��_h��@<+��`y�M�f-J!��)��1��:FfV2�5��S��s'	�@wT>��`��O��ۑ��%Bw�{R�w��%!�s���%Ug\�G��h�,/Q1��VµyH�;�،b�o	�H��l�m�3C�8F��d}�Z�%� \Gq�
؍"�g��}娹�-6�܅�@�k5s�.?���By!�C�4�!�H�!Q�`��.fx���k�����C^�@&�J�ˡ�^�V��y.DH{K�/�?c5􀵍�A�Q���f��>N������r�J�N �P��n�����{ɻw�V����Ki����55�6�L5�2֫�޵)��ΔB�Ț�fX��R!)��F�-;	A�:S$A�J//;��Π�qn�i���@��혫��"�����"�$8�� v�\^Ux���t�!T;ũ銀Bk�v��\�.�l�Z"|��4�0����¡lSًIz��Yiü���$*]v����A$g��W�O%'q��X�Ie��w5ĝQ�Ű��J�M����,��M�zD'�.��.E���8�?�Q�d��k�4�S�-��W���?��H���E��yI�
$ 0R�.�����f)ί ��g�W��CP���u���V�]���8T8|��[�'=�����҆�&�M���W���Dt���(es�PKa�ig
�U�Ό0�Q *��
�f���0�k�u��%�����'�#��k���|9\;"_$L��F�Uf�7�x���Um|�#�֓%�@G��ˎ/�;�9u�K�����cq���NEn}iׅ�AƎ	������M��|w�����Q���PE��5!6C�scgQ ����}|��Ы�ŷWަ������v�*9!���):(��d�j`z��D���@� D!v%���/���"qX�����h8�=��,���v�2wT���f�	�ŏ���e���8Ҧ�{݇��=�j�Z���s���^;+cP2@ϊ�2Az?�q��V�ՠ�}�J��Iy|�����ߚ<�^>�j�ۜ=PJ����o*2�B����Zc��DTv����}Ւ���x�q�"5΢èh����X�jF�q~�'��f���}qy��UYj�6��l�9u^\!`��������㻨����<���k�h�L�p�/h�x2��v�2� ��z�������Ԙi?�p���7z�Q��l����lN���3�\�d/�%�w�*�P���p:�!}Ï�j
��� �Lyz�4�ad<��A>�}G���?r>��OT�|�H^}�L�>ܥ��f���Z��Gp۳�9�?�9���)Y���Y�������N�0B�&s���uOzҎ+��:g��W�Y9�Yz��r+XE��)��+�feܽ
�bp�� ����o�ÍVu*8���r=b}�]���O_���x�9ߋm��q�?-p�{Xe�5������@�_��S��B�fDY}�M�|��}��d����AI��D�Ը�o�A���ͺ��Уs�V��Ya`���#�a��h�\�2��jS���o��U�~���wjZA�D�a�3���&n5RCr{�^r-�~T9�CwZ�H����}��4y���r��R�������i�Ïl����&�ZE�v��h�c1�؇t�~�n�K�͡��XK�Z�eZA�٣���L
n�@
R������ŏj\�j`�+�8��c$[�z����l*�7AS�d����^L6��X�շ�8��1��@MP�0����Mu��m�"�8�K�yQ����ܩr����'2m��GQ�3��j�~2f�ܦy�j!C�O~�Ϳ�z2��H�}�����hͷ��e����B�V~A�A}��U}V��LG����W�4M������ʸ����Ձ�Œ�^����t �����jl�q� �CX�(��H��bNޮg���[�!s��j5#���#�����ݔ�Z�_�b�w֠Ï�RύmS��7o6bh�a�Ңq�W�>���0ꇺ�=n����}Q&��0�'kl;�������9��we���tI���љX,:T��]��W>�|�JP@�S>[�ZГ�kӷ�V4��#.U���(���������Q���KL��⣖�i��Z���,�������8�5�<��[tBB��I�����:@�Mi}D�b�I�/�eP�ayF�ɐ@q�Q�*BR��ܵyY�L���v����Vb���*�,�;�u��C�vBմ�l�z��ʗt���'��Ȗ�Ȩ 	�wt����-�|!S��/k�K�t�Iu�S ά+_�d'>��48rxn/���D��v��*����	n��9���2��8�\��Ӗ�����K�G��i/q��@�������#�\��Yh~h�R���</g�}$�"a40\�!�@��o �*el��� L�@a�Op�f�����dbȉZ��k��w�yw�SG���- ���!L�B|3�����+���шR��B�^o����[���> ��vc6͂��=��+K�R��j����`g�!�R��29>�A�2�Hc��Z�m�u匽���mCY�k�y�����z;�3�f�'�2%�x�K2]��s�'�w�Te0���[w�бf.� ��T�:�]�;��}1�sYE��z�jebb}�͚3�OF;�<RXiW;�nU�,�����a$����7��Y IHJ�:���~��'\]/N�nw��!37i9N�j�  ��a�/�{����ϔg�!�s_�v�t�5,8;�ݪ�b�6L^�^'�U�ru
푁�ؒO�v`�K.ߓĳ���S#��u�:���c*m>'�(J�e�AP@;�N��!����~�R{h��eu-����m�}�-�S���hf�s�������B��l%O[K�j}JD��q`#������!�!o��-���Jsq�ȿ����M�����[��7�j@�X�*��Ō�򙱖���8���n��|y:�ʜ�s�KY-��ݙ#����<� ���!���~�*~�:���a��Ѯ�k��w�/�����I��T�8�BFL&s:��׹�6��eK=�>�_/c��r�8��X?|�9�ވ�Oy��C�p(47�	L�8�ıۑ�N;�� [�";}p�dᫌ*K1�ϭ��I�'�h�Z�ҁ.��s�YK\4��5TA�v�?�؝�=���'�h�| du����(�� 
�8E��㵕����h�ҐR�����(��fz���ݶ�Hl�������$Vdh�h���%�cz`�=e�qmm��{��H�Rl)ED�v�O��;��r����X��ϴvo{�Q�QdM��k:� d4���T^��8ǽ���������r8��|/�o`#[aVI��v��a�&EJ��xYvA�w�M�{^R8�S�p6�R��2��:��a���wg��
���qF<L>{[ l5P�	Q��`ᨬ��c*�䚇fx;���MeQ�t���6)�d�I��r/�e4?���ÒxJMu�꾯�i6(s�_}�T�yX�~I����e�h���۞�ߢ��#��y�Jd�����FvǕ19�T�ք�u��1���.�@d�V��o��,o	�I����j!c>.5I�����Lo���vDMN��4k��C
�0��3F�K��o}��p:z7����]��a1��5#�~'��d���߁�� ���?%Q�ͮF��η2 V�$Y h-�]h;�&ҥQ��Tk����G����I�򂈶O���BR�qn��|R��_"���sԛ���Y4����d Y�#O该���!v\�3�(o�6�����Z0si�b5T�5�RrM���M���2���_�g�4x��I:D!X<G���0��� ��y=Q��D�e������j�8���R7m��`�;�_�����Á;���fK}y�,���J�*s�5�~5�T��D���.�Zea C��e
b�H����{��޹��+�[u� �(�M,|k�%�1092��"K����F9��*K�o+���Ls�|���0��<���a(d�����B.f��`�$�!�5Dͣ�1`{j�	�쇏� ���v�t����=���#(R��x�7˶�l-A��ܹ?��Q\��c��=��s�����rR���r���H+j+�gɱ��ϥ�< ����J�M(rl0�Z���9V�P�\_��)E;}��k��O's��$i1P�)6��ȁ�[�O<~+���㞰A���H��>ț<V>�~���k��@X�,;�PΨNBr���J{�%��3(ӚO7����,���il�t�#�A3<�߉���Q����p�߼��@�1��?'*�΍F~�D�+��q�t�L=|++�vx�F�c������.��\"d/c'��V��u7ɼ���+���*T/g�%m졬����^S�\�L��3�8��>Ĵ��y
�G�A>9mn���\��4)�F��MgNP�
|� h�|O�~NU�U��5�UqD0�2r]ˡ�Ux��]�r��p�?ټ4�MX�~_�y��w~/�S*QiZ�:Ŧ��M��B�!MU��e<;��Mo�7�_�{�W���?q7u7�I,��7��P�`d���^��XC_�2���qUv���Ǡ
����Ǯ�,� t?/�ﯜ�:j��X��A Ї(���a����o��H��p
i��:]��Ye������͎o!��(�;��l�c�'��H=�E0��;&HD�.�|�Y�sh�ݭ/~iܯ��`=:�x��|��]��d�;��D�������ez�\����^�Uܭ��.
�r��^�8!>b�ʛ�[3,�/��
'��.����aʧ�JTu�ꬆz7I��?��|��o
�R���g��^��(�L<nV�U�I~(�+Uք~H�\;W�w�+/L-փ���A��%�u�DY��h���p&�L"̨��:M�VCC\��LY����|o`.8X��6�F�6���ù	�����[B�3�t�ĵ�ض*D��1
��	l�Ƥ0v;��j��i�*�-CB� ��l�L��Y0? ?���U󷆝~L�J6M�n����S%f�B�]ۥ�ɉ�Zz�1��v3�BM�$S�4eii����%��ç�4���hxJ��E���_�ސ�v�뺜<�T6F;Oƥ��#ߌ��N�VI� ��I����D¢ g����n�^N�~r,�}tf]�����%�q���>-]����B+Z�t)� �<�h=sc*����c�W����v�z�$
\�n��U��lQe:}���+(����'k7,���C��}5��Q E�ߖ"n��d��'C��S`�!�} `���-�k�g��b��x�sr�����!��F��V���%7{�Y�\>(�L;9ĝ�3�8������U�a��{�-C�P���A{��LI̮M6�	�Q�h����[�����8B%,Z�
��,�V����	�t�K��'īK|�N����t"9l�6v��[��Wp��\-W��4�w�g�'o�*Q���8�ݷh+�a�]���F�]�v�P_@�)^��"ݻ��	�*���4���YHA�T�p%��%��\����m��2R�\>�K���v~�Nzx�2[Y��5��^���9��ucb|��ݢ����N`�A�6�f��z�%)���#�_ȓ��8�[���&L�v�}m�ikj��e�:�i�JEd�i4C�"]3oQ��0���?����\�~ڶ'@�l�e�}�Ҿ���+�M����� �$�M�[��&�J����kA��z�a�d���	��k���-���XǨ�V=�0�톳�b��1B��g��)-��������DC/���9V"ς�>2�5K����	���>pi�P�����Znf�q���.?�Y��}^iI�R�
[����8%c0bPv�l��F@WT�͇GH�1�Q������Ɂ={��֢D1%�Y3L�n���� �h��(��nYWbG�E;��Oj$j�������L��~�T�h��2��Qu&"����(��2��u�!T[��d2���0$ò�j\�R��ِ���.�̯��}�G���Tw�F�ݟN�#����\���^M�e�O냈�Z"xި[���FsA�t�Y�R�uv�����0P�ـ�+�9�����F�@�
6v�T)���?qXW\E2[Z鸘3PG�V���a
h�c5`�1����șX�1�y�����ZB��b�"�e�xc |b�'�K:5�ٚs$�������!6EC;aF��M����A�g�s97m5.�|)}�N������'؄�v�mn�mj�
`w�:�1�@���9XI	��*k��Yr؜ �l����q}�)ʑU\+�8lr
�O͋u�l��T�����4 Z�-���?*X��[�˅��UW5�(6�A$lrNG�� �'4��� P�0����n�!̀��wLNb��6�����ʺI���q=ӭAqQ̇��V0�D�����Ɓ��{��{�7�X�D*y?����\AZP�ҐzV�L|L�'�@걚8\{W*y	�4P ~h�y�����"-�@���p߆	ۭ����Jt�һh��1���3��Sʝdq<�	�D�n��D{p�S�n���q�M\c�)�pD��״�?(,��^��D����q��{tw�o�x^�Cڃ~-�������)��b8_�����*���� c�L\������e�����5�QB���P�����*��[�ɚ:k���l�|�P�>�2����@A�*��$8��h&�~ͷOj�~��f��j%�Xj���e/���y�׷�5�w��Y�x2W��/;\(���R�(��G��k��T� *��;�?�g/�׿r%��f��h��hǑ2,���̨���������&'/&�S��Dcdl�l	ǳE�RY-�9v�����ޚ��8��.iE߇�8��W�E �E��{9�ǛTH2K�j{�t���D5H�Icג��=Q���!<�N6f������W�����̟!]<��N�E4�y�	A�0�b�&jǬvQ`MϡO
��-�#�t)�˵����0YÞ�<���d~����������:���>#2�w/}��Cփ�o�B�����^m6�4�L��ˏ����A�G����X����Ů��ȍ,�e��>L��N(a'�/RS��N�1��V��U����pd
�rėq�N93X�n*vO=��pu �̓����[��)�~�l{9�
Զn�_ܨ� �kAo�Ʊg�������P˯���ci
V�X��jg�$=U'�`JV	��?(S��"~T��=�.����ك׽3k�+�:�j|���J�5X����y��wap߉��-o^��	�l�ߓQ�Q%�I��>7=	�L�C���,�?�%a�����<����f�5��z������ �Xx�Q�C+�t���#(�1A�!�:A]��H��<R;u��	T+��)�R4L���2��*#�!g�\����r��p��N~�Ѽe���ah--V��j������I@�m|���,{Fom�aM��q��M���-�g)�H��ٞ �����N
������ r�p2�. Gp��Y;xT ����̘{4��P����f�B�zn��֙ sg����jp%�F3"�^�Y���1Yw���ΰ�o�e;�|Ru3bY]^2_���X����	�R>��@!���G��*_UԆ�~1��c�QH$�z%z���6��27�eU"�Y�ҿ&.sƦ��[��S��`�'�n݈�6/Y�́�77�Ui-#����)�'88TRk�)6&y�M8��a9JU�ʜo>ܣ�����$r ��a7[���$mԦ&9D-�����pK����B�O(S���I5	���@��lm���T��3c�>�7C+�2��]Oô;j�!t)n���zh�2GhH��`p�
u���F�D��]�.�g����7gP�>�t��N)��e%"1�+��\���	M���^�Wh֠�}�yk��'�B�K�F6:5��K4������Տ�Z�Z!8����L�,�r���%���݊gZ�n�e����"qU��ā$�o���|�- Ϩ���r����2Ɲ��&Z��"���2�� �p�!g�$�S�Oo�u�I�ﴯE���t#��f�g������Ƈ٥��"�U�*ԯ��8ݎ����1�/)1r�*��/ 
i}�y[}�?�a݌���9����r��W�@�w�)k��e�ΑZ�_�K��ȝP	���8O5��Y^�	)�41RDѲ:�V�d����ص8�&h��髦!���"@�*]>̱��H��/G	�D���~MYs#�&}rn�M����&�U�)e�9�_����(�?�F�φ�����i��9�<D�W��FOc̯�^:C��uA�A�oۡV�{���%�B+,-�o�YIn�cq���!:�����4��<˼}��6g��j��	i��E�C��qyP�C��L�;>m)]�W���@����6*B a�a@�����!
 R�2ES��w�:`\n{S���۔��$y��8M��n�5�g��j������Ĩ}�n[̸C1��wz׽�-g�]M&vA5�ՍL�V�VP8�t9s�{�>�����o��`w1*'�d�'�Ͻv�|~>y��<�Ov����;�^���D�̄��C\}Yo��Z��7I�\�J+��Fh�
�� ��ql;ugd}��ϸw�$���tY�׏��
�_)��0�M�U��1*材�S�a'Dl�9�wKm(��ʷm��'L:;�*6�Ļ��gN�Dm͗ٱ�}3 �P�s���]W�8!Rv݁`v��~L8�"�7Nͥ���'.����T� i�;�=em�3*9	+�*Bϵ�!�JQK�#8���zD��
;�e�.zީż+zL�giU���C,��ݜ��_�ӝbƙ1�:1�4+�/�,o��ÔÅI�C�c�Ԫ ��N��צ�0���,��w`�f��X&���-73�����Fk���*^�L�j�P�V��a���ovȪ"y�b�7w ��Q�W�~	�k��c��4Mf�\&��!)Ws]"df�`�*�h9]L:����:R_U�N��!��LJ)�Q/���ND;�8��~o]'*;K��s�����D�1�4(;9�Q��`� &�2i�+�f[O����wo�\�F^�.Da�x.�-I|5�W�	�s�0�����$0�A��h*L+��)̻͡�>�ڎ@�{E���찴w|��N�WĎ����M��]ڛG�X4�#;�&�l-�Ǉ��)�@��L9�-Ia@$�>I�h��n�5yJڧ�!@�^(�{)��֟ID�?�b`v�G��g4rZ��ET]�C����&;Q9'��^(
vM�}q�= ��幪�=��F�ON�&7�Ҧ%���q2�!�	��ݷ�1q�̸c���R'�%d�\o��?.���oڢb�Dg9(����bRL	�R���ˍ˰�x�0Yo���y���!��K��
Qmu�_6ۿ�N��=�]����"`F9=фWI��Y�����a����al-��X��ň*ӫǳ�o ��hy��+�B���/i#���Z�	�cd�]�~�r.}4�Z�%��h)"�:QV5F�.Q�L4�{�Q/bQɁy"���l+��2^����9K_��d�>�S�@�Ma��J�i�������Wbg��<�I8���ɚ��ƹ#�Fc�9B?�Js����%�;�4�w��WX���'S�MZ�mN�t-
�H E�C�T��������Ūg���m}9�0���&�W P�;�g$�s�$jT"��-L��<������~�x����%����K��Aj\���p�~�}m�+������ײ����I�F#�|E�C��Jx��7��r(�.T�����
4�Ky��~Nﲇ,�O��6̷�f؜F�V�I�Lň>� ����)�L��@�)�� º7�o��0�$��=*�_Q۴�m�A��hY���Ew�B���C3iM?��H�pY�k������o�/������x���n���ſ/��:��|Ȥ���_��F���& �k�0��9M�.�?�*�����"ر��E��c�2k4,�9#Z+n�\��L��9U���h��6�Am�g
T��O���`��
:p��� j��|l'O��jy	|f�KƦ� ������Ip�m��Q��� [�����bX��v�^���1�MH"v$�8W9���`�;������b��J#3h����d�5�Xk�����o�ǧ�Jr���H�Qb��8��j���i��������Qe��I�26p��H5M��R��i��Z�U�Ru0H�[�+4i]�y�k���\�+6m�lrc-Dj����Bl�0T�7�<�Z ���}Q�u��Q�)���_�9����Vp��}�͗<�әf -?i�E~�*Z�$�?�m���e�Ôc��PE���`8��`c�N ���\�`�A�(p���E8sr�z�����޿�7��,/�ifvq�ݤK���nH�a�S�%+��齼��E!V�eև�g��F��ޞvn@��1��G/�a�������s��i+��TB��EP�f38�BAS8��6Y'��S�Ќ��4A8��D87�;�.<�w܋�[j_{�!x ��a�Y�/101�Q)���6(�r�8̟�"���gKO��Q?u�Y���G��\��l����)jz_�B�3�.�x���� �wM۪Mh�� �Ѷ�S7D6��N���:�BW��,�\�F��ED�\H���v���O��B�KwRɻ���w%~B�}��3}M�9��d��[�r%t����Q��*?x��_�d�H��w��=�<n<�����_5�$��/�0'�4���1�+W�oe���D��PT�-Ū�aL0�v�h��=�<����]�'���M���P���H���ů��ʱH1��f�Is�q��[\0�M5�+o�L(	Je~Ap��'D��1��.���wC<�,(�ou�WCn�����Æ���"\����N�qp��}^9S��� ��s�gcf ;v��i��8Ć���5��7��k�������,�(�E\�ޯpN���1 j� S��8S�H�3���)��L����#d���	5��2�7��

4#��!�u�"~�h)�k����Ҧ���������H|s����Msϒ��N*��wy���:�k��N���8_pUBVp&���S���~!�T������O�G��L΄h���{E.$g"|��g���f�@�:���-Zo,�P}�kq���«��p����Z���">0E>�|���K�7 J0��(?l��#<��!�a�*?��C��.�Eu9v�j*���*#�}�7x,�u��,]rq�$eb����@���
��ËkX�n/�U|�wD�������S/�7Z�C�{C{���.���P	����k4&Kؚ���Ϲ���� �5�RΏ�U�|������%,}sU;�mn�ū��\)}Dݡ�;�o�F �q�xllЌ��VǡG������o��#i�b���,�tY��8l���o�H�2X�J#�D5W]^�����m�(A�׊����_�%B��`�W��u.M�QE�J�2�m�N �ZUXߟEٛ*��^�:X�".+�%�;��0�{[9���97k�hg.S^�K�=,#�O�_�*����ڕ��2�J�.�]r�9��u�k�z*��~��*� A�-!N����W�Bd�{�'X��Z��kkW��~ޗ�{�9�3�#^-V����)���`�d�;����f!�Z�q�pM�R�BVyzD�����{-l�ق�쪓1��֌����^�������[v����L��B�ǝ.�EP}�#��G"��'A)&��"�Z?eCZ���F��^��ݪ:���
��C�1��^y4�X:���r�T��p2Ο�b����쓭�j��7��Cʐ����L���\�I\|9�މҩT'�i�so�%���:�����XO�B��@H	a �f�e�x=��6g���Xq��e��[�WJ�����k�t��6��P*�i~Dhm	�6�L�bf�����5tZx�Nݵw�%�9n��+B�6^�;��͟���$��k1���^�!��]�1ٿN}�}��Ö��c̴��/�w��;k:X�x���E{TuN���ex�^�Bp��5��U�)dT"8 �W�v����B ~�v	����1LL~�}Cv��=�`Uz	�	�}V��5ɡ��8!��G=�M�"��%���7�3�y()h�7L�i9b����,w��V��������-A�J��@/�j�8�B���¼Gs�e�M-ie^�#g�K@朗~�7�V@C%0\XH��`�ݙ�H���'����$��U�R���$2o w�d[���H�S�ID%�]�mk�Jed��6���,���.���;�O����͠u���E��|vG���Tt�_z�
������1�}GI��4���iܖ%��Θ������U���;ein��H���6?��������M��n&Y�>m���4}���z�� ?�K|��AǞ[cݒ����j�nA`�������7�<���)��sw}���}I}��;Bf�����S��&H��p(W�Q��~��*��m�ݘ6�S̹��5s� �h�y��?#���+i-�]}<3W	ȃ!ٝ�����a�l�m/ճ�1�〲{���Tõ�m5��!4ln��;����$mCi@��l�����+hW;d0u�L8;Ha��(�����ɇ����fc�C ���5�#K�b���@h��wk}��Φ&��v}0�'zv�֛j�|��]�z�YX,��hRiw~^�X�����#`����޾���q8�*��u(kF'�!r��CA�F���ڷ[�}d*싡.v4nU�����K'�B��BT��E��I7��a�a;E��.r_��`b���{]Y���6kVM�~8(?2���*�l'`�cД�� ��|��c��0�$�,���E`{8~o��V�P8�����%>���җ�P��]=1�^�-wc����f\?#9yj%UIwũ��o��t-��p?+��B�*Ic��W��w��͈T�|f�͝w]�;x�M����W<�v�E��P�����[]U�H2'����5���8��?�B��� �A�W���E��n`\���,ec<ک黕�Xjj{o�V"@��Lsoa�Sc�HZ��3�dD�b�
o������7�H��NX-hܩz�]
i�a��d�:����{�ݞP�#K��3�C�2�_o���A_1�(-hg�B�k�)#X�	Rt(h¥oȊ�
i��:�V�Q^��L�AY�_�Z}uZ�+�f�e�f�����L�{1H�7備-h1��ٟ%���?�3��g������MrR��#��Kb��~�`��Eo�kz�-�v^z[�sD��&:�M�y3|�F�%�~�	NA����d��/�	�\�d�������F6�ݨ�� �r'��tD�]��Q��S�Xf�ȿ�����;�00�O�T����\��&L*�&'���3CV��Dp=|�0jV+0K�>l���X�p�o%�Y�.,j�� ��h�uU���C%�"���\;'�5g'�{�-g����syT��hl�@%��d��=�my�_�M�O����C�~�ّ��]��v�&��{n��P�i[��cȁ&��ꗝg����Ɂ�h0�8�hT]gRF��p��׿��GW��[�l�z��#a�7�y����	�̈k#�Z5g�2��H
����=���3����8I��B'�LH��������i���5-ؒ�%�x~\T�?����<�(f��q�"hSd�8�N�l��ý�:�B����4�n0��i����4H��v��v4C�����i'��(X�%9��:Gp++�h��u�N�׎/����|���71�����=�O�[�n`&���蠰�����jo,�f6��Ё�;}���p��'[�y�l���-̒�6T���^� ������a��i�����gWIZ�Л���呎N��Ӂ�+
&."7V�i�ucD�b�ؓQ��5jb)Et	Y�}K�ɎF�p�S�j��<�	�W�$^C���Ӓq��R��Q� B�*��

�+�1Ю���%���i�6��kv<ߚ|��_�(�����0�WŁ�v��4��)��q9��?���,�3`�"���^^��.�W�U�x��"��`�ES�bZ��׶�E��--:$�S�U��pp��a�++a��� ��@��2���^�*��-�fw�-z�V@	��Io��[ �\��WH8Of�=C�(P���ON�n~/�՞���* ��uH�(����~�m�n�L���!`$� y���7o�����^�B�/�`������Ӳҵ<;�"<��3g�`7'� ���ܘ@�wfͮ�E.���	h�I��Ű �Qձ�OM��5^���n0ŕ��ziĚ=)��3ȱ�D�������`�,Fw�*z��=ص)b��(�(d��"_י�O�H�?Ms�I��^���a�FӋ奢�T0ګ��$ȋ �ܡn���0l����7�qh�T�@��T>y{���}�?UOg�rC^c5��$�G���q��~�uw���-�q	��������4)m�	!�N��ٷ���nEG,�����=��9yQ�	�!���L.��;B4d�rʷ�t���?彮懞v5�{K4]P���gJ���%�ȟ���J�Q����m�ڙнg1�R�u.8�
��蜕�$9p@�{�H�G�&�H�Y�׋��Q���ۜV�l}��u�3f34�O�Ύe����w_KB����Y�����9��oT�N�����^og҅���A��o�i8�]t����4���"F��>���Q��.Rrj҈�^ގ޵<nD;
*j����F��~�{ ѱ0J�?B6oc`#��zM�)4��y��Z���!'��}�S�[7X���;���=��?�*�I
��~�xFwӀ�u�/ft���H}�Yʠ�&NT�ԕ��ⱇ��~H���KBV�kȲ�L# t�f�`��M�� ���������0���2��نz
��R
jpz���9�JjT)R�P�#�g.$3;�t=�J��� �l�[����d�_�޻�	����.Ij�k�
���`?_  �hmN(ޛ!�Q�1]�]u��V1��d-8y�4XS��n[jL��!�����h��l2Q��ʭt�� |ӽh��*0pL�SOU�mGU�Z�p�|k��`�Ȗ1�N���`a��x�az���� �D��r�V�u�v^�8?<���oX}�ҳ/_c�����a%Q��,���Y�J�
���ϙԜ�óK��o������N��������
�v�����A�Ά�oR��=ġ�6�fNn����2�KJ� ,�V������O�gu�V���d����=7�,V>��\�sv	�N����p�f���8g�BE9����E�y����Iw��+�������W-��V{�X!
�Xx�)�������c����EvJEk>h	�Iϟ��;\G�s�Ý�k��xk���ګ�V:3L���w�.���&?�% ݕ���E�6��z@���i���7>"���&��G~ӕ�	�����_�}��|�:��+��6v�ډ���jDx��;�r��G0
�n��c'��=�����V�e�#'h'��m�����u�Lt���Y� ж�牶B{���|��A]�^�tq��	e�	�2ۣ��[A��o�栋��G�.e���v��~nӿ��d5L���5�G|������EP�"��h"�z*�X@<�G�����cЫ#:�]��yoO�x5`���h��y��z 8RT��ߺ[Rӝ��j����9��BGOCp8)9i "U,�A�P�n�c;��L.�}x9O��3���+���E�����CI�G��m�'4�A��!F���|��ȝ��3�����ӿd�1����ލ���a{�8��<IS���D�_��)��"�V��Dy�hè��Ǥ�S�!oEN��Zb%)`X-4�������������M0\�n�h�YFeS��69���R�4ݒ��WR��K��4K{�]���-��D�/޻I��3��D���m�|��3�̎��7�Q���M!��l0Iv�Kמ�[�#����ح���d�QEO�Í�~䎎i��ɋi���V�.���05�PT�P��ȹ�ӊ%ԴrB׺j|x0ڳ��40n�r�?lrծ����?�Zs-�sZ���`Q�����0a}���Uq���ϡ�'�����K��`Φ��뫗¤Zg1����%���Y�Eü���lW��}o��z�UW_�Vo�ק9k�p��/�
�ѢT�>�0�Ɠߙg5��;��bގl0�me�j�*ĥy Wؽm��~u�Ҵ�����sH��������/e �=�̾B YH�wb�.�?�T,����BO-��w{�x�Z���������Z0�����m>՞X�
���ɖĻj��z��\�z��uZCb|���ϬA��~^�|��v�8�q�,��ٸ@�Ym)C��a�D��`_���>J~�@
>0�r�$ s������B�Q����ln�HDn=���?��OP+���PUZ
��NS����<N�o]y���ça~�����O<5� ��s5|ލH��5���c�.���k:�tQ�{����$	���d��^�H!v����fǻ� ��*���x��[����q�^�sK/�x���#�eg�i���Q
:@M5�݌��.�\(�Z_�]�a�n	:���3���f�5� 0��k'B*��U~5�H�S��͙�_�[|#n͡*/_�FDG�����H�h���`����@���++P�3(�1��ѽ])a�d�X���P���QΣ�|�#@��dNIA�0{y��s�Y`H(.~��~(�U���	�3"��C���7��H�*Cנ%g��c�s!�pc7Ń��r�����q�҄H��{�P�F���z=�Y

<}.1�=�� u��}x�xQ�N��8i��es�|m�3*�G��<J��HV޾P��삠3/�|i��گ�����<��[������.���
�"�մ:%�L$��^��#��_�]��7�TGO=�_�y_9�pj���j�j�I�=X�y,*Q8�!�;&6�5�.���p�V6߇�U�d�jj�h�g�%O:lO�r�^8�����9��D1c���]�_�;�V�P��ۀ(%8$`*#'^��b�N�
K�1� m��f~�tN9�6(ư���n��s�e��!21��H�J=�]��H.1�Qv���M�o�Dp��N�&�Dhء�ڃ�Mg^��(h(�$��YGg��g�MV�%��T~�<Kԓm���Y��0��~mH���*��}y��lC�z�Jh�9@�#m�!�w������?ƕ��<S�}���HHZ� �=#|2YN�-H%`Ϫ���;V�ݭ���ܥU1�K��IE��;�7.�TK�h�6$���3����C�5��������5Q�t�p6�n��}V�*'&��$���mq�,(�͆�֋�TO��m޸J����s6�qPI�M\X)�
��^s�_6�%�gU�Ӈ������L5E����*@X)�&��G��$X�U4oe����8(tom"�V�$蛲�|��-�ۍ~b��&�z9��̷�����X#*�38g�u�d1-�UP�i�� F�\BI��e+F��(�� �[k��t$��'�{B�B�����N��,�p��X���N�b���3�r�^#L��I�F]��XoS�(`G�'TDZBc�Z'n�ٔ� ~EJS@����2�hQ��7�&�N~2BF����|&��d�aµ��3��l`��+Y2��^EY��&]�}��j�/�(T��\B��0��,+	��,��`!�{[C�6ܘ6�����̛$��'d�b،��[(C���&q�c�Mc:S�p�(C�\�'��JF�b��?q�[�q��F�|N琊H��WNd�F \��Q��C�Q�؆�����mÚ?����q��ǣ�^�W�D��W��Y�&k�L9���I���~f`8�F#�57�.[ժ[��*f���_Q�	g�
�s�/�{C��M�w�}�6r��Hpe��ԥK�Cd��@?�֭� W�Gm00u�DO]�{ʎi���ޙ^�YԲ�0��ln�M�A�I
�q���]+2 3�>���.y�b,|�0��u$�[�M�I�1��A5~�E)�ġ)����Q��;�%��,�������'Tm�l�odߺI�F7\�t$�V�z"�!��<d��`K�S�Q[��8��"�A&�4\xZD���e���x��)�B�v��Oe��<*گ���R^e�R�S&!�DR]j����du!re�E�"���e�bx�:��H��)�sI��I�H/���-�+Lf�F�b�($�j�l��#��!IΙ�9�4[�!)=B�zm_b��b����7fXs4FP��H��[9|9���[5��e��Q�)��O�GbUF2�2)=�ܵu`���<t�=�~����=���Ʋ�ek�������[7T�.rܸ=��dq!'��H��{E���;������B w k��	�X�>�D:ǽε��s��"�$Q��n"�+����<�Il{�y�xg�I��A����20�����<��ƺP��%�G�<}�4�;J��6Z�f���:�=/[���\�!����ʰ�;����b���PQ����2d���3����,������#�ɹ����B��r��d�iUV����"ND��=��!O�J�<a�8lSG.r���j,���,0(�]f\�}�R�����w����Ier�(�l[�a���u4�܆�#�� b�7�tFBm�*ť&�p�22�w&��`�����͹�Y��sM=�"S��
�1A�V�T�?���<!X=���M $��p�;�k�/�&��4h�B��>�^�F���.A)�P�%Q��CD��p��q��W=������_�c�&	� ��+G؋�y�}�J�p�#t����ByL�!3Wo&��gB,�8s;�̽{���ɂ�3�'�=���3)d�ޖʊY
O1��'Z��H�jm�S��o�\�o����apH�����*ɲX@a+t��[(1ƞ����N�9ZJg�vK1�^�u���o�d���Z[�X \=������,"xr�+�-��B�6��������]Թ�-�c�i�,��e�x�@s@=禼�Iiѧ!v�${��F[�̶��5�����\�c�(C}o����8.���y���ͷh��o	L��iq��A�佝�z3�v�|vʊ�JϞ�s��2B��>���T�榓z�;��=!;5��Ë�j��=�d-�jr+U[L������`wV,��Q��<2��YB�u�5�u�J���cL��' ~Ɇ���Q��U�2���n��@g=��	K|���@�L]>I���L�vY�l�1<VV���~��K�����jU�I�ki��h�%hg���M�.��駷�;6
!������#3�l�do�McQ��D6�IE	��!q�9v��#7�I�7K�sםn+�0@xҧ�!4�u��}�j�\��M�&z��Э�"������Ľ���n3�VnY�?vrp
�A;��R�~i��}���C��	f���� ���=��`s�J0� ��Y�;	tbc.�r "�ـn�^�U��(��=��������E��!��ᴀ�}��G}|Y%΂^Z�@��}����"��J��[�y�k��L8�V[��
6�9Nx���oU�B���H>Q��\ç)C��0��[�b�I��6"�jgѕ��HcCD�YnǸ&���LGxVW<}I&�D��4d
�/S�П���?�_Šu������������B�ѹ�2r���F�4���9cQ�U�Q/�������Ş�Rm�(!\���p���ѣ������k���X�D�_lޮ��q������A��`��F��wɐ��������PBFK������ݬB�d\�z��n���Ҫ[7ޮ�sJ����F�������0s�BT����E�wN���J�zV=~�̷Nд�$}�jT�PVV��$�@�/�~r�[Yd�����ꅍ�����@)5Jy�N�109p4�:5uAQ��w��ZM�����Ѭ|;���!q��Vwesa������E3X�0��.U�+o��Jv�a����+�f���eR��|pn�Wt��u��u�MKxw��ZHG&]�#O<���f^�����=2@��\�	Y���z�
{j�5��u�k/#����"��+R�����H�{��c�*H���]��	w�"�<�l�E+��Vk��ky�@�3�z�cY�.��A��""b������ƈ�6�9vF�b�?�E���vp�­���Y�a4B"1��䧖�NT�����l��tΜw��z/�d#�H$'K��Gm��}R����_i�^������2�#�:VZ��^e?T^	D�ra�fo����B����M�ͯnAυ��XF�e���"�S�%k�"B�UZ�l���z+a�v��G�3e�йItT(����2������b�)T�XLI����v��~Τ���5+�=B�µ���ҟl�.߯Z;��d�U��>z�E��wf�f�?�S�p�V�~fW'��6�q����bxX6�K�/f�k�%�$fU
"N9�	��f��;��"��ΫB;D�*izar`�⚠Dv%f��Xjd_ǡZna5��f�F�b_r_��@[5T�����v̄|Bl�mB��>À�[U<��H�K8�V�+���٥I�D`F;�`�Z�a5	�t�,&ozb�wza�[��� cq�6����!��M�+�>&G��`��y���t�N�ô m�����:F�⅕m�d�W�S���/��W����qA��8H
XmT��0hā�<��؟��(mLZS�!f�a�4^���J�d�P
=d�K��|@M��N��^�ď�1���v��HP�jd���i}[�P��A���\���Ԗ�>_9��8�6qM	E�z�;���y��&׺ݯ��T���pv�B^+P }�Xh�%�y�9�Ȩ�'��)�-���߽]6�����������10��e��̾��-F��Q���ri��S������f��e�4�X6�3��%xi�w�>dװ�S�F�>���ä''.��G+�q��sP�xpG�������W(	0�1c�@cw�q���)�^9 I	�#]Ȩk���`�N&���g���W#[lOG��%�!D��
��pO�3�l�@0\)��0�t���wxQ�6���L��Z1�<�5���\��1O�U2o��+_�xQH�ك��W�������� �*.�8�([n��|Y���/���W0�C�Xl�:�)�%뽞��hw�b8z�7Ï�N�O	�a׽��j�P���r�
W WKm�<K���M���ʀ��E�`ϗK��_�y��W0Q���ƺn�؇�����!aY�l��)��ˑ֢آҨs�G�@2�D�'�NX���{�/���V��\Hq�9p��XwZn^�� c�D2�+��u�2Kj���H�	T����d0(D�ze�F�2�{�#��1F䠺5R	��^
�����H.�� ��Нej��:�_�����='3߷�xǉmR%m�H�0�%��j�q/���~��]ޢ�W���i�l�ι��&VX�V�o���F�L�r�Ҕ�Q�+��a��F�-�*�:�q���e����P=���Z{�Y�!gm�?����p��I�4����;���Z��i7`�G[N�����-/J`�N���]�U����_^��-`��������-��ײ��$9FMZtîB���|�5��A�W,�������L��2>����Ӡ0I�T
�[��pU&@v�"0�3��
c�"&�rc#�����v~�Aȣ:�L�*�_�I�Vo܇��r��%)�!�M��S&�c�`��:5�oL�!�W�"�,�`�!Q��kM2�Vl����'�ٽ��z6�ѭ�z�Uu��W�i�
����k����I��!��)��[����hfٝ*���.�A�8��Ac�Qܣq����,��� ��)��g�i��S��ib�窕�!oA>��\��妭�$�Lɣ�kJ�L�u�&�Ȫ�e�i���LUrv��̥7�*�Œ7\��5L�X�»dTVVJ��6�t�O.}�x����p�Ӓ�j�!rR�����x�������S��/A�y�"��7��`���pD�/
�G?
\��q��`��D\1N=,�\�>�H�j�����巙�&EQ�Lh;�Y�*�'=��l���Ð��F�et�N��r>/x���W6�oU�#���
ء#�y}����L��W�!�n���>Ƒ�~P=Z:��2���c~��}'�&�di��]u��f���]�$��E�h���/�&/�ܸs`ˆ�ۓ7�~y��i����^j� ��w��$��E9W�Y����8r�0�����Rqx��M
�kIl�VM������ �(���g#RGJ�*Ĵw��^�~j� 
����]�� ��QɈȻ�1�ձ�d`�|�]��	�Q�b�M>�e�E:=.ӝ4����蒯D][ή��x	�NA4��P�MG�/v*c��V�a����M8���-NB����]�����%^��m�C�l�4��λ��p[�,
H��]F��H�Y�u�z�{dgK[�>�+�a��A[�2O�i���N��#�p3���VM�Z���T�r�W: ku"�
eN4�!����8�΋ �K�����}���[�c~,uq{����^ʻ��jR[��&H�T)[�/�	�G��noC��GB�e8p"��.ō<�bG� W�f� l�CÜ�}��]��6��7W k�i�h,���g�����"�W�o=��c�|! ��1�b�Ւ�|��dõN�OE�B�n�؂=�:�P*-��Pǡ�v0�_�1�7FOv�~+m�6�k�:�m'�tZ�C�b�8Ngw0�0g.u��G�he鑏�;�I����f/eDr
� ���͡.��}�A��i���:��k��z���܂4K��q��M�^����xٙ������*a�mٺ�q*O�l��~1)���<,9 ��;p�i�:?����h0�ƫLĘ�Ta~�涄���I�G4>������к����v{^Z� V=i�&�Cә$�e9K�~���4/�5�F=�r�8�;�k�0!�L̈t������(pF%��a�f�ynX ��&�f�����)����P�C� �=��Qq�$D��@t��{^L�z�}������`p�aڇZf�����f<�(P�!V?c����)�����R z��jg�!��ߺ�e�h���A� ���������"��cW)> źmo��o1���"�n�Au�1n�`��[�Y���\^#�Đ����fPZE�4�!��`��%?�Kv� À�95ݵ>�Y��꿯1���{��U��V�Pcf����E�\ƠWw�-=�G��$��Z�;�O��!G�%�pL���y���~ulv5%A}�"'�;jm��I����U�������{y��.��נ���hM��ŧ
p\�#T���Z�c��Pȑ���4-�9*/�-dt<�n����8�Ӧ�G�5�޾,T4w�_��u�,�%���C�{�J�oC^�bW�)Un
������kL�S��	���J�`l�J��qѳ�>�$	q�-���`gD����Jl(�|X5KD^Źƅ�����!BA~�fh�;��%�A[�_�׏jG�!n�t�X�	D�K�i�D�7�hf�Z9΅�[o���_�ZM(\�|C��ա��@�83��]3
����cQ��R��cҢ%U�auyzBb��3t/MkЏ{�����R����E�y#2��p�S��8֙u��Pt��76=L��G��a[ʩ��M|G�e������2D:���b_�3���:W����B�`�ل�@��jϏ�_��gM�⺇U�K��<��d���Q�`��V���8�Q.t��?y���5����潌Ow�N=p\}���$u���MΉ�MU�~�P�ֈN|޻��N6r��������>���eb4��
uYo5+� �"l\p�_?
�ZF�/�̢��e�.�+/&@��+{ӯ�Q�������x8��y( �ä��'��4��VXpI�J�Y�+�A��{>��I���BN��:kW�-��܇y6=q�Z��dpp"&@��Yz�j���TXtf�|I��Y{�j�@/G��c��m�[YoCn��/���]\�,�86�O3��'�H8s�:��Ղ�[�.�Z��(n�oٙU��6�P���-,_xp1��E'��8+�E$�В+dٹ7�0'-j�M�
ir���k�O7�l��(A����Gǵ�S)&ۧ���hXFܙ�K�Ơ��1*yz�m�+m���^R�Lv��[�յZ�k�A�X���H�����&�w��He�8D�f�$K}wg�W����E���w��F�Z�o�4,%���[v����Nk}���o;!��VV�~�ݣ���Aܝ?K�����Y����U���@���ӽ�k��oD�y���k3�F��[��y΍νv�?�{c�`U=[��Z�Ʊ?msH/����������׹���ny�M����U��A�5;~k��W�k�s���Bt0���%#f�l��ڋ�+k���6U�̗n���Wa���\\� ?c>�/��3��Ff�p͐�Y&Jzcs�qo�*m!{�Q?�'V/���va;��U�v�0�c�"{�,N���["	�cҬ���_����yST?�"Y� B�I����O�ZՊ�,q�ԩ$i~�ᤆ����_�.�Yk�-����#2ŏ�]�X[�[���eL�[����*S�<Օ6����^X��O�'p1#�e4d�<�����1�p��ؗ#�����Ŭ�:��͸CEv�7��<p�=^��$wuva�-�Эe����dg�!�m0�=�(��M���yh��u ����D�LǢ}�5F����5ε�`]����ڰ���P�IZ��d�^G�ץ�k9\?�\�|qg��!��!���uT��3}�jt�"�q�2��=�/=��<�ё�~��A^Ɍ)��u{U�Z�+���P�Sj�7��^�:�!Oૃ�@�y�ȇ�#kǑlfF�o!j�up�w{�Z�[�aa�v�5]��yR�E=�����ؿ����P�A!���5��~�V>��jyM�AV��~�����/Uҝ�o�5C�P�f���87P����{�MT������K�mmQq�~G��p���AjI
m�������	�,v�����F�����|_m\F>��p-�� D�9�q�e��K���?�'7A�1���(��	�2�ܗ���M-I�76@����+̻�R��e�\�Υe��7al��P�5r ^���X�>��ilˆѹ5���ϵDQ�$�lb�k�v��܇a�/�����S�OY��$�ޢ����Z�ˎ���4E+N�fӰ3=HO'�q�x7���s�Y襎W#S�XY���ȯJr*l��U�;V�!	�P%�w���J�Z�g�y�RB�t�k�/\���� ��ω�CN��)��ěѯ�d9��p��ap����F[BN�)�h�Z��K%�E�� qQ �y�kxL�~Jye�r�ܫObpRu�����l%�I�e ��'$�%S	��}���蜣�0Q͒1S���s�P�%'�i�	�s �x����]7#A�FТ�W ��v�ǅ�o�nk��h3rM��+�-���ʌc�V���@�	�:�+9f�U�Iƣ�*(�XV���e}�>��P�eg��N�����8��9s;���l� ż��(���Q�[x�\�����m�Ǟ����g\�Lc��I�r}7���+��e﨟ڕf<���Ԗ�βU�r>a0�m�-?�a��R�	�B�S�8}G�4�&�U���4�hT� R�2���q��D@C�ܺ�R}åi�	�z�$W�\d3�2��O�0z�2虹��b&���L6��?�M���2P	�DYpwc����7�� <�����n��G'�
V��NB�ʊ�8�K8>�|Y�(�UʴE��[���"rP���J�M�W��e���̟P�q LO���8}�x0z0��*�iMH�N�2�w����>���܌l6'���ι�J�
�W3�t��g��xs-���ݺfHh��d��C�4Vz���Rn?@&*�u�����	$и7���øx
�����6�,!�+Lm\a_��= �$,s~�L/uo��kpݽ�m���c��j���PG���������v�^"�J�1P q�[� �������GM�B�� �T*c�秩b�]0���� �;nP����`{�@�g�w��[/(�y�-�8��Sb�����^*s`��a�(o�OJӒ��J�'����E4s��5pyYڷ��#��E��BS�o"`��,x��8�o�W;��ڡ�6Eo��#��pq�<�}0����7J��>+t�V1y�Q���U�lK�xh` ���TiӬ��[j�b�#����is�����S�F�����|A
�∐�^]��Ur���㢌(:�ls�;�A ��L��1�>��~�
d����@������SP_��^U�y@�e��B�����˚K��������{���?�ċ��ޣMI����ΝKG�	���cg�8C �Rċ�R�P��ɛa��t4P��6��R�0��9�p���/��π���]����`�;�W%�i�8�|�� b�����a��=�;ߧ�o$�=oy��~��M��iJE��������@�U�k�ut(��9����b ۅכL�'k�L7������P����%M�)h�Z� �	��@]�靥�ߗ��j�>���x�¸&�S�=$� ���������X��(�"AIt�q�H i���~@u~�7yC	�@��	��1-@i�T��l,�%_�ؘ�I�X��r>p?kZY��hZG�\�R�GxT���`K��kձ^���py¢��gW�7�Ѭg���Z��h�j� �7�=��V٧�σ{�%e2��<G}�KS)Y��� ����"�YϮ
A*�\DU�l��G������ �[�Pi��m�@\r��x���"�$ʇ�]Gg^Ge�G9��3%�5b���Q#:��A^�X�A5H�h����bJgM!'YA�iO�gw��u�t�< �\'��!�v������V\��$�����i����52E,v*��`:�%M�&��g��7s�K�����F�Vo�}JZF���"�7\ 
�J�"�׳8��\b��Ek�m/$�0���l����ג�lI�j���A��
_�\SaN�S�.����q���z��	��:�ҕF�v8�U�_^W����U�*nV�Ի�D������*i&_�bؖ�'c��������S�$c7DHf�t�<�G�E�=_0�י�q��7�V�z�1vI��'�]����c�Z$Cr�}�^,�4�e�?���"O+�e�,F���-s	A���PI�_�,�_}�����8�����9�i��_L����Yֹ���*���Ĕ,L�� ̨~gĬ&8�ͻ= ��մ��X��!֑��=a�{S�>���:����(R ��D�*�x/N�f��}jp=~�긞������ƬB�ǎ�.\�t�T�a��V��S{41ͧ����#��}��e��_�]�{u���%�S�:\�f]m�eڋy+����PH��>�����:cW j�}���P�v��x�$����[(�Du�z�S,)6�Vw"ύ2�� F6ܚ��Wb8¬�c�啓���Ԝ�*_!�z��ٓ�ܱ�A��k�2 Rf�����p0����̆u��>����m�����ޢ"4m��Q�sbNl^��� ���ne�*��_��[S�Uj��*R�ǎ��-��'���e�|���Qm^U`(<�d���{	��0Q�{JoN����n
S�y� �H'���B���@j���Q��)�^�t ��KQ��N&�Pg&��D'\ S��I���5.;�`�,��;f�x��:�+�j�q�[��7��hg��<w�Οsc,��ó[���0��6��N���a�e���Oh�و^`��5fg����P�ץ�.d]�A��G��qe� �Q]�~拕�E���%BI1�<8P�)��7i����wĎ��R1ιw�<�]z%/a��$00ƫ�4��l�N�q��������hu��d�XW6_k��I\������D	@l
g��iiW�v���o�Q�}݇H����V���bQK$f�i� v��%������(�gErŏ�w��̈���P����wBj��`�mb�(��D�� �K%�޳��N��p��T���LB��'�ꃘ�UP|I{�ׅpJ����*�l?vr`��n];G#�ï�����2hBă��qc���,��!��s.4Q~�$����ؽ�*m�ؘ�/iȮ�H(e�œ���#��2�s�a�0|�AฯQ�V�2g3��j^�E��J	�R�4�Mi9�ע�E	=����ǡ��D�㟅1���Z����m������,��_�b�[�K ���N��:��J#��ᴌS�4��멘��F��Rw�V4i*q�'�'�х�u����8�_���1P|13�ł>�[���s_�T��h�7J���4�����ړRh�Du__ۜJa���9� r�z7S ���70F?�0d�m�G(y�`�F������S?��Y�:��ZC��oʈ	B|-���0R�~�S�˿�T��2o����Y�����fS'�Ÿ`ӥ��)B�4�&qD������`�1Y���1���@8�Ï+�,;M
�̞�w��}OM;5����b;c��u�/��$4�lRm�	��Ko���`�S�j,њ�`H�},ֿk��-p|��F`d)	 y�<]�!wH�mn/� ��L�rt1�Z��'�A�ǐ�N]������?�M;.˾�e1���lC��J�Qm��RN��!ll�����L^LfU�:ޑ�x��Mq���7�ţ�x~{0<�c1�*��1�M������i��
�P`c������`��E�lú)k�U����D��(Ȋ�9G^'����bL�?m�h.)��8�6_e�p4Y��{�U-�Yi6ѷK>W�ˮ���9n�t�/��i�+֜i��x���m�zT�wl�00d�7�k������E����N���F�,B���%D>"�:ƶ���Q�������(@=�\�Q�&��`����F�~�\䍱}�L]G�F��҃o�C�`�֧s�Sm��լ�S�tH~���������Nm�9�qN�js���#Y\e*lBH�&��W����jap{qc��t�@��)��lH)p��:�8�D�ڊ�,�)�I�p�(7��&�ey%$��)��v��l�' 	�Jj� �K��	���{R�Q` �=G!;�I+���{�o��5i���!jm�.�s�	�wqm��$ONTu��^�2��$��� #.�e�u�����穼4<R/C��#�K�,N�@VyF��t ��#���t�_WtKu����S�)㳉=?_��*��������\ �$�
�Ҍf3� �1Z��q�S�8�e�.��}t����qlwI��*��e���+��a�#XD3 0w��fu,��煨O��EGL�FX��Cp!w&� �~���<��:|�@��k��߫����X�n���~�>�+Ae�s�1sW֠{q�G�J'/���b�G�;.��`�R��>8c�zΥX؛�l�� �K��-��F@e�ma{�O������#!z�b��y�[ҁ<���4*�V�9����.��9� �B9l4��N��&�(�.`�G�S+��O x}?���!��Z����0
�ݍ(��u���*m(����ms7Džj�?k��w U�v�:Zs�,_Ϯƫ�8,�r��2f����X�nˁ_z�K~��5�cl�1m�&����[-3�9)��!��zJ�g�VE�J�Yՠ��8�ApǌD-2[_W�?��E�g:m2�]h&��F��+�i����48�P�;�'�r;���6�O5�L�ze�ak�����٪"��9D�/^2�q�F8�?kL%���&�]����	 ���m�
�g��ru@��ɰY��U�^Nla�&��LMd��!��L�2Q��`e��*�708�~��u��c��~:ҝn������J���͢S��r@\�Nn�E�,�	Q<.��i͠#mBY������OSR�HQ��,�	�A� �1�����v�;�R3�- ���j�l �p�.���L�Tw����]7�Լ�[S!G��E6W\�7F�c�q���#�ƹi1��ƕ\Xq�r�М�#��s8V�+��T���o�@C��kZp�7�TPLq]1'A��$)�=�\3����8t���u�&��	=@�����{+m�<¹���/���l�V@�/c�ox�BC_�Q򘊙�ƢA�||���a���uE�E&1�T�;٨�\�Z+��۩��^�lOȷ�7��Ձz#�ۻn[_���,R؟	�@�6�24�oC*:��a�l��{ha������z�՜ԋ�F_^�y���G,�
�WWd�tСJҶ3���<>l���>��"N�=�v4�G��
��A\ʇ�qnLa�/�)�Lگ���5#��,ӁYf�_�-Q���Է��$J��.6-"Y�"���$�.����wzC]�4��_��ӰV�XS���l���Û�fջ��{۔�<@k=`[?VS7{J�*�\_���C(ɵGo���uJx��e�t�����r�e]ς~68�#jHI))�M�Cٓ��Ҳ�n�Į���V��7yT�g)-���譻K��i�;Ӗ=��r9���V1,��4��$�@���t��P|�:m�:��s^e�ƘmbQJȁ������AF�N1��"E����pSK�?�*[M�E;2U��E֘��	����oW��t�d(Nb=��kRg�{��G˘z���j��	�N���|��m}���a��*��w�8��4�o͸�V#�������LP����%)#wZ�#���+70*~�w��C  ��i�,>V~CD>�v:����v����:�7�����k�2�� �`yy��2I��+��E��}��t%�QfG Ze���t;�a�G�$�����gI/֫�6R���Vfo5��� �?��F-~�);�B��5��"ŗbǙ19�L�+Z��B!�@��>QTuk+K-�b�c��o��k�G�7j�4`�&�g"u#^ q�t��X�jx�f�9uLC���?�f�� n�[���$����[iwyK�3�3l��=�`i�E�a.ۼ5��"��.��2أ��S��a<�S=��W {��"�������eA��,�ce�U\��V�[+E*�m���x�9�N�;��\���P	k8fd9i�'ˑ��r}�rFO\��uOՊg�x�_��0��k%
��j��5e�Ͻ�����g�1,�@���ޘ�_�p��2������2<�7���vX���N� ��fY֍i*ۛ�jE~��݋��l|��a��)���P	>%;�����75�6�yM���%���N�_��A��FV?=@�G�C3�L�o$�>6
����/����E��~��<l��JW��Ṫ�����:kH���"!6�`��
�����+v��)w�@#zJ��5��i�G��ͬCy����j���>v��n=-�7+�g��U7�[�wW_�aE({����O�O�tJB�e�5͉،<0?PfΜ�߳��p�T/W��ao��a�`\:k!����j�RL%Rg��!�ڀ@�C�6!� V>��A�6�NG?��UD����;�?Ղ���ZY���Ia��~��n�t�3�U���F�Cz��z�����xQoq��"6=F��dB�-:D�i3�TL�~9C
ߩ�DR�v�������e��h3j�&�'¿u,�sh��d�d���P��7a�����p�X ��O�8]�C�$k.��F��6���J*�M�s�E?i�mg;K.uV�p��p!����r�	B�YT��_����&)Ep��������4i|��J�`]�ʸ��3WN�t��0����x%U�n^l�_���|�!��u=Hİ�>� �X3ꋿ)>'%!,�`���6��|�}*Uj��C�>}ߚ����<�'D^��`��(Ϊ[�|u�S�`2�&`m���g	���Ҷ�����1�-퀙�fPą��>p?�Oau���wG)�;K�a>�%�*�C��4��~oQQ���=ބ�Y.��v<c��C�v�j�H��p�6=�ВnT�+	%{B�#��s�<t�����{���|¯e�(8�S�Gl3�Ь�/�G���'�+��W��;*�;E�+Gvt����_��P�_�N�c"Y�,�hp4���
�E������_ћ�>��N����q����xPi��j��KQ��Z��\9�1!���.��H�>?���c����HY6���rS��L�t@N�'~����B�#�y'N& ����	�WW�nt���9�c�7»�* 	+Z��1k�o�  _��	3H��wwUZAP-)a�Zg�j���6��jF>HL �e����x���[�}�)yL_eo�/�~/������+�p�Hw���S�4�&j=|�!��`#(�t�N��<��M�1�&a*��bC�ȭ�4j%���@q���^�,x+ bS�ܷ��L1r>AVȿP���)��R:��a��#����kȢY�N���+s.�PԐP��ǎ��3����p���,1`�9ȣ`�q1������~J���ꙵ��Z�/r̝:"�4)�r��:�R��"�jy�6|��O�vAC�\�� �) `>B݋sȟo!˩5�L���KQr#񧛓2㪝\y�Q��^ÔT*���c��y�W�~(�o�/L�*��:S����*�,:�ld�l?��ӨW�p�;ᷳ#�u_����֧����D��L��j��T��Pr�#ٵ*�-5	ؿY?�Fe�b{�	�ɐ�-zU�[��G�A��=�	I��WU�H8ڡ���� ��Q���]�QI"h+A�"B��r�={f�B���������y��%ȸ� �ֲu(y�zM�	��L6=��\�9!0�'
A��x�΅�F��Lo����k.�Fo�EG��1+\���P�=����:!l�����+�Ț���K����d����\�\�W+0�$�TK�^n�g��6V�SiD�҈�����i�S�x�%!B��ez�bⷔ��3�����_�����&c��|zzEP�2Z�N;���c����棁�WC�,q�t���[�����,|��ٗ��W�)�4�J�`���TUe�xp���C�_����|�m�ݦ'p��#i��l��M������u�z0��@Ss={�T�w.�`*�fSeU)�����k��oj�m���ʨ��e�<�ǽk�ح�k��	s5u�F`7oŐ19��9�W���30|��4�+��V��Zȸ�U�p�/C�W�3/L1��?����=�yl5�>ʹW��/>qfnߩ�Z��d!���i��R��s0������I�?F�]L=�_��QC��l�S��Ykt)��1��V�ƃ�8���]�d-��m[/*�%JO'�x�Ɓ2��g���R�Pb��{��� ��5�+6������wਾΚ�]�R��=��$���H���{�z?���˪����n�'q�Z7�-$#��O;�r�j��o̦6�ܯWp�T��!	�E����͹iea�|@R��Yb:Z��멽���o�I���M�gך�-���J$���@����t��shO���G����ҟ�)U���4]3}�/�֗|/L�B�!T�tҞhzQ�h>��b��R�.}[�����g�=~�}|Ǔɧ�W� ��		<�x%��;\S��������D��As�翎�X�*���&��k��#�Ws/߹���,��_
-�g�MB��Edb��@���b�L{�8q0��A�w;u�=�~�`,J�4���� �G^�z�i�b�[��ey|\ooT>�\��N+m	)K-fC����rˇġc�������`�+48`��ӷ��4�
��K�5,pr�4�U؎{ �~�A@��ϥkƁ�^"k���\���π�N��{_�"��IB��F\�?n��՜����uST�l�G���3��nu�����Bd���������W0	<M���,۶���:(��H�{��r?�T���̅�]�$=}�NO#���y5��0ɜ ̞Vqٻ@�˥�8D�-қ�X�F�Fd�Ղ��C��c��d'*��"ι>������r�I�r�c�E%�4*&��I(꩟ka�\˙k%��I�C�G���"WFM��\V���m�񷏬4У�%,tr2� L6��:ֱ�UL}$KIQ �߹�]~`��G����I���x���|T�ˎ8e���N���O{�k�ʐd6goP	q�s�K+;�;�ǃ���n����a�W�Hj��g�6	0�;K`��cK��Eez�ۨv;�;3���,Ľ���k�	�8ȩ<+���-J4UR��%��؜���u�ۍ�S�U�����Ob��=bVR�����4z���1D�G�|���8���G���T��憕��K��VJ��?�����Xxzw/����������̲�}�.R�x(�G}_r�	��D=ϰ�J�-7��>�T����g*�H��/��8�6����[�����:M��g�̊}��D�z����S'���8�v�Yi*�����,N#��v/��ΐ���n6�!^pnh�O��#�\}�Ք<����J^��@/ܔ?v.��/+�cm���;4���%"9C�� ,���՗����?y�5X�C�B	z���7k�ɸE�E��*7>IR�ձ	�^����'8�K���ܦtV�T��6S]\Y̪N�=d$}��D���%�����ͬa��C�MT�?gn	��[�2��ҌL�b�^s��v钆b�0OSxޚ�&��ό���p${d���f�Y��đ��_�I�}�~@#���s���_&{�Rv_�l�]�
W�0BO�I��SmT���x��W��a�>X;ϭJ��:����G��*�k�"V��к%�j�ȶ�b\�y�c��H���Ѯamϖ�VV/�mG+���x5�ϐ�|~ƔXI�����_V��q�Xr�6p�O����(/r��n�Q�q�9=���`1���Yg�`J+"g�}<�~VV"ɤ�
<���	5��	���de���y��	e��#ZA�NP����i��<dwF�N�G�>�#-�c��`��e�֚�G�����N�[{����7 >ȀLA�
E�\FH����UB�]y	؂���a&�t��`�L�=�/{�%�+2�a��+��'�4�T��<]�`�Q�����Z���x�\�"@�D�@e������A��Mb!�q�P��ͻ��<���?�~�[`�.����8G�:"@��M�yN��)jY��R7�)�#�.�D����Ƅ�!�Ydq-x��de��<�yy�W�ԀM�J�B�l�}�9�ޔuC�e)���ԝzhe&��ǃ"�z{�� ���Ҫ���@���.��M���Ǫ���PK}������ �O/\�>꾣a��U�/a0�[�86�����M��)�p��Ѱ	;��cIg����z:_i��4�]�+N���*�}j��G�{�� W*��!�/��?+�(�>��ּz?�NΆ�韄mu`M0b���8���ͬ��G&�ս��R�0.��E}f���������G�[��΃����(��""�[ b]�FvH<�=$�r��] �������LW������[�f��)�J�D�'���w�:��7g�+e�L#^�@����3��Ue|��k�}U�>]I���*��ϭ��_:�����i�	����L:�ҎE��V�r�\-q�Vǿa��T���|� HӘJH�tn�:�J��i���~�nlT0Ҍiz)�ߦ��G��4%Ƀp.[FBe��#��B���X`	�^(缫o����ߥJ���kF�
hr����\�
&�PN��"�FY-aIę�wˌ��{�R�2q�&��o�9��0-��Ӂ�ǻ����Մ�����h��/�H��dK�)I����}Џ�{^\J�.���F��Yh.����>����Ҫ����]���ղ���B��8�4�]�).T�
�Dε��SH;b2��+�B�x���@G ��0҈�Ч&�z%@`�V�Ɛ�n	ox�7��9?J������2��?���v�dɗP�o�UfD���b�!�E
-��7z��ꮘ�����zțLg_r:?���S��3d,��ڢ�(���jf�=O���Qo�pP��"�.�Au��i�#P�,���!�*�}��=˔��w:R������M�X��y������%��AV�Q
m���D_�֍��sIZ����PH8R��j�g��Ot��7�S���N�{qЂ�?k\"�om"�a_�S2���w�
v��t�
W�Mc�a�
�cl�9��$ ������p/L헄m�Y"sL�{���A	6�Y��B��信���v�G���jn�.��
�pN���d�j�7�t-\C�bu�l�@�����JI��#W��Ϗh��S�1%���Ĥ�X�U��{E��I(�;��"���J����*�J���}*���z�x{��*��i�p@��ԡ5���,r�ܸ��\�z:_m��A�@�!s�	�,�m_�{X6�(���Ԇէ/?��I�19��*<.���`ʕVn��
!��)��wJZ�~��w5)kպqp���ܔ���\�)F�!plv}��	w�� ���"R�%j����J����]�to���\wD��Q���|iZE�w�K�����d�qV�(�8�p]ǭ�Ɛ:.��-�N���VW�L�K;��}(���(�4��{-�H�����]g���Ȑpp�O
5_���pLL��-�@8�>�G���� �a6�����*=��pG�!��b{�{���zH��Mt�H��m6	�R�|x�2S��o�,Z�j*�G���S��sѵ�WR�<GF1����$;�E(^ЋƑ?'L�h��n�Qy�����. �2��,�|i�	��Ca�{B��:�7&�lӻ=}!d�7�	~׋4�I�j�}��jW�AX
��N4��S)�뿲Kq>���\���L)=|%�>���P`�՛��� t���ʶ8-���o�z*^�O�S�ʮ���Ư����G�:[��IB�څ�5m�B���Ԧ�5	ӧއ�όp�G�_U��|�VRa"N]S F$�[�����7�r
-��n{��m��~��ޗ��zf�T�hBy6��ZY�mޯX�~G���֋���0o�N2�Eݺ�4p�!!r�]���k�C��0�+���!rkd�c���G��J��EW�z#Kv�7HIc+O��l7���ZW�f���˦��:�c�p�>�s������x;��'xʘ���n�(0נ��[ԣ��%\x�i����o��lUqLf�W	Ӊ{�����	�! y ���"�h��'���<�� �	��JE��9�e	I����mM9����搙��}^���߇{�(�{���&�z�W�Z����5��d,�&R�n���ru�#V9ׯ��F��1�]��ܚ�Cf�);,��@�H��U1�A`�Q�M���{�-�ƱG�B��Y�	��VЪ���D��2/aq�E"(�c!%���"�/OUt=�H0�;$�-�n���].q�w�&r���R8��c�N��kX��Z�`u�&��čH����nhx<i���E!SB�gg8��A��H���3+�-�7e����dI���{n��6���dR�9)R��.�;m`E�wN�+��G�W��G��.� r6jpx�,�x���v|��� �թ4����z}� �}sZ���l��K��X���2'�&^��L�B��$�J\eD��򀀻�G��̋�Ćh��\i1�H�U9v<'dG7��<���n]$k�Ⱥq4�8�6C���'���"0d�m�0s�,"������	��)˂&Xp�TG�/78siș��`�8�

�Y���P��[l�����|@B����p�u�7��>��/Uk�yH�늟������T�#��U��.��/�[�R+ָ���ʿ�}�u8�'��}7꣌��и��:J蹟쉪7�rB�8�5B,A�[�Q�������a/� 
�-�1��y��tC�+=�U�70L�Px����Z�����Z���)�7�7�t|?�:�����kW�ް��\��^A��y2�G�-�" 4gt7d�Q���\� �"�P�vmŨ��R$0�-�R�����r��I��-X^K0����s�	���12Ѹ*|`���U�`VO��@������%�R��~������s��J�Ħ���t&l�X�M�㮜k@c�:ۃ����9�_�h����c�����9����a����:l��Q�c�_z'��lE��r4��Q'���xA���3��������R�w6.�^7vai��Wf��2P�1���}�	�ٳ�Š>���е�/R����ǣ���P2
�"�ҐhC��?$֘��S��a{}~Bk�ҁ����h�+q��D�Au��A�.
TG ���oy�o`�zM��%c]�$�f4�bO�\]�śP�ϒ��~h��`��[��\�'N3�Ѳ+�vn=�N�Jw���od�fP�_�.G-�!N5�S.���y�q��2Z�%L���b�l{FL��W��g﹏��Z���� �9����5��4�Rҝ��R���z{Z�� z��).���lT^�4I�e���*�Nؿ ��:�TP�
��n�6����*_������Cp��"��h�d�
c��& ��^%�!=6M)��='���R�1����3�RG��7��x��'�4�erX����#�iL�,�db���5)���n o4ŗ�?��hh7��b�@S����tTЫ�������s�)?��e��Ɠ��q�[Z�ι�R|�_Y�){ы'5K_�t!�%GBc�v�>����-��E�Z����8���������D뚊w��x>
�xy����� =��nҖ� �N��ƻxQ�M ���դ�-n˲}3��c1U9���<e���.�l1HqŖ���}�D�O:�ܿ *������>	f�c�Ƌy�`,2����-�/�|�&�B{�bs+ӹYc��:�$�RJ��̿�y��$��uңx�ǖ[,Lޥm��YiqH����2�^��%U!�bX���*)=�8vlb�9Rl�jR�z&�S��F2��Tr	^j��z���sx2��;E�����7�e����'"*r�Iu�-��75^���t��ì���|?"��SZ+p[W�.h�&���X0���)ԯ��]E�5��?-(equk.��2�_~^v��
[*�=t� T1�ʶkt�$�n2H��Մ���p�)ӆ�TL�@�c�Ӝ�a`-���ɦ����G4X�s�g�"fQb������n׳Luy+�	��;&�Ӓx��L;Q�GwU?bH��F�u�p�IG�]ypqQW�3����Zґ<�$f瓱~XɊ���55?�諯�п��h���E�/�ʓ4U�����p���S��ͷBƉL-�G��ͯ6��|>�]��l*�(s���A�Tfu�:�m�{$:0z�7�iV|g�tw�ؽ���l�lH��=�AuY)�W>R�S5���,V;�V��|&�-��ߠ�	���R?O:�B*P)ަ�i*@ٕ�U!9�K[��ˠ��Zǂ.�
��t�e!k�8���1j!>,�QY���Lu5�EXk��j����Ź�Sp�oXm�텏��3����U�f �l���%!��Mm�b�V� ���c������9������.{��n�]����
�ϑ�b��~��K���R�[�lE6a�������B/�Ȑo�q�h�̟��$�n�yuؖ�U�
�+� ےy�n;!N���̩JS����O�Վ�wg�[���n���O.�+WW�̤r�q��GT�)�o�'��*���O}��ʵ@�g��`@B�Nwfiͅ2n���H@����x{u����E>|��_��h_ߞ��F�"�Q*6�Ö�Ӏ�����2��S4̎�������|`�O��N91L��K�s�e�WxC�ݨ�%�s^�Tڻ�<X{5���i�{t�E� ��o8�ܖ$�O�:k1�ohҙM#U�	i�]���Mp(�|�3�j�`���
l|F���4!�/�xˋ.��Wm�K��Z�7�.�}�R�D�PO�:�dx����AC�%�J�=¼��0�2�G��v�c�4{zn��� ��]��V��_� Bc
Xܡ��q%��!���
���uU~Wp�q����m��B:巋"�֬E$�G��[��@� "���լ,î�S�D{���#���0[�f�����*�'������|�����dS���:�p��Ӎ+�����H�M7��s��Ihw�*�C2�*�Zp�h�d�����;��Ӈ��_����+�Խ�ع����G�dd��[Ёy̐�W=}�q]\�g�&�{Q#�ɨt`�nu�'�o!K���F��Fb�1٦TE�!?CO��߻'��':�����V�M��ڳ*ժ�)1/YV�4!L�O�����%�zp�In�4�x���܂�
��s��D&����R�xk�Z��.��\����[%�a�N*�~�Y��ܳ��
����G���5= �B�NϺ�Wv�"ȁ�{`(5����DD{�{J��MW�-�74��*�6
�'l[� �Ә|��Q�!��*���ؙ�����i+F9����벓=9����-+A�,���\";�ڍ�Y����U��&�`��
�oz�G�X^Y���5���2�o���q�n��n+��h����԰E��-	�@�d�A��e�.|<�B8
#���} �-ą^���XP����I�9��T!��#�C�A<4���7�#�s{L$&ߢ������ ���U�	��#c�F0���k��ZX��w��H�>q�3l���% ?rU���Co]V�	~"""����&֍�^c#�k�ż�FJ ,�
�n=�!}�I8���??�Ĕ�"��{��I��8N��ʽ#�(A�O1W�-F9����Pck�.��&�e�V�K�@tN�t��,���K:�ھ���թ��.4w�r�A��("z\μ��ey=�{ 	n�f�sf�N)����8x��ВA��}��.4�}�r-k��7G�vW#<W�PؽewD,s��z�J�䣟���N�hq9��qY뤡D'���5>l�"K��t���|c󘦼*�o�ZK9�Y��IY�@�DB�ޚr�dҕ�x�r��0U7@-�Հ���օ)V�|�U�q��N�ׇ�pڦ��B��q��G+��8���=�׀�.L�P�a��UF�"&W�>4|�ٱ�	�#�2�;��0)F�kEN�C�J�N��)�X$��������۟�r�#��ґz�x.阠�X]%F�vQ������+�߆&;�ZY����37�7Z��ٍ�t��n�`���[U��w�Q�g��D�fc^{��ҥ/�?1�ϣ��U�'�qR)CF�������M
<��#�!��]�吼W��PW�����_�|@�	�Y�0K'5��Sm��
\�{��|�,�\��2Pm�g�*gX��%�`��Y�!����j��HrV:�����6 �|\���d�r=�xS���Y��	p�Uʟ���~��rP؊T�	��e��t>���-�V&�H�
��;q�I	�������@���q�͌��-le��d�bnt�Pj��RZ_��P�:�{u$��~�SAZ9�JO	m��ǰ���yo=��!:�J�tq�f��Y�QQM']Q:R$�ȞGJ����~�Ƽ��\cex.�:����ՉD$��as� �}�a���6�~���6���h9��&���@����
@P���-@��(?eD�YO~$Y�4�1�s{�K1h�3Z�s�DI0��]K���~`��i�Bo�=�
��kO�n
��$���*���!͈���&�/m�77_�It�.�F��[3����H�<Z��<���s_����B�`�dċ<�;�kD9f`.������	��;�����r�Lu��>�.��5���PU��c��v�9B�J��[�w�X�plZ��%h�v�f���Ҟ(t����TV��*A��ia�^ٽL��%�QUA�y�\a��CdN����,I�(�:�ģ��7���Wq��ȭ���tx��Dqє�B(f��i��r�?*ι�f6,Y1�C��'�Ӎ'�ٙJ�W-����_�Lh���$��|��?B��x�+NW�j�4k�]J�� Ad�����ꈽƫ�L��;�Lwȗ�	.*�r�'���N8�� �ċ۶T�!��59|: P ע�>>ަ�(��Vd�\�0�N��Z�����f���>\�վ0�E�z��a�s
F6���O^I��S�*�����G� �7j���>7e���fx��}�=���(*N��O��=�.��d)˙���r"��.sd�E|e��MQq<'���2���}��׸OH$���pd�G� ?�b�'� �����dߧ����d!����@s>!m�N_G7������:�S�g-Qu)��s�_���˭�>]��7B���ϛ�݅��@��tD�B�`�C�]��U����hOP^��f;��@\U7�ǝr-�Ed��%@�� �%^�-C�a+���A�3���zL#;��=3�ɟ��6��XxT�y r�|�i�	^J�~|�>���AT�}�5K�l;�ԫ�'O�
B [���P2bR�vƛt}�1�W����KZ��56-ɡ�'6�{,���X��w8:$4+�����zs��?�aq�=3�R�3���ð�r�r�r �v�X�#�iO6	*dU��� �a^�R�{ k�G�۶��lA8R�8?o��M�.*��6�֥	v��[�\�) �Va@mDŶ ^���W��M�9�e��k���Ɲ~|�>{2��P�2��a���ts�7H�ɝu��b)��G1�ma��;��N7{��S����N�l��ǤG�C+ؒV�i�p��k����v�O?��X6�uM�=d�Rw�J���p3��-!���(����S[����(y�o�Ѽ&ǎ�@Ym�~��'/2"���_UۢI^)��5��f� �OF`>h��ب���r��_;���BO'��7�SeL�n����O��DI�"�@Ju.����8UNy<�c%�U��{ɞ/Ie��F8��+���jN�VD"�{��޽�=� i��=� ^3JM�6�����vg��)Hǥi��e�_��"��#��!�(V����U3��@L}$T����#�I�Z��ܮI�~��
�/���.�L>�+�ٚi�	� e�Jr>��6�_*�~�OiE�R���NM_s,��8��]y$�G�!�6�\�S��Y�N|n�y^�`+�f��ӦB�E{1R%]��{�t/�^@hy��DnɂT��_��~��ҳ��J�9x��;��+��^!2���O��,�*%M����L����O����$<�uWYQ���7)B �֡����qqO���냓8p�lJq��4���>ks��TA�?�@8z�M�����wKkp��<���{@]��Ʀ@s�m�j���U�ӓ�HD�n�QJp$#���H����b�6�}���kD[RZWU��t�(�f���?�k�j�hE~������T��J�	X���M~��6��U�Ĉ1E�<	��_Վ�s�$���f��[�y�;n��O]��|/$u�������U�ҡ����z��%-mt�~5A��?���(s�}�^�Hb
���8tw�v@6���R���-O��yRyF`g��~�jZ����f"��IJ�!)�H���
�r4��:����Vf�C/W�����i-S�b��^L|�x]zqblc_���ធ<{��Τ���sP&�/��` �\�I�GfP�3�,,��O�ls�c��w�1��{XZ3'r�hi:s��V��^���2�/o����'�0�ܷ��jb��)K�=����N��YGǎ'�%�cOk�����፻Ġ��D&���q�, c�d�L�ڜ���S*��'�4��'4y�
6"B�^�Z��n"�b��ݯ`���=0��d�a��|	S$��[�.�>��q����Y��V���?���V�ZD�A'w �ȓ�̲����+N��Y�B#C|!�U+�EGY��b�7]y�>U���~�3���H���l�څ��χ��\��X��t\��[�KX%�&�r�%8�	*ya�m��Z�k|G�����6gG������$��"E�ję3���w��N�feny�SMQ�{�>~�𹢇gJ�I�E��M&�Dq�ǥ�Ja����y� 騢����B���z�d,��{�@e�lK*w������!���6�J�B8���(?��/Eݖ�%_S(��P��������~��L� oe5!��Aq��~�N	�MVy��"�ܧ��v!��d��ֆ"͟�A�s3���LW�\%�-�ǒ����M�Iz&@h�珞��Y%�@��