��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��:W�~�_�c�hɝv���hX�z��,'>﬚qì3���
-�x���\��6�b̃��~��lqm���e�k����]͠@�% ��4��C��n���+��&LhD�~�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�P�;�{��3�OT����n/\�@���V�F�	G�V��]� z�`t���y[q����a2��;��i�t��,-��1�� pz�jI;�"<i����#{���<�G�N�3�mŬ�#�:����(U-6��K��j�'��Y�}'	T�(L��ag�=���`m%5�|Nq�Y;�:�|���Q@Y遀 ץ1X�q��j�%|�H�����la�IKA�w��H�=0z �y���Ʀ#��au��#E*��p��c��>�$0i8Y=�P���(�]hϽ�8��1���y���*��V]�t����śvrs�C�l��Z:*B�G2�2�̒8y�����
'R��9]D�"����)@����A���xu�G���z^��Z�+�)���I�v��R����^� ���QJt�rG�@[��Ó�3�}C�	]�ڄ�0M�)��2�l2-�r$�L�Q�7'�qL�����Vj��ϻ���2��s8؇I8& ���4�&FW���!�Q��%ǌ���b~��<]&����`V`H�J��J���a �o�cp�2m0��OjpPx���қ��_��E����p#��c��5��42����!�δ�XJAl,��lvֈ��5[��஘}�쫓��.T��˓*o�SM�է�p��&Ue��ƊBA46�J�x�c)������f4W}�B��,��
a㓌��t5�<�57���?�,&��	 �3	j��Y�+�5'���"�K���n��F+�|J��E��%��#.����|%ا��;�\���ۧ5-A��x�jp���z��"�7�r��d����DJ�4�^��d�c8d"���仹R�c*�)�)B"��kc��f�0�y7An��}���3�]W{�m�`���V���JK��=�5�6�l �}X��t��1���L�렖0��\�:��d��/���S�:�g��Y�G�"�u^c}I*��}�����Ū���hL�$��wz��Y)N�I�^�Grh�hX/���<��>ʬA�v�$���O�W-o�n2�̋��cܒ$�u��H�����v��f(LL���p�0��"�6>�u��{^U�_T˹�\u������.��9;��sZό~�rX�T�o����UJ~�T{����k���'a{��d`�)!ʮ�<����[��&��7Ep����*�uiP&b�km��A-e���I��ƶ������x�"�Q�
,��`r`1���)���Yh	�rB����
����Xv�?�C�*�+�eb��*R��X���_ʄ ��p��w��������P��}��BH'9�<w�4�ɂ�P����^�lj��9w�р� r��`�_�=1���5^eL:(��C'n�*!��;�_= G��ȹ��%�`�N��<����I~����p��b���>GC+Yr��	�3����8ãY�%~2�/�� S����[�v�V����6��_�^*� ����zD��D�6ϸ{�=\��v)�XZ3�f�$iǥ�2*�0S�6ZC��O����e�v���Q��qWu_�t�U��$̼���~��]�C#��Q�8`!Ԕ�/�s�=���W��4�Hձ�3;�U$l_���絸��7���<����Χ��OT��óK�W�`�R�����e��!B��/�lBk5Gp�2g��b�j�S�5����靡�/ ��g"�u��!`<�Qp��L��PM�O���W-���S��hO˸nu�����_*C�ɽ�T��h�زP��tؕ�1�a�	�}�
/�� ��ٚ����mv��U�¿�V3��"u�����_6��X���ϯ>����S��QsUt�]�x�-T܂ghd���k'(��bF�N���"'*gB����=�C�3����K��X�a=:�	���UM:?O6�%�e�4�Gc��O����O-88��\��@�4�QONp(��1g���'	������,�}Ze�w'�C��"5��}̉[�Q3�[��:j�����K*�R�\����Y����q�{��×��!���o����8�X����o��>�s��9��0jb�U�^���ƭ��<Gc;RB�&�2���̓$֜�M����G>@Z�g�SS�[)�~4��$ڑ��B~���ۖ4|�'DZ��x��b���ylccv��Ou�-�Q9�D2 㾷cJ�U�I6��D����(�^��k�������./���tE����(T2�Ԋ������Cّ��:R�R\�[m�ӿKh���6��1��=sTW;�C�e�e�3l�������9�����a\�>ܕ]�-�����)�"۹sWvm��KY�PRg���R�@Æj8�_|��F��#K���W�i�=��$u� ~��5
jg��$74��|�*���������kÅr��	)d!%��h�1��B;am�����oّTL �w#��'Me���1�y��`��[=�XE<K������k�dm����:�2�`Ju��#��I��6K��`��j�mߗ�03��RE���s�7�)�SjxSȅ��W!������_�����ϺP��L�J��׶�6w|
:����ZaH�#��B{e������ؿ�|ط1���aҖ�L׀.%���R��M_����1&�(����f���5��Tl�Z���_�
�SH� ���n`���YuX&8�b��Vu�ݸ�����?0�t�0g���J��*
���+
�;�����ppR70��@b� �TZMY.�����=�2�Ф��e�A?��0��9ж�Ďc�+�g�DQ6~�sI�"
ij5��/k3SZ3��^�Ő�hȵ1f��9]Z��θ!����8���?�z�I�oD*�D�;3
L�g�����%�zS�3W�ك#�x3�JM� �\�zqG��Q�覲��wd-"��m=�LM�xGT�e��{���X\T�L��&,�F�^y~�tr՗���ѕ?��A��H7���fo�v�y�e1�Z�v�Q�?��0�����l�8r&���k�JՎ����3������^ !P�K��Ҹ^F�?7�3{�^�)��O���-�MmL�ƺ�#W�Kv� KT~r��F�#���NV*7�Հ��M�zd,0��i�r��#�P��x$؋�t��x�~w	�~��q�/��U��F�n?�P�)�K ��-{����^Gv �%_�|j����A��*R)���c�8�x��4����O�#�H�#�"�%:��6�����h��!��hމJ�U.!w[��]>��� w��1|���1De'1�.&�^@�/�^�&8��1g����	w��z��������ͧ�צ�����������hP�`�+F�d&��T��cEv�.����2Q�2��{x���/��R�ķ԰
g�	6-� O �����0��� b+�#���W�d��t�u��	[�(JF�`q}92E��
���np��?d�JVi\h��@v�{5kH�	ا�yH�&�&9r�G �Z�f�`l��Mǅ����^��(�:\�)�@gݯ�d/@p�St젏�u:.��)��M�.e���Y�"i�赵T�nI�j�i�R�J�op��.�	J*�3u��68\�0~���k����x�,R�[�[N������K����� 5S��!�3�?G�Z���!������3���NytH}/Y;�N�����cC˙�D��VEVg���+Z�u�8��ˇj�l��:��l��4&����##K�}�%�L����J]fc���ÀH��W��13VO1��Ǭ��$����"�j+�����B���t>?�����x��s�H��h�a"Oˆ�`�W��n[|M����}�,W&z��p���s��:�A�dv>!�k�+�ovR7}���n>�+���[�Y����0��>�
���7rM~+�ݫ��l�i�PL��cX�*��fe%����-�Z�Rj�E+ր4-I�)�����y��j����zD ��!������ƌ�O�Μ�w�W��TCK�3FX��B�Qڠ6��)���e�MQ�H#��v��d|�o<�l�.�0���.f���'�y<:�ͧ&��U���O��a���|��i��r�*���᳆S��L����n�ΘCݕ��wb
����Ȱþ�t1
%ġ۔�(˙q�rN�)?��ҖM5���0F#��b3�Q5�o���E�J{�#��B̍�E�6R��]�t��1Ep�J�`�w��z�\�(nHR�K��?Wr�0%ZA�:��FY0�0���|.�S���ϸ	�Ϧ�`g��X,���9o2P-�f�>ɞ�NPVD��Z$R�@���J��ل���Ωyּ����@vP�Kso@����?j7�y�2HK+'��꣤��Ud{�#�]��<��3ۊP=v����^�0PU��5�� .�X�*�mA�������%4��TU~�w���y��mv���Z�U�.x��!�0D/�N�ݏ��V���pwb��;��tѝ��	C@"T\���N�rt���B�/N�=k]�@W|��Q&�7{��Mn�[��# 1�ǜ��a��?�z=<��:u�Mʴ}"�!�WE��эQ9jW�OA�+Dk� ƭx�<���ʻ�m.I7�+��gk�uʂw�X����0B��������9��LNȀe|w;� ;?Z��\�8h�T�����ꣾ��Bq���W P�r��[����/+��G��\�z�
��H뙸�s�W!y��n�΢�u��.�
�_�Π��6�����rsPXc���꧖y4���/�bW�C\��:�sFMK�r�ߓ9� ;�$d�j��2a���WB�*��G,���Ȣ<����M�n�m�R�<��̦��h&a���>��	���%Fܾ��9U
k�U�!�)])�M>��]�K蕃�E(�1W]C���Ԑ	�R3n���"��!��� �����q�p��*�A���E�fRYImavJ�DV	��"���lU!�R�9Z@�x����Um��޴~�?-��0����W�|�r@V�ijG<�-�+�i��Y�<��">"�����i�fCc �"�jd���L��cG?���oVlE�&�!��ˋ69�rc����5:)_����� ���F�&q�K}���X�H��Z���Ƣ?d��n� �1IO�b�X��d-��&@���t�����p71���F�0i��e/����mwB�8t���0M�IZ�T�����t�?�n������ёD��S�s�4��p0X��B1*�k���!�z_����ț{8�a�5�$֕"���EM�K����
�V)��}wGŘ	�vnz�
�8�o?�΀��( oFA]Ui_18�k^�}](����]
O/�-Fe������9�/��7�#������7�����w�e�A��菼�z��9��x\x1�8�d���Q�(E5#QSX�	� �;g@0��1R<�_c��B�dsN979��	E�RnP�ߨ�w�¹�6��[K[��@Yzދ��;�ݣ���BO��E��,���7��T�2#���g����_F|2��d��M�f9C�a�A��;V�<��5�9[Σ(�⥗����c�;
n=��#�Z:�a>t�3Q���b�:�,{��{w�� q\l��:PAo����E_"��6g�,y�>�KLfLw"S��&����}���}t=�w����*X4n%~O;���&jm��6�H �H�e���N�قN��`2�sNR	��9���p�LT�ֿj0Z��F� �Ð$�y�����#z|?AI��t�դ9+��<��h�Z�8g�{H�)��%3V���+���әT�q�c���
�3���P�߶Y9�؀^��
�F�:�O3�?pt�0�Zr�6�� ���+� �g�w�[8��$�z�EJ�u�������ҤW1���@����������+w�v��	��_���󬯥~��[D�|fG��[W�dQ��Lp݅D���I�kefl	(���jؾ�Z��}v)�A�V�ҧv�l˱!$�	6M�\����b�J�,�l�$�^�s�`p\��̑E{�mF�o�~�%�3?��j�G�b_}�u��x�}�E�!��n��y���F�#��4N��y�^�u�8�����&�{��\~(iTaX�\��r!�#��mHh6���TU���0��~O��&��$�/��:�l ȩI��|'�E/���z"T<|��m��.�|�#����|�Ơ��e�O����YM4�#�ԍ��C���,��̠�$}Z6ă0��@M,��$ƈ1�2"��+!���X���.��Գ{�C7��?�5E��<=�}�+z��F���,��p?��:輓5��#�/�NF�1�HP_/R�����
�}B)�>@܇;��h0�[��w֟k����$��R��lq��|���ʃǘ���A5?{%���!��)���z�V���T���b��7Q}~F�[�3%�w�vqIP���6����'\1#oCB��J:�ӈ�L��UO0싞���'^�1���{J���m��G�%��p����-1۷Q|2�� � ��� �8<p��������!��|�+Mk,���E�3c��\j�sib�Ɓ{��`ۿ$��d�Q���oE��b�b^i~��%R�XO���*�-��бZ=�G�n�m�by�c+�����'��h!5��J�����)[s��f�GO���:��4<�9�[Ërw�79���>�a���i��������<�q
ٻ&Q�vC8�@����6�?e,%]N?�ɲ��K஌�n�HO�8��[����@g����z����Ӭ��/�a�3!��K�4G�-àt�����Q2�{k�T��(M0�[Կ-�e��p�J7驴GNi( 8W������u�iפ+01�xX�e1��ygR�K�Y�	$U�s�}��P�8� ��2�f5aw�3q0FC��_Sq�]vx�a<l���o��7\�񻲁�s�RT59q��*hNFo� �
�z�X��0}�:���&�ʰ��5��;�(3Ori��C�񊇈"��UG'�Оe��wON'%)���˖��LN�����+��=�)������U_0qd0��\�	��`Y�/K����מC'M��l�"37k�����V�B�?��`��B"�������X�jT�����SK>Z:�5�yiq60���6��PcZN�7Y�-�a(�G%�J��ӳ~ݡ�z����v���z!	�e���(Ҷ���Z�=8YW��߹�3Q]PY�4b�������{;4|n��)�Gi���L��b�*��L���M�Ae�pP3�6�]	H%��u����G蔔ħ͆�;�s��l�h�  L2S�i@˄Q�)x�9�7հ�z\	��Ud�8@��W�q_c�w �	��;��=�Q�9��Al�R�Q�ȟ����l�M6�v��1� /���T'_��$����Z�����A��-��H�Je���gB�zia�j�t��}���2��c�+ޕ�Qf ��$�����d,~�Yk��w��Nԫ��BTT� §�c\�	ѿ��8<����N�G�TsѷԎ0�f�-�Qz�7�]�h���U���3�x#��&N�����vì)A-��
0Z�M=����馟Ek��&�-�����}n%ԵЕ(qv{��>m%�?R����\�7�B����>�8bׁ�Y�M*"���ޓ��Gm�B� b��gW�"��<����	�A������mb���/]h�<+򇫿i�5|mk���_=ˏ�Uko/l\�Ŧ,e^08SReJ9qZ:t�</'{�UeBW��5�UW]A�d�v�V�ɿxv5uKfO������ �Pj��������{�Ў�`#��>���c���%P�O-3�,U�B0De�]%�'��J-S��3��V<�L�½��X��:�c�f�Ȼ({k],����T�zJ���T�����ۯ7��$��Sc�,���h|iUp~.���	Z�S�Br20a'��/��?nq�doab:s��
����^QO�9�=��O���F/�i���&�$�i�Cp$�Z�2|>S�&���2������j{����g&2��?��pas��g�'�^oR���Ԏo2�R%�r�{��^6L��8��E��Fn:� a�	�#�g�Ho��$��*^NO��m�?�~X�!��B����'�=R�9�����Q�<V���Bd��%�W�\,�+$n��FIP�|�%aX�9㺲�8ȳsF�s�Y�=s����+_���q�4�M�$���e��������Q�ԏ��A�O��+�z�ZLҐ[�h�s|�sP������ t��KJ��5��#�b��X���kCC6A&ό���VG�I��'�/]v�f�J�F��w�sI����݀�eT5�����4�6�_ⲥ��93�(�6��+�{�(�Q�
;��r�@K�f�D:��XG2��K���m�,�����.�+�9�)>-��Q�2��R�K���k	J	@K����
����J�bC�3� �(�-�G�Y^(�V�d-=�)ǂ�8qː�|I���J\���Z���`DÃ��O��I3+���*>���j�y�Ps�a��������MvY�
Ĵ�9�ϴ9�*��X�
�<b���g)�rP)�l��-�Խ3ґ,�ӱ��3�}�ul{b���aku�G`��ΎKHB���
�;G��;��-{��0X��2�*�'K�{�gm ��� �F�����>h�:�e4�[�����9Ͽ�/�oܠM�f�f���^`dJ/�ڦ�t�4�I[����NFK��䟶lmwh�`c��z��$�e�� y��#�?�j�eA!l�P��A���ǔ'�8���I�o�zo��p��]����Up5��r�X{�AF���)֔ �U�^�����m `a��"4WR��Z �4KO�{�nؤ��e�.5�o�J��
�jZ�]~$�b+|��+�ÿ˸̧'��B�l��f��
S�z� ~"��2�F��M��l�P�Z�"rTN��b3�]�/	_-����������;�]�%4��K�
�e��70���9;��Z��a�Gĳ�k���;n�c<0*����^ȕE@� �]���c�0`�u�:zE'*.og?�yX뉣~r���84��q��˳���2XBꬔ�:f�����9������L�\"y`���������x�,�`��2�6]~^9�C���A�/JH�>�k��~�Y��S7��E犰n���d�6vzB���ݞ���[����:O�F�5{ �"V7E�ۖ�N�Eq`]4ڷ̜GL[\Ⱥ�6�7��b��4Yrk*u���'����=g�8Yd7��W_�H�	�p�����Q�P�Yj2�s����d�2Ѭ��ø����huQɱ�D_u��'��s'���r��2r���:ov�g�&U���s��`��QǖF8}hb���$��_�;���(cW�Bm"J���u�������x�X�K�颒�'d���(�����o�0�!�;�uY$��6�Hʫ�E/=�[��=fs,g0��4�ZW�Mjg�v�T�~&H���� j��$i�efq�Q�~*�Iف�{5b���㸃M��&\�~l7�\x=���6�c�7T�Y2Gs�J��Ӷ��*e a 4��l(v'��
��OY͒�7�Qu��>H�!�(��M2�79�z������������Bx����1Q[��t�B*Ӻٯ"�wvΨ���kj�Ɯ�Q>R��֭`��>wf��A`�"J�:.+���7�c���?�c�_���2;rP��kX-n�叭�;��.F�Hӂ',�*�����]��q�,-��C8 Oe=�A��}7�	`��a|����Ƽ�X���=Z<�L��O' �3P�Ʌ��9���#�N����"����9�2=���?g@�@�X쟲vu��!H�D�	�.$���xk��Լ��vg�I#������h�UK�$X�eqY=�ϵ%^\[Z橇˭����?�����%P�S���	���ϖ�%.�&���r][�C����Et"����8x$�N(2RBA�_P�54�;���;N��@��cHׁ׵i�y���N��es&y��Ӻ��E����c���LI�T︸/:�"�@9����R�Y͑W�)�#0�|EbqS�_�0vYYb6g�8��_����W��(C�N�Ee���n����S4J�Bq��tݔ�Y>mKe���R �f������@ę���֘IN�\�`W��a+^�3�}��Y��%�_�E�L��.'�6K�GAH3�<S����8�J��kc&�(�:կ׍i^CI5�DF_�Z6��Q_�����;����ń�T2�q���ƥ�z��U�;��j�;�k���*5;�>��K�?:l���H�6&�4��l��`уx[jy�d���u��T�,!i�ЏU��̧����!�ָ����g��ޭ���Ҋ1�I>ٮ��P�FE�P8O5-�#���]`�{��M%�?J+�^J�_p�����@��a��P�K��K��:h!*�n+����q���jRfi玽쪏}f�\s
�Fۆ:bF�>���X@B�۩�'4ae��mB�K6C�:�2�1�Ӕ�d2S��Hے6������qD��"d���A6^	����ƐN��-�I���������y/�Ƭ�}��<�qCi�ħ6V�j�e�x8-
C�����c��1�^�zLG}ym2�g���`JJO����È�!6�wu�
6����K�P8��h�݌}�(�\ߑϹ� ��j}:����̶�$����`���ҫ��79�n��8�J�R��q�X�ԧ�I�����m�v�����b���]��{��G ��_�C)�}Z���V�K���>��c�	�vh��L��^�q�|��b�����
"�I5����[�	5�!80����$��ӳ& r;�GX>�
�8o��D���|)܇~��lʟ�;�w���zþ���ʫ�D����so,<�t+h�u"~�+P}
]��v#�Y��Pj�/JyI�-:5-��%�'�[]?0�J�deF(]���A&���ƕ��;{IJ�T�O�b�����T���S4�P';�u�(�+�P+E}�dv�v�������r�o��w��"�:V�c�&�'m��3wsx��Xi��s$��B�}-�?m�vv-�$M�,�q^�\l,�F̯��+�Ay!F1�}���5ȼY���5!�|�b�AY��.G�:�b��$IHܬ]�8��'@�k�2��e���͵um�X;�w��@=ÂΈˎH�枧S�a}���
�Z4	�(� S+�Ӝ���:;�J�^L�W�a@f0����./�G���o��)��c-�8�=x��Z&d'�?v���s��z��E��x�z��*/�����0XH�q��=>�I�K����7ɚ^U���=��_�������N�=x��u���Φ.��U$}�jN�7���2��u��_D���\ⷫ&�п���?���Ĥ��W���c��~��>dґ?9[�N��9~�_/�9�d�����x���Yj"���Kg�<��tR�����Y�z��m[[b���~�u\ۣ7�sLwD ͦ	ꙸ�"�U3��<�o�L��l��q�&ëTV:S�g�*�tpN]��G�STk�y �fm�f:��+��r������z��x�fki��^��,�:�#[��XY�����G/�@n[��ul��[hg^~	
�@��T�^-9`|�:%*�Qv���ƫ����wF����'�e�L���2�Љ;V�6l�Z���I���{32��������L$�*��ڎߤ6xNu���۠�a���U�y����e◖���Y(?�/����/<z���~�Ca�#�aߕl=�@ش����r��H�7ga�i�#v��+�W��_�3�P0X_��͠Ӡ�&`�;���� �Oby��Co?�Ɯ��&�"0og[�=w�.g��@�ᩎ�`�!Tbf��͉n�F�nڃ��ˍ����l�jShl��y��;�
�wfS�r�hp��<�������>�E�ߓ\�����)]u�
,����v���O��5���С7ߨ�^z91-�%d$L�C�O���1m;7�c}G���l"J���y�>aG���p��C�*C��� ���{R�V�y�f��p����S���k$B��}�����J�B��Sp(k���$�7()}���A�=��ۑ��KG�������څqݖ��Q<�2e%��[�g�Ȏ54%fZ�w���H���C�@f��;�bf��LI���\$��0�I�^��.l�������Si�fz�H����65��r��`�ʙx8/:����ry������l��2ůR#hɜq��t�oW���u��~��ZVYu��>�ՅN�N��q�R}���T�e���	���N{�R]����juD���q���eT5��>�V�����*�&��D������]1',�DZ�>�������4�������i�U1�	#�s� ����tó���ja��m�U⳽!��e�^����a�*�B�vls�G�L��yܱ�?�Otn>roɒU��땁���z,�Q|k�f���$��yMt�x��q�9׌A�C����~��?�`r��q��8AǶtCߵ�V:�hi��3��St��A?h�	�㉙�4,�L_Â�|�1��p��	��Hо�%�B�������_�]����\����5~������R��E$�=��>������!]Un��,׊�Kd����[h"��+��$�k>oda�P7�-ܒ���GM�lB�S�������~''���y���,��vr!>U#32t�x6<?��c��NgA��f���	������V��c����	�LM{���Ggj}��xb��hY��� �j�d���~�]%�L���-��������R ����v�ͣ����x���C���cS���;�=	�E����r&��`���>ϐ����y��ڑ�)%T�.�(}?����� �m�x�9��cN�v�W��*)�|)�}/W��(����ȹp�^
����h}�8�e��v�\�z6a �Uc�b/P)*���m��h�� �^�2��K(�C�hr�(��.�&7�̿8�D�Y~'�l�ٔ@S+�{�\��@r�MDԵG7kc�$6_��F³c��1�ݤ^�}�'&�Y��6�k���������B#`�#�b��r�tP�mo�����Q��n*���>��ki��S���ƅE,��ڢ�LŴ�7{�IV&g�oI�=��+�Ӟ)��[�8�����־*~'�պt���`�F�!4�]��"��3��qUO�b�K����LN,����vF�ʷ8��r9fB�dr�hgi�S3��I����hM�ȗ�'��9��Y�e)�DD�=V�A�E���_��q#�H�@Ól�|HN,1i0"8=`�!n�	�.�&F�KT��Q�U��>(4`0~"��>�{���D-��ӷgG��R��Qs�~n�������a��s��e��GKcT?MJ� ���/���#7��j2���M�-h��;Pdo��$]( ����V1���� ��^&��80�\��2�i1'�dt�j�a�|�;K�A�yZ�u�y�S��qŏ�,r��*c�T	��U��q��d�Lm ��Y��m�t����2�7�����ꢻk1���6֤]%E�-T]n��yE�r�?�&(�+��D�p�G^�����[�G�1IĞ�YoD�q�z� !9U�e�d׻��d�o31+[4�-E�؅l�oL$��O}D�!���������m�׏a�=����k�7T{Ȳ	1��f@�Fҁ����4j�x��zӿ���* t4��Ov�3�O�����Cğ��pτ�a���ӊ_4�=���a*R3�z���6���T�α�V�l�UA�!0NBo�v�$����e�T�{f��4�(���*���$^.�G9C㉸�y�o4%������a=в�#d�tY"�����[wp��r�v��*S^U�G"��7���'�~�z�)s�y�"�_/Zd?��@�O�!��s�`���B�B����M����AI1���Gó��x�h1�R���9 v�o1x�d�
V�D|���dun�Ut�Y��R�[or���P�s@P�/!��y@������p����"L��ڝ�*K����Qػ�!��
�yL�� ��Ǎ|�k'"�m�{�!|�X�Vwa���
RV�7�3��汚a[�{F#�2�y�X���1k��b�C�dIؾY!{�#���z�����t?�l�\� s�ɢ����� _�<v�N-� ��~������8��G�U.�j�E�5�K�Z�e.�\��^�����3�!t+�4�S�q�-{h���Xj`��ø�LR=o`m��B�L�Į����^<Ų�|~�"�jp��r�葵����e��cTA��QU+�^��)�P�)I���<��w��b
��P@�n1tӑ�,!p�8HfwC���b�]4�w�Q9R1�F�0��D�?i��sS��"ںܔ=w�Ɔ<г���'��GV__@�e�c}����a=�o8�k�<��pi�J���^C���W�V��vU+�u�C3����zq����)�J�G���Mt�a4��Pm=��oR!΂�cu���U�\h�6��L�{�]������C��W��-��!������-6��&~2����<1� )��=IC�z��;���7�ݡ��\cH�=K��sxu�l��&�t��zGg�/z�`�a�m�z���-3�zs�$4;��`;�b�i�%1�
����Ƶ�EvZ *�=�+ �β���_�'�*�f� Zs�p�=�`���e���g��VN-<�%Wjw�hwz;
833h�B���!�]iC��r=���9J×A���F-�k�Uk����"�r�wL�ħ�ʦ�"%O�8�T�խ�E�_��\�;��=>����Y�4AL��zԫ�Z2Ts�}r��'邝Y�j%f�sA:Q�P���L����o��y�RL�QL�-����%��d}4\}�L�)��xE�5o����<�3X:��Ss
����|��j=@7�0`B�C��5�+sW�=��_� �^��cZJ=o�t.�eB < ��0��Z`d�4��8�ŇA��8�}����	�v���[J�@���xԞr��:�nO��C#�ߠ���<�,���ExƑX�&OG���^�+5�}h�Z�S��m��PDc �TJ�H���v����љ��Ŝ��bތ�Z��`>,�[�!����:� �^9j�k�@8i%�(ە����k��	��ôvHC�j��������m؀}̔�<�]qQ�mi��CK�T�V����`�C��+�n��$u�"^x.����H](���x��~4�S��|'v\�Vx`�{��D����&\�&�'\�Ef�'9s��@dퟡ.q�2�<ra3 ,)D�4�g(t�?te�Ex0��?+H�SJ��oTz�*U���]��!�pAz�3� �3��U� k��h��:��w7���s�$D�cɟ�\�����͑�'��YpȸzS12^��������<��n��N�{]�����M�_�1=(��P�I��ŀ��F4_$�x3��F�C���߁X����s�q��ܨ��@َư�G>U��P�a�^J���uZF�*`rd�@��}�u#ļ$L�7Q*ڛ&��0~^��1��Ȏ��~"su����(8�z�V�JJ-9x]���q� ^��.��o��$C��`���DFUQX�Elt�������G �|�����㛍 ��t�������v�k:�T����Q%�۽����ٚ黑�*v�䡍���'2@�S�YS��\�����|��1I;��Pǳ*�m38y�k�(7^��?��I��<�=�b��>�6��eJ���� پ[�]I������[^�9s�}�὘O؀fҿ������NX�43���~0i } �B@m��9�*b�BD�}��}f��W�9-a��QV��umu�u�ʟQDb߂��"Wgk�d��w��r�l�s��rؘ�=����(�Q�N�K"�05��3+��;xNh�o�r�,6����0�QH���^d[}e&,�ۊ�!M ��ш�e��4���2ޏ�V ���#��h�G�O�Pw��(۲��F^
CR�"��Ә������'��6�UQ�5\ru�d<ț7)�ϰ?A��!��(�] {�%���h#IuNqS�x�.!PΎ�PP���i"B�ܛV.L;�<[�1�}C&BJ�B�5Rl����)�" �G���Lb�5�Q�8fi]Ԣ!\�+C��o�t��կ��:$�A�EIW��l&e�*�����a�db���j��.�*)Pz&�6�y#��V��W�>�1��+ �B��i�$-- ��p��jB�0	/2B��+2j�&���@3�p$5.�
��]v>��S�  �]5�S�����|%oA���``��gp%Yt� '�ڎp�u���v��?�������7��AvU�q鴜#4(��\�.Zҳ�x����*����h��j��\pw�����7�<(�L��D���!π��`$,;��w�M� ]^�CSX�T��!��Xp���	Ş�ݟ��5�<�ު�A�����y��(�I�O�h(�z�qK6Rou|b@6�QX�-A��ao{k�ET�}�\zA�n�sD����9�񥪃恉��D,����`#b3�����6�?^��*�D�܁�[�pc��/�;�y��;K�����IJ��2�����`f����=�9 K$,6�v�3��`lq��P)pU"߰�@L�*����${>��f�`�Ie�1޳sz�qt���-����=��XT�;FƘY� x���@Ev��*�l��ۤ_��T��=?D-ȸ��S��F��	sUiU�v�,d?i�|�D�˯�|vKB>�;�����P�J�!���V���л!�4�1���>c~���:GnY����ٳ�w�|~ℭ�}B��l��Y��iAV}��_0�G�����V���^E�Ԧ�z��@&��*���QB�~\r�cV��+k���n�IF�����TQ�]�gS�.�ܯ�D�I{�yp��������Q�b�,r��<��p;��iq#Q���T���a\_R�{�gJw��:�̦�A8�5h�ŋ	�7��<�Ԭw�o@�@� {.�\�@t+I(XL��`Kb�%}[L�K�?�]��VStBԶ�/�I��  �q���'�W=[a�� ��w�Z:]�,��郳� �T�)')���G���L��[q�;mA�0��Y��I�#�`;�1�gtV�B�|�R�]/�R6A�"�9�/�E�����w���t�C_�m��������s"}�H�z��M�~@��EØ,�0A�"j�����c�·/g��s5�@�C�*�]M�BkN�C��VF5RUᴪ.믇��z@h��f�#�?h݊0�)-��_�668I
�
j������]��_N���Q{���
b�>�F%�z-�t��@�ԕ	��d��E5I���7Xhb�Qn[��mhnQõ+�?�~Q�޹�m� ���f)���}���������#���AR������Q&����cD��T�r��r��&|�,��ʺ#�]��j��5ӆg�7���ô����-?{'�AA����x%hhv�!C�߃�6� m���Uz����D�V���$e��v���݄�]$i��H�v�f�yhف�-n��-�Nn�����'���U�&#��.�N܀��h9=qBi}j��C�y��s	}C�U��A�œ��#��EI�U� 0M����O����l>��t(9�F6Fm��.,&x�r�0ύ;V�q��[F6�Eq���@i� �AΫ�[]��")��a��	%3Q�����jH���h��Y�6qA�T!�3�6]�Rr�¹�����R��/ǩ\��������Pf�	�h�yXI�K��4��w@c��дfc�G6�b�<׼�-%�"W�i"��t�Y�е�v�`�cHO%�S8C΍z>�������������Be'��C+m6X���n�� 6��<&��勢2����{��e"�`���e���2E��}��f�C(i�允*橙���h7y~<�P_[DOO�E�>�1��x�K�>��W�DlW��#p�"�J�������l�A��!�Tn\i#,؎�x�j!��1�L;Ĭ���`MFw�bwNd`�XzV"����L2n���J"#�ul����)����0����n��qɔ��5	�=}��}F�kI�A���juZPr�D�e �e��-�nm-���}���~�e�c���?��+�;��b`\-?DP[���S7��]�7���Ʉ�i�܃��W�_��w ��1K��,k烬	�T�N,L%�MNN�t�_*�^A�g� U58����ާ��?�W2U��Z�1�v)�;�0���=��$��	��f�S�3|�M�¿v�A?�[W�v���V��\���,���#���6�޷�l��u���N��K=
m���Rw��-3�=��R�;�r�c��Z. �������Q����������v�-Uv�7�/�e�>�ڄ/�K�����^��Q�������p���VNM��Z���v�����I�KKhh�D����S]a<�:��#>g�oJ�g��W�־Q��	�a:���ҶN
��B��`,~%8m��a"&�sk0���U��Ğ�w�J��c:�'��t�:�o����e�c���D`��'�QT՘Wr܄���M��?̓�E��rRs7{����g�!H1�'.-�Qdr"qV����|$Cn��˵y��02ق��ʵ�:��񾱉�ɤ,F=tV�F�PM$g��H�'}N�=1WjЖ�xWS�Տ��Y�"�����bM%/ol	����M���!4��1/�/~�-H��;}�m/�Z�ٓ~z��-]:4<�J
 �@4��{t�=Z9��c�E8�v�"
�qć��<��gAϯG$Q{D�gd��ת�V>ײq�n�
�!`8����Պ%�".���O5��
b��`�Qv�ZJ�Y4�)iX�����F�,�Α�8��1��cl�T�4ŷ�^w���ǣ���.�t��X���!�Ao�Hތ�e�)�|c��k�U#bN�� ��""S�U��7e�z`	�kM�6i�����w0�l����HzD��J���"���6��Ra�����W��
���3�ZG��c�32-[n�����A��0Dl��{��w�ݕe�E���X:@�^�=��#C�4LN�|G��4k�0E2�{%@�}�5���cĬ��g��4��� pu�u�;pA��t�h�M����-`,�V�v��Y"x�+Wz��_'6���4z{+�M1�z[��%v���T�L�eF!U��)ځ��!��LA��u���C1���g!D�oU���u#��
��t���}7���'_�S���p@o�P{G4���'�Ls��C8�d�$��.&�@��'���~N��%����8�y�*�s�}�śCT!p؈��n��lAz�cO^Ι4���(V���%(Q���3
���&��� V;�k�ט���γ���z�E��=�\T~�C6>w�W��|�#|je�ȝ.���ɦ�P���1޾���9U瀈u�_��P�vUr{��e��\f颐~#k�-����d�����gy��F~��({B��{$��u����-C�uL�}%ji��m�ˢ�{����t�]ZW8�N�p�e�[OF���d�Uj��J�/�X���!�T�̣6U�L��K6z=���"[当��v$��� �c�O�����2�Զ�mL�i� f��Y��I�FMJkb�Z�S�N�U�\B\ۀ��v��C#V
����Ӑ����F��R�d��v��.�7�y�ًT����6@Q�Wk(���J��S�ͯ�G��#1|,������~�2���@�%ӽp;��I��7���	˹;�*j6��p�T{�-�T��p�e�A�K��.�?`e�U�?�g��%y4n�9SD�hD^QМTu*�����[=��#���K��S�ɇ�1�2��B��d�F�8��S���`$�俩�܅���	�བ0�������ٚ"�v,54�*��#~���`�{�c/�w�'j�>0���S��I��d���ޣ]�f�z�l�ҪY�$*�
�%�ɶ����� .�We2��M�k�3э#��k��e#�Ơt��E�\�-�K�7�̨���?V��c٭9cې2$�irKL,���!I F����@�H���Ig�K�>�X�p'�$7��g��O:����|OU����2S#�5u��oh^���������W���0�^��p��p�K�2d�Giu�F/!nD���	4��NAG ?'׃�χ��k2������n�.��,="����v��	��}P��]�R�_�>���y��:�z��%o�;/+]-���=7z��b>�:L��tZڝB9�jO�/$>E���B���[-:�LK�\�Pz0S�3�<f�ڢ�a�DU�r�
uH&Ψ�1,����C���d�� c�R�7�6��]���LJ����\yx��� ��d�y������̤F���5��fpg��x��9�7�mN�Q�������ܱD��7�R/�2Ҵ1Q����_�ig�`e(��o.W ��`f��<p�"�����'�.g��&�'�|�e2O ��Tv��L�H���`�X�Q� �S;��T�DGK�#���җr�5�Q�ңa����S��MJu���*	�^��@;2�yj�'d��D&��������9b��ݨ�0F��V&n&�5c»I�2��J��!��b�*p��)��rՋq0�t�Ih��pA�	�[�~���o�lf� R#����R�cQ2�3Y�"�r��
�����aIlBL�B_�����u�Zx�,Pŷy�*�u��	|��ǯ��&f6�h�v@���f�<�B��O�=f�|��N��Tj�����0�5�|w����t�[�ZA$�\C ���Xw�NխN��,=
,��5�{l������r�Ɖc�����>��0��:۲��������ｲ��ʑ.T����&Ax�1���}}T���|�[��P���]*D'y����.��³��\|o�uW.5�==�qC�FQ��$&���{C������Hj���*�����������QP�9r�R?]��̴NYvʥ�2G������$��|�B�
�z_F� f�Fja�����-o�d�ֺU�M8(���aEA�[B��-	|�S�P)��K1+�5��bV���9�-v�@m���w�,�?�qS�'t����c���nSd�X�^Ij��)a�i�cf	/��i	��眑~g����Q��L����0ʃ&ˣ��O2*����=�{���KFuh3l���2��|7���51�e��('�����v�0���Y�1����w��#�|ES�C\�m���0G���!Ĥ3��vuG�E4�����O�}��J���65�-g��ɀ��'�/F�WR�6���K���۴ș��~��;+_�R*O�QOYa�*P��
��D��D�|��-�T
�BWA�~(�Q���%������-�t�~���������Yxh��Y[�g�Hr4�௄k�K%eY!�V,+Q�}G�'�a}���{X�i�\�U
*_P���if}���HPϡ3��V��}����a�D��n��&���� .E$fY�y����9,}r����b	�xs���]^�r��V��WW�!L���P�sw�qD&�4��3v��Y 7��O�;�6��w��Z4zqHY	���T��H"�:�T1�,����}���Ɇ%�2��Y����9Ja��#�T+��ŋH(�_�Zj�:bq�ߓ�x��(����V3I�q�`0��Г��ֹ�-����J�è/N�|��bɋ�hz��)�����'K*C:�S	�TZu��T��!)!Z�D�^�T�I)h:�+�C�zk�����&�*l��Ă^����9�P�E�|�<�x9m����$�F@�	
�ʼ��+}9"�
�jM^�v��j��o���ι�/)b����W ��N�ft�M���57�_9�D\�~����l׺�v���#(fx����I�fJ�:�M˞t���R8k��"5��Hji�uE9j6�f+@�܉z����p�	meX�_���e,�<P'����A�����U��8(W�^�M��=N+�!�O�$�e� Y��|T;�;x�Zn1�O@��Ed��>>�d&�i�2��Z�[���~��k�p��(z����I���8�4ꡒ�yg:~�������i���F�#�\�H�B���^�%�!��K�&=fk6������A�.�hC�J���T���74KJ��SaڀH"b�l����_HF�4=�*ê�F63n���k
4(���:�3�E� ��X$�?H�;�&�N�&2��U�@�+�F��~pr���7@G�����)�Q��������7����.>�F*̵�q5���	JE�4C*���JəRZ�(2��5��r��5�a�������_�H�}�
�6����"ȧWvI�����666�bj<�	���:��P���}W�U,d[tM8���^t�J&(*�����SjGǢ��&t�W�si0	4�X�|��0�{F|9QU3z��8�,�x������;��nP�h�pҟ��e������9KT]@1k���H�s[)��wj�K��^X�|������8yb�<�Y��U|f&E��]E4�0ɣΘ�ʢ��E1���OW��&���A��G�;��;���%/P���S�E��5��$Ol����QVÔ�~m���SKM�Ea%����Ĕ�C�5��*�)��Q�o���ĺ��CT)�B����\8�BǤ),t�ۃ�Ͻ�����d�g|*z+
�"dE�D@�͆|�*�B����kZ��U~?^ ^�>�c1�6A�ŭ�����B���K��N�^k��]{|�]�]g��+9F�8��ّ�u(� ��������3�d����3((�D����x*_1��0�e�"G�{
y�B��n�V�eשO��� 3z���	�����ՙ����=��ަ� i�R`A�5h����Mr���udb4F�Ϭ���'���١�8�)#�c=�_.���/��;̜�u�D��$y���],7�x�b�c�"�=<�S��!�a��0Qj���g����ʘ�NԤ'T�"�-Ap�>�q�s��x�*���G�y>g�ʄl��� �u]��3W�J�}iW7�'�.L�O����p�����V?�Y�6B�{n��3	*W��dY1#��@�lq<�Z<�S;��!$O�׾��-L��O�t-5�I��x0I�mj(�"����`�Q:~����	�"��J
[��N>̅'q��(�yU����:Ql�٩�V��~�1���R��T���)��)��]�J��^N>H��M>5�d���k95�Y�&�J������6;�F�c�_EA5w���$ҷ�NWp��'WH�|<L� 5T�d���i��xs����?<ڶ<,Y�χ�+/��N�&�����+#T3�,��]��w�d���{������W���+w��m8o��1��[^6����8���Mib�]���N���m������7#s<ۜϸ1p�j�\&�Mi�
Ӳ�ul��P���`���	�;�<�&C��Sh�wKk����o���|��&��FpT����/H��3�o.�����ݴ���Ր=|AaK�סݑ�"�������PJ��N'�(8���]���=����^��i�}o^�)�� =];�g�ن㦜j�_��Hvd�y�aƻ�i,t��~���G�10�ܥ�)9�;0FP���.�?| �u�S������[a�4bA�>��D	�`�7%K�͆�;"0h�"�q�mp6zr�|K����/7ԭa�@�Z���
�c���a!|̌�5��y@3��D>2$�Tdi�0��NhFgYx���{8D4C{��5t���n:�=A��gq!�+<'��E9��X_�"��2��u�u�/_�o?�챼V;��S��{\��3�HQu�yf��)�Xrz��N�R�&�"
pM;�-�؏���y���s�o�LffB��
��	�D�V��cS{z�7 �|���GGg�@S�#��b��]g.�S�\IC�Y�v��a��,D��uz$�;�.%A�k��+w�u�Y܂P\�)HG{9�68iX��6��"MN �q�a`P�=�=��C�֡aT ��R�5k�ewn%(�t�M�B�M��\���!����$�o����cx��/���1⑹�/�i���rs���ڸ��ށ��:���j�Uo��"����j}�*��I�ܘ���<=�H��K�X��ג_w#�,>_��¶b);#�(&�p�X_�������ʼ]j���)ux��
�|؂8u_I�@��g�c�Q�?�y�t������#�v��� �mT����ʢ+�2��������H����84�������F]-v�5���~��J�1Či�8]���]P&\��	]���m��ۡ�N�Xu���m��T���q�X������b�sǬU��[̨��������Zű�5 ���P�d��.�(���(��t��Iw�#Bh���!F'���M�/�.^e���1�3��b}����G
�{�� �<)��
����u���Nt��N3�r�+�����o��d5l��G߹�q�f����B��p�����Qł����z�\�$��1�0��'���k*	���ց�~ ,������ڞsvwW/&1�F���Mmp��)�Q����D^�F�y�u�,����H�T��.��n���@�ԝ�=�2��D����_��/-hY
6�[{L�h�9�79�I��4���&-͔}G��<������A���A���A^�N����M��r��20_��P�@������c����f�[x��6m����r�ϰq4�řQ=�nͮ,�X��X����W��c<Ԗ�[ ���R�!q}��h��Y}�j�f�s��
҆��[�Z ��=�L;�#����*�dKd�'���إ%��T8�
�h��^�-�A	QS	�������(X��u4�
������og�D[���p��k��2�I8��w�d���F������(����$a�r�0�������%��',��uS|��va��2Tw�8NP���n:�6~5���H%p��������ݵ?I�R��. ����Q<8�פ�DwYM��]�٨ظ�rY�£�{J�������
��!7 �E	)dp/��R��U�%A*��p��� î+��^F�J2�������y�C�Q'�&\��[5�TŌ�0��,�v�g-����au�����1YcS�3�2�L�<lnW���E1�9�m�H�e@�,]�E�0��t٪��x�l���^ջy��Y7<Z��-Ca��K���@D-Y)�6��s#N_��a&"Q+�{E��"�nf�8_ߎ	�#��4��0T�����c�L7��rA@�А��܊���Y4n��2���gN�Kg��Nպ?E۝���B���ID��W� ��i��^�7��ኩ~�D�LK(��̚~
X�S��{t�g-9�#�L�:e��]����o?�UeL��V{n^���41d+bm��膆�Ҍ���L���r�6��4GL��E���uin��&�?�����$8�=la~Z*��9�B��Pl�)k5t_����+����/���:��4~3!
w(�a#{�*��ܒ���hlȫ��*������ q�vGGC���� -�\S�Cڅ]PB[�d��wJ��\�F�.5���~�*q��m�@��\ق^�~� FQ,?^��q;�4S�yNAؒ�\��&D�����y7� i��Ey���C���[�Jqe2rL���T�Æa'&���`'D�.��HQ��}YG�bS��v<�7�c:���*�E���
+6=�'�� �xې�J(����p��f�4m��R�Y�`?<#n�N�)�)� �(-�¬ �D�)*d�����Ӧ\[U��#��]����!̴����0���)����&n�`,�������5{�-2ZWk|�yʑ}5� PE�`����[v�"B�т�e�:m���qLm��-D:#F[�����(ӻ��M���s���Ҟ�{?�=��a#4H�w���	pಋ+�#���1
�j�Xw;=:���G��|=��!��7��L���k�+���1�^���{[%]�=Bw�<円I���t��z��S�)���f�-��'�]|���]�S`�\@�1�fZ1�_;�J>{��̯Ֆ g�6�i�����{���?<�A�j���<)>M\���-d��p@�L��;/ &H��� ����W#|XH�R
�����V�K�9F��t%B�n�y��Ǌߗ~��C��u��M��M^|�lf��_3R�/q���):zј�e�����m) ��Z�6|�>���S"�f	�'Z���P����zh�� �]u���G�q�sЩ^��ip�>�E���ٔ��W��*F�P��9%G��o�z-�\��1/��l�¿As��Z�z%S����\�E!h��W��P�v6����Q��N#+�"(�|\�үA6?�)���9Sݚ�墤�	-66r�I��Ѓ�Zc+2�N�h��o����=;6ް�n粔��X)�	#iLi /��d�Fϱ1 )ơ�W2x��2�G�6��)��C��a/�ʢ�U�	�6*�׀gW�X�ֻ�v2)|/��5���}r��N�N[��qe� ����M�;6Fc�'}#�F^`z���9M��Z�=0ثQ��;�|�R��4��� 1�܇!����)'��j��kR0Ã�(�U(I8b9��?���z>m�Ƅ��7Ը��ž��X�<~�	6��Կ�Хd���t��j��#J����{V u"��-9���������Pu¥/����(s�.@qb��Wo{����1t��s*��|p���Tгd���f^����|G~W+F�~�����%����-k�>�p�E �et�9Z�� t�Xn��=��~�C Y5�>�(1�/����_X����-p�IeJ��-Q6��EK���H�ߒ���HWHY��<��6��E>���+�k>�WBd����eյ�DL�{z*�e XZ���,�l�e�I!�0i�|1�v��E�
%�u%�ͧM��(@���{Z��x�S���e�	7��Ë�|��PF��t���X���H<�!b�
4��I+!n5����xD�Ɂ�ω��<c�pv_W�ey��㏺�C�ԒH	
��J�2���g#�q)Ǫ�je���\Py���ٶ3
�8�;ڍ������O��*�O���;�"r٠H#n7�!VߦƏ4���7@p���J�E5��Q��7��q�2�s/I�Ӵ�v� :��B�Ѫ�J\��fB�1rl�! ������]NzJ~�l��~���ы�~!���Ǣ��	��҄���<G���4��*�����q{耾���s�2s[�Z3:Q������-L�A�/��7Q�1��u��]�����Յ�[6t��ğ�Nc��.]ʧ<dʜ*���.�k�y"b�a��;�?�\�[IԍXu̫*���j�P+��h������V��ߴ0�3�#�5�2��a�Ͷm.O�[k�{6{��R�譔�=�$ذ�v��¢Ba�;��z����Q����-t�-��#�IE�����''c�c&��< �}*�'���?P�A��Wf��8{����B�K<����Q8�V�aNo<dm��p3q0��И"�q�ۨ����jj�����zB�����]��&`6�׎�4L�2�s���!GKe=�b�4�~�����*�dV��)�r#s��*���w��q�k�B���/&���ҰQo�7ߘ���nD����J6C`�eRـ$�HvZ��{/��H�:�LZTS����Y9�����Sz!��%K�Gh=s�RU�U@PXs_�󘖙�.XO�ץ�\%~f����l��#�>�aٜ�o���� x	%���S��j�>Da)�m�q�]�Js�^
�j]Y1ʗ�f�"����UG�Jg�Ɛ:��e�M��Ў���X7�4�= �Bٌ�$��15\U\)%pG�?vP�fmV���s��7}�n���Х�cߊ��Q���uxI+r"���	gk�&oTѿ�?��2l�߶>ɺ���X������4������TkC#�ְܨ�jR��X}�r��<X���0��W��p}Q곝�<���7L2�ZF�7;�r�}�Y��7V&����z�`]I��d�ᶎ�LF�K�H�a����O�
��&�G(�+<�1��d�$�
�C�#���8q.��q��x���*Hm��9� i�G�ʁ�GY#;x�r���dCgQ+�&�$�m�
�9+���80��Hɻ*��Ս,qS7���l=�Td��$-e����5�2l8x��e��`N��_ILS�q�M��̼����	���CtN�Q�Κ��D@���f�m1��Q l���Mӱ��nP��i�ѡp��2$��|S��J�o�o
��dn���:T	=K�q�y|2��ԙ����Ƒ �B���b�?C���
N�R��G�s\���^'����X��C�<��+Ig���$�L8�����jn�gE�o�`SDb�F��Ȉr�Bz�-��Ub

��� �/���P��j��Ę=5�S^��$ Tܙ7���������rЧ���D�!�7.��!, �!�������5-t ��.�Sֵ_�y�����<�
a�V�����&`	|��� ���w~~���r3[�g��e� C�dﺷ<Љ;�hh�'�WQwͰf;��)���z�(̝D�`@��V���z8��1 �����.�]�$0���������b6�=��Fн��[ZQo���LU��g���	3pJ�*�C>;������o�#+���X	t�����\7V��έj�٢Ӱ-��?Pp=+�C�i�#
��VK�QƮ"�!DE-cq���ˎh@�U����ɰ��7Н.���an�>���o��f�)�sx�� #:�IS��J�ʦ��Ѐ�zYw�K��m���Gt4'9��_�`�۱��W��&j��\I6�V�"*�%�*|�R�}]���4#�|6�m��O�@�LdpTN�y	���y�i�?�ƽ�SQ	�c>�Ba���,�t�U�w�j#B�,`�e��RC+��(����f �>������i��V�����b��(`�:��=�:#��� ���KL�EzU������-0B0<i��''a�CG?���B� 7������h�hO��q	��Kرb���# ?D�C0�%�s���� �㸧�^����>��_��Cs�j������/��]!��$�	��`Z	��G��m��S?�~ч ͭ��f
���:ϐ_��G"�g��'XP�O{|����q�PZڼ��t�}go@vZ=b�����t��*N�ut�����\��n�ʓ�9�Y�;:�	�9�n�y7����]b���i��n�� 2����g�T�>���`�f��ٟ���|yʶ{7؅�Qd��8��<� V!* �|�&��{5�?��
iO`ȔĠ���|`层������(Akڋ��'�*e2V�H�@䐬�	A�az�T����s<'��<�}�"����M�tzp�r��y��N�6L!6E��bŀON�ɚ���
�-�Hr��f�H���!�;���b��N�7�I��=7އ��ow�hJ^?�``�O���Y��D�����te߻���Yh��z���^�:��
ɷǁ&��|<&�{O�*�¯�U�-c0�ΝT�w�"A
�j����zG;�ol�Q�ٟ>M������F�P6�q'��z.��;�!�`�Vٖ��A5H �?��)4�X��{�]2��t�:�x��8���W�Ů�r�a��tu>����.G�vx�+��܆3�&R̮�W] �q��$er*?l��ޕ�ɟJA��_��+@�gv
l��f�i���Q�U"-���g$>[1Ȑ�O]oڔ��>���O�Ò��T��6�"���gGc�#�M��pU���""��P
C���c!C䔰'�;Ғ�r���WVVi��h�â���{Y��������A�D��>���������!d�f<ă� �j�=J*�&�f�wp�&��5���R���J��ɐw��w�Y	�ҕ���x�c4��9v4ψ	���,�+ꙏ����@��B��N�ю����cu	5�R�5��P
9���y�WwB�04h3w�Qq.�J��֏��c�A+iwס	O��5�:X��w[CI��z�R���a��������<�f��VRg�Xg�N������*���g��F0��_��D��M�O���x�i�q�=l��i^9�ae,����e���SB�)�.7a!�육�uN�з@';�Pw�ɜ�P�xx\�;��M����-��l���P�ӗ�2$�o�j�v�t�n;���Ħj�����`�V���o��T����>W�N�%���b]H��W���I �RT��ƾv_t"�p*��q�=P��cg`EJCQ�n�w-��>�c䆚�c�g�?�k�+?��|���`f�K7��E���g��7��*�ў}U+#����^X�dz/�]������vVd�˧1��j�)��o���-iԍh���̣���G��_e��A�ձ9n�hjf�w��bd�GX�H􊺙���9;�W��L�E��l���àd	6�J�W6%=��U���=�D̽��������7D���	L~� �te�5J9��$�|�q 8�����G�g:��~�k֍Ki
�,����ki;p�ɿ�W���n٠-��x(���� �C_���F���}�&D-�Fd14?�o����|���fi�[\>ĵȩV���!ٳ��Ao�A6�	��G����ѣ��w��:�ʌ��H��p8x��B�����¿�cl���/̣v��*�s�қ��!�~,ˀ>��+�Q˔�v.�C��@u �x��x�z[��[A't;����ϒ�=d�����	^E7�X�t?�C�^Sq4O���d��w�[g>�]}H����E$�4�0+����I�>G��
�>QjU�F��5pz\(��:�����Yi���(p�=��U
rW��L��^]&�K���(�CI�[�>i�kzF��;~��s�H,H����������"���N���t�nn�ڶ`����,�ƀy�ߨ��^I���ޤ+�#�ޕ[��܆������j�i�o�s��Dz���n*�Jۗ�H����?���[r���;Á!�P���q���!�Z}����BU�$nZD�
���x��|S;Eu�4\(�&S��'@�@#����!�������w��Vm@�{��~�4�锛J�!�����,����Y�V����b�vh5)[`QM"��-͑��x�:Su5�XP��ܵ�FP��I�i��w0�������Av��;S������x���h�A��>b"VX��X)v�qNCL`��z���`�Ex��t���5#2���%!8?� �\��h��	�H�x|/�fMH8i��"q��s��jpC��̀U��Zx�����Fq���(��
�ru6Pi�+���v��a���:�(`B�n��'��_�		��8��.�pkɇ�,�:ƞ�I��z���d�2=4$����M��,獢���g	���g|�f�e��$��!�xO&/؞Ҕ�I�s	e�F���#IEf'�1�b ��b�'[��j8LW�4���.���I6��@1�Ք ?l}���lT�>�޷������a��K2+�QL��o1|[���ܣ���7L�ՒBK�M[ձ'�Ôu�7�A�2˜k�}Ǜ���\ӷ�m��
Z�����`2r���|2���?�I��V�OIcN�f�@�Ua7'4���,JC�L87��ԵLt�p��� ���9�m������ۆ]�LJ:���%V@��'����������У�C�${�d$��H��9%�9����
�V�9G3DA��'�	g�+ݏF��q3{����!��oɘ�������=�Gg#As
��_t���1rTї���������Ujf��,7��	+Ǹ�J�ں�j���w�\u�ٿQAb~FB8*-��EA��6��f諸O���
�@Ы%�_���|��>�hahX��ᨐ��e	* �v����n��a�Fɳ���$yn)�����,��Ws
6S��-��)}į!�nc����O������H�R�>���2Z%��I��s�*���8��!B*�|v���p�P�]�FQj��.qd-3Z�1�
�����vX��J�Ú�B5.�Uϙ�t�^��C�(��
0/����l�i.��D��{��f_��}T��~I�*����c�fU��A)���s�+bMbj����Ӆ��9��f�3P&�A��-"l�@���nG��-���>�@K5i�{YRa���>��%��m�/�92�Y�2����<�:p�m�#W��DF��)]�]��c0�_���0�Q��P%�@���e���d�����Rfq����F�����A"<YC k��uUL� ��Tk%�5-H4�%k8�^���R�QvV�ϻp��e�wS����@4�ptE��3����d���KN������6��_�� (�JLG�bZt��P_��9-|7�5�/�]�(2���h�-?+5�Sa.�f�gh�;{?޳)8�:¡��Qt�a!��a�W&�(�v�O����m�ۭ:S-��V鼚΅#�������)<5|�-_t&b.�Zջ"��/mc�HՁ(��_�Q���݁�����|X��}���N�dd�}@q�J�l	��>W�����?m��6.����I��)]��s�����1�?��4����癵v��u�d��ma�?1@��o7�9**h��	/�Zr��2��|൤z��[pĉ�'|`�)�Ա�fΊp
yq��ZBDL���c�=A��YiFF�KP��Y��u}x�r���|V%�g���f���p(��+�V��oƻ�	#���({�5�����v5��vIS���O"�����q���K��g>Y��.L����6K�� ��=P����v��S�X��?f3���������D	@vx�����o`���h�٭�XlcS�/N�=�)� *T�}3���.z����)3ua��r�E���uhm�`x�ӧ�Q��(ɭ�`7����Q��I�B�Ö�p���c����4�*��Z��"�{�,��8�$[��_�����[Үs%E���z���v~Tm|�nÔ"c���q#vP޲�sXO�͞+��3�y�NȦ��9m1�GiYg��P��3=ۊT�掫Ar�P��K����j�/�o�b��7w!|�� �*/.��f�\��U�H��A�W��G=���	��l:K���}u���g~&����ԁ����U�����k�`�۰ᵶm����2g,f@����W y��ʂ�+��H��ԓ����6sǶ�cJ֧���J#�c���.�&3�ʚZ����׍o`v���v�y\̵�$7�zp�Y �g	�UU���t�]B����˒n\�����*�!��6���R ������ӿ��P�I5�:Zc�}]�6o-�Ŏ���NbܱNh�j�[�����s�'�oG��=�n�U|��X�B�w��:Uu4V,�L�,nd��O��U��x�&�_�m��;ߚ�;+"��T�N�=���fd�����9��ؼ��%0��p�g�\�\s�l+�AH��ë�G�Q��qj�2�W���
2fDфik�|�*���G�a����iS�)�S0�)��pl��)���g�S�����Y9����0��]�o�a��|�siC�;@s�1¯�Y���YMM����HG��)X���*lz��$�t�U��_U���,�F���>�9�fO\5,�t�2�	���2[�15܂@��xp/O��t�WᑏT"}�,
�ި��0�t�V5�C�������&F���~z{�o�5/z8f�y��C�xa��R�Rk�e����W�%g���Vo��ު&�(S��-:Y^��i�LD;��}��#9(AY�5���/��XPt@�W�%��}4v�E{u�3v��u�~������M:)uM-����s�vc�'��X�\a�����[�f1�������~��߿�EԾ�O�F�Y}�9����L�>[���^�����⏗�P�L�=l"FP'���˧���L��d*IA���H��,:M��KA��� RYc�i�0E�����g�����m��(Q�V���}ʟ.]0�5����^g;ż��F��~�P�6�_�&ͻ��e�h�P�I8�R����O��!��-�yX���������xN�Z$,��~�v�������wcr��{������p��Iv����akQ�k)�S��
�I���Z�����SgʲR�H?��Jb���.k;�*t��
u��nX[61��pYi��[��fvW΂D�c��ln,���#�Kkv^&oƂ2�o}J�s��9����+]vxo�پ5�`.�J)�H4@)��ۛ=��+�X��U�,[�H8�s�+g'�Ҷ1g�6eg�Zc�ehy]��q��X<�^TH Fu`�LYl�ߘ�V͖��j����z�$�W֤�[d����P�U��	A5��ȿ�v�jD�V�,��:�7�~Őʹ_(��ٌZX�m��c^��a�,1��w������툟����~��v;.{R�u�*��ZEF�*D�HX��e$�ɑ%�O�C�i72���,������Q����	ܶXL'����Z�S_{���b��K���5RyƴhV�UՊ���Ʒ�@0)BNZ�0��kh�x�_�L&>��pU�UwOa�L����g��F#F>�Y����&��V`0�as3��	sxW���P6l�ǠEal��Q�Ëq���e]��d})2i���Fm�<�i_e�H�qAR1�F^�kb�"g��9����%̥o�������r\G��v��"-3��K��,B\S �lp��Կ8���!��*<�\�D�J�&,Q>�6g��yvoV��u��!��1/�;��[���i���ap})��N�D��C�Z���7���Y���`����������f��n1�M�FQ�